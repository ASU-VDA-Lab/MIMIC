module fake_jpeg_1690_n_657 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_657);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_657;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_646;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_419;
wire n_378;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx10_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_3),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

BUFx6f_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_8),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_2),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_7),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_16),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_12),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_0),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_3),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_45),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_58),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g132 ( 
.A(n_59),
.Y(n_132)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_17),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_61),
.B(n_65),
.Y(n_140)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_62),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_63),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_64),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

HB1xp67_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_66),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_40),
.Y(n_67)
);

NAND2xp33_ASAP7_75t_SL g225 ( 
.A(n_67),
.B(n_121),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_68),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_69),
.Y(n_202)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_SL g200 ( 
.A(n_70),
.Y(n_200)
);

INVx11_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx11_ASAP7_75t_L g156 ( 
.A(n_71),
.Y(n_156)
);

INVx6_ASAP7_75t_SL g72 ( 
.A(n_40),
.Y(n_72)
);

BUFx4f_ASAP7_75t_SL g213 ( 
.A(n_72),
.Y(n_213)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_73),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_18),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_74),
.B(n_79),
.Y(n_141)
);

BUFx10_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g139 ( 
.A(n_75),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_37),
.B(n_15),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_76),
.B(n_78),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g207 ( 
.A(n_77),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_34),
.B(n_15),
.Y(n_78)
);

AND2x2_ASAP7_75t_SL g79 ( 
.A(n_56),
.B(n_0),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_24),
.Y(n_80)
);

INVx5_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_24),
.Y(n_81)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_82),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_83),
.Y(n_137)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_84),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

BUFx10_ASAP7_75t_L g208 ( 
.A(n_85),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

INVx4_ASAP7_75t_SL g218 ( 
.A(n_86),
.Y(n_218)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_87),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_45),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_89),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_38),
.B(n_14),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_43),
.B(n_14),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_90),
.B(n_93),
.Y(n_160)
);

INVx8_ASAP7_75t_L g91 ( 
.A(n_52),
.Y(n_91)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_91),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_52),
.Y(n_92)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_92),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_38),
.B(n_14),
.Y(n_93)
);

HB1xp67_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_94),
.Y(n_157)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_95),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_50),
.B(n_15),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_96),
.B(n_101),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_13),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_97),
.B(n_105),
.Y(n_174)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_25),
.Y(n_98)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_98),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx8_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_45),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_102),
.Y(n_164)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_45),
.Y(n_103)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_103),
.Y(n_185)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx6_ASAP7_75t_L g177 ( 
.A(n_104),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_51),
.B(n_0),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_27),
.Y(n_106)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_28),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_111),
.Y(n_189)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_22),
.Y(n_108)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_108),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_28),
.Y(n_109)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_27),
.Y(n_110)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_110),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_51),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_41),
.B(n_3),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_112),
.B(n_113),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_21),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_26),
.Y(n_114)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_114),
.Y(n_201)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_19),
.Y(n_116)
);

INVx6_ASAP7_75t_L g194 ( 
.A(n_116),
.Y(n_194)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_31),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_117),
.Y(n_147)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_26),
.Y(n_118)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_118),
.Y(n_205)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_19),
.Y(n_119)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_119),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_31),
.Y(n_120)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_120),
.Y(n_221)
);

OR2x2_ASAP7_75t_L g121 ( 
.A(n_21),
.B(n_3),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_122),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_31),
.Y(n_123)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_123),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_41),
.B(n_21),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_124),
.B(n_23),
.Y(n_212)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_125),
.Y(n_199)
);

BUFx12f_ASAP7_75t_L g126 ( 
.A(n_19),
.Y(n_126)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_126),
.Y(n_155)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_42),
.Y(n_127)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_127),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_46),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx1_ASAP7_75t_SL g129 ( 
.A(n_20),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_129),
.B(n_57),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g130 ( 
.A(n_90),
.B(n_39),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_130),
.B(n_133),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_72),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_106),
.A2(n_39),
.B1(n_55),
.B2(n_47),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_138),
.B(n_20),
.Y(n_232)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_67),
.Y(n_144)
);

INVx1_ASAP7_75t_SL g292 ( 
.A(n_144),
.Y(n_292)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_128),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g243 ( 
.A(n_153),
.Y(n_243)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_70),
.Y(n_158)
);

BUFx2_ASAP7_75t_L g298 ( 
.A(n_158),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_58),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_161),
.B(n_167),
.Y(n_252)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_71),
.Y(n_163)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_163),
.Y(n_253)
);

AOI21xp33_ASAP7_75t_L g167 ( 
.A1(n_121),
.A2(n_57),
.B(n_46),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_169),
.B(n_180),
.Y(n_257)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_110),
.Y(n_172)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_172),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_126),
.A2(n_35),
.B1(n_54),
.B2(n_44),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_173),
.A2(n_29),
.B1(n_54),
.B2(n_44),
.Y(n_259)
);

CKINVDCx14_ASAP7_75t_R g240 ( 
.A(n_175),
.Y(n_240)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_126),
.Y(n_176)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_116),
.Y(n_178)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_178),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_109),
.Y(n_180)
);

INVx4_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_182),
.Y(n_235)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_183),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_87),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_184),
.B(n_204),
.Y(n_305)
);

INVx3_ASAP7_75t_L g186 ( 
.A(n_80),
.Y(n_186)
);

BUFx12f_ASAP7_75t_L g245 ( 
.A(n_186),
.Y(n_245)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_98),
.Y(n_188)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_188),
.Y(n_226)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_115),
.Y(n_193)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_193),
.Y(n_241)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_81),
.Y(n_196)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_196),
.Y(n_250)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_95),
.Y(n_197)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_197),
.Y(n_271)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_129),
.Y(n_203)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_203),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_100),
.Y(n_204)
);

INVx11_ASAP7_75t_L g209 ( 
.A(n_85),
.Y(n_209)
);

INVx11_ASAP7_75t_L g282 ( 
.A(n_209),
.Y(n_282)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_120),
.Y(n_210)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_210),
.Y(n_289)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_104),
.Y(n_211)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_211),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_212),
.B(n_224),
.Y(n_231)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_59),
.Y(n_214)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_214),
.Y(n_297)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_123),
.Y(n_215)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_215),
.Y(n_300)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_85),
.Y(n_216)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx4_ASAP7_75t_L g220 ( 
.A(n_86),
.Y(n_220)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_220),
.Y(n_302)
);

INVx3_ASAP7_75t_L g222 ( 
.A(n_86),
.Y(n_222)
);

INVx5_ASAP7_75t_L g276 ( 
.A(n_222),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_79),
.Y(n_224)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_132),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_227),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_224),
.A2(n_79),
.B1(n_55),
.B2(n_32),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_228),
.A2(n_139),
.B(n_162),
.Y(n_325)
);

INVx6_ASAP7_75t_L g230 ( 
.A(n_132),
.Y(n_230)
);

INVx5_ASAP7_75t_L g344 ( 
.A(n_230),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_232),
.B(n_292),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_165),
.B(n_174),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g345 ( 
.A(n_233),
.B(n_238),
.Y(n_345)
);

INVx6_ASAP7_75t_L g234 ( 
.A(n_146),
.Y(n_234)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_234),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g236 ( 
.A1(n_173),
.A2(n_64),
.B1(n_99),
.B2(n_92),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_236),
.A2(n_199),
.B1(n_208),
.B2(n_291),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_140),
.B(n_32),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_146),
.Y(n_239)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_239),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_147),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_242),
.B(n_247),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_140),
.B(n_23),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_244),
.B(n_251),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_198),
.B(n_33),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_191),
.A2(n_33),
.B1(n_47),
.B2(n_35),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_248),
.A2(n_277),
.B1(n_278),
.B2(n_280),
.Y(n_348)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_159),
.Y(n_249)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_198),
.B(n_29),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g254 ( 
.A(n_213),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_254),
.B(n_256),
.Y(n_349)
);

INVx8_ASAP7_75t_L g255 ( 
.A(n_194),
.Y(n_255)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_255),
.Y(n_312)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_175),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_225),
.B(n_125),
.Y(n_258)
);

AND2x4_ASAP7_75t_L g359 ( 
.A(n_258),
.B(n_266),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_259),
.A2(n_260),
.B1(n_263),
.B2(n_265),
.Y(n_333)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_157),
.A2(n_29),
.B1(n_54),
.B2(n_44),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_143),
.B(n_30),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_261),
.B(n_262),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_160),
.B(n_143),
.Y(n_262)
);

AOI22xp33_ASAP7_75t_SL g263 ( 
.A1(n_189),
.A2(n_30),
.B1(n_20),
.B2(n_91),
.Y(n_263)
);

A2O1A1Ixp33_ASAP7_75t_L g264 ( 
.A1(n_141),
.A2(n_30),
.B(n_75),
.C(n_19),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g361 ( 
.A1(n_264),
.A2(n_237),
.B(n_243),
.Y(n_361)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_189),
.A2(n_77),
.B1(n_69),
.B2(n_68),
.Y(n_265)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_135),
.B(n_149),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_160),
.B(n_4),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_270),
.B(n_274),
.Y(n_313)
);

CKINVDCx12_ASAP7_75t_R g272 ( 
.A(n_213),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_272),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_152),
.Y(n_273)
);

INVx8_ASAP7_75t_L g314 ( 
.A(n_273),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_170),
.B(n_63),
.Y(n_274)
);

CKINVDCx12_ASAP7_75t_R g275 ( 
.A(n_171),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_275),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_201),
.A2(n_19),
.B1(n_53),
.B2(n_75),
.Y(n_277)
);

AOI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_205),
.A2(n_53),
.B1(n_5),
.B2(n_6),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_170),
.B(n_4),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_279),
.B(n_281),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_206),
.A2(n_53),
.B1(n_6),
.B2(n_7),
.Y(n_280)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_187),
.Y(n_281)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_164),
.Y(n_283)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_283),
.Y(n_318)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_152),
.Y(n_284)
);

INVx8_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_141),
.B(n_195),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_285),
.B(n_200),
.Y(n_319)
);

INVx8_ASAP7_75t_L g287 ( 
.A(n_219),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_287),
.Y(n_354)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_137),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_290),
.A2(n_294),
.B1(n_307),
.B2(n_218),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_223),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_291),
.A2(n_207),
.B1(n_202),
.B2(n_131),
.Y(n_317)
);

INVx5_ASAP7_75t_L g293 ( 
.A(n_181),
.Y(n_293)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_293),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_148),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_294)
);

INVx6_ASAP7_75t_L g295 ( 
.A(n_179),
.Y(n_295)
);

INVx2_ASAP7_75t_L g350 ( 
.A(n_295),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_171),
.B(n_9),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_296),
.B(n_303),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_179),
.Y(n_299)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_151),
.B(n_9),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_136),
.B(n_12),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_304),
.B(n_218),
.Y(n_340)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_187),
.Y(n_306)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_306),
.Y(n_330)
);

OAI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_223),
.A2(n_168),
.B1(n_202),
.B2(n_207),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_310),
.B(n_361),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_317),
.A2(n_323),
.B1(n_329),
.B2(n_337),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_319),
.B(n_325),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_258),
.A2(n_154),
.B(n_155),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_320),
.A2(n_365),
.B(n_298),
.Y(n_376)
);

OAI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_232),
.A2(n_150),
.B1(n_156),
.B2(n_185),
.Y(n_323)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_328),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_228),
.A2(n_190),
.B1(n_177),
.B2(n_145),
.Y(n_329)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_297),
.Y(n_331)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_331),
.Y(n_390)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_334),
.Y(n_400)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_266),
.Y(n_336)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_336),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_240),
.A2(n_221),
.B1(n_134),
.B2(n_181),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_340),
.B(n_355),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g341 ( 
.A1(n_258),
.A2(n_134),
.B1(n_217),
.B2(n_166),
.Y(n_341)
);

AO22x1_ASAP7_75t_L g391 ( 
.A1(n_341),
.A2(n_282),
.B1(n_293),
.B2(n_226),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_285),
.B(n_139),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_342),
.B(n_343),
.C(n_356),
.Y(n_371)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_231),
.B(n_200),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_264),
.B(n_217),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_346),
.B(n_362),
.Y(n_368)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_257),
.Y(n_347)
);

INVx2_ASAP7_75t_SL g378 ( 
.A(n_347),
.Y(n_378)
);

OAI22xp33_ASAP7_75t_SL g351 ( 
.A1(n_252),
.A2(n_208),
.B1(n_192),
.B2(n_142),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_351),
.B(n_241),
.Y(n_392)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_305),
.Y(n_353)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_353),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_246),
.B(n_208),
.C(n_199),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_243),
.Y(n_357)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_357),
.Y(n_381)
);

INVx2_ASAP7_75t_L g358 ( 
.A(n_300),
.Y(n_358)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_358),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_360),
.A2(n_282),
.B1(n_239),
.B2(n_273),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_250),
.B(n_271),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_300),
.Y(n_363)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

OA22x2_ASAP7_75t_L g364 ( 
.A1(n_236),
.A2(n_268),
.B1(n_229),
.B2(n_250),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_367),
.Y(n_413)
);

AOI21xp5_ASAP7_75t_L g365 ( 
.A1(n_235),
.A2(n_226),
.B(n_241),
.Y(n_365)
);

INVx2_ASAP7_75t_L g366 ( 
.A(n_229),
.Y(n_366)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_366),
.Y(n_408)
);

NAND2xp33_ASAP7_75t_SL g367 ( 
.A(n_268),
.B(n_298),
.Y(n_367)
);

INVx13_ASAP7_75t_L g369 ( 
.A(n_315),
.Y(n_369)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_369),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_309),
.B(n_292),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_372),
.B(n_388),
.Y(n_425)
);

INVx13_ASAP7_75t_L g373 ( 
.A(n_327),
.Y(n_373)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_373),
.Y(n_440)
);

INVx13_ASAP7_75t_L g375 ( 
.A(n_367),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_375),
.Y(n_453)
);

AND2x2_ASAP7_75t_L g445 ( 
.A(n_376),
.B(n_391),
.Y(n_445)
);

INVxp67_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

BUFx2_ASAP7_75t_L g451 ( 
.A(n_380),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_346),
.B(n_271),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_382),
.B(n_397),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_312),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_401),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_333),
.A2(n_287),
.B1(n_255),
.B2(n_230),
.Y(n_384)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_384),
.A2(n_386),
.B1(n_410),
.B2(n_317),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_360),
.A2(n_295),
.B1(n_284),
.B2(n_234),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_316),
.B(n_235),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_345),
.B(n_267),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g444 ( 
.A(n_389),
.B(n_399),
.Y(n_444)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_392),
.A2(n_382),
.B1(n_368),
.B2(n_406),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_343),
.B(n_286),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_393),
.B(n_359),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_330),
.Y(n_394)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_394),
.Y(n_420)
);

INVx13_ASAP7_75t_L g396 ( 
.A(n_366),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g441 ( 
.A1(n_396),
.A2(n_403),
.B1(n_354),
.B2(n_335),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_342),
.B(n_289),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_321),
.B(n_267),
.Y(n_399)
);

AND2x6_ASAP7_75t_L g401 ( 
.A(n_361),
.B(n_276),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_308),
.B(n_318),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g455 ( 
.A(n_402),
.B(n_409),
.Y(n_455)
);

INVx13_ASAP7_75t_L g403 ( 
.A(n_365),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_332),
.B(n_289),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g434 ( 
.A(n_404),
.B(n_405),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_311),
.B(n_286),
.Y(n_405)
);

BUFx16f_ASAP7_75t_L g407 ( 
.A(n_354),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_407),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_313),
.B(n_276),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_320),
.Y(n_411)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_411),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_349),
.B(n_301),
.Y(n_412)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_412),
.B(n_414),
.Y(n_430)
);

INVxp67_ASAP7_75t_L g414 ( 
.A(n_356),
.Y(n_414)
);

AND2x6_ASAP7_75t_L g415 ( 
.A(n_325),
.B(n_245),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_393),
.Y(n_452)
);

A2O1A1Ixp33_ASAP7_75t_SL g416 ( 
.A1(n_413),
.A2(n_374),
.B(n_403),
.C(n_368),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_422),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_376),
.A2(n_355),
.B(n_348),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_417),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g419 ( 
.A1(n_411),
.A2(n_355),
.B(n_341),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g464 ( 
.A(n_419),
.B(n_428),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_L g422 ( 
.A1(n_379),
.A2(n_364),
.B(n_336),
.C(n_334),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_369),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_423),
.B(n_443),
.Y(n_471)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_424),
.B(n_431),
.Y(n_478)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_377),
.Y(n_427)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_427),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_429),
.B(n_397),
.Y(n_459)
);

NOR2x1_ASAP7_75t_L g431 ( 
.A(n_374),
.B(n_359),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_377),
.Y(n_432)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_432),
.Y(n_458)
);

AOI22xp33_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_364),
.B1(n_319),
.B2(n_335),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g484 ( 
.A1(n_433),
.A2(n_454),
.B1(n_408),
.B2(n_381),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_371),
.B(n_359),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_436),
.B(n_439),
.C(n_429),
.Y(n_472)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_390),
.Y(n_437)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_437),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_374),
.A2(n_414),
.B1(n_385),
.B2(n_413),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_438),
.A2(n_449),
.B1(n_410),
.B2(n_391),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_371),
.B(n_359),
.Y(n_439)
);

INVx13_ASAP7_75t_L g491 ( 
.A(n_441),
.Y(n_491)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_390),
.Y(n_442)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_442),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_386),
.A2(n_329),
.B1(n_337),
.B2(n_364),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g465 ( 
.A1(n_446),
.A2(n_400),
.B1(n_406),
.B2(n_405),
.Y(n_465)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_398),
.Y(n_447)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_SL g448 ( 
.A1(n_379),
.A2(n_310),
.B(n_363),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_448),
.B(n_395),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g449 ( 
.A1(n_385),
.A2(n_312),
.B1(n_338),
.B2(n_339),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_452),
.B(n_395),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_SL g454 ( 
.A1(n_384),
.A2(n_339),
.B1(n_338),
.B2(n_358),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_L g456 ( 
.A1(n_417),
.A2(n_413),
.B1(n_380),
.B2(n_401),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_L g512 ( 
.A1(n_456),
.A2(n_460),
.B1(n_465),
.B2(n_474),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_459),
.B(n_472),
.C(n_439),
.Y(n_495)
);

OAI22xp5_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_446),
.B1(n_421),
.B2(n_452),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_SL g510 ( 
.A1(n_461),
.A2(n_416),
.B1(n_422),
.B2(n_442),
.Y(n_510)
);

AND2x2_ASAP7_75t_L g520 ( 
.A(n_463),
.B(n_449),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g466 ( 
.A(n_440),
.B(n_409),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_SL g517 ( 
.A(n_466),
.B(n_477),
.Y(n_517)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_438),
.Y(n_470)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_470),
.Y(n_515)
);

CKINVDCx20_ASAP7_75t_R g493 ( 
.A(n_471),
.Y(n_493)
);

OAI22xp5_ASAP7_75t_SL g474 ( 
.A1(n_426),
.A2(n_400),
.B1(n_415),
.B2(n_378),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_476),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_378),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g479 ( 
.A(n_455),
.B(n_378),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_479),
.B(n_482),
.Y(n_498)
);

INVx3_ASAP7_75t_L g480 ( 
.A(n_420),
.Y(n_480)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_480),
.Y(n_494)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_427),
.Y(n_481)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_481),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_451),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_383),
.Y(n_483)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_483),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_445),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_444),
.B(n_404),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_485),
.B(n_434),
.Y(n_497)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_425),
.Y(n_486)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_486),
.B(n_492),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_426),
.B(n_370),
.Y(n_487)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_487),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_434),
.B(n_370),
.Y(n_488)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_488),
.Y(n_523)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_432),
.Y(n_489)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_489),
.Y(n_525)
);

AOI22xp5_ASAP7_75t_L g490 ( 
.A1(n_445),
.A2(n_391),
.B1(n_375),
.B2(n_381),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_SL g500 ( 
.A1(n_490),
.A2(n_445),
.B1(n_419),
.B2(n_453),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_420),
.B(n_324),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_495),
.B(n_527),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_497),
.B(n_499),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g499 ( 
.A(n_483),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_500),
.A2(n_501),
.B1(n_520),
.B2(n_473),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_472),
.B(n_436),
.C(n_431),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g534 ( 
.A(n_502),
.B(n_507),
.C(n_464),
.Y(n_534)
);

OR2x2_ASAP7_75t_L g504 ( 
.A(n_475),
.B(n_435),
.Y(n_504)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_504),
.Y(n_528)
);

CKINVDCx16_ASAP7_75t_R g505 ( 
.A(n_465),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_505),
.B(n_526),
.Y(n_545)
);

OAI21xp5_ASAP7_75t_L g506 ( 
.A1(n_469),
.A2(n_416),
.B(n_453),
.Y(n_506)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_506),
.A2(n_521),
.B(n_524),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_459),
.B(n_448),
.C(n_435),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_482),
.B(n_450),
.Y(n_508)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_508),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_486),
.B(n_418),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g550 ( 
.A(n_509),
.B(n_514),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_SL g554 ( 
.A1(n_510),
.A2(n_491),
.B1(n_350),
.B2(n_344),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_485),
.B(n_328),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_488),
.B(n_487),
.Y(n_516)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_516),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_447),
.Y(n_518)
);

INVxp67_ASAP7_75t_SL g553 ( 
.A(n_518),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g521 ( 
.A1(n_469),
.A2(n_416),
.B(n_437),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_468),
.B(n_408),
.Y(n_522)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_522),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_475),
.A2(n_407),
.B(n_387),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_478),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_474),
.B(n_387),
.Y(n_527)
);

INVxp67_ASAP7_75t_L g529 ( 
.A(n_518),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g561 ( 
.A(n_529),
.B(n_531),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_521),
.A2(n_456),
.B(n_464),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_495),
.B(n_476),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g559 ( 
.A(n_532),
.B(n_540),
.Y(n_559)
);

AOI21xp5_ASAP7_75t_L g533 ( 
.A1(n_501),
.A2(n_478),
.B(n_460),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_533),
.B(n_549),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g578 ( 
.A(n_534),
.B(n_548),
.Y(n_578)
);

OA21x2_ASAP7_75t_L g535 ( 
.A1(n_504),
.A2(n_464),
.B(n_463),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_535),
.B(n_541),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_502),
.B(n_470),
.C(n_490),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g565 ( 
.A(n_536),
.B(n_537),
.C(n_544),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_507),
.B(n_468),
.C(n_473),
.Y(n_537)
);

OAI22xp5_ASAP7_75t_SL g580 ( 
.A1(n_539),
.A2(n_513),
.B1(n_523),
.B2(n_508),
.Y(n_580)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_512),
.B(n_458),
.Y(n_540)
);

AND2x6_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_407),
.Y(n_541)
);

AO22x1_ASAP7_75t_L g543 ( 
.A1(n_500),
.A2(n_458),
.B1(n_489),
.B2(n_481),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_543),
.B(n_499),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_505),
.B(n_467),
.C(n_457),
.Y(n_544)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_512),
.B(n_467),
.C(n_457),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_546),
.B(n_552),
.C(n_494),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_510),
.B(n_462),
.Y(n_548)
);

NOR3xp33_ASAP7_75t_SL g549 ( 
.A(n_503),
.B(n_462),
.C(n_373),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_503),
.A2(n_493),
.B1(n_517),
.B2(n_526),
.Y(n_551)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_551),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_497),
.B(n_331),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g562 ( 
.A1(n_554),
.A2(n_515),
.B1(n_520),
.B2(n_498),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_SL g557 ( 
.A(n_506),
.B(n_491),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_557),
.B(n_515),
.Y(n_566)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_545),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g582 ( 
.A(n_560),
.B(n_552),
.Y(n_582)
);

OAI22xp5_ASAP7_75t_SL g585 ( 
.A1(n_562),
.A2(n_570),
.B1(n_530),
.B2(n_542),
.Y(n_585)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_538),
.Y(n_564)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_564),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_SL g600 ( 
.A1(n_566),
.A2(n_525),
.B1(n_496),
.B2(n_522),
.Y(n_600)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_567),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g583 ( 
.A(n_568),
.B(n_576),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_529),
.B(n_498),
.Y(n_569)
);

CKINVDCx14_ASAP7_75t_R g592 ( 
.A(n_569),
.Y(n_592)
);

AOI22xp5_ASAP7_75t_L g570 ( 
.A1(n_540),
.A2(n_511),
.B1(n_520),
.B2(n_527),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_549),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_L g588 ( 
.A(n_571),
.B(n_575),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g572 ( 
.A(n_550),
.B(n_493),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_L g597 ( 
.A(n_572),
.B(n_573),
.C(n_579),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_556),
.B(n_517),
.Y(n_573)
);

FAx1_ASAP7_75t_SL g575 ( 
.A(n_534),
.B(n_504),
.CI(n_524),
.CON(n_575),
.SN(n_575)
);

AOI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_528),
.A2(n_511),
.B(n_523),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_553),
.Y(n_577)
);

NOR3xp33_ASAP7_75t_L g589 ( 
.A(n_577),
.B(n_544),
.C(n_546),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g579 ( 
.A(n_537),
.B(n_494),
.Y(n_579)
);

AOI22xp5_ASAP7_75t_L g593 ( 
.A1(n_580),
.A2(n_543),
.B1(n_570),
.B2(n_548),
.Y(n_593)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_547),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g598 ( 
.A(n_581),
.Y(n_598)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_582),
.Y(n_612)
);

MAJIxp5_ASAP7_75t_L g584 ( 
.A(n_565),
.B(n_559),
.C(n_578),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_584),
.B(n_590),
.Y(n_608)
);

AOI22xp5_ASAP7_75t_L g610 ( 
.A1(n_585),
.A2(n_587),
.B1(n_594),
.B2(n_564),
.Y(n_610)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_574),
.A2(n_513),
.B1(n_555),
.B2(n_541),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_589),
.B(n_593),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g590 ( 
.A(n_567),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_563),
.A2(n_531),
.B1(n_535),
.B2(n_516),
.Y(n_594)
);

AOI22xp5_ASAP7_75t_L g595 ( 
.A1(n_563),
.A2(n_535),
.B1(n_536),
.B2(n_532),
.Y(n_595)
);

OAI22xp5_ASAP7_75t_L g604 ( 
.A1(n_595),
.A2(n_561),
.B1(n_558),
.B2(n_562),
.Y(n_604)
);

BUFx12_ASAP7_75t_L g596 ( 
.A(n_568),
.Y(n_596)
);

CKINVDCx20_ASAP7_75t_R g603 ( 
.A(n_596),
.Y(n_603)
);

MAJIxp5_ASAP7_75t_L g599 ( 
.A(n_565),
.B(n_557),
.C(n_525),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g609 ( 
.A(n_599),
.B(n_600),
.Y(n_609)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_584),
.B(n_559),
.C(n_578),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_601),
.B(n_602),
.Y(n_622)
);

MAJIxp5_ASAP7_75t_L g602 ( 
.A(n_599),
.B(n_561),
.C(n_580),
.Y(n_602)
);

AOI22xp5_ASAP7_75t_L g621 ( 
.A1(n_604),
.A2(n_592),
.B1(n_586),
.B2(n_598),
.Y(n_621)
);

INVxp33_ASAP7_75t_L g605 ( 
.A(n_597),
.Y(n_605)
);

OR2x2_ASAP7_75t_L g618 ( 
.A(n_605),
.B(n_610),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g606 ( 
.A(n_595),
.B(n_581),
.C(n_569),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_606),
.B(n_607),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_583),
.B(n_576),
.C(n_571),
.Y(n_607)
);

NOR2xp67_ASAP7_75t_L g611 ( 
.A(n_588),
.B(n_496),
.Y(n_611)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_611),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_587),
.B(n_575),
.Y(n_613)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_613),
.Y(n_625)
);

XOR2xp5_ASAP7_75t_L g615 ( 
.A(n_594),
.B(n_575),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g629 ( 
.A(n_615),
.B(n_616),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_588),
.B(n_326),
.Y(n_616)
);

MAJIxp5_ASAP7_75t_L g617 ( 
.A(n_585),
.B(n_350),
.C(n_352),
.Y(n_617)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_617),
.B(n_602),
.C(n_603),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g620 ( 
.A1(n_614),
.A2(n_591),
.B(n_593),
.Y(n_620)
);

OR2x2_ASAP7_75t_L g638 ( 
.A(n_620),
.B(n_322),
.Y(n_638)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_621),
.Y(n_633)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_623),
.Y(n_639)
);

OAI22xp5_ASAP7_75t_SL g624 ( 
.A1(n_605),
.A2(n_600),
.B1(n_598),
.B2(n_596),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_624),
.A2(n_615),
.B1(n_614),
.B2(n_610),
.Y(n_631)
);

MAJIxp5_ASAP7_75t_L g627 ( 
.A(n_601),
.B(n_596),
.C(n_352),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_627),
.B(n_628),
.Y(n_637)
);

MAJIxp5_ASAP7_75t_L g628 ( 
.A(n_608),
.B(n_322),
.C(n_227),
.Y(n_628)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_607),
.B(n_326),
.Y(n_630)
);

NOR2xp33_ASAP7_75t_SL g636 ( 
.A(n_630),
.B(n_344),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_631),
.B(n_634),
.Y(n_643)
);

INVxp67_ASAP7_75t_L g632 ( 
.A(n_629),
.Y(n_632)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_632),
.B(n_636),
.Y(n_641)
);

XNOR2xp5_ASAP7_75t_L g634 ( 
.A(n_627),
.B(n_606),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g635 ( 
.A1(n_625),
.A2(n_612),
.B1(n_609),
.B2(n_617),
.Y(n_635)
);

XNOR2xp5_ASAP7_75t_L g646 ( 
.A(n_635),
.B(n_640),
.Y(n_646)
);

XOR2xp5_ASAP7_75t_L g644 ( 
.A(n_638),
.B(n_628),
.Y(n_644)
);

OAI21xp5_ASAP7_75t_L g640 ( 
.A1(n_618),
.A2(n_314),
.B(n_396),
.Y(n_640)
);

MAJIxp5_ASAP7_75t_L g642 ( 
.A(n_639),
.B(n_622),
.C(n_626),
.Y(n_642)
);

A2O1A1O1Ixp25_ASAP7_75t_L g648 ( 
.A1(n_642),
.A2(n_619),
.B(n_621),
.C(n_632),
.D(n_618),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_SL g647 ( 
.A1(n_644),
.A2(n_623),
.B(n_637),
.Y(n_647)
);

NAND2x1p5_ASAP7_75t_R g645 ( 
.A(n_633),
.B(n_620),
.Y(n_645)
);

AO21x1_ASAP7_75t_L g650 ( 
.A1(n_645),
.A2(n_301),
.B(n_302),
.Y(n_650)
);

OR2x2_ASAP7_75t_L g652 ( 
.A(n_647),
.B(n_648),
.Y(n_652)
);

OAI21xp5_ASAP7_75t_SL g649 ( 
.A1(n_643),
.A2(n_638),
.B(n_299),
.Y(n_649)
);

AOI322xp5_ASAP7_75t_L g651 ( 
.A1(n_649),
.A2(n_650),
.A3(n_641),
.B1(n_245),
.B2(n_645),
.C1(n_314),
.C2(n_646),
.Y(n_651)
);

OA21x2_ASAP7_75t_L g653 ( 
.A1(n_651),
.A2(n_269),
.B(n_253),
.Y(n_653)
);

OR2x2_ASAP7_75t_L g654 ( 
.A(n_653),
.B(n_644),
.Y(n_654)
);

XOR2xp5_ASAP7_75t_L g655 ( 
.A(n_654),
.B(n_652),
.Y(n_655)
);

NOR4xp25_ASAP7_75t_L g656 ( 
.A(n_655),
.B(n_302),
.C(n_245),
.D(n_253),
.Y(n_656)
);

XNOR2xp5_ASAP7_75t_L g657 ( 
.A(n_656),
.B(n_269),
.Y(n_657)
);


endmodule