module fake_jpeg_15719_n_85 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_85);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_85;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_82;

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_8),
.B(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_19),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_18),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_35),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_48),
.Y(n_59)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_46),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_0),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_53),
.B(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_41),
.B(n_1),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_34),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_3),
.Y(n_65)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_61),
.B(n_6),
.Y(n_68)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_62),
.Y(n_67)
);

O2A1O1Ixp33_ASAP7_75t_L g63 ( 
.A1(n_60),
.A2(n_39),
.B(n_43),
.C(n_45),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_58),
.B(n_42),
.C(n_4),
.Y(n_64)
);

HAxp5_ASAP7_75t_SL g70 ( 
.A(n_64),
.B(n_7),
.CON(n_70),
.SN(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_59),
.B1(n_55),
.B2(n_10),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_69),
.B(n_12),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_9),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

OA21x2_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_75),
.B(n_71),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_66),
.Y(n_75)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_76),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_77),
.B1(n_15),
.B2(n_17),
.Y(n_79)
);

NOR3xp33_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_13),
.C(n_20),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_80),
.B(n_23),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_24),
.C(n_25),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_82),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g84 ( 
.A1(n_83),
.A2(n_27),
.A3(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_31),
.Y(n_85)
);


endmodule