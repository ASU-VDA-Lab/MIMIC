module fake_aes_7264_n_26 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_8, n_0, n_26);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_8;
input n_0;
output n_26;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
INVx1_ASAP7_75t_L g10 ( .A(n_9), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_6), .Y(n_11) );
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
CKINVDCx20_ASAP7_75t_R g14 ( .A(n_2), .Y(n_14) );
AOI21xp5_ASAP7_75t_L g15 ( .A1(n_10), .A2(n_5), .B(n_8), .Y(n_15) );
AOI21x1_ASAP7_75t_L g16 ( .A1(n_11), .A2(n_0), .B(n_3), .Y(n_16) );
A2O1A1Ixp33_ASAP7_75t_SL g17 ( .A1(n_13), .A2(n_4), .B(n_12), .C(n_14), .Y(n_17) );
CKINVDCx20_ASAP7_75t_R g18 ( .A(n_15), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_16), .B(n_13), .Y(n_19) );
HB1xp67_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NOR2x1_ASAP7_75t_L g22 ( .A(n_21), .B(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
BUFx2_ASAP7_75t_L g25 ( .A(n_23), .Y(n_25) );
AOI222xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_4), .B1(n_13), .B2(n_17), .C1(n_19), .C2(n_24), .Y(n_26) );
endmodule