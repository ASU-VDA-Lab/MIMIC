module real_aes_16653_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_254;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_260;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1382;
wire n_1225;
wire n_875;
wire n_951;
wire n_1199;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_805;
wire n_619;
wire n_1095;
wire n_1284;
wire n_1250;
wire n_360;
wire n_859;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_1351;
wire n_972;
wire n_1209;
wire n_411;
wire n_498;
wire n_1397;
wire n_765;
wire n_648;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_712;
wire n_266;
wire n_422;
wire n_861;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_258;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_337;
wire n_264;
wire n_480;
wire n_684;
wire n_1178;
wire n_821;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_635;
wire n_792;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1368;
wire n_994;
wire n_384;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_746;
wire n_656;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_651;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1386;
wire n_406;
wire n_617;
wire n_1404;
wire n_733;
wire n_402;
wire n_602;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_255;
wire n_286;
wire n_1011;
wire n_416;
wire n_895;
wire n_799;
wire n_490;
wire n_261;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_557;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_701;
wire n_809;
wire n_520;
wire n_679;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_689;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1431;
wire n_721;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1162;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_253;
wire n_459;
wire n_1172;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_257;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_773;
wire n_353;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1373;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_467;
wire n_1213;
wire n_1053;
wire n_263;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_324;
wire n_664;
wire n_367;
wire n_267;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1414;
wire n_1241;
wire n_502;
wire n_434;
wire n_769;
wire n_250;
wire n_1212;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_251;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1028;
wire n_366;
wire n_1083;
wire n_727;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_262;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_252;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_1343;
wire n_719;
wire n_1156;
wire n_988;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1151;
wire n_1254;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_319;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_466;
wire n_1049;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_655;
wire n_654;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_969;
wire n_256;
wire n_1009;
wire n_1202;
wire n_302;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_385;
wire n_275;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1043;
wire n_435;
wire n_511;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1087;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_338;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_803;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1352;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1369;
wire n_1097;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_342;
wire n_348;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_259;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AOI22xp33_ASAP7_75t_SL g816 ( .A1(n_0), .A2(n_58), .B1(n_401), .B2(n_813), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_0), .A2(n_231), .B1(n_585), .B2(n_611), .Y(n_829) );
AOI22xp33_ASAP7_75t_L g1143 ( .A1(n_1), .A2(n_5), .B1(n_1144), .B2(n_1147), .Y(n_1143) );
AOI22xp33_ASAP7_75t_L g1345 ( .A1(n_2), .A2(n_181), .B1(n_585), .B2(n_638), .Y(n_1345) );
AOI22xp33_ASAP7_75t_L g1363 ( .A1(n_2), .A2(n_49), .B1(n_546), .B2(n_1364), .Y(n_1363) );
INVx1_ASAP7_75t_L g821 ( .A(n_3), .Y(n_821) );
OAI211xp5_ASAP7_75t_L g909 ( .A1(n_4), .A2(n_910), .B(n_911), .C(n_921), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g931 ( .A(n_4), .B(n_525), .Y(n_931) );
AOI22xp33_ASAP7_75t_SL g1418 ( .A1(n_6), .A2(n_234), .B1(n_585), .B2(n_1419), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g1426 ( .A1(n_6), .A2(n_161), .B1(n_1081), .B2(n_1427), .Y(n_1426) );
INVx1_ASAP7_75t_L g1354 ( .A(n_7), .Y(n_1354) );
OAI22xp33_ASAP7_75t_L g1369 ( .A1(n_7), .A2(n_52), .B1(n_671), .B2(n_892), .Y(n_1369) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_8), .A2(n_59), .B1(n_813), .B2(n_1081), .Y(n_1080) );
AOI22xp33_ASAP7_75t_L g1105 ( .A1(n_8), .A2(n_39), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g637 ( .A1(n_9), .A2(n_193), .B1(n_585), .B2(n_638), .Y(n_637) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_9), .A2(n_236), .B1(n_531), .B2(n_546), .Y(n_662) );
AOI22xp33_ASAP7_75t_SL g1414 ( .A1(n_10), .A2(n_214), .B1(n_583), .B2(n_585), .Y(n_1414) );
AOI22xp33_ASAP7_75t_L g1429 ( .A1(n_10), .A2(n_194), .B1(n_380), .B2(n_1430), .Y(n_1429) );
INVx1_ASAP7_75t_L g971 ( .A(n_11), .Y(n_971) );
AO22x1_ASAP7_75t_L g994 ( .A1(n_11), .A2(n_120), .B1(n_577), .B2(n_918), .Y(n_994) );
INVx1_ASAP7_75t_L g259 ( .A(n_12), .Y(n_259) );
AND2x2_ASAP7_75t_L g311 ( .A(n_12), .B(n_203), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g330 ( .A(n_12), .B(n_269), .Y(n_330) );
AND2x2_ASAP7_75t_L g344 ( .A(n_12), .B(n_345), .Y(n_344) );
INVx1_ASAP7_75t_L g979 ( .A(n_13), .Y(n_979) );
AOI22xp33_ASAP7_75t_L g993 ( .A1(n_13), .A2(n_81), .B1(n_484), .B2(n_915), .Y(n_993) );
XNOR2xp5_ASAP7_75t_L g1333 ( .A(n_14), .B(n_1334), .Y(n_1333) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_15), .A2(n_121), .B1(n_390), .B2(n_810), .C(n_815), .Y(n_814) );
AOI22xp33_ASAP7_75t_L g832 ( .A1(n_15), .A2(n_44), .B1(n_585), .B2(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g1140 ( .A(n_16), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1142 ( .A(n_16), .B(n_86), .Y(n_1142) );
AND2x2_ASAP7_75t_L g1148 ( .A(n_16), .B(n_1146), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g553 ( .A(n_17), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g653 ( .A1(n_18), .A2(n_73), .B1(n_525), .B2(n_654), .Y(n_653) );
CKINVDCx5p33_ASAP7_75t_R g807 ( .A(n_19), .Y(n_807) );
INVx1_ASAP7_75t_L g561 ( .A(n_20), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g1165 ( .A1(n_21), .A2(n_207), .B1(n_1144), .B2(n_1147), .Y(n_1165) );
OAI211xp5_ASAP7_75t_L g922 ( .A1(n_22), .A2(n_603), .B(n_712), .C(n_923), .Y(n_922) );
INVx1_ASAP7_75t_L g952 ( .A(n_22), .Y(n_952) );
OAI22xp5_ASAP7_75t_L g1357 ( .A1(n_23), .A2(n_79), .B1(n_525), .B2(n_654), .Y(n_1357) );
OAI22xp5_ASAP7_75t_L g742 ( .A1(n_24), .A2(n_240), .B1(n_743), .B2(n_747), .Y(n_742) );
OAI22xp33_ASAP7_75t_L g781 ( .A1(n_24), .A2(n_240), .B1(n_782), .B2(n_785), .Y(n_781) );
AOI22xp5_ASAP7_75t_L g1153 ( .A1(n_25), .A2(n_239), .B1(n_1137), .B2(n_1154), .Y(n_1153) );
NAND2xp5_ASAP7_75t_SL g1035 ( .A(n_26), .B(n_1036), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_26), .A2(n_133), .B1(n_378), .B2(n_1058), .Y(n_1057) );
XNOR2xp5_ASAP7_75t_L g622 ( .A(n_27), .B(n_623), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g1040 ( .A1(n_28), .A2(n_133), .B1(n_577), .B2(n_584), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_28), .A2(n_224), .B1(n_378), .B2(n_533), .Y(n_1052) );
INVx1_ASAP7_75t_L g1340 ( .A(n_29), .Y(n_1340) );
XOR2x2_ASAP7_75t_L g840 ( .A(n_30), .B(n_841), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g644 ( .A1(n_31), .A2(n_141), .B1(n_585), .B2(n_645), .Y(n_644) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_31), .A2(n_101), .B1(n_401), .B2(n_572), .Y(n_665) );
INVx1_ASAP7_75t_L g445 ( .A(n_32), .Y(n_445) );
AO22x1_ASAP7_75t_L g1162 ( .A1(n_32), .A2(n_40), .B1(n_1137), .B2(n_1141), .Y(n_1162) );
AOI22xp5_ASAP7_75t_L g1158 ( .A1(n_33), .A2(n_219), .B1(n_1144), .B2(n_1147), .Y(n_1158) );
AOI22xp33_ASAP7_75t_L g912 ( .A1(n_34), .A2(n_51), .B1(n_584), .B2(n_913), .Y(n_912) );
AOI22xp33_ASAP7_75t_SL g934 ( .A1(n_34), .A2(n_245), .B1(n_380), .B2(n_935), .Y(n_934) );
AOI22xp33_ASAP7_75t_SL g1086 ( .A1(n_35), .A2(n_110), .B1(n_539), .B2(n_1087), .Y(n_1086) );
INVxp67_ASAP7_75t_SL g1121 ( .A(n_35), .Y(n_1121) );
INVx1_ASAP7_75t_L g1383 ( .A(n_36), .Y(n_1383) );
INVx1_ASAP7_75t_L g368 ( .A(n_37), .Y(n_368) );
INVx1_ASAP7_75t_L g376 ( .A(n_37), .Y(n_376) );
INVx1_ASAP7_75t_L g1023 ( .A(n_38), .Y(n_1023) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_39), .A2(n_113), .B1(n_813), .B2(n_1084), .Y(n_1083) );
INVx1_ASAP7_75t_L g253 ( .A(n_41), .Y(n_253) );
INVx2_ASAP7_75t_L g388 ( .A(n_42), .Y(n_388) );
INVx1_ASAP7_75t_L g1013 ( .A(n_43), .Y(n_1013) );
AOI221xp5_ASAP7_75t_L g809 ( .A1(n_44), .A2(n_55), .B1(n_669), .B2(n_810), .C(n_811), .Y(n_809) );
AOI221xp5_ASAP7_75t_L g847 ( .A1(n_45), .A2(n_98), .B1(n_642), .B2(n_643), .C(n_848), .Y(n_847) );
INVx1_ASAP7_75t_L g891 ( .A(n_45), .Y(n_891) );
INVx1_ASAP7_75t_L g1091 ( .A(n_46), .Y(n_1091) );
INVx1_ASAP7_75t_L g803 ( .A(n_47), .Y(n_803) );
AOI22xp5_ASAP7_75t_L g1159 ( .A1(n_48), .A2(n_156), .B1(n_1137), .B2(n_1141), .Y(n_1159) );
AOI221xp5_ASAP7_75t_L g1349 ( .A1(n_49), .A2(n_172), .B1(n_580), .B2(n_581), .C(n_1350), .Y(n_1349) );
INVx1_ASAP7_75t_L g802 ( .A(n_50), .Y(n_802) );
AOI22xp33_ASAP7_75t_SL g939 ( .A1(n_51), .A2(n_80), .B1(n_380), .B2(n_940), .Y(n_939) );
INVx1_ASAP7_75t_L g1353 ( .A(n_52), .Y(n_1353) );
AO221x2_ASAP7_75t_L g1229 ( .A1(n_53), .A2(n_191), .B1(n_1144), .B2(n_1147), .C(n_1230), .Y(n_1229) );
AOI22xp33_ASAP7_75t_L g855 ( .A1(n_54), .A2(n_109), .B1(n_611), .B2(n_851), .Y(n_855) );
INVx1_ASAP7_75t_L g878 ( .A(n_54), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g825 ( .A1(n_55), .A2(n_121), .B1(n_580), .B2(n_826), .C(n_828), .Y(n_825) );
INVx1_ASAP7_75t_L g1060 ( .A(n_56), .Y(n_1060) );
AOI22xp33_ASAP7_75t_SL g530 ( .A1(n_57), .A2(n_160), .B1(n_378), .B2(n_531), .Y(n_530) );
AOI22xp33_ASAP7_75t_SL g610 ( .A1(n_57), .A2(n_211), .B1(n_611), .B2(n_613), .Y(n_610) );
AOI221xp5_ASAP7_75t_L g834 ( .A1(n_58), .A2(n_62), .B1(n_483), .B2(n_608), .C(n_826), .Y(n_834) );
INVx1_ASAP7_75t_L g1116 ( .A(n_59), .Y(n_1116) );
INVx1_ASAP7_75t_L g474 ( .A(n_60), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g492 ( .A1(n_60), .A2(n_105), .B1(n_483), .B2(n_486), .C(n_493), .Y(n_492) );
AOI21xp33_ASAP7_75t_L g1343 ( .A1(n_61), .A2(n_857), .B(n_1344), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1365 ( .A1(n_61), .A2(n_148), .B1(n_401), .B2(n_664), .Y(n_1365) );
AOI22xp33_ASAP7_75t_SL g812 ( .A1(n_62), .A2(n_231), .B1(n_401), .B2(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g1395 ( .A(n_63), .Y(n_1395) );
OAI221xp5_ASAP7_75t_L g1403 ( .A1(n_63), .A2(n_220), .B1(n_1404), .B2(n_1405), .C(n_1406), .Y(n_1403) );
OAI222xp33_ASAP7_75t_L g984 ( .A1(n_64), .A2(n_183), .B1(n_417), .B2(n_421), .C1(n_985), .C2(n_987), .Y(n_984) );
INVx1_ASAP7_75t_L g997 ( .A(n_64), .Y(n_997) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_65), .Y(n_688) );
INVx1_ASAP7_75t_L g1073 ( .A(n_66), .Y(n_1073) );
OAI222xp33_ASAP7_75t_L g1110 ( .A1(n_66), .A2(n_103), .B1(n_845), .B2(n_1111), .C1(n_1117), .C2(n_1124), .Y(n_1110) );
OAI22xp5_ASAP7_75t_SL g1031 ( .A1(n_67), .A2(n_84), .B1(n_716), .B2(n_718), .Y(n_1031) );
OAI21xp33_ASAP7_75t_L g1042 ( .A1(n_67), .A2(n_671), .B(n_1043), .Y(n_1042) );
INVx1_ASAP7_75t_L g860 ( .A(n_68), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g1338 ( .A1(n_69), .A2(n_626), .B(n_1339), .C(n_1341), .Y(n_1338) );
INVx1_ASAP7_75t_L g1361 ( .A(n_69), .Y(n_1361) );
OAI22xp5_ASAP7_75t_L g1396 ( .A1(n_70), .A2(n_134), .B1(n_1397), .B2(n_1398), .Y(n_1396) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_70), .A2(n_134), .B1(n_784), .B2(n_786), .Y(n_1402) );
INVx1_ASAP7_75t_L g630 ( .A(n_71), .Y(n_630) );
CKINVDCx5p33_ASAP7_75t_R g974 ( .A(n_72), .Y(n_974) );
OAI211xp5_ASAP7_75t_L g639 ( .A1(n_73), .A2(n_575), .B(n_640), .C(n_647), .Y(n_639) );
INVx1_ASAP7_75t_L g327 ( .A(n_74), .Y(n_327) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_74), .A2(n_192), .B1(n_390), .B2(n_392), .C(n_395), .Y(n_389) );
HB1xp67_ASAP7_75t_L g255 ( .A(n_75), .Y(n_255) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_75), .B(n_253), .Y(n_1138) );
AOI22xp33_ASAP7_75t_SL g534 ( .A1(n_76), .A2(n_248), .B1(n_371), .B2(n_535), .Y(n_534) );
AOI21xp33_ASAP7_75t_L g605 ( .A1(n_76), .A2(n_606), .B(n_608), .Y(n_605) );
CKINVDCx5p33_ASAP7_75t_R g965 ( .A(n_77), .Y(n_965) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_78), .Y(n_806) );
OAI211xp5_ASAP7_75t_SL g1346 ( .A1(n_79), .A2(n_1347), .B(n_1348), .C(n_1352), .Y(n_1346) );
AOI221xp5_ASAP7_75t_SL g919 ( .A1(n_80), .A2(n_245), .B1(n_484), .B2(n_828), .C(n_920), .Y(n_919) );
INVx1_ASAP7_75t_L g975 ( .A(n_81), .Y(n_975) );
OAI22xp5_ASAP7_75t_L g562 ( .A1(n_82), .A2(n_237), .B1(n_563), .B2(n_569), .Y(n_562) );
INVx1_ASAP7_75t_L g588 ( .A(n_82), .Y(n_588) );
OAI211xp5_ASAP7_75t_L g1025 ( .A1(n_83), .A2(n_1026), .B(n_1027), .C(n_1028), .Y(n_1025) );
INVxp33_ASAP7_75t_SL g1044 ( .A(n_83), .Y(n_1044) );
INVxp67_ASAP7_75t_SL g1063 ( .A(n_84), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g1067 ( .A(n_85), .Y(n_1067) );
AND2x2_ASAP7_75t_L g1139 ( .A(n_86), .B(n_1140), .Y(n_1139) );
INVx1_ASAP7_75t_L g1146 ( .A(n_86), .Y(n_1146) );
OAI22xp33_ASAP7_75t_L g429 ( .A1(n_87), .A2(n_208), .B1(n_430), .B2(n_433), .Y(n_429) );
INVxp67_ASAP7_75t_SL g439 ( .A(n_87), .Y(n_439) );
CKINVDCx5p33_ASAP7_75t_R g927 ( .A(n_88), .Y(n_927) );
INVx1_ASAP7_75t_L g863 ( .A(n_89), .Y(n_863) );
CKINVDCx5p33_ASAP7_75t_R g706 ( .A(n_90), .Y(n_706) );
INVx1_ASAP7_75t_L g386 ( .A(n_91), .Y(n_386) );
INVx2_ASAP7_75t_L g397 ( .A(n_91), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_91), .B(n_388), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_92), .A2(n_127), .B1(n_372), .B2(n_400), .Y(n_479) );
INVx1_ASAP7_75t_L g494 ( .A(n_92), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g634 ( .A1(n_93), .A2(n_635), .B(n_636), .Y(n_634) );
AOI22xp33_ASAP7_75t_L g663 ( .A1(n_93), .A2(n_141), .B1(n_401), .B2(n_664), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g1136 ( .A1(n_94), .A2(n_187), .B1(n_1137), .B2(n_1141), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g752 ( .A1(n_95), .A2(n_151), .B1(n_753), .B2(n_754), .Y(n_752) );
OAI22xp33_ASAP7_75t_L g760 ( .A1(n_95), .A2(n_151), .B1(n_761), .B2(n_764), .Y(n_760) );
INVx1_ASAP7_75t_L g349 ( .A(n_96), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_97), .A2(n_123), .B1(n_281), .B2(n_288), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g398 ( .A1(n_97), .A2(n_180), .B1(n_399), .B2(n_401), .Y(n_398) );
INVx1_ASAP7_75t_L g879 ( .A(n_98), .Y(n_879) );
NOR2xp33_ASAP7_75t_L g898 ( .A(n_99), .B(n_549), .Y(n_898) );
OAI22xp5_ASAP7_75t_L g930 ( .A1(n_100), .A2(n_116), .B1(n_633), .B2(n_712), .Y(n_930) );
INVx1_ASAP7_75t_L g943 ( .A(n_100), .Y(n_943) );
INVxp67_ASAP7_75t_SL g632 ( .A(n_101), .Y(n_632) );
INVx1_ASAP7_75t_L g982 ( .A(n_102), .Y(n_982) );
NAND2xp33_ASAP7_75t_SL g1006 ( .A(n_102), .B(n_484), .Y(n_1006) );
INVx1_ASAP7_75t_L g1071 ( .A(n_103), .Y(n_1071) );
INVx1_ASAP7_75t_L g652 ( .A(n_104), .Y(n_652) );
AOI221xp5_ASAP7_75t_L g467 ( .A1(n_105), .A2(n_222), .B1(n_379), .B2(n_468), .C(n_469), .Y(n_467) );
XNOR2xp5_ASAP7_75t_L g446 ( .A(n_106), .B(n_447), .Y(n_446) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_107), .Y(n_691) );
OAI211xp5_ASAP7_75t_SL g730 ( .A1(n_108), .A2(n_725), .B(n_731), .C(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g780 ( .A(n_108), .Y(n_780) );
INVx1_ASAP7_75t_L g887 ( .A(n_109), .Y(n_887) );
AOI221xp5_ASAP7_75t_L g1100 ( .A1(n_110), .A2(n_241), .B1(n_643), .B2(n_1101), .C(n_1104), .Y(n_1100) );
INVx1_ASAP7_75t_L g649 ( .A(n_111), .Y(n_649) );
OAI22xp33_ASAP7_75t_L g670 ( .A1(n_111), .A2(n_157), .B1(n_563), .B2(n_671), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g701 ( .A(n_112), .Y(n_701) );
INVx1_ASAP7_75t_L g1112 ( .A(n_113), .Y(n_1112) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_114), .Y(n_523) );
OAI211xp5_ASAP7_75t_L g574 ( .A1(n_114), .A2(n_575), .B(n_578), .C(n_587), .Y(n_574) );
AOI22xp33_ASAP7_75t_SL g537 ( .A1(n_115), .A2(n_230), .B1(n_371), .B2(n_535), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_115), .A2(n_248), .B1(n_583), .B2(n_585), .Y(n_582) );
INVx1_ASAP7_75t_L g950 ( .A(n_116), .Y(n_950) );
CKINVDCx16_ASAP7_75t_R g986 ( .A(n_117), .Y(n_986) );
OAI22xp33_ASAP7_75t_L g454 ( .A1(n_118), .A2(n_243), .B1(n_430), .B2(n_433), .Y(n_454) );
INVxp33_ASAP7_75t_SL g504 ( .A(n_118), .Y(n_504) );
NAND5xp2_ASAP7_75t_L g907 ( .A(n_119), .B(n_908), .C(n_932), .D(n_944), .E(n_948), .Y(n_907) );
INVx1_ASAP7_75t_L g956 ( .A(n_119), .Y(n_956) );
AOI21xp5_ASAP7_75t_L g983 ( .A1(n_120), .A2(n_385), .B(n_400), .Y(n_983) );
INVx1_ASAP7_75t_L g1008 ( .A(n_122), .Y(n_1008) );
AOI22xp33_ASAP7_75t_SL g363 ( .A1(n_123), .A2(n_233), .B1(n_364), .B2(n_371), .Y(n_363) );
AO22x1_ASAP7_75t_L g1163 ( .A1(n_124), .A2(n_205), .B1(n_1144), .B2(n_1147), .Y(n_1163) );
INVx1_ASAP7_75t_L g514 ( .A(n_125), .Y(n_514) );
OAI221xp5_ASAP7_75t_L g592 ( .A1(n_125), .A2(n_128), .B1(n_593), .B2(n_597), .C(n_601), .Y(n_592) );
BUFx3_ASAP7_75t_L g370 ( .A(n_126), .Y(n_370) );
INVx1_ASAP7_75t_L g488 ( .A(n_127), .Y(n_488) );
INVx1_ASAP7_75t_L g518 ( .A(n_128), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g704 ( .A(n_129), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g457 ( .A(n_130), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_131), .A2(n_211), .B1(n_378), .B2(n_539), .Y(n_538) );
AOI221xp5_ASAP7_75t_L g579 ( .A1(n_131), .A2(n_160), .B1(n_486), .B2(n_580), .C(n_581), .Y(n_579) );
INVx1_ASAP7_75t_L g461 ( .A(n_132), .Y(n_461) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_132), .A2(n_175), .B1(n_483), .B2(n_486), .C(n_487), .Y(n_482) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_135), .A2(n_236), .B1(n_580), .B2(n_642), .C(n_643), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_135), .A2(n_193), .B1(n_539), .B2(n_669), .Y(n_668) );
INVx1_ASAP7_75t_L g867 ( .A(n_136), .Y(n_867) );
OAI21xp33_ASAP7_75t_L g1089 ( .A1(n_137), .A2(n_559), .B(n_1090), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1190 ( .A1(n_138), .A2(n_150), .B1(n_1144), .B2(n_1147), .Y(n_1190) );
BUFx6f_ASAP7_75t_L g266 ( .A(n_139), .Y(n_266) );
INVx1_ASAP7_75t_L g449 ( .A(n_140), .Y(n_449) );
INVx1_ASAP7_75t_L g822 ( .A(n_142), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_143), .A2(n_179), .B1(n_913), .B2(n_918), .Y(n_917) );
AOI22xp33_ASAP7_75t_L g937 ( .A1(n_143), .A2(n_173), .B1(n_401), .B2(n_938), .Y(n_937) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_144), .Y(n_738) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_145), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g322 ( .A1(n_146), .A2(n_180), .B1(n_288), .B2(n_323), .C(n_325), .Y(n_322) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_146), .A2(n_186), .B1(n_378), .B2(n_380), .C(n_385), .Y(n_377) );
AOI22xp33_ASAP7_75t_SL g1416 ( .A1(n_147), .A2(n_194), .B1(n_857), .B2(n_1417), .Y(n_1416) );
AOI22xp33_ASAP7_75t_L g1421 ( .A1(n_147), .A2(n_214), .B1(n_399), .B2(n_1422), .Y(n_1421) );
AOI22xp33_ASAP7_75t_L g1351 ( .A1(n_148), .A2(n_228), .B1(n_585), .B2(n_645), .Y(n_1351) );
OAI21xp5_ASAP7_75t_SL g835 ( .A1(n_149), .A2(n_654), .B(n_836), .Y(n_835) );
INVx1_ASAP7_75t_L g472 ( .A(n_152), .Y(n_472) );
INVx1_ASAP7_75t_L g1093 ( .A(n_153), .Y(n_1093) );
CKINVDCx5p33_ASAP7_75t_R g685 ( .A(n_154), .Y(n_685) );
INVx1_ASAP7_75t_L g966 ( .A(n_155), .Y(n_966) );
NOR2xp33_ASAP7_75t_L g968 ( .A(n_155), .B(n_430), .Y(n_968) );
INVx1_ASAP7_75t_L g648 ( .A(n_157), .Y(n_648) );
AOI22xp5_ASAP7_75t_L g1166 ( .A1(n_158), .A2(n_218), .B1(n_1137), .B2(n_1141), .Y(n_1166) );
INVx1_ASAP7_75t_L g1076 ( .A(n_159), .Y(n_1076) );
AOI22xp33_ASAP7_75t_L g1415 ( .A1(n_161), .A2(n_226), .B1(n_580), .B2(n_857), .Y(n_1415) );
AOI21xp33_ASAP7_75t_L g1039 ( .A1(n_162), .A2(n_486), .B(n_636), .Y(n_1039) );
INVx1_ASAP7_75t_L g1049 ( .A(n_162), .Y(n_1049) );
INVx1_ASAP7_75t_L g739 ( .A(n_163), .Y(n_739) );
OAI211xp5_ASAP7_75t_L g767 ( .A1(n_163), .A2(n_768), .B(n_770), .C(n_772), .Y(n_767) );
XOR2x2_ASAP7_75t_L g674 ( .A(n_164), .B(n_675), .Y(n_674) );
OAI211xp5_ASAP7_75t_L g844 ( .A1(n_165), .A2(n_845), .B(n_846), .C(n_852), .Y(n_844) );
INVx1_ASAP7_75t_L g895 ( .A(n_165), .Y(n_895) );
AOI221xp5_ASAP7_75t_L g856 ( .A1(n_166), .A2(n_232), .B1(n_580), .B2(n_857), .C(n_859), .Y(n_856) );
INVx1_ASAP7_75t_L g870 ( .A(n_166), .Y(n_870) );
INVx1_ASAP7_75t_L g947 ( .A(n_167), .Y(n_947) );
INVx1_ASAP7_75t_L g1382 ( .A(n_168), .Y(n_1382) );
INVx1_ASAP7_75t_L g865 ( .A(n_169), .Y(n_865) );
OAI332xp33_ASAP7_75t_SL g868 ( .A1(n_169), .A2(n_667), .A3(n_869), .B1(n_875), .B2(n_876), .B3(n_882), .C1(n_886), .C2(n_892), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g1189 ( .A1(n_170), .A2(n_215), .B1(n_1137), .B2(n_1141), .Y(n_1189) );
BUFx6f_ASAP7_75t_L g265 ( .A(n_171), .Y(n_265) );
AOI22xp33_ASAP7_75t_L g1366 ( .A1(n_172), .A2(n_181), .B1(n_669), .B2(n_1364), .Y(n_1366) );
AOI221xp5_ASAP7_75t_L g914 ( .A1(n_173), .A2(n_221), .B1(n_484), .B2(n_636), .C(n_915), .Y(n_914) );
INVx1_ASAP7_75t_L g1392 ( .A(n_174), .Y(n_1392) );
AOI21xp33_ASAP7_75t_L g478 ( .A1(n_175), .A2(n_394), .B(n_395), .Y(n_478) );
XOR2x2_ASAP7_75t_L g1018 ( .A(n_176), .B(n_1019), .Y(n_1018) );
AOI22xp33_ASAP7_75t_SL g1034 ( .A1(n_177), .A2(n_235), .B1(n_577), .B2(n_833), .Y(n_1034) );
INVx1_ASAP7_75t_L g1051 ( .A(n_177), .Y(n_1051) );
INVxp67_ASAP7_75t_SL g1342 ( .A(n_178), .Y(n_1342) );
AOI22xp33_ASAP7_75t_SL g1367 ( .A1(n_178), .A2(n_228), .B1(n_572), .B2(n_1368), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_179), .A2(n_221), .B1(n_401), .B2(n_813), .Y(n_936) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_182), .B(n_510), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g554 ( .A1(n_182), .A2(n_555), .B1(n_556), .B2(n_617), .Y(n_554) );
INVx1_ASAP7_75t_L g619 ( .A(n_182), .Y(n_619) );
NOR2xp33_ASAP7_75t_R g999 ( .A(n_183), .B(n_1000), .Y(n_999) );
AO22x1_ASAP7_75t_L g1179 ( .A1(n_184), .A2(n_206), .B1(n_1137), .B2(n_1180), .Y(n_1179) );
CKINVDCx16_ASAP7_75t_R g1231 ( .A(n_185), .Y(n_1231) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_186), .A2(n_192), .B1(n_292), .B2(n_296), .C(n_300), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g682 ( .A(n_188), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g850 ( .A1(n_189), .A2(n_212), .B1(n_611), .B2(n_851), .Y(n_850) );
INVx1_ASAP7_75t_L g885 ( .A(n_189), .Y(n_885) );
INVx1_ASAP7_75t_L g961 ( .A(n_190), .Y(n_961) );
AOI222xp33_ASAP7_75t_L g1331 ( .A1(n_191), .A2(n_1332), .B1(n_1370), .B2(n_1372), .C1(n_1377), .C2(n_1434), .Y(n_1331) );
OA22x2_ASAP7_75t_L g1378 ( .A1(n_191), .A2(n_1379), .B1(n_1432), .B2(n_1433), .Y(n_1378) );
INVxp67_ASAP7_75t_SL g1433 ( .A(n_191), .Y(n_1433) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_195), .Y(n_353) );
OAI221xp5_ASAP7_75t_L g416 ( .A1(n_195), .A2(n_198), .B1(n_417), .B2(n_421), .C(n_424), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g1079 ( .A1(n_196), .A2(n_241), .B1(n_390), .B2(n_531), .Y(n_1079) );
INVxp67_ASAP7_75t_SL g1118 ( .A(n_196), .Y(n_1118) );
OAI211xp5_ASAP7_75t_SL g455 ( .A1(n_197), .A2(n_411), .B(n_424), .C(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g499 ( .A(n_197), .Y(n_499) );
OAI221xp5_ASAP7_75t_L g306 ( .A1(n_198), .A2(n_210), .B1(n_307), .B2(n_315), .C(n_320), .Y(n_306) );
OAI211xp5_ASAP7_75t_L g625 ( .A1(n_199), .A2(n_626), .B(n_627), .C(n_631), .Y(n_625) );
INVx1_ASAP7_75t_L g659 ( .A(n_199), .Y(n_659) );
INVx1_ASAP7_75t_L g862 ( .A(n_200), .Y(n_862) );
CKINVDCx5p33_ASAP7_75t_R g1030 ( .A(n_201), .Y(n_1030) );
AOI22xp5_ASAP7_75t_L g1152 ( .A1(n_202), .A2(n_227), .B1(n_1144), .B2(n_1147), .Y(n_1152) );
BUFx3_ASAP7_75t_L g269 ( .A(n_203), .Y(n_269) );
INVx1_ASAP7_75t_L g345 ( .A(n_203), .Y(n_345) );
CKINVDCx20_ASAP7_75t_R g1233 ( .A(n_204), .Y(n_1233) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_208), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g924 ( .A(n_209), .Y(n_924) );
OAI22xp5_ASAP7_75t_L g402 ( .A1(n_210), .A2(n_213), .B1(n_403), .B2(n_407), .Y(n_402) );
INVx1_ASAP7_75t_L g872 ( .A(n_212), .Y(n_872) );
INVxp67_ASAP7_75t_SL g355 ( .A(n_213), .Y(n_355) );
CKINVDCx5p33_ASAP7_75t_R g698 ( .A(n_216), .Y(n_698) );
INVx1_ASAP7_75t_L g305 ( .A(n_217), .Y(n_305) );
INVx2_ASAP7_75t_L g310 ( .A(n_217), .Y(n_310) );
INVx1_ASAP7_75t_L g335 ( .A(n_217), .Y(n_335) );
XNOR2x1_ASAP7_75t_L g798 ( .A(n_218), .B(n_799), .Y(n_798) );
OAI211xp5_ASAP7_75t_L g1385 ( .A1(n_220), .A2(n_1386), .B(n_1387), .C(n_1390), .Y(n_1385) );
INVx1_ASAP7_75t_L g489 ( .A(n_222), .Y(n_489) );
INVx1_ASAP7_75t_L g972 ( .A(n_223), .Y(n_972) );
AOI22xp33_ASAP7_75t_L g1005 ( .A1(n_223), .A2(n_247), .B1(n_913), .B2(n_918), .Y(n_1005) );
NAND2xp5_ASAP7_75t_SL g1033 ( .A(n_224), .B(n_486), .Y(n_1033) );
AO22x1_ASAP7_75t_L g1181 ( .A1(n_225), .A2(n_242), .B1(n_1144), .B2(n_1147), .Y(n_1181) );
AOI22xp33_ASAP7_75t_L g1423 ( .A1(n_226), .A2(n_234), .B1(n_1424), .B2(n_1425), .Y(n_1423) );
INVx1_ASAP7_75t_L g1356 ( .A(n_229), .Y(n_1356) );
INVx1_ASAP7_75t_L g602 ( .A(n_230), .Y(n_602) );
INVxp67_ASAP7_75t_SL g883 ( .A(n_232), .Y(n_883) );
INVx1_ASAP7_75t_L g326 ( .A(n_233), .Y(n_326) );
INVxp67_ASAP7_75t_SL g1056 ( .A(n_235), .Y(n_1056) );
INVx1_ASAP7_75t_L g590 ( .A(n_237), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g466 ( .A(n_238), .Y(n_466) );
INVx1_ASAP7_75t_L g1125 ( .A(n_239), .Y(n_1125) );
INVxp67_ASAP7_75t_SL g452 ( .A(n_243), .Y(n_452) );
CKINVDCx5p33_ASAP7_75t_R g1029 ( .A(n_244), .Y(n_1029) );
INVx1_ASAP7_75t_L g1038 ( .A(n_246), .Y(n_1038) );
INVx1_ASAP7_75t_L g980 ( .A(n_247), .Y(n_980) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_250), .A2(n_270), .B(n_1128), .Y(n_249) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_256), .Y(n_250) );
INVx1_ASAP7_75t_L g1437 ( .A(n_251), .Y(n_1437) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
NOR2xp33_ASAP7_75t_L g1371 ( .A(n_252), .B(n_255), .Y(n_1371) );
INVx1_ASAP7_75t_L g1373 ( .A(n_252), .Y(n_1373) );
HB1xp67_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g1376 ( .A(n_255), .B(n_1373), .Y(n_1376) );
NAND2xp5_ASAP7_75t_L g256 ( .A(n_257), .B(n_260), .Y(n_256) );
INVx1_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
AND2x4_ASAP7_75t_L g757 ( .A(n_258), .B(n_758), .Y(n_757) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_258), .B(n_1437), .Y(n_1436) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x4_ASAP7_75t_L g302 ( .A(n_259), .B(n_269), .Y(n_302) );
AND2x4_ASAP7_75t_L g609 ( .A(n_259), .B(n_268), .Y(n_609) );
INVx1_ASAP7_75t_L g753 ( .A(n_260), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g1381 ( .A1(n_260), .A2(n_755), .B1(n_1382), .B2(n_1383), .Y(n_1381) );
AND2x4_ASAP7_75t_SL g1435 ( .A(n_260), .B(n_1436), .Y(n_1435) );
INVx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OR2x6_ASAP7_75t_L g261 ( .A(n_262), .B(n_267), .Y(n_261) );
OR2x6_ASAP7_75t_L g745 ( .A(n_262), .B(n_746), .Y(n_745) );
OR2x2_ASAP7_75t_L g1397 ( .A(n_262), .B(n_746), .Y(n_1397) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g290 ( .A(n_263), .Y(n_290) );
BUFx4f_ASAP7_75t_L g713 ( .A(n_263), .Y(n_713) );
INVx3_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
OR2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g287 ( .A(n_265), .Y(n_287) );
INVx2_ASAP7_75t_L g295 ( .A(n_265), .Y(n_295) );
NAND2x1_ASAP7_75t_L g299 ( .A(n_265), .B(n_266), .Y(n_299) );
INVx1_ASAP7_75t_L g318 ( .A(n_265), .Y(n_318) );
AND2x2_ASAP7_75t_L g443 ( .A(n_265), .B(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g485 ( .A(n_265), .B(n_266), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_266), .B(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g294 ( .A(n_266), .B(n_295), .Y(n_294) );
BUFx2_ASAP7_75t_L g314 ( .A(n_266), .Y(n_314) );
INVx1_ASAP7_75t_L g339 ( .A(n_266), .Y(n_339) );
AND2x2_ASAP7_75t_L g348 ( .A(n_266), .B(n_287), .Y(n_348) );
INVx2_ASAP7_75t_L g444 ( .A(n_266), .Y(n_444) );
INVxp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx1_ASAP7_75t_L g733 ( .A(n_268), .Y(n_733) );
INVx2_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g737 ( .A(n_269), .Y(n_737) );
AND2x4_ASAP7_75t_L g741 ( .A(n_269), .B(n_317), .Y(n_741) );
OAI22xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_272), .B1(n_900), .B2(n_901), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
XNOR2xp5_ASAP7_75t_L g272 ( .A(n_273), .B(n_795), .Y(n_272) );
XOR2xp5_ASAP7_75t_L g273 ( .A(n_274), .B(n_506), .Y(n_273) );
INVxp67_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
XNOR2x1_ASAP7_75t_L g275 ( .A(n_276), .B(n_446), .Y(n_275) );
XNOR2x1_ASAP7_75t_L g276 ( .A(n_277), .B(n_445), .Y(n_276) );
OR2x2_ASAP7_75t_L g277 ( .A(n_278), .B(n_361), .Y(n_277) );
NAND3xp33_ASAP7_75t_SL g278 ( .A(n_279), .B(n_331), .C(n_354), .Y(n_278) );
AOI211xp5_ASAP7_75t_SL g279 ( .A1(n_280), .A2(n_291), .B(n_306), .C(n_322), .Y(n_279) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g490 ( .A(n_284), .Y(n_490) );
INVx4_ASAP7_75t_L g716 ( .A(n_284), .Y(n_716) );
BUFx6f_ASAP7_75t_L g1123 ( .A(n_284), .Y(n_1123) );
INVx8_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
BUFx2_ASAP7_75t_L g324 ( .A(n_285), .Y(n_324) );
OR2x2_ASAP7_75t_L g751 ( .A(n_285), .B(n_737), .Y(n_751) );
OR2x2_ASAP7_75t_L g1398 ( .A(n_285), .B(n_733), .Y(n_1398) );
BUFx6f_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
BUFx6f_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
OAI22xp5_ASAP7_75t_L g487 ( .A1(n_290), .A2(n_488), .B1(n_489), .B2(n_490), .Y(n_487) );
OAI22x1_ASAP7_75t_SL g493 ( .A1(n_290), .A2(n_466), .B1(n_490), .B2(n_494), .Y(n_493) );
INVx2_ASAP7_75t_SL g724 ( .A(n_290), .Y(n_724) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g325 ( .A1(n_293), .A2(n_297), .B1(n_326), .B2(n_327), .C(n_328), .Y(n_325) );
BUFx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
BUFx2_ASAP7_75t_L g718 ( .A(n_294), .Y(n_718) );
INVx1_ASAP7_75t_L g1004 ( .A(n_294), .Y(n_1004) );
BUFx2_ASAP7_75t_L g1115 ( .A(n_294), .Y(n_1115) );
AND2x2_ASAP7_75t_L g338 ( .A(n_295), .B(n_339), .Y(n_338) );
HB1xp67_ASAP7_75t_L g926 ( .A(n_295), .Y(n_926) );
INVxp67_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
OAI221xp5_ASAP7_75t_L g1111 ( .A1(n_297), .A2(n_609), .B1(n_1112), .B2(n_1113), .C(n_1116), .Y(n_1111) );
BUFx4f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g320 ( .A(n_298), .B(n_321), .Y(n_320) );
INVx4_ASAP7_75t_L g604 ( .A(n_298), .Y(n_604) );
BUFx4f_ASAP7_75t_L g633 ( .A(n_298), .Y(n_633) );
BUFx6f_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
BUFx3_ASAP7_75t_L g352 ( .A(n_299), .Y(n_352) );
OAI21xp5_ASAP7_75t_L g1001 ( .A1(n_300), .A2(n_320), .B(n_1002), .Y(n_1001) );
INVx2_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AOI33xp33_ASAP7_75t_L g1412 ( .A1(n_301), .A2(n_1413), .A3(n_1414), .B1(n_1415), .B2(n_1416), .B3(n_1418), .Y(n_1412) );
AND2x2_ASAP7_75t_SL g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x4_ASAP7_75t_L g495 ( .A(n_302), .B(n_496), .Y(n_495) );
INVx4_ASAP7_75t_L g581 ( .A(n_302), .Y(n_581) );
INVx1_ASAP7_75t_SL g643 ( .A(n_302), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_302), .B(n_496), .Y(n_728) );
INVx4_ASAP7_75t_L g828 ( .A(n_302), .Y(n_828) );
NAND4xp25_ASAP7_75t_L g1032 ( .A(n_302), .B(n_1033), .C(n_1034), .D(n_1035), .Y(n_1032) );
INVx1_ASAP7_75t_L g497 ( .A(n_303), .Y(n_497) );
OR2x2_ASAP7_75t_L g551 ( .A(n_303), .B(n_406), .Y(n_551) );
OR2x2_ASAP7_75t_L g680 ( .A(n_303), .B(n_396), .Y(n_680) );
HB1xp67_ASAP7_75t_L g792 ( .A(n_303), .Y(n_792) );
INVx2_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx2_ASAP7_75t_L g319 ( .A(n_304), .Y(n_319) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g500 ( .A(n_307), .Y(n_500) );
INVx2_ASAP7_75t_SL g998 ( .A(n_307), .Y(n_998) );
NAND2x2_ASAP7_75t_L g307 ( .A(n_308), .B(n_312), .Y(n_307) );
INVx1_ASAP7_75t_L g321 ( .A(n_308), .Y(n_321) );
INVx2_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_310), .B(n_311), .Y(n_309) );
BUFx2_ASAP7_75t_L g329 ( .A(n_310), .Y(n_329) );
INVx2_ASAP7_75t_L g437 ( .A(n_310), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g316 ( .A(n_311), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_311), .B(n_338), .Y(n_337) );
AND2x6_ASAP7_75t_L g586 ( .A(n_311), .B(n_484), .Y(n_586) );
INVx1_ASAP7_75t_L g600 ( .A(n_311), .Y(n_600) );
AND2x2_ASAP7_75t_L g628 ( .A(n_311), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_SL g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_L g599 ( .A(n_314), .Y(n_599) );
BUFx2_ASAP7_75t_L g629 ( .A(n_314), .Y(n_629) );
AND2x4_ASAP7_75t_L g736 ( .A(n_314), .B(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_314), .B(n_733), .Y(n_1391) );
INVx1_ASAP7_75t_SL g996 ( .A(n_315), .Y(n_996) );
OR2x2_ASAP7_75t_L g315 ( .A(n_316), .B(n_319), .Y(n_315) );
OR2x2_ASAP7_75t_L g502 ( .A(n_316), .B(n_319), .Y(n_502) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx1_ASAP7_75t_L g359 ( .A(n_319), .Y(n_359) );
INVxp67_ASAP7_75t_L g526 ( .A(n_319), .Y(n_526) );
INVx1_ASAP7_75t_L g758 ( .A(n_319), .Y(n_758) );
CKINVDCx5p33_ASAP7_75t_R g505 ( .A(n_320), .Y(n_505) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_328), .Y(n_491) );
INVx4_ASAP7_75t_L g708 ( .A(n_328), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g992 ( .A(n_328), .B(n_993), .Y(n_992) );
AND2x4_ASAP7_75t_L g328 ( .A(n_329), .B(n_330), .Y(n_328) );
INVx1_ASAP7_75t_L g616 ( .A(n_329), .Y(n_616) );
OR2x6_ASAP7_75t_L g667 ( .A(n_329), .B(n_385), .Y(n_667) );
OR2x2_ASAP7_75t_L g811 ( .A(n_329), .B(n_385), .Y(n_811) );
AOI222xp33_ASAP7_75t_L g331 ( .A1(n_332), .A2(n_340), .B1(n_341), .B2(n_349), .C1(n_350), .C2(n_353), .Y(n_331) );
AOI21xp33_ASAP7_75t_SL g503 ( .A1(n_332), .A2(n_504), .B(n_505), .Y(n_503) );
AND2x4_ASAP7_75t_L g332 ( .A(n_333), .B(n_336), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
AND2x4_ASAP7_75t_L g517 ( .A(n_334), .B(n_414), .Y(n_517) );
OR2x2_ASAP7_75t_L g552 ( .A(n_334), .B(n_337), .Y(n_552) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_335), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g543 ( .A(n_335), .Y(n_543) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
AND2x2_ASAP7_75t_L g360 ( .A(n_338), .B(n_344), .Y(n_360) );
BUFx6f_ASAP7_75t_L g584 ( .A(n_338), .Y(n_584) );
INVx3_ASAP7_75t_L g612 ( .A(n_338), .Y(n_612) );
AOI222xp33_ASAP7_75t_L g498 ( .A1(n_341), .A2(n_457), .B1(n_472), .B2(n_499), .C1(n_500), .C2(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g1011 ( .A(n_341), .Y(n_1011) );
AND2x4_ASAP7_75t_L g341 ( .A(n_342), .B(n_346), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
OR2x2_ASAP7_75t_L g351 ( .A(n_343), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g1000 ( .A(n_343), .B(n_352), .Y(n_1000) );
AND2x2_ASAP7_75t_L g441 ( .A(n_344), .B(n_442), .Y(n_441) );
AND2x4_ASAP7_75t_L g576 ( .A(n_344), .B(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g591 ( .A(n_344), .B(n_442), .Y(n_591) );
AND2x4_ASAP7_75t_SL g596 ( .A(n_344), .B(n_484), .Y(n_596) );
AND2x2_ASAP7_75t_L g824 ( .A(n_344), .B(n_346), .Y(n_824) );
BUFx2_ASAP7_75t_L g929 ( .A(n_344), .Y(n_929) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_345), .Y(n_746) );
INVx3_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g613 ( .A(n_347), .Y(n_613) );
INVx2_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_348), .Y(n_577) );
BUFx3_ASAP7_75t_L g585 ( .A(n_348), .Y(n_585) );
BUFx3_ASAP7_75t_L g913 ( .A(n_348), .Y(n_913) );
AOI211xp5_ASAP7_75t_L g409 ( .A1(n_349), .A2(n_410), .B(n_416), .C(n_429), .Y(n_409) );
AOI222xp33_ASAP7_75t_L g481 ( .A1(n_350), .A2(n_458), .B1(n_482), .B2(n_491), .C1(n_492), .C2(n_495), .Y(n_481) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_SL g720 ( .A(n_352), .Y(n_720) );
BUFx2_ASAP7_75t_SL g725 ( .A(n_352), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_355), .B(n_356), .Y(n_354) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g1061 ( .A(n_357), .B(n_892), .Y(n_1061) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
HB1xp67_ASAP7_75t_L g448 ( .A(n_358), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g964 ( .A1(n_358), .A2(n_440), .B1(n_965), .B2(n_966), .Y(n_964) );
AND2x4_ASAP7_75t_L g358 ( .A(n_359), .B(n_360), .Y(n_358) );
AND2x4_ASAP7_75t_L g440 ( .A(n_359), .B(n_441), .Y(n_440) );
BUFx6f_ASAP7_75t_L g589 ( .A(n_360), .Y(n_589) );
INVx1_ASAP7_75t_L g1098 ( .A(n_360), .Y(n_1098) );
A2O1A1Ixp33_ASAP7_75t_L g361 ( .A1(n_362), .A2(n_409), .B(n_435), .C(n_438), .Y(n_361) );
AOI221xp5_ASAP7_75t_L g362 ( .A1(n_363), .A2(n_377), .B1(n_389), .B2(n_398), .C(n_402), .Y(n_362) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x6_ASAP7_75t_SL g430 ( .A(n_365), .B(n_431), .Y(n_430) );
INVx3_ASAP7_75t_L g664 ( .A(n_365), .Y(n_664) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
BUFx6f_ASAP7_75t_L g394 ( .A(n_366), .Y(n_394) );
BUFx8_ASAP7_75t_L g572 ( .A(n_366), .Y(n_572) );
BUFx6f_ASAP7_75t_L g690 ( .A(n_366), .Y(n_690) );
AND2x4_ASAP7_75t_L g366 ( .A(n_367), .B(n_369), .Y(n_366) );
INVxp67_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g384 ( .A(n_368), .Y(n_384) );
AND2x4_ASAP7_75t_L g382 ( .A(n_369), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_370), .Y(n_373) );
AND2x4_ASAP7_75t_L g379 ( .A(n_370), .B(n_375), .Y(n_379) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_370), .B(n_376), .Y(n_465) );
OR2x2_ASAP7_75t_L g566 ( .A(n_370), .B(n_384), .Y(n_566) );
BUFx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx12f_ASAP7_75t_L g401 ( .A(n_372), .Y(n_401) );
AND2x4_ASAP7_75t_L g434 ( .A(n_372), .B(n_432), .Y(n_434) );
INVx5_ASAP7_75t_L g1082 ( .A(n_372), .Y(n_1082) );
BUFx3_ASAP7_75t_L g1368 ( .A(n_372), .Y(n_1368) );
AND2x4_ASAP7_75t_L g372 ( .A(n_373), .B(n_374), .Y(n_372) );
INVx2_ASAP7_75t_L g420 ( .A(n_373), .Y(n_420) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_373), .B(n_427), .Y(n_426) );
BUFx2_ASAP7_75t_L g776 ( .A(n_373), .Y(n_776) );
INVx1_ASAP7_75t_L g423 ( .A(n_374), .Y(n_423) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g427 ( .A(n_376), .Y(n_427) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g391 ( .A(n_379), .Y(n_391) );
AND2x2_ASAP7_75t_L g408 ( .A(n_379), .B(n_405), .Y(n_408) );
BUFx2_ASAP7_75t_L g546 ( .A(n_379), .Y(n_546) );
BUFx2_ASAP7_75t_L g669 ( .A(n_379), .Y(n_669) );
AND2x4_ASAP7_75t_L g771 ( .A(n_379), .B(n_387), .Y(n_771) );
BUFx2_ASAP7_75t_L g935 ( .A(n_379), .Y(n_935) );
BUFx2_ASAP7_75t_L g1430 ( .A(n_379), .Y(n_1430) );
INVx8_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g468 ( .A(n_381), .Y(n_468) );
INVx3_ASAP7_75t_L g539 ( .A(n_381), .Y(n_539) );
INVx2_ASAP7_75t_L g810 ( .A(n_381), .Y(n_810) );
INVx2_ASAP7_75t_L g838 ( .A(n_381), .Y(n_838) );
INVx8_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
BUFx3_ASAP7_75t_L g400 ( .A(n_382), .Y(n_400) );
AND2x2_ASAP7_75t_L g404 ( .A(n_382), .B(n_405), .Y(n_404) );
NAND2x1p5_ASAP7_75t_L g413 ( .A(n_382), .B(n_414), .Y(n_413) );
BUFx3_ASAP7_75t_L g533 ( .A(n_382), .Y(n_533) );
HB1xp67_ASAP7_75t_L g1058 ( .A(n_382), .Y(n_1058) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx3_ASAP7_75t_L g470 ( .A(n_385), .Y(n_470) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
NAND3x1_ASAP7_75t_L g542 ( .A(n_386), .B(n_387), .C(n_543), .Y(n_542) );
AND2x4_ASAP7_75t_L g414 ( .A(n_387), .B(n_415), .Y(n_414) );
OR2x4_ASAP7_75t_L g763 ( .A(n_387), .B(n_566), .Y(n_763) );
INVx1_ASAP7_75t_L g766 ( .A(n_387), .Y(n_766) );
OR2x6_ASAP7_75t_L g786 ( .A(n_387), .B(n_787), .Y(n_786) );
INVx3_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
NAND2xp33_ASAP7_75t_SL g396 ( .A(n_388), .B(n_397), .Y(n_396) );
BUFx3_ASAP7_75t_L g529 ( .A(n_388), .Y(n_529) );
INVx2_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx2_ASAP7_75t_L g940 ( .A(n_391), .Y(n_940) );
INVx1_ASAP7_75t_L g1422 ( .A(n_391), .Y(n_1422) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g460 ( .A1(n_393), .A2(n_461), .B1(n_462), .B2(n_466), .C(n_467), .Y(n_460) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_393), .A2(n_425), .B1(n_974), .B2(n_975), .C(n_976), .Y(n_973) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
INVx2_ASAP7_75t_SL g536 ( .A(n_394), .Y(n_536) );
INVx5_ASAP7_75t_L g697 ( .A(n_394), .Y(n_697) );
INVx2_ASAP7_75t_SL g978 ( .A(n_394), .Y(n_978) );
BUFx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx1_ASAP7_75t_L g415 ( .A(n_397), .Y(n_415) );
AND3x4_ASAP7_75t_L g528 ( .A(n_397), .B(n_437), .C(n_529), .Y(n_528) );
HB1xp67_ASAP7_75t_L g790 ( .A(n_397), .Y(n_790) );
AND2x2_ASAP7_75t_L g976 ( .A(n_397), .B(n_529), .Y(n_976) );
BUFx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx2_ASAP7_75t_L g1084 ( .A(n_401), .Y(n_1084) );
INVx2_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
AOI22xp5_ASAP7_75t_L g471 ( .A1(n_404), .A2(n_408), .B1(n_449), .B2(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_L g432 ( .A(n_406), .Y(n_432) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
OR2x6_ASAP7_75t_L g525 ( .A(n_413), .B(n_526), .Y(n_525) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_413), .B(n_526), .Y(n_1010) );
AND2x6_ASAP7_75t_L g418 ( .A(n_414), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g422 ( .A(n_414), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g428 ( .A(n_414), .Y(n_428) );
INVx4_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g456 ( .A1(n_418), .A2(n_422), .B1(n_457), .B2(n_458), .Y(n_456) );
NAND2x1_ASAP7_75t_L g516 ( .A(n_419), .B(n_517), .Y(n_516) );
AND2x4_ASAP7_75t_SL g658 ( .A(n_419), .B(n_517), .Y(n_658) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_419), .B(n_517), .Y(n_1072) );
INVx3_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g521 ( .A(n_423), .Y(n_521) );
OAI221xp5_ASAP7_75t_L g969 ( .A1(n_424), .A2(n_970), .B1(n_973), .B2(n_977), .C(n_981), .Y(n_969) );
OR2x6_ASAP7_75t_L g424 ( .A(n_425), .B(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g890 ( .A(n_425), .Y(n_890) );
BUFx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx6f_ASAP7_75t_L g477 ( .A(n_426), .Y(n_477) );
BUFx3_ASAP7_75t_L g700 ( .A(n_426), .Y(n_700) );
BUFx2_ASAP7_75t_L g779 ( .A(n_427), .Y(n_779) );
INVx2_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
HB1xp67_ASAP7_75t_L g988 ( .A(n_432), .Y(n_988) );
INVx3_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g1015 ( .A(n_434), .B(n_616), .Y(n_1015) );
HB1xp67_ASAP7_75t_L g1041 ( .A(n_435), .Y(n_1041) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
AOI21x1_ASAP7_75t_L g908 ( .A1(n_436), .A2(n_909), .B(n_931), .Y(n_908) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
OAI31xp33_ASAP7_75t_SL g453 ( .A1(n_437), .A2(n_454), .A3(n_455), .B(n_459), .Y(n_453) );
OAI31xp33_ASAP7_75t_L g967 ( .A1(n_437), .A2(n_968), .A3(n_969), .B(n_984), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_440), .B(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g946 ( .A(n_440), .Y(n_946) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_442), .Y(n_635) );
INVx2_ASAP7_75t_L g827 ( .A(n_442), .Y(n_827) );
INVx1_ASAP7_75t_L g858 ( .A(n_442), .Y(n_858) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
BUFx3_ASAP7_75t_L g486 ( .A(n_443), .Y(n_486) );
AND2x4_ASAP7_75t_L g755 ( .A(n_443), .B(n_746), .Y(n_755) );
INVx2_ASAP7_75t_L g916 ( .A(n_443), .Y(n_916) );
AOI211x1_ASAP7_75t_L g447 ( .A1(n_448), .A2(n_449), .B(n_450), .C(n_480), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_453), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g459 ( .A(n_460), .B(n_471), .C(n_473), .Y(n_459) );
OAI22xp5_ASAP7_75t_L g882 ( .A1(n_462), .A2(n_883), .B1(n_884), .B2(n_885), .Y(n_882) );
OAI221xp5_ASAP7_75t_L g1055 ( .A1(n_462), .A2(n_697), .B1(n_1038), .B2(n_1056), .C(n_1057), .Y(n_1055) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g550 ( .A(n_463), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g874 ( .A(n_463), .Y(n_874) );
INVx1_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
BUFx6f_ASAP7_75t_L g693 ( .A(n_464), .Y(n_693) );
INVx1_ASAP7_75t_L g464 ( .A(n_465), .Y(n_464) );
BUFx2_ASAP7_75t_L g787 ( .A(n_465), .Y(n_787) );
INVx3_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
OAI211xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_478), .C(n_479), .Y(n_473) );
OAI21xp5_ASAP7_75t_SL g981 ( .A1(n_475), .A2(n_982), .B(n_983), .Y(n_981) );
INVx3_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g686 ( .A(n_476), .Y(n_686) );
INVx3_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
OR2x2_ASAP7_75t_L g560 ( .A(n_477), .B(n_551), .Y(n_560) );
INVx4_ASAP7_75t_L g881 ( .A(n_477), .Y(n_881) );
BUFx6f_ASAP7_75t_L g1404 ( .A(n_477), .Y(n_1404) );
NAND3xp33_ASAP7_75t_L g480 ( .A(n_481), .B(n_498), .C(n_503), .Y(n_480) );
BUFx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g580 ( .A(n_484), .Y(n_580) );
AND2x2_ASAP7_75t_L g732 ( .A(n_484), .B(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g849 ( .A(n_484), .Y(n_849) );
BUFx3_ASAP7_75t_L g1036 ( .A(n_484), .Y(n_1036) );
BUFx3_ASAP7_75t_L g1417 ( .A(n_484), .Y(n_1417) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx1_ASAP7_75t_L g1103 ( .A(n_485), .Y(n_1103) );
INVx1_ASAP7_75t_L g607 ( .A(n_486), .Y(n_607) );
HB1xp67_ASAP7_75t_L g1350 ( .A(n_486), .Y(n_1350) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
INVx2_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
AND2x4_ASAP7_75t_L g559 ( .A(n_502), .B(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g654 ( .A(n_502), .B(n_560), .Y(n_654) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_507), .A2(n_620), .B1(n_793), .B2(n_794), .Y(n_506) );
INVx1_ASAP7_75t_L g793 ( .A(n_507), .Y(n_793) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2x1p5_ASAP7_75t_L g508 ( .A(n_509), .B(n_554), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_511), .B(n_547), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
NOR2xp33_ASAP7_75t_SL g617 ( .A(n_512), .B(n_618), .Y(n_617) );
NAND4xp25_ASAP7_75t_SL g512 ( .A(n_513), .B(n_522), .C(n_527), .D(n_544), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_514), .A2(n_515), .B1(n_518), .B2(n_519), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_515), .A2(n_519), .B1(n_860), .B2(n_895), .Y(n_894) );
AOI221x1_ASAP7_75t_L g1045 ( .A1(n_515), .A2(n_519), .B1(n_1023), .B2(n_1029), .C(n_1046), .Y(n_1045) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x4_ASAP7_75t_L g519 ( .A(n_517), .B(n_520), .Y(n_519) );
AND2x4_ASAP7_75t_L g545 ( .A(n_517), .B(n_546), .Y(n_545) );
AND2x4_ASAP7_75t_SL g660 ( .A(n_517), .B(n_520), .Y(n_660) );
AO22x1_ASAP7_75t_L g1070 ( .A1(n_519), .A2(n_1071), .B1(n_1072), .B2(n_1073), .Y(n_1070) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_523), .B(n_524), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g896 ( .A(n_524), .B(n_863), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_524), .B(n_1063), .Y(n_1062) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_524), .B(n_1076), .Y(n_1075) );
INVx5_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx3_ASAP7_75t_L g801 ( .A(n_525), .Y(n_801) );
AOI33xp33_ASAP7_75t_L g527 ( .A1(n_528), .A2(n_530), .A3(n_534), .B1(n_537), .B2(n_538), .B3(n_540), .Y(n_527) );
AOI33xp33_ASAP7_75t_L g661 ( .A1(n_528), .A2(n_662), .A3(n_663), .B1(n_665), .B2(n_666), .B3(n_668), .Y(n_661) );
INVx1_ASAP7_75t_L g815 ( .A(n_528), .Y(n_815) );
AOI33xp33_ASAP7_75t_L g933 ( .A1(n_528), .A2(n_934), .A3(n_936), .B1(n_937), .B2(n_939), .B3(n_941), .Y(n_933) );
BUFx3_ASAP7_75t_L g1078 ( .A(n_528), .Y(n_1078) );
AOI33xp33_ASAP7_75t_L g1362 ( .A1(n_528), .A2(n_666), .A3(n_1363), .B1(n_1365), .B2(n_1366), .B3(n_1367), .Y(n_1362) );
AOI33xp33_ASAP7_75t_L g1420 ( .A1(n_528), .A2(n_1421), .A3(n_1423), .B1(n_1426), .B2(n_1429), .B3(n_1431), .Y(n_1420) );
INVx3_ASAP7_75t_L g775 ( .A(n_529), .Y(n_775) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_SL g532 ( .A(n_533), .Y(n_532) );
BUFx3_ASAP7_75t_L g1364 ( .A(n_533), .Y(n_1364) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g702 ( .A(n_540), .Y(n_702) );
BUFx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
BUFx2_ASAP7_75t_L g1085 ( .A(n_541), .Y(n_1085) );
INVx3_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
INVx3_ASAP7_75t_L g1054 ( .A(n_542), .Y(n_1054) );
NAND4xp25_ASAP7_75t_L g893 ( .A(n_544), .B(n_894), .C(n_896), .D(n_897), .Y(n_893) );
NAND2xp5_ASAP7_75t_SL g1074 ( .A(n_544), .B(n_1075), .Y(n_1074) );
INVx3_ASAP7_75t_L g544 ( .A(n_545), .Y(n_544) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_545), .Y(n_673) );
INVx3_ASAP7_75t_L g817 ( .A(n_545), .Y(n_817) );
AOI221xp5_ASAP7_75t_L g942 ( .A1(n_545), .A2(n_658), .B1(n_660), .B2(n_924), .C(n_943), .Y(n_942) );
NOR3xp33_ASAP7_75t_L g1358 ( .A(n_545), .B(n_1359), .C(n_1369), .Y(n_1358) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_547), .B(n_619), .Y(n_618) );
NAND2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_553), .Y(n_547) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_548), .A2(n_652), .B(n_653), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g800 ( .A1(n_548), .A2(n_801), .B1(n_802), .B2(n_803), .C(n_804), .Y(n_800) );
AOI211x1_ASAP7_75t_L g1066 ( .A1(n_548), .A2(n_1067), .B(n_1068), .C(n_1089), .Y(n_1066) );
AOI21xp5_ASAP7_75t_L g1355 ( .A1(n_548), .A2(n_1356), .B(n_1357), .Y(n_1355) );
INVx8_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x4_ASAP7_75t_L g549 ( .A(n_550), .B(n_552), .Y(n_549) );
INVx1_ASAP7_75t_L g951 ( .A(n_550), .Y(n_951) );
INVx1_ASAP7_75t_L g568 ( .A(n_551), .Y(n_568) );
INVx1_ASAP7_75t_L g571 ( .A(n_551), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g1014 ( .A(n_552), .B(n_1015), .Y(n_1014) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_573), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_562), .Y(n_557) );
AOI21xp5_ASAP7_75t_L g866 ( .A1(n_558), .A2(n_867), .B(n_868), .Y(n_866) );
INVx2_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx2_ASAP7_75t_L g949 ( .A(n_560), .Y(n_949) );
OR2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_567), .Y(n_563) );
OR2x6_ASAP7_75t_L g892 ( .A(n_564), .B(n_567), .Y(n_892) );
INVx2_ASAP7_75t_SL g564 ( .A(n_565), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
BUFx4f_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
OR2x4_ASAP7_75t_L g784 ( .A(n_566), .B(n_766), .Y(n_784) );
BUFx3_ASAP7_75t_L g877 ( .A(n_566), .Y(n_877) );
BUFx3_ASAP7_75t_L g888 ( .A(n_566), .Y(n_888) );
INVxp67_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
AND2x2_ASAP7_75t_L g672 ( .A(n_568), .B(n_664), .Y(n_672) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_570), .B(n_862), .Y(n_897) );
AOI22xp33_ASAP7_75t_L g1090 ( .A1(n_570), .A2(n_1091), .B1(n_1092), .B2(n_1093), .Y(n_1090) );
AND2x4_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
AND2x4_ASAP7_75t_L g837 ( .A(n_571), .B(n_838), .Y(n_837) );
AND2x4_ASAP7_75t_L g1092 ( .A(n_571), .B(n_838), .Y(n_1092) );
INVx3_ASAP7_75t_L g871 ( .A(n_572), .Y(n_871) );
OAI21xp5_ASAP7_75t_L g573 ( .A1(n_574), .A2(n_592), .B(n_614), .Y(n_573) );
INVx2_ASAP7_75t_SL g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_R g1109 ( .A(n_576), .B(n_1076), .Y(n_1109) );
INVx3_ASAP7_75t_L g1347 ( .A(n_576), .Y(n_1347) );
BUFx2_ASAP7_75t_L g851 ( .A(n_577), .Y(n_851) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_582), .B(n_586), .Y(n_578) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g646 ( .A(n_584), .Y(n_646) );
INVx1_ASAP7_75t_SL g1108 ( .A(n_585), .Y(n_1108) );
AOI21xp5_ASAP7_75t_L g640 ( .A1(n_586), .A2(n_641), .B(n_644), .Y(n_640) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_586), .A2(n_802), .B1(n_824), .B2(n_825), .C(n_829), .Y(n_823) );
INVx1_ASAP7_75t_L g852 ( .A(n_586), .Y(n_852) );
AOI21xp5_ASAP7_75t_L g1099 ( .A1(n_586), .A2(n_1100), .B(n_1105), .Y(n_1099) );
AOI21xp5_ASAP7_75t_L g1348 ( .A1(n_586), .A2(n_1349), .B(n_1351), .Y(n_1348) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_590), .B2(n_591), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g647 ( .A1(n_589), .A2(n_648), .B1(n_649), .B2(n_650), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g820 ( .A1(n_589), .A2(n_591), .B1(n_821), .B2(n_822), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g864 ( .A(n_589), .B(n_865), .Y(n_864) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_591), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_591), .A2(n_824), .B1(n_862), .B2(n_863), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1096 ( .A1(n_591), .A2(n_1091), .B1(n_1093), .B2(n_1097), .Y(n_1096) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g626 ( .A(n_594), .Y(n_626) );
INVx1_ASAP7_75t_L g845 ( .A(n_594), .Y(n_845) );
INVx4_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
BUFx3_ASAP7_75t_L g831 ( .A(n_596), .Y(n_831) );
BUFx2_ASAP7_75t_L g1124 ( .A(n_597), .Y(n_1124) );
INVx2_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
NOR2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_600), .Y(n_598) );
INVx1_ASAP7_75t_L g928 ( .A(n_600), .Y(n_928) );
OAI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_603), .B(n_605), .C(n_610), .Y(n_601) );
INVx2_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
INVx2_ASAP7_75t_L g1027 ( .A(n_604), .Y(n_1027) );
INVx1_ASAP7_75t_L g1386 ( .A(n_604), .Y(n_1386) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g642 ( .A(n_607), .Y(n_642) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx3_ASAP7_75t_L g636 ( .A(n_609), .Y(n_636) );
INVx2_ASAP7_75t_L g859 ( .A(n_609), .Y(n_859) );
INVx1_ASAP7_75t_L g1344 ( .A(n_609), .Y(n_1344) );
INVx2_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g638 ( .A(n_612), .Y(n_638) );
INVx1_ASAP7_75t_L g833 ( .A(n_612), .Y(n_833) );
INVx2_ASAP7_75t_L g918 ( .A(n_612), .Y(n_918) );
INVx2_ASAP7_75t_L g1106 ( .A(n_612), .Y(n_1106) );
OAI21xp5_ASAP7_75t_SL g624 ( .A1(n_614), .A2(n_625), .B(n_639), .Y(n_624) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_614), .A2(n_819), .B(n_835), .Y(n_818) );
OAI21xp5_ASAP7_75t_L g843 ( .A1(n_614), .A2(n_844), .B(n_853), .Y(n_843) );
OAI21xp5_ASAP7_75t_L g1094 ( .A1(n_614), .A2(n_1095), .B(n_1110), .Y(n_1094) );
OAI21xp5_ASAP7_75t_SL g1337 ( .A1(n_614), .A2(n_1338), .B(n_1346), .Y(n_1337) );
INVx2_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
BUFx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g794 ( .A(n_620), .Y(n_794) );
XNOR2xp5_ASAP7_75t_L g620 ( .A(n_621), .B(n_674), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_624), .B(n_651), .C(n_655), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_628), .B(n_630), .Y(n_627) );
AOI222xp33_ASAP7_75t_L g830 ( .A1(n_628), .A2(n_806), .B1(n_807), .B2(n_831), .C1(n_832), .C2(n_834), .Y(n_830) );
AOI22xp33_ASAP7_75t_L g854 ( .A1(n_628), .A2(n_855), .B1(n_856), .B2(n_860), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_628), .B(n_1340), .Y(n_1339) );
AOI22xp5_ASAP7_75t_L g923 ( .A1(n_629), .A2(n_924), .B1(n_925), .B2(n_927), .Y(n_923) );
AOI22xp33_ASAP7_75t_L g1028 ( .A1(n_629), .A2(n_925), .B1(n_1029), .B2(n_1030), .Y(n_1028) );
AOI22xp33_ASAP7_75t_L g657 ( .A1(n_630), .A2(n_658), .B1(n_659), .B2(n_660), .Y(n_657) );
OAI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_633), .B(n_634), .C(n_637), .Y(n_631) );
OAI211xp5_ASAP7_75t_L g1341 ( .A1(n_633), .A2(n_1342), .B(n_1343), .C(n_1345), .Y(n_1341) );
BUFx3_ASAP7_75t_L g1104 ( .A(n_635), .Y(n_1104) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx2_ASAP7_75t_SL g1419 ( .A(n_646), .Y(n_1419) );
AOI22xp33_ASAP7_75t_L g1352 ( .A1(n_650), .A2(n_1097), .B1(n_1353), .B2(n_1354), .Y(n_1352) );
NOR3xp33_ASAP7_75t_L g655 ( .A(n_656), .B(n_670), .C(n_673), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_661), .Y(n_656) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_658), .A2(n_660), .B1(n_806), .B2(n_807), .Y(n_805) );
AOI22xp33_ASAP7_75t_L g1360 ( .A1(n_658), .A2(n_660), .B1(n_1340), .B2(n_1361), .Y(n_1360) );
INVx1_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g941 ( .A(n_667), .Y(n_941) );
INVx1_ASAP7_75t_L g1431 ( .A(n_667), .Y(n_1431) );
INVx1_ASAP7_75t_L g1088 ( .A(n_669), .Y(n_1088) );
NAND2x1_ASAP7_75t_L g945 ( .A(n_671), .B(n_946), .Y(n_945) );
INVx2_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g836 ( .A1(n_672), .A2(n_821), .B1(n_822), .B2(n_837), .Y(n_836) );
NAND3xp33_ASAP7_75t_L g675 ( .A(n_676), .B(n_729), .C(n_759), .Y(n_675) );
NOR2xp33_ASAP7_75t_L g676 ( .A(n_677), .B(n_707), .Y(n_676) );
OAI33xp33_ASAP7_75t_L g677 ( .A1(n_678), .A2(n_681), .A3(n_687), .B1(n_694), .B2(n_702), .B3(n_703), .Y(n_677) );
BUFx3_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
BUFx4f_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
BUFx8_ASAP7_75t_L g875 ( .A(n_680), .Y(n_875) );
BUFx2_ASAP7_75t_L g1047 ( .A(n_680), .Y(n_1047) );
OAI22xp33_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_683), .B1(n_685), .B2(n_686), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_682), .A2(n_704), .B1(n_710), .B2(n_714), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g703 ( .A1(n_683), .A2(n_704), .B1(n_705), .B2(n_706), .Y(n_703) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g970 ( .A1(n_684), .A2(n_705), .B1(n_971), .B2(n_972), .Y(n_970) );
OAI22xp5_ASAP7_75t_L g721 ( .A1(n_685), .A2(n_706), .B1(n_714), .B2(n_718), .Y(n_721) );
OAI22xp5_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_689), .B1(n_691), .B2(n_692), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g717 ( .A1(n_688), .A2(n_698), .B1(n_718), .B2(n_719), .Y(n_717) );
INVx1_ASAP7_75t_L g1424 ( .A(n_689), .Y(n_1424) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x4_ASAP7_75t_L g765 ( .A(n_690), .B(n_766), .Y(n_765) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_690), .Y(n_813) );
BUFx6f_ASAP7_75t_L g938 ( .A(n_690), .Y(n_938) );
INVx1_ASAP7_75t_L g1428 ( .A(n_690), .Y(n_1428) );
OAI22xp33_ASAP7_75t_L g722 ( .A1(n_691), .A2(n_701), .B1(n_723), .B2(n_725), .Y(n_722) );
OAI22xp5_ASAP7_75t_L g977 ( .A1(n_692), .A2(n_978), .B1(n_979), .B2(n_980), .Y(n_977) );
INVx3_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx3_ASAP7_75t_L g705 ( .A(n_693), .Y(n_705) );
INVx3_ASAP7_75t_L g1050 ( .A(n_693), .Y(n_1050) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_695), .A2(n_698), .B1(n_699), .B2(n_701), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx8_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
BUFx6f_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g769 ( .A(n_700), .Y(n_769) );
OAI33xp33_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .A3(n_717), .B1(n_721), .B2(n_722), .B3(n_726), .Y(n_707) );
INVx2_ASAP7_75t_SL g1413 ( .A(n_708), .Y(n_1413) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_SL g711 ( .A(n_712), .Y(n_711) );
INVx3_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx4_ASAP7_75t_L g1026 ( .A(n_713), .Y(n_1026) );
BUFx6f_ASAP7_75t_L g1120 ( .A(n_713), .Y(n_1120) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
OAI211xp5_ASAP7_75t_L g1037 ( .A1(n_719), .A2(n_1038), .B(n_1039), .C(n_1040), .Y(n_1037) );
INVx5_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
OAI31xp33_ASAP7_75t_SL g729 ( .A1(n_730), .A2(n_742), .A3(n_752), .B(n_756), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
AND2x2_ASAP7_75t_L g1388 ( .A(n_733), .B(n_1389), .Y(n_1388) );
AOI22xp33_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_738), .B1(n_739), .B2(n_740), .Y(n_734) );
BUFx3_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_738), .A2(n_773), .B1(n_777), .B2(n_780), .Y(n_772) );
BUFx3_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g1394 ( .A(n_741), .Y(n_1394) );
INVx1_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx2_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx2_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
INVx3_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
BUFx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
INVx1_ASAP7_75t_L g1399 ( .A(n_757), .Y(n_1399) );
OAI31xp33_ASAP7_75t_SL g759 ( .A1(n_760), .A2(n_767), .A3(n_781), .B(n_788), .Y(n_759) );
INVx1_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx2_ASAP7_75t_SL g1409 ( .A(n_763), .Y(n_1409) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
AOI22xp33_ASAP7_75t_L g1408 ( .A1(n_765), .A2(n_1382), .B1(n_1383), .B2(n_1409), .Y(n_1408) );
INVx2_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
CKINVDCx8_ASAP7_75t_R g770 ( .A(n_771), .Y(n_770) );
NOR3xp33_ASAP7_75t_L g1401 ( .A(n_771), .B(n_1402), .C(n_1403), .Y(n_1401) );
BUFx3_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AND2x2_ASAP7_75t_L g774 ( .A(n_775), .B(n_776), .Y(n_774) );
AND2x4_ASAP7_75t_L g778 ( .A(n_775), .B(n_779), .Y(n_778) );
AND2x4_ASAP7_75t_L g1407 ( .A(n_775), .B(n_776), .Y(n_1407) );
BUFx6f_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g1405 ( .A(n_778), .Y(n_1405) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
BUFx3_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
AND2x2_ASAP7_75t_L g788 ( .A(n_789), .B(n_791), .Y(n_788) );
AND2x2_ASAP7_75t_L g1411 ( .A(n_789), .B(n_791), .Y(n_1411) );
INVx1_ASAP7_75t_SL g789 ( .A(n_790), .Y(n_789) );
INVx1_ASAP7_75t_L g791 ( .A(n_792), .Y(n_791) );
HB1xp67_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
AOI22xp5_ASAP7_75t_L g796 ( .A1(n_797), .A2(n_839), .B1(n_840), .B2(n_899), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
HB1xp67_ASAP7_75t_L g899 ( .A(n_798), .Y(n_899) );
AND2x2_ASAP7_75t_L g799 ( .A(n_800), .B(n_818), .Y(n_799) );
NAND3xp33_ASAP7_75t_SL g804 ( .A(n_805), .B(n_808), .C(n_817), .Y(n_804) );
AOI22xp5_ASAP7_75t_L g808 ( .A1(n_809), .A2(n_812), .B1(n_814), .B2(n_816), .Y(n_808) );
INVx2_ASAP7_75t_L g884 ( .A(n_813), .Y(n_884) );
AND5x1_ASAP7_75t_L g1019 ( .A(n_817), .B(n_1020), .C(n_1045), .D(n_1059), .E(n_1062), .Y(n_1019) );
NAND3xp33_ASAP7_75t_L g819 ( .A(n_820), .B(n_823), .C(n_830), .Y(n_819) );
INVx2_ASAP7_75t_L g910 ( .A(n_824), .Y(n_910) );
INVx2_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_831), .B(n_1023), .Y(n_1022) );
AOI222xp33_ASAP7_75t_L g948 ( .A1(n_837), .A2(n_927), .B1(n_949), .B2(n_950), .C1(n_951), .C2(n_952), .Y(n_948) );
AOI22xp5_ASAP7_75t_L g985 ( .A1(n_838), .A2(n_940), .B1(n_965), .B2(n_986), .Y(n_985) );
INVxp67_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
NOR3xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_893), .C(n_898), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_843), .B(n_866), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g846 ( .A(n_847), .B(n_850), .Y(n_846) );
INVx1_ASAP7_75t_L g848 ( .A(n_849), .Y(n_848) );
NAND3xp33_ASAP7_75t_L g853 ( .A(n_854), .B(n_861), .C(n_864), .Y(n_853) );
INVx2_ASAP7_75t_SL g857 ( .A(n_858), .Y(n_857) );
OAI22xp5_ASAP7_75t_L g869 ( .A1(n_870), .A2(n_871), .B1(n_872), .B2(n_873), .Y(n_869) );
INVx1_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI22xp33_ASAP7_75t_L g876 ( .A1(n_877), .A2(n_878), .B1(n_879), .B2(n_880), .Y(n_876) );
INVx1_ASAP7_75t_L g880 ( .A(n_881), .Y(n_880) );
OAI22xp5_ASAP7_75t_L g886 ( .A1(n_887), .A2(n_888), .B1(n_889), .B2(n_891), .Y(n_886) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_L g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_L g901 ( .A(n_902), .Y(n_901) );
INVx1_ASAP7_75t_L g902 ( .A(n_903), .Y(n_902) );
AO22x2_ASAP7_75t_L g903 ( .A1(n_904), .A2(n_1064), .B1(n_1126), .B2(n_1127), .Y(n_903) );
INVx1_ASAP7_75t_L g1126 ( .A(n_904), .Y(n_1126) );
XNOR2xp5_ASAP7_75t_L g904 ( .A(n_905), .B(n_1018), .Y(n_904) );
OAI22xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_960), .B1(n_1016), .B2(n_1017), .Y(n_905) );
INVx1_ASAP7_75t_L g1017 ( .A(n_906), .Y(n_1017) );
NAND3xp33_ASAP7_75t_L g906 ( .A(n_907), .B(n_953), .C(n_957), .Y(n_906) );
INVx1_ASAP7_75t_L g954 ( .A(n_908), .Y(n_954) );
AOI22xp5_ASAP7_75t_L g911 ( .A1(n_912), .A2(n_914), .B1(n_917), .B2(n_919), .Y(n_911) );
INVx2_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g920 ( .A(n_916), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_922), .A2(n_928), .B1(n_929), .B2(n_930), .Y(n_921) );
INVx1_ASAP7_75t_L g925 ( .A(n_926), .Y(n_925) );
AOI22xp5_ASAP7_75t_L g1024 ( .A1(n_928), .A2(n_929), .B1(n_1025), .B2(n_1031), .Y(n_1024) );
INVx1_ASAP7_75t_L g955 ( .A(n_932), .Y(n_955) );
AND2x2_ASAP7_75t_L g932 ( .A(n_933), .B(n_942), .Y(n_932) );
INVx1_ASAP7_75t_L g959 ( .A(n_944), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_945), .B(n_947), .Y(n_944) );
INVx1_ASAP7_75t_L g958 ( .A(n_948), .Y(n_958) );
AOI22xp5_ASAP7_75t_L g1043 ( .A1(n_949), .A2(n_951), .B1(n_1030), .B2(n_1044), .Y(n_1043) );
OAI21xp5_ASAP7_75t_L g953 ( .A1(n_954), .A2(n_955), .B(n_956), .Y(n_953) );
OAI21xp33_ASAP7_75t_L g957 ( .A1(n_956), .A2(n_958), .B(n_959), .Y(n_957) );
INVx1_ASAP7_75t_L g1016 ( .A(n_960), .Y(n_1016) );
XNOR2xp5_ASAP7_75t_L g960 ( .A(n_961), .B(n_962), .Y(n_960) );
NOR2x1_ASAP7_75t_L g962 ( .A(n_963), .B(n_989), .Y(n_962) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_964), .B(n_967), .Y(n_963) );
OAI211xp5_ASAP7_75t_L g1002 ( .A1(n_974), .A2(n_1003), .B(n_1005), .C(n_1006), .Y(n_1002) );
OAI221xp5_ASAP7_75t_L g1048 ( .A1(n_978), .A2(n_1049), .B1(n_1050), .B2(n_1051), .C(n_1052), .Y(n_1048) );
AOI22xp5_ASAP7_75t_L g995 ( .A1(n_986), .A2(n_996), .B1(n_997), .B2(n_998), .Y(n_995) );
INVx1_ASAP7_75t_L g987 ( .A(n_988), .Y(n_987) );
NAND3xp33_ASAP7_75t_L g989 ( .A(n_990), .B(n_1007), .C(n_1012), .Y(n_989) );
NOR3xp33_ASAP7_75t_SL g990 ( .A(n_991), .B(n_999), .C(n_1001), .Y(n_990) );
OAI21xp5_ASAP7_75t_SL g991 ( .A1(n_992), .A2(n_994), .B(n_995), .Y(n_991) );
INVx2_ASAP7_75t_L g1003 ( .A(n_1004), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_1010), .B(n_1011), .Y(n_1009) );
NAND2xp5_ASAP7_75t_L g1012 ( .A(n_1013), .B(n_1014), .Y(n_1012) );
AOI21xp5_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1041), .B(n_1042), .Y(n_1020) );
NAND4xp25_ASAP7_75t_L g1021 ( .A(n_1022), .B(n_1024), .C(n_1032), .D(n_1037), .Y(n_1021) );
OAI22xp5_ASAP7_75t_SL g1046 ( .A1(n_1047), .A2(n_1048), .B1(n_1053), .B2(n_1055), .Y(n_1046) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
NAND2xp5_ASAP7_75t_L g1059 ( .A(n_1060), .B(n_1061), .Y(n_1059) );
INVx2_ASAP7_75t_L g1127 ( .A(n_1064), .Y(n_1127) );
XOR2x2_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1125), .Y(n_1064) );
NAND2xp5_ASAP7_75t_SL g1065 ( .A(n_1066), .B(n_1094), .Y(n_1065) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1077), .Y(n_1068) );
NOR2xp33_ASAP7_75t_L g1069 ( .A(n_1070), .B(n_1074), .Y(n_1069) );
AOI33xp33_ASAP7_75t_L g1077 ( .A1(n_1078), .A2(n_1079), .A3(n_1080), .B1(n_1083), .B2(n_1085), .B3(n_1086), .Y(n_1077) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx2_ASAP7_75t_R g1425 ( .A(n_1082), .Y(n_1425) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
NAND3xp33_ASAP7_75t_SL g1095 ( .A(n_1096), .B(n_1099), .C(n_1109), .Y(n_1095) );
INVx2_ASAP7_75t_L g1097 ( .A(n_1098), .Y(n_1097) );
INVx1_ASAP7_75t_L g1101 ( .A(n_1102), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1102 ( .A(n_1103), .Y(n_1102) );
INVx1_ASAP7_75t_L g1389 ( .A(n_1103), .Y(n_1389) );
INVx1_ASAP7_75t_SL g1107 ( .A(n_1108), .Y(n_1107) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
INVx4_ASAP7_75t_L g1114 ( .A(n_1115), .Y(n_1114) );
OAI22xp5_ASAP7_75t_L g1117 ( .A1(n_1118), .A2(n_1119), .B1(n_1121), .B2(n_1122), .Y(n_1117) );
INVx2_ASAP7_75t_L g1119 ( .A(n_1120), .Y(n_1119) );
INVx5_ASAP7_75t_L g1122 ( .A(n_1123), .Y(n_1122) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1329), .B(n_1331), .Y(n_1128) );
NOR2xp67_ASAP7_75t_SL g1129 ( .A(n_1130), .B(n_1280), .Y(n_1129) );
OAI21xp5_ASAP7_75t_L g1130 ( .A1(n_1131), .A2(n_1227), .B(n_1235), .Y(n_1130) );
NOR4xp25_ASAP7_75t_L g1131 ( .A(n_1132), .B(n_1194), .C(n_1206), .D(n_1222), .Y(n_1131) );
OAI211xp5_ASAP7_75t_L g1132 ( .A1(n_1133), .A2(n_1149), .B(n_1167), .C(n_1182), .Y(n_1132) );
CKINVDCx14_ASAP7_75t_R g1133 ( .A(n_1134), .Y(n_1133) );
OAI322xp33_ASAP7_75t_L g1206 ( .A1(n_1134), .A2(n_1151), .A3(n_1207), .B1(n_1208), .B2(n_1213), .C1(n_1218), .C2(n_1220), .Y(n_1206) );
AOI22xp33_ASAP7_75t_L g1247 ( .A1(n_1134), .A2(n_1160), .B1(n_1248), .B2(n_1249), .Y(n_1247) );
INVx3_ASAP7_75t_L g1134 ( .A(n_1135), .Y(n_1134) );
OR2x2_ASAP7_75t_L g1176 ( .A(n_1135), .B(n_1177), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1186 ( .A(n_1135), .B(n_1187), .Y(n_1186) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1135), .Y(n_1212) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1135), .B(n_1196), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1135), .B(n_1188), .Y(n_1250) );
AND2x2_ASAP7_75t_L g1257 ( .A(n_1135), .B(n_1178), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1275 ( .A(n_1135), .B(n_1177), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1299 ( .A(n_1135), .B(n_1188), .Y(n_1299) );
OR2x2_ASAP7_75t_L g1319 ( .A(n_1135), .B(n_1178), .Y(n_1319) );
AND2x4_ASAP7_75t_L g1135 ( .A(n_1136), .B(n_1143), .Y(n_1135) );
INVx2_ASAP7_75t_L g1232 ( .A(n_1137), .Y(n_1232) );
AND2x6_ASAP7_75t_L g1137 ( .A(n_1138), .B(n_1139), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_1138), .B(n_1142), .Y(n_1141) );
AND2x4_ASAP7_75t_L g1144 ( .A(n_1138), .B(n_1145), .Y(n_1144) );
AND2x6_ASAP7_75t_L g1147 ( .A(n_1138), .B(n_1148), .Y(n_1147) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_1138), .B(n_1142), .Y(n_1154) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_1138), .B(n_1142), .Y(n_1180) );
NAND2xp5_ASAP7_75t_L g1330 ( .A(n_1138), .B(n_1145), .Y(n_1330) );
AND2x2_ASAP7_75t_L g1145 ( .A(n_1140), .B(n_1146), .Y(n_1145) );
INVxp67_ASAP7_75t_L g1234 ( .A(n_1141), .Y(n_1234) );
HB1xp67_ASAP7_75t_L g1374 ( .A(n_1145), .Y(n_1374) );
OR2x2_ASAP7_75t_L g1149 ( .A(n_1150), .B(n_1155), .Y(n_1149) );
NAND2xp5_ASAP7_75t_L g1170 ( .A(n_1150), .B(n_1164), .Y(n_1170) );
AND2x2_ASAP7_75t_L g1202 ( .A(n_1150), .B(n_1203), .Y(n_1202) );
AND3x1_ASAP7_75t_L g1255 ( .A(n_1150), .B(n_1164), .C(n_1174), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1263 ( .A(n_1150), .B(n_1174), .Y(n_1263) );
AND2x2_ASAP7_75t_L g1273 ( .A(n_1150), .B(n_1156), .Y(n_1273) );
AND2x2_ASAP7_75t_L g1293 ( .A(n_1150), .B(n_1294), .Y(n_1293) );
INVx2_ASAP7_75t_L g1150 ( .A(n_1151), .Y(n_1150) );
BUFx2_ASAP7_75t_L g1172 ( .A(n_1151), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1151), .B(n_1203), .Y(n_1219) );
OR2x2_ASAP7_75t_L g1225 ( .A(n_1151), .B(n_1226), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1151), .B(n_1160), .Y(n_1259) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1151), .B(n_1294), .Y(n_1312) );
AND2x2_ASAP7_75t_L g1151 ( .A(n_1152), .B(n_1153), .Y(n_1151) );
NAND2xp5_ASAP7_75t_L g1155 ( .A(n_1156), .B(n_1160), .Y(n_1155) );
INVx1_ASAP7_75t_L g1185 ( .A(n_1156), .Y(n_1185) );
NAND2xp5_ASAP7_75t_L g1215 ( .A(n_1156), .B(n_1216), .Y(n_1215) );
NAND2xp5_ASAP7_75t_L g1251 ( .A(n_1156), .B(n_1203), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1289 ( .A(n_1156), .B(n_1211), .Y(n_1289) );
INVx2_ASAP7_75t_L g1156 ( .A(n_1157), .Y(n_1156) );
AND2x2_ASAP7_75t_L g1168 ( .A(n_1157), .B(n_1169), .Y(n_1168) );
OR2x2_ASAP7_75t_L g1192 ( .A(n_1157), .B(n_1188), .Y(n_1192) );
AND2x2_ASAP7_75t_L g1196 ( .A(n_1157), .B(n_1188), .Y(n_1196) );
INVx1_ASAP7_75t_L g1201 ( .A(n_1157), .Y(n_1201) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1157), .B(n_1178), .Y(n_1266) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1157), .B(n_1172), .Y(n_1279) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1157), .B(n_1187), .Y(n_1305) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1157), .B(n_1197), .Y(n_1317) );
OR2x2_ASAP7_75t_L g1320 ( .A(n_1157), .B(n_1321), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1157 ( .A(n_1158), .B(n_1159), .Y(n_1157) );
INVx1_ASAP7_75t_L g1226 ( .A(n_1160), .Y(n_1226) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1160), .B(n_1273), .Y(n_1315) );
AND2x2_ASAP7_75t_L g1160 ( .A(n_1161), .B(n_1164), .Y(n_1160) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1161), .Y(n_1174) );
AND2x2_ASAP7_75t_L g1203 ( .A(n_1161), .B(n_1204), .Y(n_1203) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1161), .B(n_1172), .Y(n_1321) );
NAND3xp33_ASAP7_75t_L g1322 ( .A(n_1161), .B(n_1229), .C(n_1284), .Y(n_1322) );
OR2x2_ASAP7_75t_L g1161 ( .A(n_1162), .B(n_1163), .Y(n_1161) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1164), .B(n_1174), .Y(n_1173) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1164), .Y(n_1204) );
OAI211xp5_ASAP7_75t_L g1246 ( .A1(n_1164), .A2(n_1192), .B(n_1247), .C(n_1251), .Y(n_1246) );
NOR2xp33_ASAP7_75t_L g1304 ( .A(n_1164), .B(n_1305), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1164 ( .A(n_1165), .B(n_1166), .Y(n_1164) );
OAI21xp5_ASAP7_75t_L g1167 ( .A1(n_1168), .A2(n_1171), .B(n_1175), .Y(n_1167) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1170), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1248 ( .A(n_1170), .B(n_1185), .Y(n_1248) );
OAI221xp5_ASAP7_75t_L g1301 ( .A1(n_1170), .A2(n_1225), .B1(n_1256), .B2(n_1302), .C(n_1303), .Y(n_1301) );
AOI21xp33_ASAP7_75t_L g1306 ( .A1(n_1170), .A2(n_1192), .B(n_1307), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1241 ( .A(n_1171), .B(n_1201), .Y(n_1241) );
NOR2xp33_ASAP7_75t_L g1287 ( .A(n_1171), .B(n_1202), .Y(n_1287) );
AND2x2_ASAP7_75t_L g1171 ( .A(n_1172), .B(n_1173), .Y(n_1171) );
AND2x2_ASAP7_75t_L g1193 ( .A(n_1172), .B(n_1174), .Y(n_1193) );
OR2x2_ASAP7_75t_L g1197 ( .A(n_1172), .B(n_1174), .Y(n_1197) );
OR2x2_ASAP7_75t_L g1207 ( .A(n_1173), .B(n_1203), .Y(n_1207) );
NAND3xp33_ASAP7_75t_L g1213 ( .A(n_1173), .B(n_1214), .C(n_1217), .Y(n_1213) );
AND2x2_ASAP7_75t_L g1272 ( .A(n_1173), .B(n_1273), .Y(n_1272) );
AOI221xp5_ASAP7_75t_L g1242 ( .A1(n_1174), .A2(n_1202), .B1(n_1243), .B2(n_1244), .C(n_1246), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1174), .B(n_1204), .Y(n_1294) );
AOI21xp5_ASAP7_75t_L g1303 ( .A1(n_1175), .A2(n_1304), .B(n_1306), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1308 ( .A(n_1175), .B(n_1241), .Y(n_1308) );
INVx1_ASAP7_75t_L g1175 ( .A(n_1176), .Y(n_1175) );
NOR2xp33_ASAP7_75t_L g1191 ( .A(n_1177), .B(n_1192), .Y(n_1191) );
NOR2xp33_ASAP7_75t_SL g1209 ( .A(n_1177), .B(n_1210), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1221 ( .A(n_1177), .B(n_1187), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1177), .B(n_1229), .Y(n_1237) );
NAND2xp5_ASAP7_75t_L g1260 ( .A(n_1177), .B(n_1249), .Y(n_1260) );
AND2x2_ASAP7_75t_L g1313 ( .A(n_1177), .B(n_1211), .Y(n_1313) );
CKINVDCx6p67_ASAP7_75t_R g1177 ( .A(n_1178), .Y(n_1177) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_1178), .Y(n_1205) );
OR2x2_ASAP7_75t_L g1223 ( .A(n_1178), .B(n_1224), .Y(n_1223) );
OR2x6_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1181), .Y(n_1178) );
OR2x2_ASAP7_75t_L g1217 ( .A(n_1179), .B(n_1181), .Y(n_1217) );
OAI21xp5_ASAP7_75t_L g1182 ( .A1(n_1183), .A2(n_1191), .B(n_1193), .Y(n_1182) );
INVx1_ASAP7_75t_L g1183 ( .A(n_1184), .Y(n_1183) );
NAND2xp5_ASAP7_75t_L g1184 ( .A(n_1185), .B(n_1186), .Y(n_1184) );
CKINVDCx6p67_ASAP7_75t_R g1224 ( .A(n_1186), .Y(n_1224) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1187), .Y(n_1216) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1188), .B(n_1212), .Y(n_1211) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1189), .B(n_1190), .Y(n_1188) );
CKINVDCx14_ASAP7_75t_R g1269 ( .A(n_1193), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1288 ( .A(n_1193), .B(n_1289), .Y(n_1288) );
O2A1O1Ixp33_ASAP7_75t_L g1194 ( .A1(n_1195), .A2(n_1197), .B(n_1198), .C(n_1205), .Y(n_1194) );
AOI21xp33_ASAP7_75t_L g1326 ( .A1(n_1195), .A2(n_1327), .B(n_1328), .Y(n_1326) );
CKINVDCx14_ASAP7_75t_R g1195 ( .A(n_1196), .Y(n_1195) );
INVx1_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
AND2x2_ASAP7_75t_L g1199 ( .A(n_1200), .B(n_1202), .Y(n_1199) );
AND2x2_ASAP7_75t_L g1254 ( .A(n_1200), .B(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1284 ( .A(n_1200), .Y(n_1284) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1200), .B(n_1249), .Y(n_1286) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_1200), .B(n_1293), .Y(n_1292) );
INVx2_ASAP7_75t_L g1200 ( .A(n_1201), .Y(n_1200) );
NAND2xp5_ASAP7_75t_L g1283 ( .A(n_1202), .B(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1202), .Y(n_1327) );
AND2x2_ASAP7_75t_L g1278 ( .A(n_1203), .B(n_1279), .Y(n_1278) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1203), .Y(n_1307) );
O2A1O1Ixp33_ASAP7_75t_L g1297 ( .A1(n_1205), .A2(n_1218), .B(n_1298), .C(n_1300), .Y(n_1297) );
INVx1_ASAP7_75t_L g1208 ( .A(n_1209), .Y(n_1208) );
AOI21xp33_ASAP7_75t_L g1290 ( .A1(n_1210), .A2(n_1291), .B(n_1292), .Y(n_1290) );
INVx1_ASAP7_75t_L g1210 ( .A(n_1211), .Y(n_1210) );
NAND2xp5_ASAP7_75t_L g1265 ( .A(n_1211), .B(n_1266), .Y(n_1265) );
NAND2xp5_ASAP7_75t_L g1325 ( .A(n_1214), .B(n_1219), .Y(n_1325) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx2_ASAP7_75t_L g1239 ( .A(n_1216), .Y(n_1239) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1216), .B(n_1219), .Y(n_1296) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1219), .Y(n_1218) );
OAI21xp5_ASAP7_75t_SL g1261 ( .A1(n_1219), .A2(n_1262), .B(n_1264), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1314 ( .A1(n_1220), .A2(n_1224), .B1(n_1315), .B2(n_1316), .Y(n_1314) );
INVx1_ASAP7_75t_L g1220 ( .A(n_1221), .Y(n_1220) );
NOR2xp33_ASAP7_75t_L g1222 ( .A(n_1223), .B(n_1225), .Y(n_1222) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_1224), .A2(n_1319), .B1(n_1320), .B2(n_1322), .Y(n_1318) );
OAI31xp33_ASAP7_75t_SL g1295 ( .A1(n_1227), .A2(n_1296), .A3(n_1297), .B(n_1301), .Y(n_1295) );
INVx3_ASAP7_75t_L g1227 ( .A(n_1228), .Y(n_1227) );
INVx2_ASAP7_75t_SL g1228 ( .A(n_1229), .Y(n_1228) );
INVx2_ASAP7_75t_SL g1270 ( .A(n_1229), .Y(n_1270) );
OAI22xp5_ASAP7_75t_SL g1230 ( .A1(n_1231), .A2(n_1232), .B1(n_1233), .B2(n_1234), .Y(n_1230) );
AOI211xp5_ASAP7_75t_L g1235 ( .A1(n_1236), .A2(n_1238), .B(n_1252), .C(n_1267), .Y(n_1235) );
INVx1_ASAP7_75t_L g1236 ( .A(n_1237), .Y(n_1236) );
OAI21xp5_ASAP7_75t_L g1238 ( .A1(n_1239), .A2(n_1240), .B(n_1242), .Y(n_1238) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1239), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1239), .B(n_1257), .Y(n_1256) );
NOR2xp33_ASAP7_75t_L g1276 ( .A(n_1239), .B(n_1277), .Y(n_1276) );
INVxp67_ASAP7_75t_L g1240 ( .A(n_1241), .Y(n_1240) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_1243), .Y(n_1268) );
INVx1_ASAP7_75t_L g1244 ( .A(n_1245), .Y(n_1244) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
OAI321xp33_ASAP7_75t_L g1267 ( .A1(n_1250), .A2(n_1268), .A3(n_1269), .B1(n_1270), .B2(n_1271), .C(n_1274), .Y(n_1267) );
OAI221xp5_ASAP7_75t_L g1252 ( .A1(n_1253), .A2(n_1256), .B1(n_1258), .B2(n_1260), .C(n_1261), .Y(n_1252) );
INVx1_ASAP7_75t_L g1253 ( .A(n_1254), .Y(n_1253) );
NAND2xp5_ASAP7_75t_L g1302 ( .A(n_1257), .B(n_1284), .Y(n_1302) );
OAI21xp5_ASAP7_75t_L g1323 ( .A1(n_1257), .A2(n_1324), .B(n_1326), .Y(n_1323) );
INVx1_ASAP7_75t_L g1258 ( .A(n_1259), .Y(n_1258) );
INVx1_ASAP7_75t_L g1262 ( .A(n_1263), .Y(n_1262) );
INVxp67_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1272), .Y(n_1271) );
NAND2xp5_ASAP7_75t_L g1274 ( .A(n_1275), .B(n_1276), .Y(n_1274) );
AOI211xp5_ASAP7_75t_L g1281 ( .A1(n_1275), .A2(n_1282), .B(n_1285), .C(n_1290), .Y(n_1281) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1275), .Y(n_1291) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1278), .Y(n_1277) );
NAND5xp2_ASAP7_75t_L g1280 ( .A(n_1281), .B(n_1295), .C(n_1308), .D(n_1309), .E(n_1323), .Y(n_1280) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1283), .Y(n_1282) );
OAI21xp5_ASAP7_75t_L g1285 ( .A1(n_1286), .A2(n_1287), .B(n_1288), .Y(n_1285) );
INVx1_ASAP7_75t_L g1300 ( .A(n_1293), .Y(n_1300) );
INVx2_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
NOR3xp33_ASAP7_75t_SL g1309 ( .A(n_1310), .B(n_1314), .C(n_1318), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
NAND2xp5_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1312), .Y(n_1328) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVxp67_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
BUFx2_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
INVxp67_ASAP7_75t_SL g1332 ( .A(n_1333), .Y(n_1332) );
HB1xp67_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx1_ASAP7_75t_L g1335 ( .A(n_1336), .Y(n_1335) );
NAND3xp33_ASAP7_75t_L g1336 ( .A(n_1337), .B(n_1355), .C(n_1358), .Y(n_1336) );
NAND2xp5_ASAP7_75t_L g1359 ( .A(n_1360), .B(n_1362), .Y(n_1359) );
HB1xp67_ASAP7_75t_L g1370 ( .A(n_1371), .Y(n_1370) );
OAI21xp5_ASAP7_75t_L g1372 ( .A1(n_1373), .A2(n_1374), .B(n_1375), .Y(n_1372) );
INVx1_ASAP7_75t_L g1375 ( .A(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1379), .Y(n_1432) );
NAND4xp75_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1400), .C(n_1412), .D(n_1420), .Y(n_1379) );
AO21x1_ASAP7_75t_L g1380 ( .A1(n_1381), .A2(n_1384), .B(n_1399), .Y(n_1380) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1385), .B(n_1396), .Y(n_1384) );
INVx2_ASAP7_75t_L g1387 ( .A(n_1388), .Y(n_1387) );
AOI22xp5_ASAP7_75t_L g1390 ( .A1(n_1391), .A2(n_1392), .B1(n_1393), .B2(n_1395), .Y(n_1390) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1392), .B(n_1407), .Y(n_1406) );
INVx2_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
AO21x1_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1408), .B(n_1410), .Y(n_1400) );
INVx1_ASAP7_75t_L g1410 ( .A(n_1411), .Y(n_1410) );
INVx1_ASAP7_75t_L g1427 ( .A(n_1428), .Y(n_1427) );
BUFx4f_ASAP7_75t_L g1434 ( .A(n_1435), .Y(n_1434) );
endmodule