module fake_jpeg_29723_n_396 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_396);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_396;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_8),
.B(n_11),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx12_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_8),
.Y(n_26)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_7),
.B(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_8),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_44),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_34),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_47),
.Y(n_87)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_34),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_29),
.Y(n_48)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_21),
.B(n_14),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_49),
.B(n_51),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_29),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_53),
.B(n_67),
.Y(n_107)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_54),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_17),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_30),
.B(n_0),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_56),
.B(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_59),
.Y(n_113)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_60),
.Y(n_110)
);

INVx2_ASAP7_75t_SL g61 ( 
.A(n_32),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g103 ( 
.A(n_61),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_30),
.B(n_1),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_16),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g127 ( 
.A(n_63),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_25),
.B(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_64),
.B(n_77),
.Y(n_124)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_31),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_65),
.Y(n_128)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_25),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g68 ( 
.A(n_24),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_68),
.B(n_75),
.Y(n_108)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_23),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_69),
.Y(n_111)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_20),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_71),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_39),
.Y(n_72)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_72),
.Y(n_135)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_74),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_15),
.B(n_1),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_15),
.B(n_33),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_78),
.Y(n_122)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_79),
.Y(n_123)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_32),
.Y(n_80)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_80),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

INVx4_ASAP7_75t_SL g82 ( 
.A(n_24),
.Y(n_82)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_82),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_83),
.Y(n_132)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_27),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_84),
.B(n_35),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_86),
.Y(n_134)
);

INVx5_ASAP7_75t_SL g86 ( 
.A(n_16),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_56),
.A2(n_62),
.B1(n_72),
.B2(n_55),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g150 ( 
.A1(n_94),
.A2(n_98),
.B1(n_112),
.B2(n_125),
.Y(n_150)
);

AND2x4_ASAP7_75t_L g95 ( 
.A(n_44),
.B(n_22),
.Y(n_95)
);

AND2x2_ASAP7_75t_SL g152 ( 
.A(n_95),
.B(n_44),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_58),
.A2(n_27),
.B1(n_41),
.B2(n_38),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_63),
.B(n_18),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_102),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_48),
.B(n_57),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_100),
.B(n_50),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_36),
.B1(n_22),
.B2(n_16),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_101),
.A2(n_46),
.B1(n_65),
.B2(n_76),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_63),
.B(n_38),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_61),
.A2(n_18),
.B1(n_41),
.B2(n_33),
.Y(n_105)
);

OA22x2_ASAP7_75t_L g180 ( 
.A1(n_105),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_71),
.A2(n_43),
.B1(n_26),
.B2(n_28),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_115),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g116 ( 
.A(n_52),
.B(n_26),
.CON(n_116),
.SN(n_116)
);

OR2x2_ASAP7_75t_SL g167 ( 
.A(n_116),
.B(n_13),
.Y(n_167)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_59),
.B(n_37),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_120),
.B(n_121),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_68),
.B(n_82),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_37),
.B1(n_35),
.B2(n_28),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_84),
.A2(n_36),
.B1(n_22),
.B2(n_4),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_129),
.B1(n_2),
.B2(n_3),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_60),
.A2(n_74),
.B1(n_73),
.B2(n_69),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_90),
.B(n_54),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_138),
.B(n_142),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_89),
.Y(n_139)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_139),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_83),
.B1(n_80),
.B2(n_78),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_140),
.A2(n_159),
.B1(n_163),
.B2(n_166),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_68),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_124),
.B(n_36),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_144),
.B(n_151),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_136),
.Y(n_146)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_136),
.Y(n_147)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_147),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_108),
.B(n_96),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_148),
.B(n_149),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_66),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_87),
.Y(n_151)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_152),
.B(n_95),
.Y(n_186)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_91),
.Y(n_153)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_153),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_93),
.B(n_36),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_154),
.B(n_157),
.Y(n_204)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx13_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_174),
.B1(n_175),
.B2(n_109),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_134),
.B(n_120),
.Y(n_157)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_158),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_50),
.B1(n_22),
.B2(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_171),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_115),
.B(n_24),
.C(n_3),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_161),
.B(n_130),
.C(n_103),
.Y(n_183)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_104),
.Y(n_162)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_162),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_163)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_109),
.Y(n_164)
);

BUFx5_ASAP7_75t_L g215 ( 
.A(n_164),
.Y(n_215)
);

BUFx4f_ASAP7_75t_SL g165 ( 
.A(n_127),
.Y(n_165)
);

INVx13_ASAP7_75t_L g212 ( 
.A(n_165),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_167),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_216)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_106),
.Y(n_168)
);

INVx13_ASAP7_75t_L g217 ( 
.A(n_168),
.Y(n_217)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_170),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_137),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_172),
.B(n_177),
.Y(n_192)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_173),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_116),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_174)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_118),
.A2(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_119),
.Y(n_176)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_176),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_103),
.B(n_6),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_137),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_114),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_179),
.A2(n_180),
.B1(n_131),
.B2(n_133),
.Y(n_195)
);

INVx8_ASAP7_75t_L g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_111),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_183),
.B(n_172),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_185),
.B(n_186),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_95),
.C(n_133),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_187),
.B(n_194),
.C(n_207),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_141),
.A2(n_92),
.B1(n_110),
.B2(n_132),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_197),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_169),
.A2(n_92),
.B1(n_110),
.B2(n_135),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_150),
.A2(n_114),
.B1(n_131),
.B2(n_135),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_95),
.C(n_119),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_195),
.B(n_208),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_169),
.A2(n_97),
.B1(n_117),
.B2(n_122),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_152),
.B(n_161),
.C(n_167),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_140),
.A2(n_117),
.B1(n_122),
.B2(n_111),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_208),
.A2(n_178),
.B1(n_145),
.B2(n_139),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_144),
.A2(n_128),
.B1(n_88),
.B2(n_11),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_211),
.B1(n_214),
.B2(n_163),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_152),
.B1(n_177),
.B2(n_159),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_180),
.A2(n_88),
.B1(n_9),
.B2(n_12),
.Y(n_214)
);

AO22x2_ASAP7_75t_L g218 ( 
.A1(n_152),
.A2(n_6),
.B1(n_13),
.B2(n_180),
.Y(n_218)
);

AO21x1_ASAP7_75t_L g252 ( 
.A1(n_218),
.A2(n_139),
.B(n_145),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_143),
.B(n_13),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_219),
.B(n_173),
.C(n_153),
.Y(n_243)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_184),
.Y(n_222)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_222),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_224),
.A2(n_244),
.B1(n_202),
.B2(n_183),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_192),
.B(n_143),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_226),
.B(n_232),
.Y(n_267)
);

INVx6_ASAP7_75t_L g227 ( 
.A(n_196),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_227),
.B(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_201),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_229),
.Y(n_271)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_230),
.B(n_234),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_216),
.A2(n_164),
.B(n_165),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_252),
.B(n_212),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_192),
.B(n_170),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_243),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_193),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g235 ( 
.A1(n_191),
.A2(n_151),
.A3(n_162),
.B1(n_146),
.B2(n_147),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_235),
.B(n_237),
.Y(n_273)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_220),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_199),
.B(n_165),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_238),
.B(n_239),
.Y(n_274)
);

CKINVDCx14_ASAP7_75t_R g239 ( 
.A(n_200),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_191),
.Y(n_240)
);

NAND3xp33_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_186),
.C(n_218),
.Y(n_261)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_210),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_241),
.B(n_242),
.Y(n_269)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_206),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_190),
.A2(n_158),
.B1(n_179),
.B2(n_181),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_187),
.B(n_168),
.C(n_155),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_245),
.B(n_251),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_196),
.A2(n_181),
.B1(n_182),
.B2(n_171),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g264 ( 
.A(n_246),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_247),
.A2(n_253),
.B1(n_198),
.B2(n_203),
.Y(n_275)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_206),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_248),
.Y(n_256)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_221),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_249),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_197),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_165),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_204),
.B(n_219),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_254),
.B(n_213),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_231),
.A2(n_207),
.B(n_216),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_255),
.A2(n_265),
.B(n_270),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_260),
.B1(n_268),
.B2(n_282),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_224),
.A2(n_202),
.B1(n_195),
.B2(n_194),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_261),
.B(n_252),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_236),
.A2(n_186),
.B(n_218),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_240),
.A2(n_195),
.B1(n_186),
.B2(n_214),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_251),
.A2(n_236),
.B(n_253),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g272 ( 
.A1(n_236),
.A2(n_195),
.B(n_198),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_272),
.A2(n_278),
.B(n_280),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_275),
.A2(n_277),
.B1(n_223),
.B2(n_244),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_253),
.A2(n_203),
.B1(n_221),
.B2(n_215),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_232),
.A2(n_213),
.B(n_212),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_279),
.B(n_226),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_223),
.A2(n_215),
.B1(n_205),
.B2(n_217),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_269),
.Y(n_283)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_283),
.Y(n_311)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_269),
.Y(n_284)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_284),
.Y(n_321)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_281),
.Y(n_285)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_285),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_263),
.B(n_225),
.C(n_233),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_286),
.B(n_299),
.C(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_281),
.Y(n_287)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_287),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_288),
.B(n_289),
.Y(n_316)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_262),
.Y(n_289)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_262),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_292),
.B(n_294),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_293),
.A2(n_296),
.B1(n_260),
.B2(n_259),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g294 ( 
.A(n_279),
.Y(n_294)
);

XNOR2x1_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_258),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_252),
.B1(n_235),
.B2(n_245),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_274),
.B(n_228),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_297),
.B(n_298),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_267),
.B(n_243),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_263),
.B(n_225),
.Y(n_299)
);

BUFx12f_ASAP7_75t_SL g300 ( 
.A(n_278),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_300),
.A2(n_301),
.B(n_303),
.Y(n_314)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_257),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_274),
.B(n_237),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_302),
.A2(n_230),
.B(n_229),
.Y(n_322)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_257),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_276),
.B(n_267),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_273),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_278),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_306),
.A2(n_255),
.B(n_272),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_307),
.A2(n_323),
.B1(n_305),
.B2(n_304),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_270),
.B1(n_276),
.B2(n_275),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_308),
.A2(n_320),
.B1(n_325),
.B2(n_293),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_318),
.C(n_319),
.Y(n_331)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_310),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_312),
.B(n_290),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_313),
.B(n_304),
.Y(n_333)
);

AOI322xp5_ASAP7_75t_L g315 ( 
.A1(n_288),
.A2(n_273),
.A3(n_265),
.B1(n_282),
.B2(n_261),
.C1(n_258),
.C2(n_268),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_315),
.B(n_316),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_299),
.B(n_258),
.C(n_271),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_286),
.B(n_271),
.C(n_277),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_291),
.A2(n_264),
.B1(n_256),
.B2(n_266),
.Y(n_320)
);

CKINVDCx16_ASAP7_75t_R g330 ( 
.A(n_322),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_296),
.A2(n_256),
.B1(n_266),
.B2(n_222),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_295),
.A2(n_284),
.B1(n_283),
.B2(n_306),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g358 ( 
.A(n_328),
.B(n_329),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_309),
.B(n_298),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_318),
.B(n_303),
.C(n_301),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_332),
.B(n_342),
.C(n_343),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_333),
.B(n_336),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_334),
.A2(n_300),
.B1(n_310),
.B2(n_321),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_335),
.B(n_341),
.Y(n_350)
);

INVx13_ASAP7_75t_L g336 ( 
.A(n_314),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_326),
.B(n_292),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_337),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_326),
.B(n_316),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_339),
.B(n_340),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_317),
.B(n_297),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_308),
.A2(n_325),
.B1(n_320),
.B2(n_321),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_319),
.B(n_289),
.C(n_290),
.Y(n_343)
);

CKINVDCx16_ASAP7_75t_R g344 ( 
.A(n_317),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_344),
.B(n_345),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_312),
.B(n_300),
.C(n_302),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_349),
.B(n_335),
.Y(n_364)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_334),
.A2(n_311),
.B1(n_307),
.B2(n_323),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_352),
.B(n_353),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_340),
.B(n_313),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_330),
.A2(n_311),
.B1(n_314),
.B2(n_327),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_354),
.B(n_357),
.Y(n_363)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_341),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_356),
.B(n_336),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_330),
.A2(n_327),
.B1(n_324),
.B2(n_285),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_324),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_359),
.Y(n_360)
);

BUFx24_ASAP7_75t_SL g361 ( 
.A(n_358),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_361),
.B(n_345),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_358),
.B(n_329),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_362),
.B(n_365),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_364),
.B(n_369),
.Y(n_372)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_355),
.B(n_331),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_367),
.B(n_368),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_355),
.B(n_331),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_351),
.B(n_332),
.Y(n_369)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_338),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_370),
.B(n_349),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_370),
.A2(n_347),
.B1(n_356),
.B2(n_346),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_373),
.B(n_375),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_364),
.B(n_343),
.C(n_352),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_376),
.B(n_377),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g378 ( 
.A(n_360),
.B(n_354),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_378),
.B(n_374),
.Y(n_385)
);

NAND3xp33_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_338),
.C(n_350),
.Y(n_379)
);

OAI21xp5_ASAP7_75t_L g383 ( 
.A1(n_379),
.A2(n_363),
.B(n_357),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_372),
.B(n_350),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_382),
.B(n_383),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_371),
.B(n_342),
.Y(n_384)
);

BUFx24_ASAP7_75t_SL g387 ( 
.A(n_384),
.Y(n_387)
);

AOI21xp33_ASAP7_75t_L g389 ( 
.A1(n_385),
.A2(n_381),
.B(n_380),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g386 ( 
.A(n_379),
.Y(n_386)
);

AOI322xp5_ASAP7_75t_L g390 ( 
.A1(n_386),
.A2(n_287),
.A3(n_376),
.B1(n_322),
.B2(n_227),
.C1(n_205),
.C2(n_217),
.Y(n_390)
);

AOI21x1_ASAP7_75t_L g391 ( 
.A1(n_389),
.A2(n_390),
.B(n_386),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_391),
.B(n_392),
.C(n_393),
.Y(n_394)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_388),
.Y(n_392)
);

OAI21x1_ASAP7_75t_L g393 ( 
.A1(n_387),
.A2(n_241),
.B(n_249),
.Y(n_393)
);

MAJx2_ASAP7_75t_L g395 ( 
.A(n_394),
.B(n_242),
.C(n_248),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_395),
.B(n_213),
.Y(n_396)
);


endmodule