module fake_jpeg_17146_n_80 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_80);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_80;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_0),
.B(n_4),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx4_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_8),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_7),
.B(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_11),
.B(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_26),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_27),
.B(n_29),
.Y(n_40)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_12),
.B(n_0),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

OR2x2_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_1),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_22),
.B(n_2),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_35),
.B(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_22),
.B(n_2),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_26),
.Y(n_37)
);

AO21x1_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_20),
.B(n_3),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_17),
.B1(n_19),
.B2(n_15),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_39),
.A2(n_25),
.B1(n_18),
.B2(n_16),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_30),
.A2(n_20),
.B(n_24),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_42),
.A2(n_47),
.B(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_44),
.B(n_45),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_32),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_30),
.A2(n_21),
.B(n_31),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_32),
.B(n_21),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_51),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_25),
.A2(n_18),
.B1(n_16),
.B2(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_34),
.B1(n_31),
.B2(n_2),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_27),
.B(n_23),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_35),
.C(n_31),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_41),
.B(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_56),
.A2(n_62),
.B1(n_46),
.B2(n_43),
.Y(n_65)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_48),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_4),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_61),
.B(n_38),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_45),
.A2(n_3),
.B1(n_5),
.B2(n_9),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_54),
.B(n_48),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_58),
.C(n_54),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_64),
.B(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_68),
.B(n_70),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_69),
.B(n_67),
.Y(n_73)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_67),
.B(n_60),
.C(n_57),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_63),
.Y(n_74)
);

AOI221xp5_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_65),
.B1(n_59),
.B2(n_53),
.C(n_40),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_75),
.B(n_72),
.Y(n_77)
);

AO22x1_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_43),
.B1(n_37),
.B2(n_5),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_77),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_76),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_79),
.Y(n_80)
);


endmodule