module fake_jpeg_12080_n_630 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_630);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_630;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_620;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_288;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_509;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_10),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_5),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g45 ( 
.A(n_1),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_0),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_10),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_18),
.B(n_3),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_15),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_0),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_6),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_59),
.Y(n_147)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_60),
.Y(n_165)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_61),
.Y(n_130)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_62),
.Y(n_142)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_63),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_64),
.B(n_73),
.Y(n_182)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_65),
.Y(n_129)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_47),
.Y(n_66)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_66),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g135 ( 
.A(n_67),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_69),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_70),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_29),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_74),
.Y(n_146)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_25),
.Y(n_75)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_75),
.Y(n_151)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

INVx3_ASAP7_75t_L g178 ( 
.A(n_76),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_77),
.Y(n_158)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g179 ( 
.A(n_78),
.Y(n_179)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_20),
.Y(n_79)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_79),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_19),
.B(n_17),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_80),
.B(n_88),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_81),
.Y(n_162)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_26),
.Y(n_83)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_83),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_20),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_84),
.Y(n_144)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_51),
.Y(n_85)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_85),
.Y(n_159)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_51),
.Y(n_86)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_87),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_19),
.B(n_1),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_89),
.B(n_93),
.Y(n_186)
);

BUFx5_ASAP7_75t_L g90 ( 
.A(n_53),
.Y(n_90)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_22),
.Y(n_91)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_91),
.Y(n_161)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_92),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_24),
.Y(n_94)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_24),
.Y(n_95)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_95),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_55),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_96),
.B(n_98),
.Y(n_193)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_35),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_97),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_55),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_27),
.Y(n_99)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_99),
.Y(n_183)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_100),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_20),
.Y(n_101)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_101),
.Y(n_150)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_22),
.Y(n_102)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_102),
.Y(n_205)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_31),
.Y(n_103)
);

INVx3_ASAP7_75t_L g191 ( 
.A(n_103),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_35),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_104),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_31),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_105),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_38),
.Y(n_106)
);

INVx5_ASAP7_75t_L g181 ( 
.A(n_106),
.Y(n_181)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_22),
.Y(n_107)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_107),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_35),
.Y(n_108)
);

INVx6_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_27),
.Y(n_109)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_109),
.Y(n_210)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_31),
.Y(n_110)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_23),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_111),
.B(n_32),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_112),
.B(n_123),
.Y(n_200)
);

BUFx3_ASAP7_75t_SL g113 ( 
.A(n_38),
.Y(n_113)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_113),
.Y(n_172)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_31),
.Y(n_114)
);

INVx3_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_28),
.Y(n_115)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_115),
.Y(n_214)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_40),
.Y(n_116)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_116),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_41),
.Y(n_117)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_40),
.Y(n_118)
);

INVx2_ASAP7_75t_SL g217 ( 
.A(n_118),
.Y(n_217)
);

BUFx2_ASAP7_75t_L g119 ( 
.A(n_38),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_119),
.Y(n_157)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_40),
.Y(n_120)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_41),
.Y(n_121)
);

INVx6_ASAP7_75t_L g166 ( 
.A(n_121),
.Y(n_166)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_41),
.Y(n_122)
);

INVx3_ASAP7_75t_SL g153 ( 
.A(n_122),
.Y(n_153)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_28),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_23),
.B(n_2),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_124),
.B(n_126),
.Y(n_206)
);

BUFx5_ASAP7_75t_L g125 ( 
.A(n_38),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g154 ( 
.A(n_125),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_34),
.Y(n_126)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_33),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g173 ( 
.A(n_127),
.B(n_45),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_40),
.Y(n_128)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_128),
.Y(n_212)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_68),
.Y(n_132)
);

BUFx2_ASAP7_75t_L g220 ( 
.A(n_132),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_79),
.B(n_57),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_134),
.B(n_138),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_120),
.B(n_57),
.Y(n_138)
);

AND2x2_ASAP7_75t_SL g140 ( 
.A(n_103),
.B(n_45),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_140),
.B(n_173),
.Y(n_229)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_113),
.Y(n_141)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_141),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_70),
.A2(n_42),
.B1(n_46),
.B2(n_43),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_145),
.A2(n_176),
.B1(n_166),
.B2(n_163),
.Y(n_286)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

BUFx2_ASAP7_75t_L g232 ( 
.A(n_148),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_61),
.A2(n_54),
.B1(n_44),
.B2(n_48),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_149),
.A2(n_52),
.B(n_33),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_113),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_167),
.B(n_177),
.Y(n_248)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_118),
.B(n_52),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_169),
.B(n_209),
.Y(n_222)
);

INVx6_ASAP7_75t_SL g171 ( 
.A(n_113),
.Y(n_171)
);

BUFx4f_ASAP7_75t_SL g263 ( 
.A(n_171),
.Y(n_263)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_71),
.Y(n_175)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_97),
.A2(n_42),
.B1(n_43),
.B2(n_46),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_119),
.B(n_49),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_122),
.A2(n_34),
.B(n_48),
.C(n_45),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_187),
.A2(n_110),
.B1(n_78),
.B2(n_45),
.Y(n_231)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_77),
.Y(n_192)
);

INVx6_ASAP7_75t_L g273 ( 
.A(n_192),
.Y(n_273)
);

INVx6_ASAP7_75t_L g195 ( 
.A(n_81),
.Y(n_195)
);

INVx6_ASAP7_75t_L g296 ( 
.A(n_195),
.Y(n_296)
);

INVx8_ASAP7_75t_L g199 ( 
.A(n_87),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_199),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_106),
.B(n_32),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_201),
.B(n_203),
.Y(n_261)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_92),
.Y(n_202)
);

INVx4_ASAP7_75t_L g266 ( 
.A(n_202),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_59),
.Y(n_203)
);

INVx6_ASAP7_75t_L g204 ( 
.A(n_104),
.Y(n_204)
);

INVx5_ASAP7_75t_L g246 ( 
.A(n_204),
.Y(n_246)
);

INVx13_ASAP7_75t_L g208 ( 
.A(n_84),
.Y(n_208)
);

BUFx8_ASAP7_75t_L g267 ( 
.A(n_208),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_128),
.B(n_49),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g213 ( 
.A(n_101),
.Y(n_213)
);

BUFx3_ASAP7_75t_L g226 ( 
.A(n_213),
.Y(n_226)
);

INVx5_ASAP7_75t_L g216 ( 
.A(n_72),
.Y(n_216)
);

INVx4_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_105),
.Y(n_218)
);

INVx4_ASAP7_75t_L g288 ( 
.A(n_218),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_219),
.B(n_7),
.Y(n_250)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_185),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g348 ( 
.A(n_221),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_184),
.A2(n_121),
.B1(n_117),
.B2(n_108),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_223),
.A2(n_284),
.B1(n_294),
.B2(n_197),
.Y(n_306)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_168),
.Y(n_224)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_224),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_200),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_234),
.Y(n_309)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_170),
.Y(n_227)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_227),
.Y(n_333)
);

OAI21xp33_ASAP7_75t_SL g337 ( 
.A1(n_228),
.A2(n_135),
.B(n_198),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_231),
.A2(n_247),
.B1(n_249),
.B2(n_254),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_169),
.A2(n_37),
.B(n_36),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g310 ( 
.A1(n_233),
.A2(n_197),
.B(n_205),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_200),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_184),
.A2(n_37),
.B(n_36),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_235),
.B(n_242),
.C(n_281),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_206),
.B(n_2),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_236),
.B(n_238),
.Y(n_301)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_237),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_4),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_239),
.Y(n_329)
);

BUFx3_ASAP7_75t_L g240 ( 
.A(n_213),
.Y(n_240)
);

INVx5_ASAP7_75t_L g303 ( 
.A(n_240),
.Y(n_303)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_147),
.Y(n_241)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_241),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_183),
.B(n_46),
.C(n_43),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_186),
.B(n_4),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_243),
.B(n_287),
.Y(n_302)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g354 ( 
.A(n_244),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g247 ( 
.A1(n_145),
.A2(n_42),
.B1(n_5),
.B2(n_6),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_187),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g305 ( 
.A(n_250),
.B(n_279),
.Y(n_305)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_179),
.Y(n_251)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_251),
.Y(n_345)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_153),
.Y(n_252)
);

INVx3_ASAP7_75t_L g304 ( 
.A(n_252),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_182),
.B(n_7),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_253),
.B(n_265),
.Y(n_300)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_210),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_254)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_130),
.Y(n_255)
);

INVxp33_ASAP7_75t_L g311 ( 
.A(n_255),
.Y(n_311)
);

AND2x2_ASAP7_75t_SL g256 ( 
.A(n_142),
.B(n_7),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g299 ( 
.A(n_256),
.B(n_283),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_193),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_257),
.B(n_275),
.Y(n_312)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_181),
.Y(n_258)
);

INVx4_ASAP7_75t_L g318 ( 
.A(n_258),
.Y(n_318)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_153),
.Y(n_260)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_260),
.Y(n_319)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_155),
.Y(n_262)
);

INVx3_ASAP7_75t_L g339 ( 
.A(n_262),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_130),
.A2(n_214),
.B1(n_188),
.B2(n_129),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_182),
.B(n_8),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_137),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_269),
.Y(n_350)
);

AOI22xp33_ASAP7_75t_SL g271 ( 
.A1(n_159),
.A2(n_164),
.B1(n_157),
.B2(n_178),
.Y(n_271)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_271),
.A2(n_274),
.B1(n_276),
.B2(n_154),
.Y(n_308)
);

BUFx10_ASAP7_75t_L g272 ( 
.A(n_172),
.Y(n_272)
);

INVx5_ASAP7_75t_L g334 ( 
.A(n_272),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g274 ( 
.A1(n_165),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_193),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_SL g276 ( 
.A1(n_174),
.A2(n_8),
.B1(n_11),
.B2(n_12),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_140),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_277),
.B(n_278),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_209),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_186),
.B(n_11),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g280 ( 
.A1(n_173),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_286),
.B1(n_199),
.B2(n_131),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_143),
.B(n_13),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_219),
.B(n_14),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_SL g355 ( 
.A(n_282),
.B(n_285),
.Y(n_355)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_161),
.Y(n_283)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_149),
.A2(n_14),
.B1(n_16),
.B2(n_160),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_146),
.B(n_16),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_151),
.B(n_215),
.Y(n_287)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_191),
.Y(n_289)
);

INVx5_ASAP7_75t_L g353 ( 
.A(n_289),
.Y(n_353)
);

CKINVDCx12_ASAP7_75t_R g290 ( 
.A(n_172),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_290),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_133),
.B(n_211),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_291),
.B(n_292),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_141),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_207),
.B(n_180),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_293),
.B(n_190),
.Y(n_325)
);

OAI22xp33_ASAP7_75t_L g294 ( 
.A1(n_136),
.A2(n_156),
.B1(n_194),
.B2(n_162),
.Y(n_294)
);

INVx3_ASAP7_75t_L g295 ( 
.A(n_132),
.Y(n_295)
);

INVx6_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_194),
.B1(n_189),
.B2(n_139),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_321),
.B1(n_327),
.B2(n_347),
.Y(n_357)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_306),
.B(n_246),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_308),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_310),
.B(n_338),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_272),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_314),
.B(n_331),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_229),
.B(n_208),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_315),
.B(n_237),
.C(n_239),
.Y(n_383)
);

AOI22xp33_ASAP7_75t_L g322 ( 
.A1(n_223),
.A2(n_131),
.B1(n_196),
.B2(n_139),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_L g377 ( 
.A1(n_322),
.A2(n_273),
.B1(n_260),
.B2(n_252),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_256),
.B(n_158),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_323),
.B(n_324),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_256),
.B(n_158),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_325),
.B(n_330),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_231),
.A2(n_152),
.B1(n_196),
.B2(n_162),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_235),
.B(n_152),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_328),
.B(n_335),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_261),
.B(n_144),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_272),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g332 ( 
.A(n_272),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_332),
.B(n_336),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_189),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_230),
.B(n_150),
.Y(n_336)
);

NAND2xp33_ASAP7_75t_SL g356 ( 
.A(n_337),
.B(n_229),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_248),
.B(n_154),
.Y(n_338)
);

CKINVDCx16_ASAP7_75t_R g340 ( 
.A(n_255),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_340),
.B(n_341),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_245),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_243),
.B(n_281),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_343),
.B(n_352),
.Y(n_381)
);

INVx8_ASAP7_75t_L g344 ( 
.A(n_259),
.Y(n_344)
);

INVx3_ASAP7_75t_SL g386 ( 
.A(n_344),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_SL g347 ( 
.A1(n_233),
.A2(n_222),
.B1(n_242),
.B2(n_269),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_236),
.A2(n_238),
.B1(n_228),
.B2(n_224),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_349),
.A2(n_262),
.B1(n_270),
.B2(n_246),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_281),
.B(n_229),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_356),
.A2(n_370),
.B(n_263),
.Y(n_435)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_313),
.Y(n_358)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_358),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_328),
.A2(n_227),
.B1(n_294),
.B2(n_296),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_359),
.A2(n_360),
.B1(n_362),
.B2(n_377),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_306),
.A2(n_259),
.B1(n_273),
.B2(n_296),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_346),
.A2(n_335),
.B1(n_302),
.B2(n_352),
.Y(n_362)
);

INVx3_ASAP7_75t_L g363 ( 
.A(n_351),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g408 ( 
.A(n_363),
.Y(n_408)
);

INVx5_ASAP7_75t_L g364 ( 
.A(n_344),
.Y(n_364)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_364),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_320),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_367),
.B(n_369),
.Y(n_415)
);

INVx4_ASAP7_75t_L g368 ( 
.A(n_351),
.Y(n_368)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_368),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g369 ( 
.A(n_310),
.Y(n_369)
);

AOI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_346),
.A2(n_263),
.B(n_283),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_241),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_371),
.B(n_315),
.C(n_324),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g372 ( 
.A(n_309),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_372),
.B(n_394),
.Y(n_439)
);

INVx5_ASAP7_75t_L g373 ( 
.A(n_318),
.Y(n_373)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_373),
.Y(n_413)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_374),
.Y(n_418)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_333),
.Y(n_378)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_378),
.Y(n_427)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_297),
.A2(n_270),
.B(n_288),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g425 ( 
.A1(n_380),
.A2(n_356),
.B(n_334),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_299),
.B(n_251),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_382),
.B(n_398),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_383),
.B(n_345),
.Y(n_426)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_384),
.A2(n_395),
.B1(n_311),
.B2(n_331),
.Y(n_404)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_333),
.Y(n_385)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

INVx13_ASAP7_75t_L g387 ( 
.A(n_307),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_387),
.Y(n_411)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_312),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_388),
.B(n_396),
.Y(n_431)
);

AOI22xp33_ASAP7_75t_L g390 ( 
.A1(n_298),
.A2(n_220),
.B1(n_268),
.B2(n_295),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g416 ( 
.A1(n_390),
.A2(n_392),
.B1(n_314),
.B2(n_348),
.Y(n_416)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_342),
.Y(n_391)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_391),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_341),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_323),
.A2(n_220),
.B1(n_268),
.B2(n_289),
.Y(n_395)
);

INVxp67_ASAP7_75t_L g396 ( 
.A(n_354),
.Y(n_396)
);

CKINVDCx12_ASAP7_75t_R g397 ( 
.A(n_334),
.Y(n_397)
);

CKINVDCx16_ASAP7_75t_R g421 ( 
.A(n_397),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_299),
.B(n_288),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_342),
.Y(n_399)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_399),
.B(n_400),
.Y(n_428)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_345),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_299),
.B(n_266),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_350),
.Y(n_420)
);

AO21x2_ASAP7_75t_L g402 ( 
.A1(n_375),
.A2(n_327),
.B(n_297),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_402),
.B(n_417),
.Y(n_462)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_404),
.Y(n_468)
);

XNOR2x1_ASAP7_75t_L g473 ( 
.A(n_405),
.B(n_426),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_362),
.B(n_316),
.C(n_343),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_410),
.B(n_412),
.C(n_383),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_301),
.C(n_350),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g446 ( 
.A(n_416),
.Y(n_446)
);

OAI32xp33_ASAP7_75t_L g417 ( 
.A1(n_375),
.A2(n_355),
.A3(n_301),
.B1(n_305),
.B2(n_317),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_357),
.A2(n_355),
.B1(n_305),
.B2(n_300),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_419),
.A2(n_395),
.B1(n_358),
.B2(n_385),
.Y(n_459)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_420),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_SL g422 ( 
.A(n_372),
.B(n_263),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_422),
.B(n_389),
.Y(n_440)
);

NAND2x1_ASAP7_75t_SL g423 ( 
.A(n_369),
.B(n_267),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g442 ( 
.A1(n_423),
.A2(n_429),
.B(n_401),
.Y(n_442)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_393),
.Y(n_424)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

OAI21xp5_ASAP7_75t_SL g460 ( 
.A1(n_425),
.A2(n_435),
.B(n_423),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_379),
.A2(n_348),
.B(n_354),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_371),
.B(n_339),
.Y(n_430)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_430),
.Y(n_453)
);

CKINVDCx16_ASAP7_75t_R g432 ( 
.A(n_376),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_365),
.Y(n_447)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_379),
.Y(n_433)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_433),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_394),
.B(n_339),
.Y(n_436)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_436),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_361),
.B(n_348),
.Y(n_437)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_437),
.Y(n_470)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_440),
.B(n_461),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_435),
.A2(n_380),
.B(n_366),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_SL g487 ( 
.A1(n_441),
.A2(n_448),
.B(n_460),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_442),
.B(n_460),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g479 ( 
.A(n_444),
.B(n_423),
.Y(n_479)
);

OAI22xp5_ASAP7_75t_SL g445 ( 
.A1(n_402),
.A2(n_357),
.B1(n_366),
.B2(n_361),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_445),
.A2(n_451),
.B1(n_457),
.B2(n_438),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_SL g492 ( 
.A(n_447),
.B(n_411),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_SL g448 ( 
.A(n_412),
.B(n_381),
.C(n_384),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_381),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g484 ( 
.A(n_450),
.B(n_452),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_402),
.A2(n_392),
.B1(n_382),
.B2(n_384),
.Y(n_451)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_318),
.Y(n_452)
);

NOR4xp25_ASAP7_75t_L g454 ( 
.A(n_417),
.B(n_433),
.C(n_437),
.D(n_403),
.Y(n_454)
);

AOI322xp5_ASAP7_75t_SL g482 ( 
.A1(n_454),
.A2(n_414),
.A3(n_428),
.B1(n_434),
.B2(n_427),
.C1(n_418),
.C2(n_406),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_436),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_455),
.B(n_463),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_303),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_456),
.B(n_471),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_402),
.A2(n_398),
.B1(n_359),
.B2(n_360),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_459),
.A2(n_467),
.B1(n_391),
.B2(n_400),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_424),
.B(n_378),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_428),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_464),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_426),
.B(n_410),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_472),
.C(n_420),
.Y(n_476)
);

AND2x6_ASAP7_75t_L g466 ( 
.A(n_419),
.B(n_387),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_466),
.B(n_474),
.Y(n_499)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_402),
.A2(n_377),
.B1(n_374),
.B2(n_386),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_431),
.B(n_303),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_405),
.B(n_430),
.C(n_403),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_428),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_440),
.B(n_421),
.Y(n_475)
);

NOR2xp33_ASAP7_75t_SL g531 ( 
.A(n_475),
.B(n_483),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_476),
.B(n_479),
.C(n_495),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g480 ( 
.A(n_473),
.B(n_429),
.Y(n_480)
);

XOR2xp5_ASAP7_75t_L g518 ( 
.A(n_480),
.B(n_490),
.Y(n_518)
);

FAx1_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_425),
.CI(n_402),
.CON(n_481),
.SN(n_481)
);

OAI21xp5_ASAP7_75t_L g509 ( 
.A1(n_481),
.A2(n_505),
.B(n_507),
.Y(n_509)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_482),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_461),
.B(n_458),
.Y(n_483)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_458),
.Y(n_485)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_485),
.Y(n_528)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_470),
.Y(n_488)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_488),
.Y(n_535)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_470),
.Y(n_489)
);

INVx1_ASAP7_75t_SL g511 ( 
.A(n_489),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_414),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_449),
.B(n_411),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_491),
.B(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_449),
.B(n_407),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_494),
.B(n_496),
.Y(n_520)
);

XNOR2xp5_ASAP7_75t_L g495 ( 
.A(n_444),
.B(n_434),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_472),
.B(n_459),
.Y(n_496)
);

NOR2x1_ASAP7_75t_L g497 ( 
.A(n_443),
.B(n_427),
.Y(n_497)
);

NOR2xp33_ASAP7_75t_L g529 ( 
.A(n_497),
.B(n_464),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_462),
.A2(n_406),
.B1(n_418),
.B2(n_438),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_498),
.A2(n_501),
.B1(n_451),
.B2(n_445),
.Y(n_523)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_500),
.A2(n_453),
.B1(n_467),
.B2(n_446),
.Y(n_512)
);

OAI22xp5_ASAP7_75t_L g502 ( 
.A1(n_446),
.A2(n_409),
.B1(n_413),
.B2(n_408),
.Y(n_502)
);

HB1xp67_ASAP7_75t_L g526 ( 
.A(n_502),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_455),
.B(n_409),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g534 ( 
.A(n_503),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_443),
.B(n_399),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_504),
.B(n_506),
.Y(n_516)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_469),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_442),
.B(n_386),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_505),
.A2(n_441),
.B(n_462),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_510),
.B(n_517),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g549 ( 
.A1(n_512),
.A2(n_527),
.B1(n_506),
.B2(n_503),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_SL g513 ( 
.A(n_480),
.B(n_465),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g539 ( 
.A(n_513),
.B(n_532),
.Y(n_539)
);

OAI22xp33_ASAP7_75t_SL g515 ( 
.A1(n_493),
.A2(n_468),
.B1(n_469),
.B2(n_466),
.Y(n_515)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_515),
.Y(n_537)
);

INVx6_ASAP7_75t_L g517 ( 
.A(n_492),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_485),
.B(n_474),
.Y(n_521)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_521),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_477),
.B(n_463),
.Y(n_522)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_522),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_SL g551 ( 
.A1(n_523),
.A2(n_504),
.B1(n_497),
.B2(n_484),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_505),
.A2(n_448),
.B(n_468),
.Y(n_524)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_524),
.A2(n_396),
.B(n_373),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_476),
.B(n_453),
.Y(n_525)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_525),
.B(n_530),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g527 ( 
.A1(n_500),
.A2(n_468),
.B1(n_457),
.B2(n_464),
.Y(n_527)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_529),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g530 ( 
.A(n_495),
.B(n_413),
.Y(n_530)
);

XNOR2xp5_ASAP7_75t_SL g532 ( 
.A(n_479),
.B(n_245),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_477),
.B(n_408),
.Y(n_533)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_533),
.Y(n_553)
);

OAI22xp33_ASAP7_75t_L g536 ( 
.A1(n_534),
.A2(n_499),
.B1(n_481),
.B2(n_489),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_536),
.A2(n_550),
.B1(n_551),
.B2(n_527),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_519),
.B(n_490),
.C(n_507),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g560 ( 
.A(n_538),
.B(n_541),
.C(n_546),
.Y(n_560)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_507),
.C(n_487),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_512),
.A2(n_499),
.B1(n_498),
.B2(n_481),
.Y(n_543)
);

OAI22xp5_ASAP7_75t_SL g573 ( 
.A1(n_543),
.A2(n_549),
.B1(n_523),
.B2(n_526),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_525),
.B(n_487),
.C(n_488),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_508),
.B(n_493),
.Y(n_547)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_547),
.Y(n_564)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_522),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g552 ( 
.A1(n_514),
.A2(n_478),
.B1(n_486),
.B2(n_408),
.Y(n_552)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_552),
.Y(n_571)
);

XNOR2x1_ASAP7_75t_L g554 ( 
.A(n_518),
.B(n_486),
.Y(n_554)
);

XOR2xp5_ASAP7_75t_L g566 ( 
.A(n_554),
.B(n_509),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_530),
.B(n_363),
.C(n_386),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g563 ( 
.A(n_555),
.B(n_557),
.C(n_511),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g576 ( 
.A(n_556),
.Y(n_576)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_513),
.B(n_329),
.C(n_326),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_521),
.B(n_364),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_533),
.Y(n_561)
);

AO221x1_ASAP7_75t_L g559 ( 
.A1(n_548),
.A2(n_520),
.B1(n_537),
.B2(n_542),
.C(n_544),
.Y(n_559)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_559),
.Y(n_586)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_561),
.Y(n_589)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_540),
.B(n_518),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_562),
.B(n_572),
.Y(n_580)
);

XNOR2xp5_ASAP7_75t_L g579 ( 
.A(n_563),
.B(n_567),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_551),
.B(n_531),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g588 ( 
.A(n_565),
.B(n_569),
.Y(n_588)
);

XOR2xp5_ASAP7_75t_L g581 ( 
.A(n_566),
.B(n_574),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g567 ( 
.A(n_540),
.B(n_524),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g585 ( 
.A1(n_568),
.A2(n_553),
.B1(n_556),
.B2(n_516),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_SL g569 ( 
.A(n_546),
.B(n_517),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_SL g570 ( 
.A(n_543),
.B(n_509),
.Y(n_570)
);

NOR2xp67_ASAP7_75t_L g577 ( 
.A(n_570),
.B(n_549),
.Y(n_577)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_558),
.Y(n_572)
);

AOI22xp5_ASAP7_75t_L g578 ( 
.A1(n_573),
.A2(n_536),
.B1(n_545),
.B2(n_558),
.Y(n_578)
);

XNOR2xp5_ASAP7_75t_L g574 ( 
.A(n_554),
.B(n_510),
.Y(n_574)
);

XOR2xp5_ASAP7_75t_L g575 ( 
.A(n_538),
.B(n_539),
.Y(n_575)
);

XOR2xp5_ASAP7_75t_L g582 ( 
.A(n_575),
.B(n_560),
.Y(n_582)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_577),
.Y(n_600)
);

OAI22xp5_ASAP7_75t_SL g594 ( 
.A1(n_578),
.A2(n_590),
.B1(n_592),
.B2(n_589),
.Y(n_594)
);

XNOR2xp5_ASAP7_75t_L g593 ( 
.A(n_582),
.B(n_583),
.Y(n_593)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_541),
.Y(n_583)
);

NAND3xp33_ASAP7_75t_SL g584 ( 
.A(n_576),
.B(n_516),
.C(n_558),
.Y(n_584)
);

OAI21xp5_ASAP7_75t_SL g601 ( 
.A1(n_584),
.A2(n_587),
.B(n_578),
.Y(n_601)
);

XOR2xp5_ASAP7_75t_L g604 ( 
.A(n_585),
.B(n_311),
.Y(n_604)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_576),
.A2(n_535),
.B(n_511),
.Y(n_587)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_587),
.A2(n_590),
.B1(n_586),
.B2(n_581),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g590 ( 
.A1(n_571),
.A2(n_535),
.B1(n_528),
.B2(n_555),
.Y(n_590)
);

OAI22xp5_ASAP7_75t_L g591 ( 
.A1(n_564),
.A2(n_557),
.B1(n_532),
.B2(n_539),
.Y(n_591)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_591),
.B(n_575),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_561),
.Y(n_592)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_592),
.B(n_560),
.Y(n_595)
);

XNOR2xp5_ASAP7_75t_SL g608 ( 
.A(n_594),
.B(n_603),
.Y(n_608)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_595),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_596),
.B(n_599),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_588),
.B(n_563),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_597),
.B(n_598),
.Y(n_613)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_579),
.B(n_566),
.C(n_574),
.Y(n_598)
);

XNOR2xp5_ASAP7_75t_L g599 ( 
.A(n_579),
.B(n_570),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g609 ( 
.A1(n_601),
.A2(n_582),
.B(n_226),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g602 ( 
.A(n_580),
.B(n_368),
.Y(n_602)
);

CKINVDCx14_ASAP7_75t_R g611 ( 
.A(n_602),
.Y(n_611)
);

MAJIxp5_ASAP7_75t_L g607 ( 
.A(n_604),
.B(n_581),
.C(n_583),
.Y(n_607)
);

AOI22xp5_ASAP7_75t_SL g615 ( 
.A1(n_607),
.A2(n_598),
.B1(n_594),
.B2(n_593),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_609),
.A2(n_610),
.B(n_612),
.Y(n_618)
);

MAJIxp5_ASAP7_75t_L g610 ( 
.A(n_593),
.B(n_304),
.C(n_319),
.Y(n_610)
);

AOI21xp33_ASAP7_75t_L g612 ( 
.A1(n_600),
.A2(n_267),
.B(n_226),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_611),
.B(n_595),
.Y(n_614)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_614),
.Y(n_623)
);

XNOR2xp5_ASAP7_75t_L g622 ( 
.A(n_615),
.B(n_616),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_613),
.B(n_599),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_605),
.A2(n_604),
.B(n_240),
.Y(n_617)
);

INVxp67_ASAP7_75t_L g620 ( 
.A(n_617),
.Y(n_620)
);

AOI322xp5_ASAP7_75t_L g619 ( 
.A1(n_606),
.A2(n_353),
.A3(n_329),
.B1(n_326),
.B2(n_258),
.C1(n_221),
.C2(n_244),
.Y(n_619)
);

O2A1O1Ixp33_ASAP7_75t_SL g621 ( 
.A1(n_619),
.A2(n_267),
.B(n_353),
.C(n_610),
.Y(n_621)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_621),
.A2(n_266),
.B1(n_232),
.B2(n_304),
.Y(n_625)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_623),
.B(n_607),
.Y(n_624)
);

AOI21x1_ASAP7_75t_SL g626 ( 
.A1(n_624),
.A2(n_625),
.B(n_618),
.Y(n_626)
);

AO21x1_ASAP7_75t_L g627 ( 
.A1(n_626),
.A2(n_620),
.B(n_622),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_627),
.B(n_608),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g629 ( 
.A(n_628),
.B(n_608),
.Y(n_629)
);

AOI21xp5_ASAP7_75t_L g630 ( 
.A1(n_629),
.A2(n_319),
.B(n_232),
.Y(n_630)
);


endmodule