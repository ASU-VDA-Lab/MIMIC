module fake_netlist_5_516_n_96 (n_29, n_16, n_0, n_12, n_9, n_36, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_28, n_21, n_40, n_34, n_38, n_4, n_32, n_35, n_11, n_17, n_19, n_7, n_37, n_15, n_26, n_30, n_20, n_5, n_33, n_14, n_2, n_31, n_23, n_13, n_3, n_6, n_39, n_96);

input n_29;
input n_16;
input n_0;
input n_12;
input n_9;
input n_36;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_28;
input n_21;
input n_40;
input n_34;
input n_38;
input n_4;
input n_32;
input n_35;
input n_11;
input n_17;
input n_19;
input n_7;
input n_37;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_14;
input n_2;
input n_31;
input n_23;
input n_13;
input n_3;
input n_6;
input n_39;

output n_96;

wire n_91;
wire n_82;
wire n_86;
wire n_83;
wire n_61;
wire n_90;
wire n_75;
wire n_65;
wire n_78;
wire n_74;
wire n_57;
wire n_66;
wire n_60;
wire n_43;
wire n_58;
wire n_69;
wire n_42;
wire n_45;
wire n_46;
wire n_94;
wire n_80;
wire n_73;
wire n_92;
wire n_84;
wire n_79;
wire n_47;
wire n_53;
wire n_44;
wire n_62;
wire n_71;
wire n_85;
wire n_95;
wire n_59;
wire n_55;
wire n_49;
wire n_54;
wire n_67;
wire n_76;
wire n_87;
wire n_64;
wire n_77;
wire n_81;
wire n_89;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_41;
wire n_56;
wire n_51;
wire n_63;
wire n_48;
wire n_50;
wire n_52;
wire n_88;

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22x1_ASAP7_75t_SL g42 ( 
.A1(n_38),
.A2(n_22),
.B1(n_24),
.B2(n_14),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_13),
.B(n_32),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

AND2x4_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_21),
.Y(n_50)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_19),
.Y(n_51)
);

AND2x2_ASAP7_75t_SL g52 ( 
.A(n_3),
.B(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_5),
.B(n_20),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_27),
.B(n_16),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_8),
.B(n_31),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_6),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_25),
.Y(n_60)
);

NOR3xp33_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_0),
.C(n_1),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_1),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_2),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_60),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

BUFx6f_ASAP7_75t_SL g68 ( 
.A(n_50),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

OR2x2_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_53),
.Y(n_70)
);

AO31x2_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_45),
.A3(n_44),
.B(n_43),
.Y(n_71)
);

AOI21x1_ASAP7_75t_L g72 ( 
.A1(n_66),
.A2(n_58),
.B(n_56),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_65),
.A2(n_49),
.B(n_55),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_67),
.A2(n_46),
.B(n_52),
.Y(n_74)
);

AO21x2_ASAP7_75t_L g75 ( 
.A1(n_73),
.A2(n_61),
.B(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_68),
.B1(n_60),
.B2(n_48),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_48),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_75),
.B(n_68),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_78),
.B(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_77),
.B(n_72),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_79),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_83),
.Y(n_85)
);

AND2x4_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_82),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_76),
.B(n_42),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_85),
.A2(n_80),
.B(n_87),
.Y(n_88)
);

OAI32xp33_ASAP7_75t_L g89 ( 
.A1(n_86),
.A2(n_9),
.A3(n_11),
.B1(n_15),
.B2(n_17),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_88),
.Y(n_90)
);

NOR3xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_89),
.C(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_90),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_18),
.B1(n_26),
.B2(n_29),
.Y(n_93)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_91),
.Y(n_94)
);

NOR2xp67_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_33),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_93),
.B(n_37),
.Y(n_96)
);


endmodule