module real_jpeg_20256_n_17 (n_5, n_4, n_8, n_0, n_12, n_306, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_306;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_286;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_237;
wire n_174;
wire n_87;
wire n_255;
wire n_40;
wire n_173;
wire n_243;
wire n_105;
wire n_299;
wire n_115;
wire n_197;
wire n_98;
wire n_27;
wire n_56;
wire n_293;
wire n_48;
wire n_164;
wire n_184;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_18;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_298;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_296;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_205;
wire n_110;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_70;
wire n_80;
wire n_41;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_240;
wire n_125;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_187;
wire n_97;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_244;
wire n_167;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_213;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_206;
wire n_210;
wire n_127;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_0),
.A2(n_27),
.B1(n_36),
.B2(n_96),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_0),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g133 ( 
.A1(n_0),
.A2(n_48),
.B1(n_51),
.B2(n_96),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_0),
.A2(n_65),
.B1(n_66),
.B2(n_96),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_0),
.A2(n_33),
.B1(n_34),
.B2(n_96),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_27),
.B1(n_36),
.B2(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_1),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_1),
.A2(n_65),
.B1(n_66),
.B2(n_117),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g183 ( 
.A1(n_1),
.A2(n_48),
.B1(n_51),
.B2(n_117),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_1),
.A2(n_33),
.B1(n_34),
.B2(n_117),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_2),
.A2(n_33),
.B1(n_34),
.B2(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_2),
.A2(n_48),
.B1(n_51),
.B2(n_57),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_2),
.A2(n_57),
.B1(n_65),
.B2(n_66),
.Y(n_109)
);

A2O1A1O1Ixp25_ASAP7_75t_L g130 ( 
.A1(n_3),
.A2(n_51),
.B(n_61),
.C(n_131),
.D(n_132),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_3),
.B(n_51),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_3),
.B(n_47),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_3),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g171 ( 
.A1(n_3),
.A2(n_84),
.B(n_150),
.Y(n_171)
);

A2O1A1O1Ixp25_ASAP7_75t_L g184 ( 
.A1(n_3),
.A2(n_33),
.B(n_44),
.C(n_185),
.D(n_186),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_33),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_3),
.B(n_119),
.Y(n_211)
);

AOI21xp33_ASAP7_75t_L g227 ( 
.A1(n_3),
.A2(n_32),
.B(n_34),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_3),
.A2(n_27),
.B1(n_36),
.B2(n_166),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g35 ( 
.A1(n_4),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_4),
.A2(n_33),
.B1(n_34),
.B2(n_37),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g196 ( 
.A1(n_4),
.A2(n_37),
.B1(n_65),
.B2(n_66),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_4),
.A2(n_37),
.B1(n_48),
.B2(n_51),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_5),
.A2(n_48),
.B1(n_51),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_5),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_5),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_7),
.Y(n_85)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_7),
.B(n_151),
.Y(n_150)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_9),
.A2(n_48),
.B1(n_51),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_9),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_9),
.A2(n_65),
.B1(n_66),
.B2(n_145),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_9),
.A2(n_33),
.B1(n_34),
.B2(n_145),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_9),
.A2(n_27),
.B1(n_36),
.B2(n_145),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_10),
.A2(n_33),
.B1(n_34),
.B2(n_54),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_10),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_10),
.A2(n_48),
.B1(n_51),
.B2(n_54),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g230 ( 
.A1(n_10),
.A2(n_54),
.B1(n_65),
.B2(n_66),
.Y(n_230)
);

BUFx12_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g38 ( 
.A1(n_12),
.A2(n_27),
.B1(n_36),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_12),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_12),
.A2(n_33),
.B1(n_34),
.B2(n_39),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_12),
.A2(n_39),
.B1(n_48),
.B2(n_51),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_12),
.A2(n_39),
.B1(n_65),
.B2(n_66),
.Y(n_210)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_16),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_122),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_120),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_98),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_20),
.B(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_80),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_72),
.B2(n_73),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_40),
.B2(n_41),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_25),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_31),
.B1(n_35),
.B2(n_38),
.Y(n_25)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_26),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_26),
.A2(n_116),
.B(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_26),
.A2(n_31),
.B1(n_116),
.B2(n_252),
.Y(n_272)
);

A2O1A1Ixp33_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_27),
.B(n_29),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g226 ( 
.A1(n_27),
.A2(n_29),
.B(n_166),
.C(n_227),
.Y(n_226)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_31)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_29),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_31),
.A2(n_35),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_31),
.Y(n_119)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_31),
.A2(n_94),
.B(n_252),
.Y(n_251)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g44 ( 
.A1(n_34),
.A2(n_45),
.B(n_46),
.C(n_47),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_34),
.B(n_45),
.Y(n_46)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_58),
.B1(n_59),
.B2(n_71),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_42),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_43),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_43),
.A2(n_55),
.B1(n_205),
.B2(n_240),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_43),
.A2(n_240),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_44),
.A2(n_47),
.B1(n_53),
.B2(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_44),
.A2(n_47),
.B1(n_75),
.B2(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_44),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_45),
.A2(n_48),
.B1(n_50),
.B2(n_51),
.Y(n_47)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_46),
.Y(n_193)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g61 ( 
.A1(n_48),
.A2(n_62),
.B(n_63),
.C(n_64),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_48),
.B(n_62),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_48),
.B(n_50),
.Y(n_192)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_51),
.A2(n_185),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_55),
.B(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_55),
.A2(n_205),
.B(n_206),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_55),
.A2(n_206),
.B(n_270),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

AOI21xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_68),
.B(n_69),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_60),
.A2(n_68),
.B1(n_78),
.B2(n_91),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_60),
.A2(n_68),
.B1(n_91),
.B2(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_60),
.A2(n_68),
.B1(n_144),
.B2(n_183),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_60),
.A2(n_183),
.B(n_218),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_60),
.A2(n_68),
.B1(n_111),
.B2(n_237),
.Y(n_260)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_64),
.B1(n_77),
.B2(n_79),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_61),
.B(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g67 ( 
.A(n_62),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_62),
.B(n_66),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_63),
.A2(n_65),
.B1(n_136),
.B2(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_85),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_66),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_68),
.B(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_68),
.A2(n_144),
.B(n_146),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g165 ( 
.A(n_68),
.B(n_166),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g236 ( 
.A1(n_68),
.A2(n_146),
.B(n_237),
.Y(n_236)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_69),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_73),
.A2(n_74),
.B(n_76),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_76),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_92),
.B(n_93),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_82),
.B1(n_100),
.B2(n_102),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_83),
.Y(n_92)
);

AOI22x1_ASAP7_75t_SL g100 ( 
.A1(n_83),
.A2(n_92),
.B1(n_93),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_83),
.A2(n_90),
.B1(n_92),
.B2(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_86),
.B(n_89),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_84),
.A2(n_85),
.B1(n_89),
.B2(n_109),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_84),
.A2(n_149),
.B(n_150),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_84),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_84),
.B(n_152),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_84),
.A2(n_85),
.B1(n_196),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_84),
.A2(n_88),
.B1(n_210),
.B2(n_230),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_84),
.A2(n_86),
.B1(n_109),
.B2(n_230),
.Y(n_259)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_85),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_85),
.A2(n_157),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_85),
.B(n_166),
.Y(n_173)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g194 ( 
.A1(n_87),
.A2(n_169),
.B(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_90),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_93),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_95),
.B(n_119),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_97),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.C(n_105),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_292),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_99),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_100),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_105),
.A2(n_106),
.B1(n_290),
.B2(n_291),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.C(n_114),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_107),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_110),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_108),
.B(n_110),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_112),
.A2(n_114),
.B1(n_115),
.B2(n_285),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_112),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_113),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_118),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI321xp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_280),
.A3(n_293),
.B1(n_299),
.B2(n_304),
.C(n_306),
.Y(n_122)
);

NOR3xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_246),
.C(n_276),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_220),
.B(n_245),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_199),
.B(n_219),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_177),
.B(n_198),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_128),
.A2(n_153),
.B(n_176),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_138),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_129),
.B(n_138),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_130),
.B(n_134),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g162 ( 
.A(n_130),
.Y(n_162)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_132),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_148),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_142),
.B2(n_143),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_140),
.B(n_143),
.C(n_148),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_149),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_163),
.B(n_175),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_161),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_155),
.B(n_161),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_164),
.A2(n_170),
.B(n_174),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_167),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_165),
.B(n_167),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_178),
.B(n_179),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_190),
.B2(n_197),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_184),
.B1(n_188),
.B2(n_189),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_182),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_184),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_184),
.B(n_189),
.C(n_197),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g207 ( 
.A(n_187),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_190),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_200),
.B(n_201),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_215),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_216),
.C(n_217),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_208),
.B2(n_214),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_203),
.B(n_211),
.C(n_212),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_208),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_212),
.B2(n_213),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_209),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_211),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_221),
.B(n_222),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_231),
.B1(n_232),
.B2(n_233),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_224),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_224),
.B(n_233),
.C(n_234),
.Y(n_277)
);

AOI22x1_ASAP7_75t_SL g224 ( 
.A1(n_225),
.A2(n_226),
.B1(n_228),
.B2(n_229),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_229),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_226),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g233 ( 
.A(n_231),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_242),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_238),
.B1(n_239),
.B2(n_241),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_236),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_241),
.C(n_242),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g300 ( 
.A1(n_247),
.A2(n_301),
.B(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_262),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_248),
.B(n_262),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_258),
.C(n_261),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_279),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_257),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_253),
.B1(n_254),
.B2(n_256),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_253),
.B(n_256),
.C(n_257),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_258),
.B(n_261),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_260),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_274),
.B2(n_275),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_265),
.B(n_266),
.C(n_275),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_267),
.B(n_271),
.C(n_273),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_269),
.A2(n_271),
.B1(n_272),
.B2(n_273),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_269),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_272),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_274),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_277),
.B(n_278),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_289),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_281),
.B(n_289),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_286),
.C(n_288),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_283),
.B1(n_286),
.B2(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_286),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_294),
.A2(n_300),
.B(n_303),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_295),
.B(n_296),
.Y(n_303)
);


endmodule