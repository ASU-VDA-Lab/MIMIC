module real_jpeg_6011_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_288;
wire n_78;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_412;
wire n_155;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_487;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_375;
wire n_196;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

INVx8_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_1),
.B(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_1),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_1),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_1),
.B(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_1),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_1),
.B(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_1),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_2),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_259),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_2),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_2),
.B(n_307),
.Y(n_306)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_2),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_2),
.B(n_288),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_2),
.B(n_431),
.Y(n_430)
);

AND2x2_ASAP7_75t_L g233 ( 
.A(n_3),
.B(n_234),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_3),
.A2(n_280),
.B(n_282),
.Y(n_279)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_3),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_3),
.B(n_352),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_3),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_3),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_3),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_3),
.B(n_440),
.Y(n_439)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_4),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_4),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_4),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_5),
.B(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_218),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_5),
.B(n_241),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_5),
.B(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_5),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_5),
.B(n_413),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_5),
.B(n_454),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_6),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_6),
.B(n_312),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_6),
.B(n_368),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_6),
.B(n_399),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_6),
.B(n_303),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_6),
.B(n_288),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_6),
.B(n_436),
.Y(n_435)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_8),
.Y(n_145)
);

INVx8_ASAP7_75t_L g232 ( 
.A(n_8),
.Y(n_232)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_8),
.Y(n_286)
);

BUFx5_ASAP7_75t_L g440 ( 
.A(n_8),
.Y(n_440)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_9),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_9),
.Y(n_281)
);

AND2x2_ASAP7_75t_SL g25 ( 
.A(n_10),
.B(n_26),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_10),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_10),
.B(n_64),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_10),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g132 ( 
.A(n_10),
.B(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_10),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_10),
.B(n_193),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_10),
.B(n_229),
.Y(n_228)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_12),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g183 ( 
.A(n_12),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_12),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_12),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_13),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_13),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_13),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_13),
.B(n_196),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_13),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_13),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_13),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_13),
.B(n_349),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g21 ( 
.A(n_14),
.B(n_22),
.Y(n_21)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_14),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_14),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_14),
.B(n_112),
.Y(n_111)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_14),
.B(n_145),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g149 ( 
.A(n_15),
.Y(n_149)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_15),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_15),
.Y(n_288)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

O2A1O1Ixp33_ASAP7_75t_SL g17 ( 
.A1(n_18),
.A2(n_101),
.B(n_117),
.C(n_495),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_31),
.Y(n_18)
);

FAx1_ASAP7_75t_SL g92 ( 
.A(n_19),
.B(n_93),
.CI(n_94),
.CON(n_92),
.SN(n_92)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_25),
.C(n_27),
.Y(n_19)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_20),
.A2(n_21),
.B1(n_27),
.B2(n_71),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_20),
.A2(n_21),
.B1(n_97),
.B2(n_99),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g495 ( 
.A(n_20),
.B(n_39),
.C(n_97),
.Y(n_495)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_21),
.B(n_178),
.C(n_182),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_21),
.B(n_224),
.Y(n_223)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_24),
.Y(n_76)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_24),
.Y(n_155)
);

BUFx5_ASAP7_75t_L g219 ( 
.A(n_24),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_24),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_25),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_25),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_25),
.A2(n_83),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_25),
.B(n_132),
.C(n_135),
.Y(n_161)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_26),
.Y(n_343)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_36),
.B1(n_71),
.B2(n_72),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_27),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_27),
.B(n_227),
.C(n_233),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_27),
.A2(n_71),
.B1(n_315),
.B2(n_316),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_29),
.Y(n_27)
);

OR2x2_ASAP7_75t_L g36 ( 
.A(n_28),
.B(n_37),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_30),
.Y(n_65)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_30),
.Y(n_131)
);

INVx3_ASAP7_75t_L g307 ( 
.A(n_30),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_92),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_78),
.C(n_79),
.Y(n_32)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_33),
.B(n_493),
.Y(n_492)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_57),
.C(n_68),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_34),
.B(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_35),
.B(n_52),
.C(n_55),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.C(n_42),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_36),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_71),
.C(n_77),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_36),
.A2(n_72),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_36),
.A2(n_72),
.B1(n_257),
.B2(n_258),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_38),
.Y(n_122)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_38),
.Y(n_134)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_38),
.Y(n_238)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_38),
.Y(n_305)
);

BUFx3_ASAP7_75t_L g395 ( 
.A(n_38),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_39),
.A2(n_95),
.B1(n_96),
.B2(n_100),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_39),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_39),
.A2(n_42),
.B1(n_43),
.B2(n_100),
.Y(n_160)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_41),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_42),
.A2(n_43),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_42),
.B(n_111),
.C(n_118),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_42),
.A2(n_43),
.B1(n_306),
.B2(n_364),
.Y(n_363)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_43),
.B(n_302),
.C(n_306),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_47),
.A2(n_52),
.B1(n_55),
.B2(n_56),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_47),
.Y(n_55)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g242 ( 
.A(n_51),
.Y(n_242)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_51),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_52),
.Y(n_56)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_57),
.B(n_68),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_58),
.B(n_62),
.C(n_66),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_58),
.A2(n_62),
.B1(n_63),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_58),
.Y(n_139)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_62),
.A2(n_63),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_63),
.B(n_144),
.C(n_192),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_65),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_66),
.B(n_138),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_69),
.A2(n_70),
.B1(n_73),
.B2(n_77),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_72),
.B(n_257),
.C(n_262),
.Y(n_256)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_73),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_73),
.B(n_118),
.C(n_120),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_73),
.A2(n_77),
.B1(n_120),
.B2(n_176),
.Y(n_175)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_78),
.B(n_79),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_84),
.B1(n_85),
.B2(n_91),
.Y(n_79)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_86),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_87),
.B(n_88),
.C(n_91),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g496 ( 
.A(n_92),
.Y(n_496)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_97),
.Y(n_99)
);

MAJx2_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_191),
.C(n_195),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_97),
.A2(n_99),
.B1(n_152),
.B2(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_97),
.A2(n_99),
.B1(n_195),
.B2(n_245),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_99),
.B(n_142),
.C(n_152),
.Y(n_141)
);

AO21x1_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_490),
.B(n_494),
.Y(n_101)
);

OAI21xp33_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_247),
.B(n_487),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_203),
.Y(n_103)
);

AOI21xp33_ASAP7_75t_SL g487 ( 
.A1(n_104),
.A2(n_488),
.B(n_489),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_165),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_105),
.B(n_165),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_156),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_106),
.B(n_157),
.C(n_163),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_137),
.C(n_140),
.Y(n_106)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_107),
.B(n_167),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_119),
.C(n_123),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_108),
.B(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_113),
.B1(n_117),
.B2(n_118),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g117 ( 
.A(n_111),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_113),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_113),
.A2(n_118),
.B1(n_174),
.B2(n_175),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_113),
.B(n_228),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_113),
.A2(n_118),
.B1(n_227),
.B2(n_228),
.Y(n_455)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_114),
.Y(n_222)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_119),
.B(n_123),
.Y(n_208)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_120),
.Y(n_176)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_132),
.B1(n_135),
.B2(n_136),
.Y(n_125)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_126),
.Y(n_135)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx8_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_130),
.Y(n_272)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_131),
.Y(n_400)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_132),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_132),
.B(n_217),
.Y(n_255)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_136),
.B(n_216),
.C(n_220),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_137),
.A2(n_140),
.B1(n_141),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_137),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

OA22x2_ASAP7_75t_L g199 ( 
.A1(n_142),
.A2(n_143),
.B1(n_200),
.B2(n_202),
.Y(n_199)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_146),
.C(n_150),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_144),
.A2(n_150),
.B1(n_186),
.B2(n_187),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_144),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_144),
.A2(n_186),
.B1(n_192),
.B2(n_214),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_144),
.A2(n_186),
.B1(n_412),
.B2(n_414),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_144),
.B(n_414),
.Y(n_456)
);

INVx4_ASAP7_75t_L g432 ( 
.A(n_145),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_146),
.A2(n_185),
.B1(n_188),
.B2(n_189),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_146),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_146),
.B(n_269),
.C(n_273),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_146),
.A2(n_188),
.B1(n_269),
.B2(n_339),
.Y(n_338)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_152),
.Y(n_201)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_155),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_163),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_161),
.C(n_162),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_162),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.C(n_171),
.Y(n_165)
);

FAx1_ASAP7_75t_SL g246 ( 
.A(n_166),
.B(n_169),
.CI(n_171),
.CON(n_246),
.SN(n_246)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_190),
.C(n_199),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_172),
.B(n_206),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_177),
.C(n_184),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_173),
.B(n_177),
.Y(n_323)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_182),
.Y(n_224)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_181),
.Y(n_420)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_184),
.B(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_185),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_199),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_191),
.B(n_244),
.Y(n_243)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_192),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_192),
.B(n_310),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_192),
.A2(n_214),
.B1(n_310),
.B2(n_311),
.Y(n_378)
);

BUFx2_ASAP7_75t_L g405 ( 
.A(n_193),
.Y(n_405)
);

INVx8_ASAP7_75t_L g429 ( 
.A(n_193),
.Y(n_429)
);

BUFx8_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

BUFx5_ASAP7_75t_L g438 ( 
.A(n_194),
.Y(n_438)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_195),
.Y(n_245)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_200),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_246),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_204),
.B(n_246),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_207),
.C(n_209),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_205),
.B(n_207),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_209),
.B(n_330),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_225),
.C(n_243),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_210),
.B(n_325),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_215),
.C(n_223),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_211),
.Y(n_295)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_215),
.B(n_223),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_220),
.B(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_225),
.B(n_243),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_235),
.C(n_239),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_226),
.B(n_292),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_227),
.A2(n_228),
.B1(n_233),
.B2(n_317),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

INVx3_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_232),
.Y(n_349)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_232),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_233),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_235),
.A2(n_239),
.B1(n_240),
.B2(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx6_ASAP7_75t_L g372 ( 
.A(n_238),
.Y(n_372)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

BUFx24_ASAP7_75t_SL g497 ( 
.A(n_246),
.Y(n_497)
);

AOI221xp5_ASAP7_75t_L g247 ( 
.A1(n_248),
.A2(n_384),
.B1(n_480),
.B2(n_485),
.C(n_486),
.Y(n_247)
);

NOR3xp33_ASAP7_75t_SL g248 ( 
.A(n_249),
.B(n_327),
.C(n_331),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g480 ( 
.A1(n_249),
.A2(n_481),
.B(n_484),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_320),
.Y(n_249)
);

OR2x2_ASAP7_75t_L g484 ( 
.A(n_250),
.B(n_320),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_294),
.C(n_297),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_251),
.B(n_294),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_252),
.B(n_277),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_252),
.B(n_278),
.C(n_291),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_256),
.C(n_267),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_254),
.B(n_268),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_256),
.B(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_261),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_262),
.B(n_300),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_266),
.Y(n_413)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_269),
.Y(n_339)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_273),
.B(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_275),
.Y(n_273)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_291),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_287),
.C(n_289),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_279),
.B(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g340 ( 
.A1(n_279),
.A2(n_282),
.B(n_341),
.Y(n_340)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

INVx5_ASAP7_75t_L g284 ( 
.A(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g319 ( 
.A(n_287),
.B(n_289),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_297),
.B(n_356),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_314),
.C(n_318),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g334 ( 
.A(n_298),
.B(n_335),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_301),
.C(n_308),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_299),
.B(n_380),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_301),
.A2(n_308),
.B1(n_309),
.B2(n_381),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_301),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_SL g362 ( 
.A(n_302),
.B(n_363),
.Y(n_362)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx4_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_306),
.Y(n_364)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_311),
.Y(n_310)
);

INVx6_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_326),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_322),
.B(n_324),
.C(n_326),
.Y(n_328)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_327),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_329),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_328),
.B(n_329),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_332),
.B(n_357),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_332),
.A2(n_482),
.B(n_483),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_355),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_333),
.B(n_355),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_336),
.C(n_353),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_383),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_336),
.B(n_353),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.C(n_344),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_337),
.B(n_340),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_342),
.B(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_344),
.B(n_360),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_347),
.C(n_350),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g467 ( 
.A1(n_345),
.A2(n_346),
.B1(n_468),
.B2(n_469),
.Y(n_467)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g468 ( 
.A1(n_347),
.A2(n_348),
.B1(n_350),
.B2(n_351),
.Y(n_468)
);

CKINVDCx14_ASAP7_75t_R g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_358),
.B(n_382),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_358),
.B(n_382),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.C(n_379),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g477 ( 
.A(n_359),
.B(n_478),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g478 ( 
.A(n_361),
.B(n_379),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.C(n_377),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_SL g470 ( 
.A(n_362),
.B(n_471),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_365),
.A2(n_377),
.B1(n_378),
.B2(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_365),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_370),
.C(n_373),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_366),
.A2(n_367),
.B1(n_373),
.B2(n_374),
.Y(n_460)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_370),
.B(n_460),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_372),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_371),
.B(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_378),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_385),
.A2(n_475),
.B(n_479),
.Y(n_384)
);

AOI21xp5_ASAP7_75t_L g385 ( 
.A1(n_386),
.A2(n_462),
.B(n_474),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_L g386 ( 
.A1(n_387),
.A2(n_449),
.B(n_461),
.Y(n_386)
);

AOI21xp5_ASAP7_75t_L g387 ( 
.A1(n_388),
.A2(n_423),
.B(n_448),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_389),
.B(n_415),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g448 ( 
.A(n_389),
.B(n_415),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_L g389 ( 
.A(n_390),
.B(n_401),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_390),
.B(n_402),
.C(n_411),
.Y(n_450)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_391),
.B(n_396),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_391),
.B(n_397),
.C(n_398),
.Y(n_458)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_398),
.Y(n_396)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_411),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_403),
.B(n_406),
.Y(n_416)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_407),
.B(n_408),
.Y(n_406)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_409),
.Y(n_408)
);

INVx8_ASAP7_75t_L g409 ( 
.A(n_410),
.Y(n_409)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_412),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.C(n_421),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_416),
.B(n_445),
.Y(n_444)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_417),
.A2(n_421),
.B1(n_422),
.B2(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_417),
.Y(n_446)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_420),
.Y(n_419)
);

INVx3_ASAP7_75t_L g454 ( 
.A(n_420),
.Y(n_454)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_442),
.B(n_447),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g424 ( 
.A1(n_425),
.A2(n_434),
.B(n_441),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_433),
.Y(n_425)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_426),
.B(n_433),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_430),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_427),
.B(n_430),
.Y(n_443)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx3_ASAP7_75t_SL g431 ( 
.A(n_432),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_439),
.Y(n_434)
);

INVx1_ASAP7_75t_SL g436 ( 
.A(n_437),
.Y(n_436)
);

INVx3_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_443),
.B(n_444),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_443),
.B(n_444),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_451),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_450),
.B(n_451),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_452),
.A2(n_465),
.B1(n_466),
.B2(n_467),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_452),
.B(n_458),
.C(n_459),
.Y(n_473)
);

FAx1_ASAP7_75t_SL g452 ( 
.A(n_453),
.B(n_455),
.CI(n_456),
.CON(n_452),
.SN(n_452)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_463),
.B(n_473),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_463),
.B(n_473),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_470),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g476 ( 
.A(n_465),
.B(n_467),
.C(n_470),
.Y(n_476)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_468),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_476),
.B(n_477),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_476),
.B(n_477),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_491),
.B(n_492),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g494 ( 
.A(n_491),
.B(n_492),
.Y(n_494)
);


endmodule