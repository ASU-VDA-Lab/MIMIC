module fake_ariane_1508_n_800 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_800);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_800;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_374;
wire n_345;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_665;
wire n_336;
wire n_731;
wire n_754;
wire n_779;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_381;
wire n_344;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_271;
wire n_465;
wire n_507;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_248;
wire n_277;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_780;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_658;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_772;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_745;
wire n_613;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_742;
wire n_716;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_697;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_548;
wire n_542;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_531;
wire n_783;
wire n_675;

INVx2_ASAP7_75t_SL g168 ( 
.A(n_111),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_3),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_64),
.Y(n_170)
);

BUFx10_ASAP7_75t_L g171 ( 
.A(n_43),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_28),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_97),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_104),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_9),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_47),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_164),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_9),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_147),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_77),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_93),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_4),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_131),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_133),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_145),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_0),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_152),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_101),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_2),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_165),
.Y(n_192)
);

INVx2_ASAP7_75t_SL g193 ( 
.A(n_159),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_67),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_83),
.Y(n_195)
);

BUFx5_ASAP7_75t_L g196 ( 
.A(n_23),
.Y(n_196)
);

BUFx3_ASAP7_75t_L g197 ( 
.A(n_72),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_137),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_15),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_4),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_142),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_0),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_80),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_87),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_130),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_48),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_82),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_30),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_78),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_117),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_119),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_128),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_70),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_109),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_108),
.Y(n_216)
);

NOR2xp67_ASAP7_75t_L g217 ( 
.A(n_106),
.B(n_57),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_41),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_126),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_91),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

BUFx2_ASAP7_75t_L g222 ( 
.A(n_102),
.Y(n_222)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_160),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_25),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_136),
.Y(n_225)
);

BUFx10_ASAP7_75t_L g226 ( 
.A(n_11),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_90),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_139),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_174),
.Y(n_229)
);

BUFx12f_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

OAI22x1_ASAP7_75t_SL g232 ( 
.A1(n_169),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_176),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

AND2x4_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_1),
.Y(n_235)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_171),
.Y(n_236)
);

OAI21x1_ASAP7_75t_L g237 ( 
.A1(n_185),
.A2(n_75),
.B(n_166),
.Y(n_237)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_184),
.Y(n_238)
);

BUFx8_ASAP7_75t_L g239 ( 
.A(n_222),
.Y(n_239)
);

OA21x2_ASAP7_75t_L g240 ( 
.A1(n_178),
.A2(n_5),
.B(n_6),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_181),
.B(n_5),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_188),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_185),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_187),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

BUFx6f_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_182),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_226),
.Y(n_249)
);

BUFx2_ASAP7_75t_L g250 ( 
.A(n_191),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_221),
.Y(n_252)
);

INVx5_ASAP7_75t_L g253 ( 
.A(n_168),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_196),
.Y(n_254)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_223),
.Y(n_255)
);

AND2x6_ASAP7_75t_L g256 ( 
.A(n_190),
.B(n_194),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_195),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_205),
.B(n_6),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_186),
.A2(n_7),
.B1(n_8),
.B2(n_10),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_200),
.Y(n_260)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_196),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_201),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_183),
.B(n_7),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_208),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_196),
.Y(n_265)
);

AND2x4_ASAP7_75t_L g266 ( 
.A(n_193),
.B(n_8),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_211),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g268 ( 
.A(n_204),
.Y(n_268)
);

INVx5_ASAP7_75t_L g269 ( 
.A(n_196),
.Y(n_269)
);

AND2x6_ASAP7_75t_L g270 ( 
.A(n_212),
.B(n_18),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_170),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_218),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_224),
.Y(n_273)
);

BUFx6f_ASAP7_75t_L g274 ( 
.A(n_172),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_236),
.B(n_183),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_229),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_229),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_233),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_234),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_245),
.Y(n_280)
);

AND2x4_ASAP7_75t_L g281 ( 
.A(n_236),
.B(n_255),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_245),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_268),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_230),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_239),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_230),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_239),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_246),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_239),
.Y(n_289)
);

INVx3_ASAP7_75t_L g290 ( 
.A(n_252),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_274),
.Y(n_291)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_252),
.Y(n_292)
);

NOR2xp67_ASAP7_75t_L g293 ( 
.A(n_236),
.B(n_173),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_274),
.Y(n_294)
);

HB1xp67_ASAP7_75t_L g295 ( 
.A(n_250),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_241),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_264),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g298 ( 
.A(n_255),
.B(n_199),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_274),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_264),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_264),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_R g303 ( 
.A(n_255),
.B(n_209),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_262),
.B(n_202),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_R g305 ( 
.A(n_260),
.B(n_215),
.Y(n_305)
);

INVx5_ASAP7_75t_L g306 ( 
.A(n_270),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_271),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_260),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_271),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_271),
.Y(n_310)
);

INVx2_ASAP7_75t_L g311 ( 
.A(n_244),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_264),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_248),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_263),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_244),
.Y(n_315)
);

NOR2x1p5_ASAP7_75t_L g316 ( 
.A(n_249),
.B(n_175),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_244),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_248),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_272),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_244),
.Y(n_320)
);

OR2x6_ASAP7_75t_L g321 ( 
.A(n_251),
.B(n_217),
.Y(n_321)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_247),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_272),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_231),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_247),
.Y(n_325)
);

NOR2xp67_ASAP7_75t_L g326 ( 
.A(n_284),
.B(n_286),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_278),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_307),
.B(n_263),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_275),
.B(n_266),
.Y(n_329)
);

BUFx6f_ASAP7_75t_SL g330 ( 
.A(n_281),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_279),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_313),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_L g333 ( 
.A(n_304),
.B(n_266),
.C(n_235),
.Y(n_333)
);

NAND2x1_ASAP7_75t_L g334 ( 
.A(n_288),
.B(n_270),
.Y(n_334)
);

INVxp33_ASAP7_75t_L g335 ( 
.A(n_295),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_309),
.B(n_266),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_310),
.B(n_235),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g338 ( 
.A(n_317),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_287),
.B(n_289),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_281),
.B(n_235),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_291),
.B(n_253),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_318),
.B(n_253),
.Y(n_342)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_290),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_296),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

INVxp67_ASAP7_75t_L g346 ( 
.A(n_295),
.Y(n_346)
);

BUFx6f_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

NAND2x1_ASAP7_75t_L g348 ( 
.A(n_288),
.B(n_270),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_319),
.B(n_253),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_292),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_317),
.Y(n_351)
);

INVx2_ASAP7_75t_SL g352 ( 
.A(n_323),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g353 ( 
.A(n_317),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g354 ( 
.A(n_298),
.B(n_231),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_294),
.B(n_253),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_299),
.B(n_300),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_256),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_293),
.B(n_256),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_311),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_292),
.B(n_256),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_315),
.Y(n_361)
);

NAND2xp33_ASAP7_75t_L g362 ( 
.A(n_316),
.B(n_270),
.Y(n_362)
);

INVx4_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_321),
.B(n_253),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_297),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_320),
.Y(n_366)
);

NOR2xp33_ASAP7_75t_L g367 ( 
.A(n_321),
.B(n_276),
.Y(n_367)
);

AO221x1_ASAP7_75t_L g368 ( 
.A1(n_305),
.A2(n_232),
.B1(n_238),
.B2(n_243),
.C(n_252),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_301),
.B(n_256),
.Y(n_369)
);

NAND2x1_ASAP7_75t_L g370 ( 
.A(n_325),
.B(n_270),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_256),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_321),
.B(n_257),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_305),
.B(n_242),
.Y(n_373)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_277),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_280),
.B(n_267),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_312),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_322),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_306),
.B(n_273),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_306),
.B(n_247),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_306),
.B(n_247),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g381 ( 
.A(n_282),
.B(n_258),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_283),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_314),
.Y(n_383)
);

INVx3_ASAP7_75t_L g384 ( 
.A(n_303),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_303),
.B(n_238),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_308),
.B(n_238),
.Y(n_386)
);

BUFx5_ASAP7_75t_L g387 ( 
.A(n_285),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_SL g388 ( 
.A(n_313),
.B(n_259),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_278),
.Y(n_389)
);

INVx2_ASAP7_75t_SL g390 ( 
.A(n_313),
.Y(n_390)
);

NOR2xp67_ASAP7_75t_L g391 ( 
.A(n_284),
.B(n_269),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_SL g392 ( 
.A(n_313),
.B(n_219),
.Y(n_392)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_333),
.A2(n_228),
.B1(n_240),
.B2(n_206),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g394 ( 
.A1(n_327),
.A2(n_240),
.B1(n_265),
.B2(n_261),
.Y(n_394)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_328),
.A2(n_216),
.B1(n_179),
.B2(n_189),
.Y(n_395)
);

NOR3xp33_ASAP7_75t_SL g396 ( 
.A(n_381),
.B(n_227),
.C(n_192),
.Y(n_396)
);

BUFx6f_ASAP7_75t_L g397 ( 
.A(n_338),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_331),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_375),
.A2(n_220),
.B1(n_198),
.B2(n_207),
.Y(n_400)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_374),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_329),
.B(n_177),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_336),
.A2(n_213),
.B1(n_214),
.B2(n_225),
.Y(n_403)
);

AOI22xp33_ASAP7_75t_L g404 ( 
.A1(n_344),
.A2(n_240),
.B1(n_265),
.B2(n_261),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_382),
.Y(n_405)
);

INVx1_ASAP7_75t_SL g406 ( 
.A(n_332),
.Y(n_406)
);

INVxp67_ASAP7_75t_L g407 ( 
.A(n_386),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_337),
.B(n_210),
.Y(n_408)
);

INVx3_ASAP7_75t_L g409 ( 
.A(n_359),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_343),
.Y(n_410)
);

O2A1O1Ixp5_ASAP7_75t_L g411 ( 
.A1(n_334),
.A2(n_246),
.B(n_254),
.C(n_237),
.Y(n_411)
);

AOI21xp33_ASAP7_75t_L g412 ( 
.A1(n_357),
.A2(n_254),
.B(n_237),
.Y(n_412)
);

AND2x2_ASAP7_75t_L g413 ( 
.A(n_335),
.B(n_10),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_340),
.B(n_269),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_269),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_354),
.B(n_269),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_382),
.Y(n_417)
);

HB1xp67_ASAP7_75t_L g418 ( 
.A(n_346),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_389),
.B(n_269),
.Y(n_419)
);

NOR3xp33_ASAP7_75t_SL g420 ( 
.A(n_383),
.B(n_11),
.C(n_12),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_343),
.B(n_196),
.Y(n_421)
);

NAND2x1p5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_12),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_13),
.Y(n_423)
);

AND2x4_ASAP7_75t_L g424 ( 
.A(n_352),
.B(n_13),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_345),
.B(n_14),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_350),
.Y(n_426)
);

BUFx12f_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_338),
.Y(n_428)
);

AND2x4_ASAP7_75t_L g429 ( 
.A(n_390),
.B(n_14),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_L g430 ( 
.A1(n_388),
.A2(n_372),
.B1(n_373),
.B2(n_365),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_376),
.B(n_360),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_362),
.A2(n_86),
.B(n_163),
.Y(n_432)
);

INVx2_ASAP7_75t_SL g433 ( 
.A(n_384),
.Y(n_433)
);

NOR2xp67_ASAP7_75t_L g434 ( 
.A(n_326),
.B(n_167),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_377),
.Y(n_435)
);

BUFx3_ASAP7_75t_L g436 ( 
.A(n_387),
.Y(n_436)
);

BUFx3_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_358),
.A2(n_85),
.B(n_161),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_361),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_367),
.B(n_15),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_359),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_364),
.B(n_16),
.Y(n_442)
);

AOI21x1_ASAP7_75t_L g443 ( 
.A1(n_348),
.A2(n_84),
.B(n_158),
.Y(n_443)
);

NOR2xp33_ASAP7_75t_R g444 ( 
.A(n_339),
.B(n_19),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_351),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_366),
.Y(n_447)
);

AOI22xp33_ASAP7_75t_L g448 ( 
.A1(n_368),
.A2(n_16),
.B1(n_17),
.B2(n_20),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_366),
.Y(n_449)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_338),
.Y(n_450)
);

HB1xp67_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_366),
.Y(n_452)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_SL g454 ( 
.A(n_391),
.B(n_17),
.Y(n_454)
);

NOR2x1p5_ASAP7_75t_L g455 ( 
.A(n_370),
.B(n_162),
.Y(n_455)
);

NOR2x2_ASAP7_75t_L g456 ( 
.A(n_387),
.B(n_21),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_347),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_378),
.B(n_22),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g459 ( 
.A(n_392),
.B(n_24),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_341),
.B(n_26),
.Y(n_460)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_342),
.B(n_27),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_347),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_439),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_407),
.B(n_349),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_399),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_406),
.B(n_355),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_418),
.Y(n_467)
);

AOI21xp5_ASAP7_75t_L g468 ( 
.A1(n_431),
.A2(n_363),
.B(n_371),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g469 ( 
.A1(n_431),
.A2(n_369),
.B(n_379),
.Y(n_469)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_401),
.A2(n_380),
.B1(n_353),
.B2(n_347),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_406),
.B(n_417),
.Y(n_471)
);

INVx3_ASAP7_75t_L g472 ( 
.A(n_397),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_453),
.B(n_353),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_402),
.B(n_353),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_414),
.A2(n_29),
.B(n_31),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_435),
.Y(n_476)
);

BUFx3_ASAP7_75t_L g477 ( 
.A(n_427),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_421),
.A2(n_32),
.B(n_33),
.Y(n_478)
);

AO22x1_ASAP7_75t_L g479 ( 
.A1(n_459),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_479)
);

BUFx3_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_433),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_410),
.B(n_157),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_436),
.B(n_40),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_426),
.Y(n_484)
);

NOR3xp33_ASAP7_75t_SL g485 ( 
.A(n_440),
.B(n_425),
.C(n_442),
.Y(n_485)
);

AOI22xp33_ASAP7_75t_L g486 ( 
.A1(n_393),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_430),
.B(n_46),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_408),
.B(n_49),
.Y(n_489)
);

O2A1O1Ixp33_ASAP7_75t_L g490 ( 
.A1(n_425),
.A2(n_423),
.B(n_429),
.C(n_424),
.Y(n_490)
);

A2O1A1Ixp33_ASAP7_75t_L g491 ( 
.A1(n_424),
.A2(n_50),
.B(n_51),
.C(n_52),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g492 ( 
.A1(n_415),
.A2(n_53),
.B(n_54),
.Y(n_492)
);

BUFx2_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_429),
.B(n_55),
.Y(n_494)
);

INVx3_ASAP7_75t_L g495 ( 
.A(n_397),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_416),
.A2(n_56),
.B(n_58),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_400),
.B(n_59),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_441),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g499 ( 
.A1(n_416),
.A2(n_60),
.B(n_61),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_395),
.B(n_62),
.Y(n_500)
);

BUFx6f_ASAP7_75t_L g501 ( 
.A(n_397),
.Y(n_501)
);

OR2x6_ASAP7_75t_L g502 ( 
.A(n_437),
.B(n_63),
.Y(n_502)
);

O2A1O1Ixp33_ASAP7_75t_L g503 ( 
.A1(n_454),
.A2(n_65),
.B(n_66),
.C(n_68),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_SL g504 ( 
.A(n_403),
.B(n_69),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_413),
.B(n_156),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_428),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_457),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_449),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_422),
.A2(n_71),
.B1(n_73),
.B2(n_74),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_462),
.B(n_409),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_422),
.A2(n_76),
.B1(n_81),
.B2(n_88),
.Y(n_511)
);

AOI21xp5_ASAP7_75t_L g512 ( 
.A1(n_419),
.A2(n_89),
.B(n_92),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_448),
.B(n_94),
.Y(n_513)
);

A2O1A1Ixp33_ASAP7_75t_L g514 ( 
.A1(n_432),
.A2(n_95),
.B(n_96),
.C(n_98),
.Y(n_514)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_419),
.A2(n_99),
.B(n_100),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_SL g516 ( 
.A(n_420),
.B(n_103),
.C(n_107),
.Y(n_516)
);

A2O1A1Ixp33_ASAP7_75t_L g517 ( 
.A1(n_461),
.A2(n_110),
.B(n_112),
.C(n_113),
.Y(n_517)
);

O2A1O1Ixp33_ASAP7_75t_L g518 ( 
.A1(n_396),
.A2(n_114),
.B(n_115),
.C(n_116),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_469),
.A2(n_411),
.B(n_468),
.Y(n_519)
);

CKINVDCx11_ASAP7_75t_R g520 ( 
.A(n_477),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_489),
.A2(n_412),
.B(n_458),
.Y(n_521)
);

AND2x2_ASAP7_75t_L g522 ( 
.A(n_467),
.B(n_444),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_465),
.B(n_409),
.Y(n_523)
);

AOI21xp5_ASAP7_75t_L g524 ( 
.A1(n_474),
.A2(n_458),
.B(n_460),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_476),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_484),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_463),
.Y(n_527)
);

AO21x2_ASAP7_75t_L g528 ( 
.A1(n_488),
.A2(n_412),
.B(n_497),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_490),
.B(n_485),
.Y(n_529)
);

AOI22xp33_ASAP7_75t_L g530 ( 
.A1(n_513),
.A2(n_447),
.B1(n_446),
.B2(n_394),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_487),
.Y(n_531)
);

INVx2_ASAP7_75t_SL g532 ( 
.A(n_493),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_501),
.Y(n_533)
);

OAI21x1_ASAP7_75t_L g534 ( 
.A1(n_492),
.A2(n_443),
.B(n_438),
.Y(n_534)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_501),
.Y(n_535)
);

INVx6_ASAP7_75t_SL g536 ( 
.A(n_502),
.Y(n_536)
);

OAI21x1_ASAP7_75t_L g537 ( 
.A1(n_496),
.A2(n_404),
.B(n_455),
.Y(n_537)
);

INVx6_ASAP7_75t_L g538 ( 
.A(n_501),
.Y(n_538)
);

BUFx6f_ASAP7_75t_L g539 ( 
.A(n_472),
.Y(n_539)
);

BUFx3_ASAP7_75t_L g540 ( 
.A(n_480),
.Y(n_540)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_505),
.A2(n_434),
.B1(n_452),
.B2(n_450),
.Y(n_541)
);

AOI21xp5_ASAP7_75t_L g542 ( 
.A1(n_464),
.A2(n_398),
.B(n_428),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_500),
.A2(n_398),
.B(n_428),
.Y(n_543)
);

AND2x4_ASAP7_75t_L g544 ( 
.A(n_472),
.B(n_398),
.Y(n_544)
);

OR2x2_ASAP7_75t_L g545 ( 
.A(n_507),
.B(n_471),
.Y(n_545)
);

OAI21x1_ASAP7_75t_L g546 ( 
.A1(n_499),
.A2(n_398),
.B(n_456),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_498),
.Y(n_547)
);

BUFx2_ASAP7_75t_L g548 ( 
.A(n_494),
.Y(n_548)
);

INVxp67_ASAP7_75t_SL g549 ( 
.A(n_473),
.Y(n_549)
);

OA21x2_ASAP7_75t_L g550 ( 
.A1(n_514),
.A2(n_118),
.B(n_120),
.Y(n_550)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_510),
.Y(n_551)
);

BUFx3_ASAP7_75t_L g552 ( 
.A(n_495),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_494),
.Y(n_553)
);

OAI21x1_ASAP7_75t_L g554 ( 
.A1(n_478),
.A2(n_121),
.B(n_122),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_502),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_508),
.Y(n_556)
);

INVx6_ASAP7_75t_L g557 ( 
.A(n_494),
.Y(n_557)
);

OAI21x1_ASAP7_75t_L g558 ( 
.A1(n_512),
.A2(n_123),
.B(n_124),
.Y(n_558)
);

OAI21x1_ASAP7_75t_L g559 ( 
.A1(n_515),
.A2(n_125),
.B(n_127),
.Y(n_559)
);

CKINVDCx20_ASAP7_75t_R g560 ( 
.A(n_483),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_495),
.Y(n_561)
);

OAI21x1_ASAP7_75t_L g562 ( 
.A1(n_475),
.A2(n_129),
.B(n_132),
.Y(n_562)
);

AND2x2_ASAP7_75t_L g563 ( 
.A(n_516),
.B(n_466),
.Y(n_563)
);

INVx1_ASAP7_75t_SL g564 ( 
.A(n_494),
.Y(n_564)
);

CKINVDCx6p67_ASAP7_75t_R g565 ( 
.A(n_520),
.Y(n_565)
);

INVx3_ASAP7_75t_L g566 ( 
.A(n_557),
.Y(n_566)
);

INVx1_ASAP7_75t_SL g567 ( 
.A(n_540),
.Y(n_567)
);

AOI21xp33_ASAP7_75t_L g568 ( 
.A1(n_529),
.A2(n_486),
.B(n_504),
.Y(n_568)
);

NAND2x1p5_ASAP7_75t_L g569 ( 
.A(n_548),
.B(n_506),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_525),
.Y(n_570)
);

INVx2_ASAP7_75t_L g571 ( 
.A(n_556),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g572 ( 
.A(n_526),
.B(n_549),
.Y(n_572)
);

AO21x2_ASAP7_75t_L g573 ( 
.A1(n_521),
.A2(n_491),
.B(n_482),
.Y(n_573)
);

AOI22xp5_ASAP7_75t_L g574 ( 
.A1(n_560),
.A2(n_470),
.B1(n_509),
.B2(n_511),
.Y(n_574)
);

AOI21x1_ASAP7_75t_L g575 ( 
.A1(n_519),
.A2(n_479),
.B(n_518),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_519),
.A2(n_534),
.B(n_524),
.Y(n_576)
);

BUFx3_ASAP7_75t_L g577 ( 
.A(n_540),
.Y(n_577)
);

AOI222xp33_ASAP7_75t_L g578 ( 
.A1(n_522),
.A2(n_517),
.B1(n_506),
.B2(n_481),
.C1(n_503),
.C2(n_141),
.Y(n_578)
);

BUFx3_ASAP7_75t_L g579 ( 
.A(n_533),
.Y(n_579)
);

CKINVDCx5p33_ASAP7_75t_R g580 ( 
.A(n_520),
.Y(n_580)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_534),
.A2(n_134),
.B(n_135),
.Y(n_581)
);

CKINVDCx16_ASAP7_75t_R g582 ( 
.A(n_560),
.Y(n_582)
);

INVx8_ASAP7_75t_L g583 ( 
.A(n_544),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_557),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_527),
.Y(n_585)
);

BUFx12f_ASAP7_75t_L g586 ( 
.A(n_532),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_531),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_547),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_523),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_557),
.Y(n_590)
);

AOI21xp5_ASAP7_75t_L g591 ( 
.A1(n_521),
.A2(n_138),
.B(n_140),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_543),
.A2(n_143),
.B(n_144),
.Y(n_592)
);

AO21x1_ASAP7_75t_SL g593 ( 
.A1(n_541),
.A2(n_146),
.B(n_148),
.Y(n_593)
);

CKINVDCx14_ASAP7_75t_R g594 ( 
.A(n_545),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_551),
.Y(n_595)
);

AND2x2_ASAP7_75t_L g596 ( 
.A(n_549),
.B(n_149),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_561),
.Y(n_597)
);

BUFx4f_ASAP7_75t_SL g598 ( 
.A(n_536),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_537),
.A2(n_150),
.B(n_151),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_561),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_558),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_558),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_538),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_563),
.B(n_153),
.Y(n_604)
);

HB1xp67_ASAP7_75t_L g605 ( 
.A(n_533),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_594),
.B(n_555),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_572),
.B(n_553),
.Y(n_607)
);

AND2x2_ASAP7_75t_L g608 ( 
.A(n_594),
.B(n_552),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_570),
.Y(n_609)
);

CKINVDCx16_ASAP7_75t_R g610 ( 
.A(n_582),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_587),
.Y(n_611)
);

OR2x2_ASAP7_75t_L g612 ( 
.A(n_572),
.B(n_552),
.Y(n_612)
);

INVx6_ASAP7_75t_L g613 ( 
.A(n_583),
.Y(n_613)
);

NOR3xp33_ASAP7_75t_SL g614 ( 
.A(n_580),
.B(n_542),
.C(n_536),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_589),
.B(n_564),
.Y(n_615)
);

CKINVDCx20_ASAP7_75t_R g616 ( 
.A(n_565),
.Y(n_616)
);

AOI22xp33_ASAP7_75t_L g617 ( 
.A1(n_568),
.A2(n_536),
.B1(n_530),
.B2(n_528),
.Y(n_617)
);

HB1xp67_ASAP7_75t_L g618 ( 
.A(n_601),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_596),
.B(n_530),
.Y(n_619)
);

BUFx2_ASAP7_75t_L g620 ( 
.A(n_586),
.Y(n_620)
);

AO31x2_ASAP7_75t_L g621 ( 
.A1(n_601),
.A2(n_528),
.A3(n_550),
.B(n_537),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_R g622 ( 
.A(n_580),
.B(n_538),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_579),
.B(n_535),
.Y(n_623)
);

BUFx2_ASAP7_75t_SL g624 ( 
.A(n_577),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_585),
.B(n_588),
.Y(n_625)
);

NOR3xp33_ASAP7_75t_SL g626 ( 
.A(n_565),
.B(n_591),
.C(n_603),
.Y(n_626)
);

NAND2xp33_ASAP7_75t_SL g627 ( 
.A(n_596),
.B(n_539),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_577),
.B(n_567),
.Y(n_628)
);

BUFx3_ASAP7_75t_L g629 ( 
.A(n_586),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_539),
.Y(n_630)
);

AND2x2_ASAP7_75t_L g631 ( 
.A(n_605),
.B(n_604),
.Y(n_631)
);

HB1xp67_ASAP7_75t_L g632 ( 
.A(n_579),
.Y(n_632)
);

OAI22xp5_ASAP7_75t_L g633 ( 
.A1(n_574),
.A2(n_550),
.B1(n_539),
.B2(n_538),
.Y(n_633)
);

NAND2xp33_ASAP7_75t_R g634 ( 
.A(n_604),
.B(n_550),
.Y(n_634)
);

AND2x2_ASAP7_75t_L g635 ( 
.A(n_595),
.B(n_539),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_598),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_583),
.Y(n_637)
);

OR2x6_ASAP7_75t_L g638 ( 
.A(n_583),
.B(n_546),
.Y(n_638)
);

AND2x2_ASAP7_75t_L g639 ( 
.A(n_566),
.B(n_535),
.Y(n_639)
);

CKINVDCx16_ASAP7_75t_R g640 ( 
.A(n_590),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_571),
.Y(n_641)
);

AND2x4_ASAP7_75t_L g642 ( 
.A(n_566),
.B(n_535),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_583),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_571),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_600),
.B(n_535),
.Y(n_645)
);

HB1xp67_ASAP7_75t_L g646 ( 
.A(n_569),
.Y(n_646)
);

INVx1_ASAP7_75t_SL g647 ( 
.A(n_590),
.Y(n_647)
);

AOI21xp33_ASAP7_75t_L g648 ( 
.A1(n_578),
.A2(n_559),
.B(n_554),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_566),
.B(n_544),
.Y(n_649)
);

BUFx2_ASAP7_75t_L g650 ( 
.A(n_590),
.Y(n_650)
);

AND2x4_ASAP7_75t_L g651 ( 
.A(n_584),
.B(n_544),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_609),
.B(n_576),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_641),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_611),
.Y(n_654)
);

NOR2x1p5_ASAP7_75t_L g655 ( 
.A(n_629),
.B(n_584),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_625),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_632),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_631),
.B(n_569),
.Y(n_658)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_607),
.B(n_576),
.Y(n_659)
);

AND2x4_ASAP7_75t_L g660 ( 
.A(n_638),
.B(n_590),
.Y(n_660)
);

OAI21x1_ASAP7_75t_L g661 ( 
.A1(n_633),
.A2(n_599),
.B(n_575),
.Y(n_661)
);

INVx2_ASAP7_75t_SL g662 ( 
.A(n_612),
.Y(n_662)
);

HB1xp67_ASAP7_75t_L g663 ( 
.A(n_607),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_635),
.B(n_569),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_618),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_644),
.Y(n_666)
);

HB1xp67_ASAP7_75t_L g667 ( 
.A(n_615),
.Y(n_667)
);

AND2x4_ASAP7_75t_L g668 ( 
.A(n_638),
.B(n_646),
.Y(n_668)
);

OR2x2_ASAP7_75t_L g669 ( 
.A(n_619),
.B(n_602),
.Y(n_669)
);

AND2x2_ASAP7_75t_L g670 ( 
.A(n_619),
.B(n_573),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_615),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_645),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_610),
.B(n_584),
.Y(n_673)
);

AND2x2_ASAP7_75t_L g674 ( 
.A(n_608),
.B(n_573),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_628),
.B(n_590),
.Y(n_675)
);

HB1xp67_ASAP7_75t_L g676 ( 
.A(n_645),
.Y(n_676)
);

OR2x2_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_602),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_638),
.B(n_599),
.Y(n_678)
);

OAI221xp5_ASAP7_75t_L g679 ( 
.A1(n_634),
.A2(n_575),
.B1(n_592),
.B2(n_593),
.C(n_581),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_621),
.B(n_639),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_630),
.Y(n_681)
);

AND2x2_ASAP7_75t_L g682 ( 
.A(n_630),
.B(n_593),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_L g683 ( 
.A(n_663),
.B(n_650),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_L g684 ( 
.A(n_667),
.B(n_606),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_671),
.B(n_623),
.Y(n_685)
);

NAND3xp33_ASAP7_75t_L g686 ( 
.A(n_657),
.B(n_626),
.C(n_614),
.Y(n_686)
);

INVx2_ASAP7_75t_SL g687 ( 
.A(n_677),
.Y(n_687)
);

HB1xp67_ASAP7_75t_L g688 ( 
.A(n_662),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_662),
.B(n_623),
.Y(n_689)
);

HB1xp67_ASAP7_75t_L g690 ( 
.A(n_665),
.Y(n_690)
);

AND2x4_ASAP7_75t_L g691 ( 
.A(n_668),
.B(n_614),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_674),
.B(n_633),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_654),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_656),
.B(n_617),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_674),
.B(n_626),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_676),
.Y(n_696)
);

BUFx3_ASAP7_75t_L g697 ( 
.A(n_675),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_659),
.B(n_649),
.Y(n_698)
);

HB1xp67_ASAP7_75t_L g699 ( 
.A(n_665),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_669),
.B(n_640),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_677),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_653),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_666),
.Y(n_703)
);

INVxp33_ASAP7_75t_L g704 ( 
.A(n_673),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_668),
.B(n_651),
.Y(n_705)
);

OR2x2_ASAP7_75t_L g706 ( 
.A(n_669),
.B(n_627),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_696),
.B(n_659),
.Y(n_707)
);

AND2x4_ASAP7_75t_L g708 ( 
.A(n_687),
.B(n_691),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_687),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_697),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_690),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_702),
.Y(n_712)
);

INVx1_ASAP7_75t_L g713 ( 
.A(n_699),
.Y(n_713)
);

AND2x2_ASAP7_75t_L g714 ( 
.A(n_698),
.B(n_652),
.Y(n_714)
);

INVx2_ASAP7_75t_SL g715 ( 
.A(n_701),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_698),
.B(n_652),
.Y(n_716)
);

NOR3xp33_ASAP7_75t_SL g717 ( 
.A(n_686),
.B(n_636),
.C(n_679),
.Y(n_717)
);

HB1xp67_ASAP7_75t_L g718 ( 
.A(n_688),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_695),
.B(n_678),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_693),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_695),
.B(n_668),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_701),
.B(n_678),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_711),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_711),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_713),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_707),
.B(n_683),
.Y(n_726)
);

NAND4xp75_ASAP7_75t_L g727 ( 
.A(n_717),
.B(n_692),
.C(n_694),
.D(n_682),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_713),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_SL g729 ( 
.A1(n_719),
.A2(n_692),
.B1(n_691),
.B2(n_670),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_720),
.B(n_701),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_707),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_712),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_723),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_732),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_724),
.Y(n_735)
);

OAI211xp5_ASAP7_75t_SL g736 ( 
.A1(n_725),
.A2(n_728),
.B(n_730),
.C(n_718),
.Y(n_736)
);

OAI22xp5_ASAP7_75t_L g737 ( 
.A1(n_733),
.A2(n_727),
.B1(n_729),
.B2(n_708),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_735),
.B(n_730),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_736),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_734),
.B(n_731),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_736),
.Y(n_741)
);

HB1xp67_ASAP7_75t_L g742 ( 
.A(n_739),
.Y(n_742)
);

INVx2_ASAP7_75t_SL g743 ( 
.A(n_738),
.Y(n_743)
);

NOR3x1_ASAP7_75t_L g744 ( 
.A(n_737),
.B(n_620),
.C(n_721),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_741),
.B(n_719),
.Y(n_745)
);

NOR3x1_ASAP7_75t_L g746 ( 
.A(n_745),
.B(n_740),
.C(n_715),
.Y(n_746)
);

AOI21xp5_ASAP7_75t_SL g747 ( 
.A1(n_742),
.A2(n_655),
.B(n_708),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_743),
.A2(n_704),
.B(n_616),
.Y(n_748)
);

NOR4xp25_ASAP7_75t_L g749 ( 
.A(n_746),
.B(n_744),
.C(n_684),
.D(n_715),
.Y(n_749)
);

NOR2x1_ASAP7_75t_L g750 ( 
.A(n_748),
.B(n_622),
.Y(n_750)
);

NOR2xp67_ASAP7_75t_L g751 ( 
.A(n_747),
.B(n_709),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_750),
.Y(n_752)
);

AND3x4_ASAP7_75t_L g753 ( 
.A(n_749),
.B(n_708),
.C(n_691),
.Y(n_753)
);

NOR4xp25_ASAP7_75t_L g754 ( 
.A(n_751),
.B(n_726),
.C(n_648),
.D(n_722),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_750),
.Y(n_755)
);

INVxp33_ASAP7_75t_SL g756 ( 
.A(n_750),
.Y(n_756)
);

NOR4xp25_ASAP7_75t_L g757 ( 
.A(n_749),
.B(n_648),
.C(n_722),
.D(n_685),
.Y(n_757)
);

NOR4xp75_ASAP7_75t_SL g758 ( 
.A(n_756),
.B(n_704),
.C(n_658),
.D(n_689),
.Y(n_758)
);

INVx2_ASAP7_75t_L g759 ( 
.A(n_753),
.Y(n_759)
);

NAND5xp2_ASAP7_75t_L g760 ( 
.A(n_752),
.B(n_682),
.C(n_714),
.D(n_716),
.E(n_664),
.Y(n_760)
);

INVx2_ASAP7_75t_L g761 ( 
.A(n_755),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_754),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_757),
.B(n_714),
.Y(n_763)
);

OAI211xp5_ASAP7_75t_SL g764 ( 
.A1(n_752),
.A2(n_706),
.B(n_700),
.C(n_643),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_759),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_761),
.B(n_710),
.Y(n_766)
);

XNOR2xp5_ASAP7_75t_L g767 ( 
.A(n_762),
.B(n_637),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_763),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_758),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_764),
.Y(n_770)
);

INVxp67_ASAP7_75t_L g771 ( 
.A(n_760),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_762),
.B(n_716),
.Y(n_772)
);

NOR2xp33_ASAP7_75t_L g773 ( 
.A(n_765),
.B(n_710),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_772),
.Y(n_774)
);

XOR2xp5_ASAP7_75t_L g775 ( 
.A(n_767),
.B(n_700),
.Y(n_775)
);

INVxp67_ASAP7_75t_SL g776 ( 
.A(n_766),
.Y(n_776)
);

INVx2_ASAP7_75t_L g777 ( 
.A(n_770),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_771),
.B(n_613),
.Y(n_778)
);

INVxp67_ASAP7_75t_L g779 ( 
.A(n_768),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_769),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_765),
.Y(n_781)
);

INVx1_ASAP7_75t_L g782 ( 
.A(n_772),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_780),
.A2(n_651),
.B1(n_613),
.B2(n_670),
.Y(n_783)
);

OAI22xp33_ASAP7_75t_L g784 ( 
.A1(n_777),
.A2(n_706),
.B1(n_672),
.B2(n_712),
.Y(n_784)
);

AOI22xp5_ASAP7_75t_L g785 ( 
.A1(n_774),
.A2(n_613),
.B1(n_642),
.B2(n_672),
.Y(n_785)
);

AOI22xp33_ASAP7_75t_L g786 ( 
.A1(n_778),
.A2(n_782),
.B1(n_779),
.B2(n_781),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_779),
.A2(n_775),
.B1(n_773),
.B2(n_776),
.Y(n_787)
);

INVxp67_ASAP7_75t_SL g788 ( 
.A(n_781),
.Y(n_788)
);

AOI22x1_ASAP7_75t_L g789 ( 
.A1(n_788),
.A2(n_642),
.B1(n_647),
.B2(n_660),
.Y(n_789)
);

HB1xp67_ASAP7_75t_L g790 ( 
.A(n_787),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_786),
.A2(n_681),
.B1(n_660),
.B2(n_680),
.Y(n_791)
);

AOI22x1_ASAP7_75t_L g792 ( 
.A1(n_783),
.A2(n_785),
.B1(n_784),
.B2(n_660),
.Y(n_792)
);

OA22x2_ASAP7_75t_L g793 ( 
.A1(n_787),
.A2(n_705),
.B1(n_681),
.B2(n_581),
.Y(n_793)
);

XOR2x2_ASAP7_75t_L g794 ( 
.A(n_790),
.B(n_697),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_793),
.Y(n_795)
);

CKINVDCx20_ASAP7_75t_R g796 ( 
.A(n_791),
.Y(n_796)
);

OAI21xp5_ASAP7_75t_L g797 ( 
.A1(n_795),
.A2(n_792),
.B(n_789),
.Y(n_797)
);

AOI22xp5_ASAP7_75t_L g798 ( 
.A1(n_797),
.A2(n_796),
.B1(n_794),
.B2(n_562),
.Y(n_798)
);

OR2x6_ASAP7_75t_L g799 ( 
.A(n_798),
.B(n_705),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_799),
.A2(n_661),
.B1(n_680),
.B2(n_703),
.Y(n_800)
);


endmodule