module fake_jpeg_8092_n_339 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_339);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_339;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

BUFx24_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_SL g28 ( 
.A(n_0),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_12),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_37),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_41),
.Y(n_62)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g47 ( 
.A(n_22),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g49 ( 
.A(n_47),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_48),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_29),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_51),
.A2(n_45),
.B1(n_26),
.B2(n_46),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_68),
.Y(n_75)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_47),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_63),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

INVx1_ASAP7_75t_SL g86 ( 
.A(n_59),
.Y(n_86)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_19),
.B1(n_18),
.B2(n_29),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_61),
.A2(n_60),
.B1(n_45),
.B2(n_20),
.Y(n_94)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_64),
.B(n_63),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_41),
.B(n_32),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_66),
.B(n_32),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_43),
.B(n_19),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_40),
.A2(n_29),
.B1(n_25),
.B2(n_26),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_69),
.A2(n_32),
.B1(n_26),
.B2(n_25),
.Y(n_79)
);

OAI31xp33_ASAP7_75t_L g105 ( 
.A1(n_71),
.A2(n_57),
.A3(n_38),
.B(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_74),
.B(n_76),
.Y(n_109)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_62),
.Y(n_76)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_78),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_79),
.A2(n_92),
.B1(n_36),
.B2(n_30),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_80),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_81),
.A2(n_88),
.B1(n_89),
.B2(n_93),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_70),
.Y(n_84)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_84),
.Y(n_126)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_85),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_67),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_87),
.B(n_90),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_66),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g89 ( 
.A(n_66),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_67),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_68),
.A2(n_45),
.B1(n_30),
.B2(n_36),
.Y(n_92)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_62),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_96),
.B1(n_20),
.B2(n_33),
.Y(n_114)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_52),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_95),
.Y(n_111)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_56),
.Y(n_98)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_98),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_58),
.C(n_55),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_99),
.B(n_121),
.Y(n_147)
);

NAND2xp33_ASAP7_75t_SL g101 ( 
.A(n_84),
.B(n_38),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_101),
.A2(n_105),
.B(n_72),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_96),
.A2(n_56),
.B1(n_64),
.B2(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_102),
.A2(n_87),
.B1(n_90),
.B2(n_95),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_106),
.A2(n_114),
.B1(n_125),
.B2(n_126),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_112),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_75),
.B(n_59),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_79),
.A2(n_55),
.B1(n_67),
.B2(n_48),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_74),
.B1(n_73),
.B2(n_97),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_78),
.A2(n_21),
.B1(n_25),
.B2(n_50),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_116),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_93),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_118),
.B(n_123),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_77),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_124),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_71),
.A2(n_38),
.B(n_59),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_121),
.A2(n_38),
.B(n_86),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_71),
.B(n_59),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_72),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_128),
.B(n_132),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_129),
.A2(n_136),
.B(n_111),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_117),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_130),
.A2(n_143),
.B1(n_100),
.B2(n_117),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_131),
.A2(n_151),
.B(n_119),
.Y(n_159)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_122),
.Y(n_132)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_148),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_108),
.A2(n_91),
.B1(n_82),
.B2(n_81),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_134),
.A2(n_138),
.B1(n_141),
.B2(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_109),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_135),
.B(n_145),
.Y(n_184)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx4_ASAP7_75t_L g177 ( 
.A(n_137),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_120),
.A2(n_91),
.B1(n_82),
.B2(n_85),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_140),
.A2(n_146),
.B1(n_149),
.B2(n_154),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_102),
.A2(n_86),
.B1(n_98),
.B2(n_80),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_126),
.A2(n_83),
.B1(n_44),
.B2(n_42),
.Y(n_142)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_104),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_109),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_123),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_147),
.B(n_124),
.C(n_111),
.Y(n_162)
);

INVx13_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_99),
.A2(n_44),
.B1(n_42),
.B2(n_39),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_105),
.A2(n_118),
.B(n_110),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_153),
.B(n_106),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_125),
.A2(n_39),
.B1(n_37),
.B2(n_21),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_112),
.A2(n_119),
.B1(n_113),
.B2(n_101),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_155),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_158),
.A2(n_160),
.B1(n_163),
.B2(n_164),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_159),
.A2(n_174),
.B(n_186),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_152),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_144),
.B1(n_145),
.B2(n_135),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_162),
.B(n_173),
.C(n_178),
.Y(n_191)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_152),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_138),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_128),
.B(n_38),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g207 ( 
.A(n_166),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_142),
.Y(n_167)
);

OAI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_167),
.A2(n_168),
.B1(n_170),
.B2(n_179),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_129),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_169),
.A2(n_171),
.B(n_27),
.Y(n_196)
);

OA21x2_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_100),
.B(n_103),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_136),
.A2(n_127),
.B(n_37),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_172),
.Y(n_190)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_147),
.B(n_37),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g174 ( 
.A1(n_151),
.A2(n_27),
.B(n_31),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_139),
.B(n_115),
.Y(n_176)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_176),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_131),
.B(n_24),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_150),
.B(n_24),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_180),
.B(n_185),
.C(n_31),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_150),
.B(n_115),
.Y(n_181)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_17),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_155),
.B(n_24),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_144),
.A2(n_27),
.B(n_107),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_156),
.A2(n_168),
.B1(n_179),
.B2(n_183),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_187),
.A2(n_195),
.B1(n_207),
.B2(n_208),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_188),
.A2(n_189),
.B1(n_203),
.B2(n_214),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_156),
.A2(n_149),
.B1(n_146),
.B2(n_134),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_130),
.Y(n_193)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_193),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_165),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_194),
.B(n_202),
.Y(n_232)
);

O2A1O1Ixp33_ASAP7_75t_L g195 ( 
.A1(n_160),
.A2(n_154),
.B(n_133),
.C(n_35),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_195),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_196),
.B(n_186),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_137),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_209),
.C(n_210),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_169),
.A2(n_143),
.B(n_27),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_200),
.B(n_27),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_213),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_184),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_17),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_176),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_208),
.B(n_211),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_148),
.C(n_104),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_159),
.B(n_148),
.C(n_104),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_181),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_31),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_213),
.C(n_216),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_23),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_164),
.A2(n_23),
.B1(n_34),
.B2(n_35),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_182),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_215),
.B(n_167),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_180),
.B(n_35),
.C(n_34),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_202),
.B(n_177),
.Y(n_218)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_218),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_204),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_222),
.B(n_224),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_215),
.B(n_163),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_226),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_191),
.B(n_174),
.C(n_171),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_227),
.C(n_230),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_175),
.C(n_166),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_194),
.B(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_228),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_197),
.B(n_175),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_229),
.B(n_233),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_157),
.C(n_161),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_192),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_231),
.A2(n_234),
.B(n_206),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_201),
.B(n_157),
.C(n_170),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_35),
.C(n_34),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_236),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_210),
.B(n_23),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_187),
.B(n_10),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_190),
.B(n_34),
.C(n_17),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_1),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_16),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_196),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_241),
.A2(n_242),
.B1(n_214),
.B2(n_206),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_232),
.A2(n_200),
.B1(n_188),
.B2(n_203),
.Y(n_244)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_244),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_190),
.B1(n_205),
.B2(n_198),
.Y(n_245)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_245),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_246),
.B(n_265),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_248),
.B(n_250),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_230),
.A2(n_205),
.B1(n_198),
.B2(n_199),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_257),
.B1(n_260),
.B2(n_263),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_255),
.A2(n_219),
.B(n_223),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_233),
.A2(n_189),
.B1(n_216),
.B2(n_10),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_258),
.B(n_223),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_227),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_261),
.B(n_240),
.C(n_235),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_217),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_262),
.B(n_264),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_241),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_12),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_252),
.B(n_220),
.Y(n_267)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_267),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_268),
.B(n_271),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_247),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_225),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_273),
.A2(n_276),
.B(n_281),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_236),
.C(n_221),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_274),
.B(n_265),
.C(n_3),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_238),
.B(n_12),
.Y(n_276)
);

BUFx24_ASAP7_75t_SL g278 ( 
.A(n_258),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_278),
.B(n_283),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_252),
.B(n_11),
.Y(n_279)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_279),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_253),
.B(n_1),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_251),
.B(n_2),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_282),
.A2(n_261),
.B(n_3),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_245),
.B(n_2),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_275),
.A2(n_257),
.B1(n_246),
.B2(n_255),
.Y(n_284)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_284),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_270),
.B(n_256),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_285),
.B(n_287),
.C(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_277),
.B(n_254),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_291),
.B(n_297),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_280),
.A2(n_255),
.B1(n_263),
.B2(n_247),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_292),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_293),
.B(n_298),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_274),
.B(n_254),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_273),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_2),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_268),
.B(n_271),
.C(n_272),
.Y(n_298)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_289),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_299),
.B(n_306),
.Y(n_316)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_288),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_300),
.B(n_310),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_290),
.B(n_266),
.Y(n_305)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_305),
.Y(n_313)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_285),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_291),
.B(n_269),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_307),
.B(n_309),
.C(n_5),
.Y(n_320)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_287),
.A2(n_272),
.B(n_276),
.Y(n_308)
);

AOI21xp5_ASAP7_75t_L g315 ( 
.A1(n_308),
.A2(n_298),
.B(n_297),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_295),
.B(n_3),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g317 ( 
.A(n_311),
.B(n_5),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_299),
.B(n_296),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_314),
.B(n_317),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_320),
.Y(n_324)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_304),
.B(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_321),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_303),
.B(n_286),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_319),
.B(n_301),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_302),
.B(n_6),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g323 ( 
.A(n_313),
.B(n_300),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_316),
.B(n_312),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_327),
.C(n_328),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_318),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_322),
.A2(n_306),
.B(n_304),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_325),
.Y(n_333)
);

OAI21x1_ASAP7_75t_L g332 ( 
.A1(n_324),
.A2(n_307),
.B(n_7),
.Y(n_332)
);

AO21x1_ASAP7_75t_L g334 ( 
.A1(n_332),
.A2(n_6),
.B(n_7),
.Y(n_334)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_334),
.C(n_330),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_331),
.C(n_8),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_6),
.B(n_8),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_9),
.B(n_322),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_9),
.Y(n_339)
);


endmodule