module real_aes_11983_n_375 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_357, n_64, n_254, n_207, n_10, n_83, n_181, n_362, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_355, n_239, n_100, n_54, n_112, n_319, n_364, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_353, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_374, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_356, n_184, n_28, n_372, n_202, n_56, n_370, n_34, n_98, n_121, n_352, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_369, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_345, n_304, n_311, n_324, n_25, n_278, n_236, n_367, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_363, n_323, n_199, n_350, n_142, n_223, n_67, n_368, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_360, n_58, n_165, n_361, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_351, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_366, n_346, n_193, n_293, n_162, n_358, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_354, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_373, n_60, n_233, n_290, n_365, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_344, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_349, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_359, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_371, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_347, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_348, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_375);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_357;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_362;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_355;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_364;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_353;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_374;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_356;
input n_184;
input n_28;
input n_372;
input n_202;
input n_56;
input n_370;
input n_34;
input n_98;
input n_121;
input n_352;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_369;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_345;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_367;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_363;
input n_323;
input n_199;
input n_350;
input n_142;
input n_223;
input n_67;
input n_368;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_360;
input n_58;
input n_165;
input n_361;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_351;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_366;
input n_346;
input n_193;
input n_293;
input n_162;
input n_358;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_354;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_373;
input n_60;
input n_233;
input n_290;
input n_365;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_344;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_349;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_359;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_371;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_347;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_348;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_375;
wire n_476;
wire n_599;
wire n_887;
wire n_1279;
wire n_2014;
wire n_2003;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_1797;
wire n_933;
wire n_485;
wire n_822;
wire n_1641;
wire n_750;
wire n_503;
wire n_1781;
wire n_1762;
wire n_1591;
wire n_1903;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_1929;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1888;
wire n_1423;
wire n_571;
wire n_549;
wire n_1328;
wire n_1034;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_1972;
wire n_593;
wire n_2029;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_2006;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1936;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1873;
wire n_1835;
wire n_1871;
wire n_1468;
wire n_1713;
wire n_1967;
wire n_1920;
wire n_870;
wire n_1248;
wire n_2021;
wire n_1602;
wire n_548;
wire n_1859;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1845;
wire n_1415;
wire n_1160;
wire n_1849;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1805;
wire n_744;
wire n_1367;
wire n_1994;
wire n_1325;
wire n_1225;
wire n_1441;
wire n_875;
wire n_951;
wire n_1199;
wire n_1382;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1833;
wire n_1477;
wire n_1944;
wire n_595;
wire n_1893;
wire n_1960;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_2016;
wire n_962;
wire n_1599;
wire n_1959;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_874;
wire n_796;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_1771;
wire n_1809;
wire n_682;
wire n_1745;
wire n_1820;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_1883;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_2022;
wire n_885;
wire n_950;
wire n_381;
wire n_1981;
wire n_1196;
wire n_1013;
wire n_1905;
wire n_808;
wire n_1694;
wire n_1224;
wire n_1639;
wire n_1872;
wire n_688;
wire n_1042;
wire n_1588;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_527;
wire n_1676;
wire n_1342;
wire n_2018;
wire n_1440;
wire n_1966;
wire n_552;
wire n_1346;
wire n_1383;
wire n_1890;
wire n_1675;
wire n_1954;
wire n_590;
wire n_1293;
wire n_1880;
wire n_432;
wire n_1882;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1865;
wire n_1600;
wire n_805;
wire n_619;
wire n_1284;
wire n_1250;
wire n_1583;
wire n_1095;
wire n_1465;
wire n_859;
wire n_1987;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_1658;
wire n_1866;
wire n_954;
wire n_702;
wire n_1874;
wire n_1007;
wire n_1906;
wire n_898;
wire n_1926;
wire n_562;
wire n_1897;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_2004;
wire n_1201;
wire n_997;
wire n_2000;
wire n_1105;
wire n_1768;
wire n_1243;
wire n_1846;
wire n_1003;
wire n_749;
wire n_1870;
wire n_914;
wire n_1837;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1813;
wire n_1978;
wire n_1628;
wire n_1587;
wire n_1821;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1825;
wire n_1615;
wire n_1763;
wire n_928;
wire n_1384;
wire n_789;
wire n_2024;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1956;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_1940;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_1814;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_1921;
wire n_422;
wire n_861;
wire n_2007;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_1914;
wire n_440;
wire n_1945;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_1793;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1751;
wire n_1765;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_1787;
wire n_424;
wire n_877;
wire n_802;
wire n_1876;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1999;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1979;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1828;
wire n_1860;
wire n_2012;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_1973;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_667;
wire n_991;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_1951;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_1606;
wire n_1129;
wire n_1760;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1770;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_1750;
wire n_1852;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1830;
wire n_1594;
wire n_2020;
wire n_1864;
wire n_537;
wire n_1767;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1991;
wire n_1776;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_1499;
wire n_948;
wire n_399;
wire n_700;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1839;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1881;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1884;
wire n_1182;
wire n_872;
wire n_1401;
wire n_2017;
wire n_1946;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1210;
wire n_1741;
wire n_1456;
wire n_1879;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_860;
wire n_748;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_1853;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_2009;
wire n_925;
wire n_1389;
wire n_1393;
wire n_1977;
wire n_1930;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_2005;
wire n_508;
wire n_1141;
wire n_1769;
wire n_1812;
wire n_1985;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_1971;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_1854;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_1856;
wire n_531;
wire n_1848;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_1993;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_985;
wire n_777;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1773;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1766;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_2002;
wire n_734;
wire n_1623;
wire n_1907;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_1857;
wire n_1984;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_1234;
wire n_1915;
wire n_622;
wire n_1634;
wire n_1353;
wire n_1002;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_1862;
wire n_1965;
wire n_850;
wire n_720;
wire n_2023;
wire n_1026;
wire n_1756;
wire n_1803;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_1699;
wire n_1794;
wire n_1748;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_1970;
wire n_526;
wire n_1513;
wire n_2015;
wire n_1983;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_1934;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1784;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1806;
wire n_1829;
wire n_1133;
wire n_1775;
wire n_1593;
wire n_1976;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1807;
wire n_459;
wire n_1172;
wire n_998;
wire n_1689;
wire n_1625;
wire n_1910;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1957;
wire n_1184;
wire n_583;
wire n_1998;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1961;
wire n_1413;
wire n_1783;
wire n_1759;
wire n_1266;
wire n_497;
wire n_911;
wire n_1904;
wire n_450;
wire n_1578;
wire n_473;
wire n_1779;
wire n_967;
wire n_1709;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1908;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_1840;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_1795;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1451;
wire n_1069;
wire n_842;
wire n_1788;
wire n_1938;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_2019;
wire n_1816;
wire n_1952;
wire n_1811;
wire n_1066;
wire n_1917;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_1928;
wire n_943;
wire n_977;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1995;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_852;
wire n_1268;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_1980;
wire n_2013;
wire n_1446;
wire n_1778;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1932;
wire n_1707;
wire n_594;
wire n_856;
wire n_1146;
wire n_1685;
wire n_1810;
wire n_1435;
wire n_1800;
wire n_932;
wire n_958;
wire n_1755;
wire n_775;
wire n_763;
wire n_1093;
wire n_1990;
wire n_427;
wire n_1540;
wire n_519;
wire n_1878;
wire n_1116;
wire n_709;
wire n_1834;
wire n_388;
wire n_1913;
wire n_1470;
wire n_816;
wire n_1899;
wire n_625;
wire n_953;
wire n_1565;
wire n_1953;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_584;
wire n_896;
wire n_1817;
wire n_2008;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_1663;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1923;
wire n_2025;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1850;
wire n_1332;
wire n_1927;
wire n_1263;
wire n_1411;
wire n_1922;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1827;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1949;
wire n_1029;
wire n_1989;
wire n_1207;
wire n_1555;
wire n_1962;
wire n_664;
wire n_1017;
wire n_1942;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_1939;
wire n_609;
wire n_1743;
wire n_1752;
wire n_1792;
wire n_1006;
wire n_1869;
wire n_1259;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1895;
wire n_1670;
wire n_1941;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_1986;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_1786;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1764;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_1948;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1749;
wire n_1158;
wire n_1886;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_1832;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_1855;
wire n_1802;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1774;
wire n_1785;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1782;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1798;
wire n_1038;
wire n_1085;
wire n_2027;
wire n_845;
wire n_1838;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1753;
wire n_1244;
wire n_1581;
wire n_1863;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_628;
wire n_487;
wire n_831;
wire n_1772;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_2028;
wire n_1693;
wire n_1791;
wire n_418;
wire n_771;
wire n_1496;
wire n_524;
wire n_1378;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1824;
wire n_1933;
wire n_1270;
wire n_1988;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_1761;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_1790;
wire n_644;
wire n_1150;
wire n_1861;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_2011;
wire n_1757;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1799;
wire n_640;
wire n_1176;
wire n_1691;
wire n_1721;
wire n_1931;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_1804;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_1964;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1844;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1937;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_1841;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_1789;
wire n_987;
wire n_1596;
wire n_1982;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_2030;
wire n_1822;
wire n_718;
wire n_1955;
wire n_669;
wire n_1091;
wire n_1969;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_1777;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1819;
wire n_1887;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1902;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_1889;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_1896;
wire n_767;
wire n_889;
wire n_1398;
wire n_1911;
wire n_379;
wire n_1847;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1912;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_1747;
wire n_573;
wire n_1654;
wire n_1099;
wire n_626;
wire n_539;
wire n_1919;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_1754;
wire n_578;
wire n_892;
wire n_938;
wire n_774;
wire n_466;
wire n_1584;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1950;
wire n_984;
wire n_726;
wire n_517;
wire n_931;
wire n_780;
wire n_1851;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1360;
wire n_1082;
wire n_468;
wire n_1916;
wire n_532;
wire n_1025;
wire n_1875;
wire n_1826;
wire n_1836;
wire n_1909;
wire n_924;
wire n_1264;
wire n_1858;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1901;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1678;
wire n_1198;
wire n_1943;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1063;
wire n_1135;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_1818;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1780;
wire n_1974;
wire n_1547;
wire n_1823;
wire n_1867;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1891;
wire n_1267;
wire n_790;
wire n_1262;
wire n_1843;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1885;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1416;
wire n_1249;
wire n_387;
wire n_1239;
wire n_1796;
wire n_1662;
wire n_1992;
wire n_1963;
wire n_1958;
wire n_969;
wire n_1535;
wire n_2010;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1801;
wire n_1925;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_1968;
wire n_430;
wire n_1647;
wire n_1252;
wire n_1132;
wire n_1947;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_1996;
wire n_536;
wire n_851;
wire n_470;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_2001;
wire n_965;
wire n_1894;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1808;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1758;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_1877;
wire n_1900;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1842;
wire n_1536;
wire n_1746;
wire n_1898;
wire n_1711;
wire n_482;
wire n_633;
wire n_1892;
wire n_971;
wire n_1052;
wire n_1071;
wire n_2026;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_1573;
wire n_1130;
wire n_1918;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_1831;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_1997;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1815;
wire n_1924;
wire n_1412;
wire n_1868;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1975;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_394;
wire n_1280;
wire n_729;
wire n_1352;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1935;
wire n_1645;
wire n_429;
XNOR2xp5_ASAP7_75t_L g909 ( .A(n_0), .B(n_910), .Y(n_909) );
AO221x1_ASAP7_75t_L g1738 ( .A1(n_0), .A2(n_153), .B1(n_1706), .B2(n_1728), .C(n_1739), .Y(n_1738) );
CKINVDCx5p33_ASAP7_75t_R g1033 ( .A(n_1), .Y(n_1033) );
AOI22xp5_ASAP7_75t_L g1705 ( .A1(n_2), .A2(n_140), .B1(n_1706), .B2(n_1710), .Y(n_1705) );
AOI22xp33_ASAP7_75t_L g472 ( .A1(n_3), .A2(n_340), .B1(n_473), .B2(n_474), .Y(n_472) );
INVx1_ASAP7_75t_L g575 ( .A(n_3), .Y(n_575) );
INVxp33_ASAP7_75t_L g1946 ( .A(n_4), .Y(n_1946) );
AOI221xp5_ASAP7_75t_L g1976 ( .A1(n_4), .A2(n_103), .B1(n_473), .B2(n_1977), .C(n_1978), .Y(n_1976) );
INVx1_ASAP7_75t_L g1957 ( .A(n_5), .Y(n_1957) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_6), .A2(n_111), .B1(n_637), .B2(n_642), .Y(n_636) );
INVx1_ASAP7_75t_L g711 ( .A(n_6), .Y(n_711) );
CKINVDCx5p33_ASAP7_75t_R g445 ( .A(n_7), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g2021 ( .A1(n_8), .A2(n_221), .B1(n_545), .B2(n_808), .C(n_809), .Y(n_2021) );
OAI22xp33_ASAP7_75t_L g2026 ( .A1(n_8), .A2(n_337), .B1(n_422), .B2(n_969), .Y(n_2026) );
INVx1_ASAP7_75t_L g796 ( .A(n_9), .Y(n_796) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_9), .A2(n_117), .B1(n_479), .B2(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g934 ( .A(n_10), .Y(n_934) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_10), .A2(n_214), .B1(n_755), .B2(n_756), .Y(n_943) );
AOI221xp5_ASAP7_75t_L g1596 ( .A1(n_11), .A2(n_35), .B1(n_1597), .B2(n_1598), .C(n_1600), .Y(n_1596) );
INVx1_ASAP7_75t_L g1633 ( .A(n_11), .Y(n_1633) );
OAI22xp33_ASAP7_75t_L g757 ( .A1(n_12), .A2(n_110), .B1(n_517), .B2(n_558), .Y(n_757) );
AOI221xp5_ASAP7_75t_L g769 ( .A1(n_12), .A2(n_110), .B1(n_485), .B2(n_761), .C(n_770), .Y(n_769) );
AOI22xp33_ASAP7_75t_L g1505 ( .A1(n_13), .A2(n_23), .B1(n_1503), .B2(n_1506), .Y(n_1505) );
INVxp67_ASAP7_75t_SL g1511 ( .A(n_13), .Y(n_1511) );
AOI221xp5_ASAP7_75t_L g1263 ( .A1(n_14), .A2(n_289), .B1(n_744), .B2(n_747), .C(n_960), .Y(n_1263) );
OAI22xp33_ASAP7_75t_L g1269 ( .A1(n_14), .A2(n_115), .B1(n_971), .B2(n_973), .Y(n_1269) );
AOI22xp33_ASAP7_75t_L g810 ( .A1(n_15), .A2(n_124), .B1(n_811), .B2(n_813), .Y(n_810) );
AOI22xp33_ASAP7_75t_SL g821 ( .A1(n_15), .A2(n_124), .B1(n_822), .B2(n_823), .Y(n_821) );
INVx1_ASAP7_75t_L g1655 ( .A(n_16), .Y(n_1655) );
OAI211xp5_ASAP7_75t_SL g1673 ( .A1(n_16), .A2(n_517), .B(n_1674), .C(n_1680), .Y(n_1673) );
INVx1_ASAP7_75t_L g1740 ( .A(n_17), .Y(n_1740) );
AOI221xp5_ASAP7_75t_L g1137 ( .A1(n_18), .A2(n_321), .B1(n_694), .B2(n_747), .C(n_799), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1146 ( .A1(n_18), .A2(n_321), .B1(n_479), .B2(n_1147), .Y(n_1146) );
INVx1_ASAP7_75t_L g1553 ( .A(n_19), .Y(n_1553) );
AOI22xp33_ASAP7_75t_SL g1567 ( .A1(n_19), .A2(n_307), .B1(n_825), .B2(n_1568), .Y(n_1567) );
CKINVDCx5p33_ASAP7_75t_R g1650 ( .A(n_20), .Y(n_1650) );
AOI22xp33_ASAP7_75t_SL g1491 ( .A1(n_21), .A2(n_39), .B1(n_799), .B2(n_1492), .Y(n_1491) );
AOI22xp33_ASAP7_75t_L g1502 ( .A1(n_21), .A2(n_39), .B1(n_1503), .B2(n_1504), .Y(n_1502) );
CKINVDCx20_ASAP7_75t_R g1193 ( .A(n_22), .Y(n_1193) );
INVxp33_ASAP7_75t_L g1518 ( .A(n_23), .Y(n_1518) );
CKINVDCx5p33_ASAP7_75t_R g1345 ( .A(n_24), .Y(n_1345) );
INVx1_ASAP7_75t_L g1377 ( .A(n_25), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1436 ( .A1(n_25), .A2(n_243), .B1(n_1437), .B2(n_1438), .C(n_1440), .Y(n_1436) );
AOI22xp33_ASAP7_75t_L g1332 ( .A1(n_26), .A2(n_98), .B1(n_1333), .B2(n_1334), .Y(n_1332) );
INVx1_ASAP7_75t_L g1359 ( .A(n_26), .Y(n_1359) );
XNOR2xp5_ASAP7_75t_L g1167 ( .A(n_27), .B(n_1168), .Y(n_1167) );
AOI22xp33_ASAP7_75t_SL g814 ( .A1(n_28), .A2(n_106), .B1(n_811), .B2(n_815), .Y(n_814) );
INVxp67_ASAP7_75t_SL g847 ( .A(n_28), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g2003 ( .A1(n_29), .A2(n_371), .B1(n_1180), .B2(n_1284), .Y(n_2003) );
INVxp67_ASAP7_75t_SL g2016 ( .A(n_29), .Y(n_2016) );
AOI22xp33_ASAP7_75t_L g1586 ( .A1(n_30), .A2(n_148), .B1(n_1587), .B2(n_1588), .Y(n_1586) );
INVx1_ASAP7_75t_L g1614 ( .A(n_30), .Y(n_1614) );
OAI222xp33_ASAP7_75t_L g1027 ( .A1(n_31), .A2(n_77), .B1(n_161), .B2(n_836), .C1(n_839), .C2(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1043 ( .A(n_31), .Y(n_1043) );
CKINVDCx5p33_ASAP7_75t_R g1105 ( .A(n_32), .Y(n_1105) );
CKINVDCx5p33_ASAP7_75t_R g1590 ( .A(n_33), .Y(n_1590) );
OAI22xp5_ASAP7_75t_L g1277 ( .A1(n_34), .A2(n_231), .B1(n_460), .B2(n_1278), .Y(n_1277) );
INVx1_ASAP7_75t_L g1306 ( .A(n_34), .Y(n_1306) );
INVx1_ASAP7_75t_L g1629 ( .A(n_35), .Y(n_1629) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_36), .A2(n_224), .B1(n_545), .B2(n_1126), .C(n_1127), .Y(n_1125) );
INVx1_ASAP7_75t_L g1154 ( .A(n_36), .Y(n_1154) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_37), .B(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g709 ( .A(n_37), .Y(n_709) );
CKINVDCx5p33_ASAP7_75t_R g1652 ( .A(n_38), .Y(n_1652) );
CKINVDCx5p33_ASAP7_75t_R g1536 ( .A(n_40), .Y(n_1536) );
AOI22xp33_ASAP7_75t_L g1076 ( .A1(n_41), .A2(n_171), .B1(n_491), .B2(n_1077), .Y(n_1076) );
AOI22xp33_ASAP7_75t_SL g1095 ( .A1(n_41), .A2(n_171), .B1(n_947), .B2(n_1096), .Y(n_1095) );
INVx1_ASAP7_75t_L g382 ( .A(n_42), .Y(n_382) );
INVx1_ASAP7_75t_L g1935 ( .A(n_43), .Y(n_1935) );
CKINVDCx5p33_ASAP7_75t_R g1982 ( .A(n_44), .Y(n_1982) );
CKINVDCx5p33_ASAP7_75t_R g1425 ( .A(n_45), .Y(n_1425) );
AOI22xp33_ASAP7_75t_L g1122 ( .A1(n_46), .A2(n_175), .B1(n_1123), .B2(n_1124), .Y(n_1122) );
INVx1_ASAP7_75t_L g1155 ( .A(n_46), .Y(n_1155) );
CKINVDCx5p33_ASAP7_75t_R g1413 ( .A(n_47), .Y(n_1413) );
AOI22xp5_ASAP7_75t_L g1764 ( .A1(n_48), .A2(n_162), .B1(n_1706), .B2(n_1710), .Y(n_1764) );
INVxp67_ASAP7_75t_SL g800 ( .A(n_49), .Y(n_800) );
OAI22xp33_ASAP7_75t_L g835 ( .A1(n_49), .A2(n_194), .B1(n_836), .B2(n_839), .Y(n_835) );
INVx1_ASAP7_75t_L g855 ( .A(n_50), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_50), .A2(n_241), .B1(n_808), .B2(n_885), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g1283 ( .A1(n_51), .A2(n_316), .B1(n_1180), .B2(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1315 ( .A(n_51), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g884 ( .A1(n_52), .A2(n_163), .B1(n_542), .B2(n_885), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g896 ( .A1(n_52), .A2(n_163), .B1(n_761), .B2(n_825), .Y(n_896) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_53), .A2(n_266), .B1(n_479), .B2(n_480), .Y(n_478) );
INVx1_ASAP7_75t_L g566 ( .A(n_53), .Y(n_566) );
INVx1_ASAP7_75t_L g1347 ( .A(n_54), .Y(n_1347) );
INVx1_ASAP7_75t_L g1576 ( .A(n_55), .Y(n_1576) );
XNOR2xp5_ASAP7_75t_L g1640 ( .A(n_56), .B(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1241 ( .A(n_57), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1249 ( .A1(n_57), .A2(n_558), .B1(n_952), .B2(n_1250), .C(n_1255), .Y(n_1249) );
AO221x2_ASAP7_75t_L g1725 ( .A1(n_58), .A2(n_300), .B1(n_1726), .B2(n_1728), .C(n_1730), .Y(n_1725) );
INVxp33_ASAP7_75t_L g1933 ( .A(n_59), .Y(n_1933) );
AOI221xp5_ASAP7_75t_L g1966 ( .A1(n_59), .A2(n_130), .B1(n_1967), .B2(n_1969), .C(n_1970), .Y(n_1966) );
INVx1_ASAP7_75t_L g1344 ( .A(n_60), .Y(n_1344) );
AOI221xp5_ASAP7_75t_L g1352 ( .A1(n_60), .A2(n_220), .B1(n_818), .B2(n_1303), .C(n_1353), .Y(n_1352) );
AOI22xp33_ASAP7_75t_L g1487 ( .A1(n_61), .A2(n_72), .B1(n_1488), .B2(n_1489), .Y(n_1487) );
AOI22xp33_ASAP7_75t_L g1498 ( .A1(n_61), .A2(n_72), .B1(n_1499), .B2(n_1500), .Y(n_1498) );
INVx1_ASAP7_75t_L g2002 ( .A(n_62), .Y(n_2002) );
INVx1_ASAP7_75t_L g997 ( .A(n_63), .Y(n_997) );
INVx1_ASAP7_75t_L g1407 ( .A(n_64), .Y(n_1407) );
AOI221xp5_ASAP7_75t_L g1448 ( .A1(n_64), .A2(n_186), .B1(n_1437), .B2(n_1449), .C(n_1451), .Y(n_1448) );
INVx1_ASAP7_75t_L g1215 ( .A(n_65), .Y(n_1215) );
OAI22xp33_ASAP7_75t_L g1221 ( .A1(n_65), .A2(n_145), .B1(n_422), .B2(n_969), .Y(n_1221) );
INVxp33_ASAP7_75t_L g1943 ( .A(n_66), .Y(n_1943) );
AOI22xp33_ASAP7_75t_L g1980 ( .A1(n_66), .A2(n_319), .B1(n_485), .B2(n_936), .Y(n_1980) );
INVxp33_ASAP7_75t_L g1473 ( .A(n_67), .Y(n_1473) );
AOI22xp33_ASAP7_75t_SL g1493 ( .A1(n_67), .A2(n_154), .B1(n_1488), .B2(n_1494), .Y(n_1493) );
AOI22xp33_ASAP7_75t_L g1288 ( .A1(n_68), .A2(n_361), .B1(n_1289), .B2(n_1290), .Y(n_1288) );
OAI22xp5_ASAP7_75t_L g1316 ( .A1(n_68), .A2(n_361), .B1(n_583), .B2(n_588), .Y(n_1316) );
OAI221xp5_ASAP7_75t_L g1939 ( .A1(n_69), .A2(n_255), .B1(n_1395), .B2(n_1622), .C(n_1940), .Y(n_1939) );
OAI22xp5_ASAP7_75t_L g1962 ( .A1(n_69), .A2(n_255), .B1(n_1963), .B2(n_1964), .Y(n_1962) );
INVx1_ASAP7_75t_L g1046 ( .A(n_70), .Y(n_1046) );
AOI22xp33_ASAP7_75t_SL g1065 ( .A1(n_70), .A2(n_123), .B1(n_761), .B2(n_902), .Y(n_1065) );
AOI22xp33_ASAP7_75t_L g1179 ( .A1(n_71), .A2(n_374), .B1(n_1180), .B2(n_1181), .Y(n_1179) );
INVx1_ASAP7_75t_L g1201 ( .A(n_71), .Y(n_1201) );
INVx1_ASAP7_75t_L g732 ( .A(n_73), .Y(n_732) );
AOI221xp5_ASAP7_75t_L g760 ( .A1(n_73), .A2(n_274), .B1(n_761), .B2(n_763), .C(n_765), .Y(n_760) );
NOR2xp33_ASAP7_75t_L g1118 ( .A(n_74), .B(n_1119), .Y(n_1118) );
CKINVDCx5p33_ASAP7_75t_R g1648 ( .A(n_75), .Y(n_1648) );
OAI22xp33_ASAP7_75t_L g1532 ( .A1(n_76), .A2(n_338), .B1(n_583), .B2(n_588), .Y(n_1532) );
AOI22xp33_ASAP7_75t_L g1570 ( .A1(n_76), .A2(n_338), .B1(n_671), .B2(n_823), .Y(n_1570) );
AOI22xp33_ASAP7_75t_SL g1050 ( .A1(n_77), .A2(n_327), .B1(n_542), .B2(n_1051), .Y(n_1050) );
AOI22xp33_ASAP7_75t_L g1747 ( .A1(n_78), .A2(n_329), .B1(n_1706), .B2(n_1710), .Y(n_1747) );
INVx1_ASAP7_75t_L g1287 ( .A(n_79), .Y(n_1287) );
OAI211xp5_ASAP7_75t_SL g1295 ( .A1(n_79), .A2(n_517), .B(n_1296), .C(n_1304), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g882 ( .A1(n_80), .A2(n_216), .B1(n_811), .B2(n_883), .Y(n_882) );
AOI22xp33_ASAP7_75t_L g893 ( .A1(n_80), .A2(n_216), .B1(n_822), .B2(n_894), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g1693 ( .A1(n_81), .A2(n_355), .B1(n_1694), .B2(n_1702), .Y(n_1693) );
AOI22xp33_ASAP7_75t_L g1335 ( .A1(n_82), .A2(n_320), .B1(n_431), .B2(n_1336), .Y(n_1335) );
OAI221xp5_ASAP7_75t_L g1356 ( .A1(n_82), .A2(n_558), .B1(n_580), .B2(n_1357), .C(n_1362), .Y(n_1356) );
INVx1_ASAP7_75t_L g1472 ( .A(n_83), .Y(n_1472) );
CKINVDCx5p33_ASAP7_75t_R g409 ( .A(n_84), .Y(n_409) );
CKINVDCx5p33_ASAP7_75t_R g1605 ( .A(n_85), .Y(n_1605) );
OAI22xp33_ASAP7_75t_L g1662 ( .A1(n_86), .A2(n_362), .B1(n_1245), .B2(n_1246), .Y(n_1662) );
INVx1_ASAP7_75t_L g1682 ( .A(n_86), .Y(n_1682) );
AO22x1_ASAP7_75t_L g1750 ( .A1(n_87), .A2(n_283), .B1(n_1710), .B2(n_1751), .Y(n_1750) );
CKINVDCx5p33_ASAP7_75t_R g1282 ( .A(n_88), .Y(n_1282) );
OAI22xp5_ASAP7_75t_L g1591 ( .A1(n_89), .A2(n_269), .B1(n_1592), .B2(n_1593), .Y(n_1591) );
OAI221xp5_ASAP7_75t_L g1621 ( .A1(n_89), .A2(n_269), .B1(n_1395), .B2(n_1397), .C(n_1622), .Y(n_1621) );
CKINVDCx5p33_ASAP7_75t_R g985 ( .A(n_90), .Y(n_985) );
CKINVDCx5p33_ASAP7_75t_R g1415 ( .A(n_91), .Y(n_1415) );
AOI22xp33_ASAP7_75t_L g484 ( .A1(n_92), .A2(n_363), .B1(n_480), .B2(n_485), .Y(n_484) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_92), .A2(n_558), .B1(n_560), .B2(n_574), .C(n_580), .Y(n_557) );
INVx1_ASAP7_75t_L g856 ( .A(n_93), .Y(n_856) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_93), .A2(n_181), .B1(n_811), .B2(n_889), .Y(n_888) );
AO22x1_ASAP7_75t_L g1752 ( .A1(n_94), .A2(n_282), .B1(n_1694), .B2(n_1702), .Y(n_1752) );
CKINVDCx5p33_ASAP7_75t_R g1341 ( .A(n_95), .Y(n_1341) );
CKINVDCx5p33_ASAP7_75t_R g926 ( .A(n_96), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g1177 ( .A(n_97), .Y(n_1177) );
INVx1_ASAP7_75t_L g1361 ( .A(n_98), .Y(n_1361) );
INVx1_ASAP7_75t_L g988 ( .A(n_99), .Y(n_988) );
OAI221xp5_ASAP7_75t_L g1000 ( .A1(n_99), .A2(n_558), .B1(n_952), .B2(n_1001), .C(n_1004), .Y(n_1000) );
INVx1_ASAP7_75t_L g1661 ( .A(n_100), .Y(n_1661) );
OAI22xp5_ASAP7_75t_L g1666 ( .A1(n_100), .A2(n_322), .B1(n_755), .B2(n_756), .Y(n_1666) );
CKINVDCx20_ASAP7_75t_R g1997 ( .A(n_101), .Y(n_1997) );
XNOR2x2_ASAP7_75t_L g722 ( .A(n_102), .B(n_723), .Y(n_722) );
INVxp67_ASAP7_75t_L g1948 ( .A(n_103), .Y(n_1948) );
INVxp67_ASAP7_75t_SL g788 ( .A(n_104), .Y(n_788) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_104), .A2(n_280), .B1(n_822), .B2(n_831), .Y(n_830) );
CKINVDCx5p33_ASAP7_75t_R g746 ( .A(n_105), .Y(n_746) );
INVxp33_ASAP7_75t_L g846 ( .A(n_106), .Y(n_846) );
INVx1_ASAP7_75t_L g419 ( .A(n_107), .Y(n_419) );
BUFx2_ASAP7_75t_L g471 ( .A(n_107), .Y(n_471) );
BUFx2_ASAP7_75t_L g493 ( .A(n_107), .Y(n_493) );
OR2x2_ASAP7_75t_L g1394 ( .A(n_107), .B(n_511), .Y(n_1394) );
OAI22xp33_ASAP7_75t_L g995 ( .A1(n_108), .A2(n_114), .B1(n_447), .B2(n_460), .Y(n_995) );
INVx1_ASAP7_75t_L g1016 ( .A(n_108), .Y(n_1016) );
INVx1_ASAP7_75t_L g1298 ( .A(n_109), .Y(n_1298) );
OAI22xp5_ASAP7_75t_L g1319 ( .A1(n_109), .A2(n_211), .B1(n_971), .B2(n_973), .Y(n_1319) );
INVx1_ASAP7_75t_L g621 ( .A(n_111), .Y(n_621) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_112), .Y(n_730) );
INVx1_ASAP7_75t_L g429 ( .A(n_113), .Y(n_429) );
AOI221xp5_ASAP7_75t_L g539 ( .A1(n_113), .A2(n_314), .B1(n_540), .B2(n_542), .C(n_545), .Y(n_539) );
INVx1_ASAP7_75t_L g1015 ( .A(n_114), .Y(n_1015) );
INVx1_ASAP7_75t_L g1261 ( .A(n_115), .Y(n_1261) );
AOI22xp33_ASAP7_75t_L g816 ( .A1(n_116), .A2(n_227), .B1(n_808), .B2(n_817), .Y(n_816) );
INVxp67_ASAP7_75t_SL g834 ( .A(n_116), .Y(n_834) );
INVxp33_ASAP7_75t_L g791 ( .A(n_117), .Y(n_791) );
AO221x1_ASAP7_75t_L g1100 ( .A1(n_118), .A2(n_223), .B1(n_743), .B2(n_744), .C(n_818), .Y(n_1100) );
INVx1_ASAP7_75t_L g1111 ( .A(n_118), .Y(n_1111) );
AOI22xp33_ASAP7_75t_L g1602 ( .A1(n_119), .A2(n_296), .B1(n_1333), .B2(n_1603), .Y(n_1602) );
INVx1_ASAP7_75t_L g1634 ( .A(n_119), .Y(n_1634) );
INVx1_ASAP7_75t_L g1040 ( .A(n_120), .Y(n_1040) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_120), .A2(n_245), .B1(n_491), .B2(n_822), .Y(n_1066) );
AOI221xp5_ASAP7_75t_L g1302 ( .A1(n_121), .A2(n_211), .B1(n_808), .B2(n_817), .C(n_1303), .Y(n_1302) );
OAI22xp5_ASAP7_75t_L g1318 ( .A1(n_121), .A2(n_261), .B1(n_422), .B2(n_969), .Y(n_1318) );
INVxp67_ASAP7_75t_SL g1475 ( .A(n_122), .Y(n_1475) );
AOI22xp33_ASAP7_75t_SL g1495 ( .A1(n_122), .A2(n_234), .B1(n_1492), .B2(n_1496), .Y(n_1495) );
INVx1_ASAP7_75t_L g1042 ( .A(n_123), .Y(n_1042) );
AO221x1_ASAP7_75t_L g1712 ( .A1(n_125), .A2(n_141), .B1(n_1706), .B2(n_1710), .C(n_1713), .Y(n_1712) );
AOI22xp33_ASAP7_75t_L g1508 ( .A1(n_126), .A2(n_238), .B1(n_1180), .B2(n_1284), .Y(n_1508) );
INVxp33_ASAP7_75t_SL g1515 ( .A(n_126), .Y(n_1515) );
INVx1_ASAP7_75t_L g994 ( .A(n_127), .Y(n_994) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_127), .A2(n_249), .B1(n_755), .B2(n_756), .Y(n_999) );
AO22x2_ASAP7_75t_L g1022 ( .A1(n_128), .A2(n_1023), .B1(n_1024), .B2(n_1069), .Y(n_1022) );
INVxp67_ASAP7_75t_SL g1023 ( .A(n_128), .Y(n_1023) );
AO221x1_ASAP7_75t_L g1719 ( .A1(n_128), .A2(n_343), .B1(n_1706), .B2(n_1710), .C(n_1720), .Y(n_1719) );
INVx1_ASAP7_75t_L g1722 ( .A(n_129), .Y(n_1722) );
INVxp33_ASAP7_75t_L g1938 ( .A(n_130), .Y(n_1938) );
XNOR2xp5_ASAP7_75t_L g975 ( .A(n_131), .B(n_976), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_132), .A2(n_304), .B1(n_825), .B2(n_1079), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g1097 ( .A1(n_132), .A2(n_304), .B1(n_694), .B2(n_747), .C(n_960), .Y(n_1097) );
CKINVDCx5p33_ASAP7_75t_R g1326 ( .A(n_133), .Y(n_1326) );
CKINVDCx5p33_ASAP7_75t_R g1325 ( .A(n_134), .Y(n_1325) );
AOI22xp33_ASAP7_75t_L g1329 ( .A1(n_135), .A2(n_160), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx1_ASAP7_75t_L g1363 ( .A(n_135), .Y(n_1363) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_136), .A2(n_226), .B1(n_540), .B2(n_542), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_136), .A2(n_226), .B1(n_761), .B2(n_825), .Y(n_1062) );
OAI22xp33_ASAP7_75t_L g1190 ( .A1(n_137), .A2(n_215), .B1(n_460), .B2(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g1219 ( .A(n_137), .Y(n_1219) );
CKINVDCx5p33_ASAP7_75t_R g1236 ( .A(n_138), .Y(n_1236) );
INVx1_ASAP7_75t_L g1717 ( .A(n_139), .Y(n_1717) );
OA22x2_ASAP7_75t_L g599 ( .A1(n_140), .A2(n_600), .B1(n_720), .B2(n_721), .Y(n_599) );
INVxp67_ASAP7_75t_SL g721 ( .A(n_140), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g1763 ( .A1(n_142), .A2(n_167), .B1(n_1694), .B2(n_1702), .Y(n_1763) );
INVx1_ASAP7_75t_L g2019 ( .A(n_143), .Y(n_2019) );
OAI22xp33_ASAP7_75t_L g2027 ( .A1(n_143), .A2(n_221), .B1(n_971), .B2(n_973), .Y(n_2027) );
XNOR2xp5_ASAP7_75t_L g403 ( .A(n_144), .B(n_404), .Y(n_403) );
AOI221xp5_ASAP7_75t_L g1216 ( .A1(n_145), .A2(n_325), .B1(n_744), .B2(n_808), .C(n_809), .Y(n_1216) );
CKINVDCx5p33_ASAP7_75t_R g1542 ( .A(n_146), .Y(n_1542) );
XNOR2xp5_ASAP7_75t_L g1993 ( .A(n_147), .B(n_1994), .Y(n_1993) );
INVx1_ASAP7_75t_L g1619 ( .A(n_148), .Y(n_1619) );
INVx1_ASAP7_75t_L g2005 ( .A(n_149), .Y(n_2005) );
OAI221xp5_ASAP7_75t_L g2011 ( .A1(n_149), .A2(n_558), .B1(n_580), .B2(n_2012), .C(n_2014), .Y(n_2011) );
INVx1_ASAP7_75t_L g1731 ( .A(n_150), .Y(n_1731) );
INVx1_ASAP7_75t_L g874 ( .A(n_151), .Y(n_874) );
AOI22xp33_ASAP7_75t_SL g901 ( .A1(n_151), .A2(n_336), .B1(n_761), .B2(n_902), .Y(n_901) );
CKINVDCx5p33_ASAP7_75t_R g738 ( .A(n_152), .Y(n_738) );
INVxp33_ASAP7_75t_SL g1470 ( .A(n_154), .Y(n_1470) );
AOI22xp33_ASAP7_75t_L g488 ( .A1(n_155), .A2(n_219), .B1(n_489), .B2(n_491), .Y(n_488) );
OAI22xp5_ASAP7_75t_L g582 ( .A1(n_155), .A2(n_219), .B1(n_583), .B2(n_588), .Y(n_582) );
INVx1_ASAP7_75t_L g1551 ( .A(n_156), .Y(n_1551) );
AOI22xp33_ASAP7_75t_L g1565 ( .A1(n_156), .A2(n_310), .B1(n_489), .B2(n_1566), .Y(n_1565) );
CKINVDCx5p33_ASAP7_75t_R g438 ( .A(n_157), .Y(n_438) );
INVx1_ASAP7_75t_L g1211 ( .A(n_158), .Y(n_1211) );
OAI22xp33_ASAP7_75t_L g1222 ( .A1(n_158), .A2(n_325), .B1(n_971), .B2(n_973), .Y(n_1222) );
CKINVDCx5p33_ASAP7_75t_R g622 ( .A(n_159), .Y(n_622) );
INVx1_ASAP7_75t_L g1365 ( .A(n_160), .Y(n_1365) );
INVx1_ASAP7_75t_L g1044 ( .A(n_161), .Y(n_1044) );
INVx1_ASAP7_75t_L g1698 ( .A(n_164), .Y(n_1698) );
OAI22xp33_ASAP7_75t_L g1244 ( .A1(n_165), .A2(n_353), .B1(n_1245), .B2(n_1246), .Y(n_1244) );
INVx1_ASAP7_75t_L g1265 ( .A(n_165), .Y(n_1265) );
INVx1_ASAP7_75t_L g1937 ( .A(n_166), .Y(n_1937) );
INVx1_ASAP7_75t_L g1721 ( .A(n_168), .Y(n_1721) );
INVx1_ASAP7_75t_L g869 ( .A(n_169), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g903 ( .A1(n_169), .A2(n_213), .B1(n_440), .B2(n_894), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g1237 ( .A1(n_170), .A2(n_369), .B1(n_936), .B2(n_1189), .Y(n_1237) );
INVx1_ASAP7_75t_L g1252 ( .A(n_170), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1337 ( .A1(n_172), .A2(n_302), .B1(n_1180), .B2(n_1284), .Y(n_1337) );
OAI22xp5_ASAP7_75t_L g1368 ( .A1(n_172), .A2(n_302), .B1(n_583), .B2(n_756), .Y(n_1368) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_173), .A2(n_330), .B1(n_1123), .B2(n_1139), .Y(n_1138) );
AOI22xp33_ASAP7_75t_L g1144 ( .A1(n_173), .A2(n_330), .B1(n_767), .B2(n_1145), .Y(n_1144) );
INVx1_ASAP7_75t_L g1558 ( .A(n_174), .Y(n_1558) );
INVx1_ASAP7_75t_L g1151 ( .A(n_175), .Y(n_1151) );
INVx1_ASAP7_75t_L g792 ( .A(n_176), .Y(n_792) );
INVx1_ASAP7_75t_L g1699 ( .A(n_177), .Y(n_1699) );
NAND2xp5_ASAP7_75t_L g1704 ( .A(n_177), .B(n_1697), .Y(n_1704) );
INVx1_ASAP7_75t_L g1476 ( .A(n_178), .Y(n_1476) );
OAI22xp5_ASAP7_75t_L g1512 ( .A1(n_178), .A2(n_365), .B1(n_802), .B2(n_1513), .Y(n_1512) );
INVx1_ASAP7_75t_L g1242 ( .A(n_179), .Y(n_1242) );
OAI211xp5_ASAP7_75t_SL g1258 ( .A1(n_179), .A2(n_517), .B(n_1259), .C(n_1264), .Y(n_1258) );
INVx2_ASAP7_75t_L g394 ( .A(n_180), .Y(n_394) );
INVx1_ASAP7_75t_L g859 ( .A(n_181), .Y(n_859) );
OAI22xp5_ASAP7_75t_L g2008 ( .A1(n_182), .A2(n_230), .B1(n_1246), .B2(n_1278), .Y(n_2008) );
INVx1_ASAP7_75t_L g2023 ( .A(n_182), .Y(n_2023) );
AOI22xp33_ASAP7_75t_L g1056 ( .A1(n_183), .A2(n_292), .B1(n_1057), .B2(n_1058), .Y(n_1056) );
AOI22xp33_ASAP7_75t_L g1063 ( .A1(n_183), .A2(n_292), .B1(n_473), .B2(n_491), .Y(n_1063) );
CKINVDCx5p33_ASAP7_75t_R g673 ( .A(n_184), .Y(n_673) );
AOI22xp33_ASAP7_75t_L g1186 ( .A1(n_185), .A2(n_366), .B1(n_894), .B2(n_1187), .Y(n_1186) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_185), .A2(n_366), .B1(n_583), .B2(n_588), .Y(n_1195) );
INVx1_ASAP7_75t_L g1409 ( .A(n_186), .Y(n_1409) );
INVx1_ASAP7_75t_L g415 ( .A(n_187), .Y(n_415) );
BUFx3_ASAP7_75t_L g435 ( .A(n_187), .Y(n_435) );
INVx1_ASAP7_75t_L g1411 ( .A(n_188), .Y(n_1411) );
AOI22xp33_ASAP7_75t_L g1452 ( .A1(n_188), .A2(n_225), .B1(n_1145), .B2(n_1453), .Y(n_1452) );
INVx1_ASAP7_75t_L g1262 ( .A(n_189), .Y(n_1262) );
OAI22xp33_ASAP7_75t_L g1268 ( .A1(n_189), .A2(n_289), .B1(n_422), .B2(n_969), .Y(n_1268) );
INVx1_ASAP7_75t_L g1136 ( .A(n_190), .Y(n_1136) );
AOI22xp33_ASAP7_75t_L g1148 ( .A1(n_190), .A2(n_285), .B1(n_431), .B2(n_498), .Y(n_1148) );
CKINVDCx5p33_ASAP7_75t_R g654 ( .A(n_191), .Y(n_654) );
CKINVDCx5p33_ASAP7_75t_R g1103 ( .A(n_192), .Y(n_1103) );
OAI22xp33_ASAP7_75t_L g939 ( .A1(n_193), .A2(n_351), .B1(n_447), .B2(n_460), .Y(n_939) );
INVx1_ASAP7_75t_L g962 ( .A(n_193), .Y(n_962) );
INVx1_ASAP7_75t_L g803 ( .A(n_194), .Y(n_803) );
CKINVDCx5p33_ASAP7_75t_R g628 ( .A(n_195), .Y(n_628) );
CKINVDCx5p33_ASAP7_75t_R g1384 ( .A(n_196), .Y(n_1384) );
AOI221xp5_ASAP7_75t_L g959 ( .A1(n_197), .A2(n_358), .B1(n_743), .B2(n_744), .C(n_960), .Y(n_959) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_197), .A2(n_222), .B1(n_971), .B2(n_973), .Y(n_970) );
INVx1_ASAP7_75t_L g1010 ( .A(n_198), .Y(n_1010) );
OAI22xp33_ASAP7_75t_L g1019 ( .A1(n_198), .A2(n_200), .B1(n_971), .B2(n_973), .Y(n_1019) );
OAI22xp5_ASAP7_75t_L g754 ( .A1(n_199), .A2(n_342), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g772 ( .A(n_199), .Y(n_772) );
AOI221xp5_ASAP7_75t_L g1013 ( .A1(n_200), .A2(n_242), .B1(n_743), .B2(n_744), .C(n_799), .Y(n_1013) );
OAI221xp5_ASAP7_75t_L g860 ( .A1(n_201), .A2(n_273), .B1(n_839), .B2(n_861), .C(n_862), .Y(n_860) );
INVx1_ASAP7_75t_L g872 ( .A(n_201), .Y(n_872) );
INVx1_ASAP7_75t_L g2006 ( .A(n_202), .Y(n_2006) );
OAI211xp5_ASAP7_75t_SL g2017 ( .A1(n_202), .A2(n_517), .B(n_2018), .C(n_2022), .Y(n_2017) );
INVx1_ASAP7_75t_L g1953 ( .A(n_203), .Y(n_1953) );
CKINVDCx5p33_ASAP7_75t_R g1088 ( .A(n_204), .Y(n_1088) );
XNOR2xp5_ASAP7_75t_L g1320 ( .A(n_205), .B(n_1321), .Y(n_1320) );
INVx1_ASAP7_75t_L g1954 ( .A(n_206), .Y(n_1954) );
AOI22xp33_ASAP7_75t_SL g1084 ( .A1(n_207), .A2(n_372), .B1(n_440), .B2(n_823), .Y(n_1084) );
INVx1_ASAP7_75t_L g1092 ( .A(n_207), .Y(n_1092) );
AOI221xp5_ASAP7_75t_L g1582 ( .A1(n_208), .A2(n_229), .B1(n_1583), .B2(n_1584), .C(n_1585), .Y(n_1582) );
INVx1_ASAP7_75t_L g1618 ( .A(n_208), .Y(n_1618) );
AOI221xp5_ASAP7_75t_L g1679 ( .A1(n_209), .A2(n_373), .B1(n_545), .B2(n_747), .C(n_799), .Y(n_1679) );
OAI22xp33_ASAP7_75t_L g1685 ( .A1(n_209), .A2(n_313), .B1(n_971), .B2(n_973), .Y(n_1685) );
AOI22xp5_ASAP7_75t_L g1748 ( .A1(n_210), .A2(n_244), .B1(n_1694), .B2(n_1702), .Y(n_1748) );
INVx1_ASAP7_75t_L g1741 ( .A(n_212), .Y(n_1741) );
INVx1_ASAP7_75t_L g870 ( .A(n_213), .Y(n_870) );
INVx1_ASAP7_75t_L g937 ( .A(n_214), .Y(n_937) );
INVx1_ASAP7_75t_L g1218 ( .A(n_215), .Y(n_1218) );
CKINVDCx5p33_ASAP7_75t_R g1537 ( .A(n_217), .Y(n_1537) );
INVx1_ASAP7_75t_L g1733 ( .A(n_218), .Y(n_1733) );
INVx1_ASAP7_75t_L g1342 ( .A(n_220), .Y(n_1342) );
INVx1_ASAP7_75t_L g956 ( .A(n_222), .Y(n_956) );
INVx1_ASAP7_75t_L g1113 ( .A(n_223), .Y(n_1113) );
INVx1_ASAP7_75t_L g1152 ( .A(n_224), .Y(n_1152) );
INVx1_ASAP7_75t_L g1404 ( .A(n_225), .Y(n_1404) );
INVxp33_ASAP7_75t_L g841 ( .A(n_227), .Y(n_841) );
INVx1_ASAP7_75t_L g418 ( .A(n_228), .Y(n_418) );
INVx1_ASAP7_75t_L g469 ( .A(n_228), .Y(n_469) );
INVx1_ASAP7_75t_L g1616 ( .A(n_229), .Y(n_1616) );
INVx1_ASAP7_75t_L g2024 ( .A(n_230), .Y(n_2024) );
INVx1_ASAP7_75t_L g1305 ( .A(n_231), .Y(n_1305) );
CKINVDCx5p33_ASAP7_75t_R g677 ( .A(n_232), .Y(n_677) );
INVx1_ASAP7_75t_L g1133 ( .A(n_233), .Y(n_1133) );
AOI22xp33_ASAP7_75t_L g1149 ( .A1(n_233), .A2(n_277), .B1(n_767), .B2(n_895), .Y(n_1149) );
INVxp33_ASAP7_75t_SL g1469 ( .A(n_234), .Y(n_1469) );
CKINVDCx5p33_ASAP7_75t_R g1544 ( .A(n_235), .Y(n_1544) );
XOR2x2_ASAP7_75t_L g1529 ( .A(n_236), .B(n_1530), .Y(n_1529) );
AOI22xp33_ASAP7_75t_L g1080 ( .A1(n_237), .A2(n_350), .B1(n_761), .B2(n_1081), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1099 ( .A1(n_237), .A2(n_517), .B1(n_1100), .B2(n_1101), .C(n_1104), .Y(n_1099) );
INVxp67_ASAP7_75t_SL g1516 ( .A(n_238), .Y(n_1516) );
INVx1_ASAP7_75t_L g1654 ( .A(n_239), .Y(n_1654) );
OAI221xp5_ASAP7_75t_L g1667 ( .A1(n_239), .A2(n_558), .B1(n_952), .B2(n_1668), .C(n_1672), .Y(n_1667) );
INVx1_ASAP7_75t_L g1714 ( .A(n_240), .Y(n_1714) );
INVx1_ASAP7_75t_L g863 ( .A(n_241), .Y(n_863) );
OAI22xp33_ASAP7_75t_L g1018 ( .A1(n_242), .A2(n_339), .B1(n_422), .B2(n_969), .Y(n_1018) );
INVx1_ASAP7_75t_L g1386 ( .A(n_243), .Y(n_1386) );
INVx1_ASAP7_75t_L g1928 ( .A(n_244), .Y(n_1928) );
AOI22xp33_ASAP7_75t_L g1987 ( .A1(n_244), .A2(n_1988), .B1(n_1992), .B2(n_2028), .Y(n_1987) );
INVx1_ASAP7_75t_L g1039 ( .A(n_245), .Y(n_1039) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_246), .Y(n_751) );
OAI221xp5_ASAP7_75t_L g773 ( .A1(n_246), .A2(n_447), .B1(n_460), .B2(n_497), .C(n_774), .Y(n_773) );
CKINVDCx5p33_ASAP7_75t_R g1417 ( .A(n_247), .Y(n_1417) );
OAI22xp5_ASAP7_75t_L g1129 ( .A1(n_248), .A2(n_268), .B1(n_555), .B2(n_1130), .Y(n_1129) );
INVx1_ASAP7_75t_L g1158 ( .A(n_248), .Y(n_1158) );
INVx1_ASAP7_75t_L g993 ( .A(n_249), .Y(n_993) );
INVx1_ASAP7_75t_L g1159 ( .A(n_250), .Y(n_1159) );
CKINVDCx5p33_ASAP7_75t_R g1541 ( .A(n_251), .Y(n_1541) );
CKINVDCx5p33_ASAP7_75t_R g919 ( .A(n_252), .Y(n_919) );
INVx1_ASAP7_75t_L g1958 ( .A(n_253), .Y(n_1958) );
CKINVDCx5p33_ASAP7_75t_R g1381 ( .A(n_254), .Y(n_1381) );
CKINVDCx5p33_ASAP7_75t_R g858 ( .A(n_256), .Y(n_858) );
INVx1_ASAP7_75t_L g1185 ( .A(n_257), .Y(n_1185) );
OAI211xp5_ASAP7_75t_SL g1208 ( .A1(n_257), .A2(n_517), .B(n_1209), .C(n_1217), .Y(n_1208) );
CKINVDCx16_ASAP7_75t_R g780 ( .A(n_258), .Y(n_780) );
INVx1_ASAP7_75t_L g928 ( .A(n_259), .Y(n_928) );
OAI221xp5_ASAP7_75t_L g944 ( .A1(n_259), .A2(n_558), .B1(n_945), .B2(n_948), .C(n_952), .Y(n_944) );
INVx1_ASAP7_75t_L g1293 ( .A(n_260), .Y(n_1293) );
INVx1_ASAP7_75t_L g1301 ( .A(n_261), .Y(n_1301) );
INVx1_ASAP7_75t_L g1229 ( .A(n_262), .Y(n_1229) );
INVx1_ASAP7_75t_L g1184 ( .A(n_263), .Y(n_1184) );
OAI221xp5_ASAP7_75t_L g1196 ( .A1(n_263), .A2(n_558), .B1(n_952), .B2(n_1197), .C(n_1206), .Y(n_1196) );
CKINVDCx5p33_ASAP7_75t_R g1281 ( .A(n_264), .Y(n_1281) );
XNOR2xp5_ASAP7_75t_L g1372 ( .A(n_265), .B(n_1373), .Y(n_1372) );
XNOR2x1_ASAP7_75t_L g1522 ( .A(n_265), .B(n_1373), .Y(n_1522) );
INVx1_ASAP7_75t_L g570 ( .A(n_266), .Y(n_570) );
CKINVDCx5p33_ASAP7_75t_R g923 ( .A(n_267), .Y(n_923) );
INVx1_ASAP7_75t_L g1157 ( .A(n_268), .Y(n_1157) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_270), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g605 ( .A1(n_271), .A2(n_294), .B1(n_606), .B2(n_611), .Y(n_605) );
INVx1_ASAP7_75t_L g688 ( .A(n_271), .Y(n_688) );
INVx1_ASAP7_75t_L g1234 ( .A(n_272), .Y(n_1234) );
AOI21xp33_ASAP7_75t_L g1256 ( .A1(n_272), .A2(n_694), .B(n_1257), .Y(n_1256) );
INVx1_ASAP7_75t_L g873 ( .A(n_273), .Y(n_873) );
AOI21xp33_ASAP7_75t_L g734 ( .A1(n_274), .A2(n_512), .B(n_694), .Y(n_734) );
CKINVDCx5p33_ASAP7_75t_R g1176 ( .A(n_275), .Y(n_1176) );
OAI221xp5_ASAP7_75t_L g1533 ( .A1(n_276), .A2(n_517), .B1(n_1534), .B2(n_1539), .C(n_1543), .Y(n_1533) );
AOI22xp33_ASAP7_75t_SL g1569 ( .A1(n_276), .A2(n_349), .B1(n_485), .B2(n_1568), .Y(n_1569) );
INVx1_ASAP7_75t_L g1134 ( .A(n_277), .Y(n_1134) );
INVx1_ASAP7_75t_L g1609 ( .A(n_278), .Y(n_1609) );
OAI211xp5_ASAP7_75t_L g614 ( .A1(n_279), .A2(n_561), .B(n_615), .C(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g685 ( .A(n_279), .Y(n_685) );
INVx1_ASAP7_75t_L g786 ( .A(n_280), .Y(n_786) );
CKINVDCx5p33_ASAP7_75t_R g1607 ( .A(n_281), .Y(n_1607) );
XNOR2xp5_ASAP7_75t_L g1226 ( .A(n_283), .B(n_1227), .Y(n_1226) );
OAI221xp5_ASAP7_75t_L g1389 ( .A1(n_284), .A2(n_364), .B1(n_1390), .B2(n_1395), .C(n_1397), .Y(n_1389) );
OAI22xp5_ASAP7_75t_L g1430 ( .A1(n_284), .A2(n_364), .B1(n_1431), .B2(n_1434), .Y(n_1430) );
INVx1_ASAP7_75t_L g1128 ( .A(n_285), .Y(n_1128) );
AOI22xp33_ASAP7_75t_SL g1243 ( .A1(n_286), .A2(n_315), .B1(n_831), .B2(n_918), .Y(n_1243) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_286), .A2(n_315), .B1(n_583), .B2(n_588), .Y(n_1248) );
BUFx3_ASAP7_75t_L g414 ( .A(n_287), .Y(n_414) );
INVx1_ASAP7_75t_L g427 ( .A(n_287), .Y(n_427) );
XNOR2xp5_ASAP7_75t_L g1274 ( .A(n_288), .B(n_1275), .Y(n_1274) );
INVx1_ASAP7_75t_L g931 ( .A(n_290), .Y(n_931) );
OAI211xp5_ASAP7_75t_L g953 ( .A1(n_290), .A2(n_517), .B(n_954), .C(n_961), .Y(n_953) );
CKINVDCx5p33_ASAP7_75t_R g1087 ( .A(n_291), .Y(n_1087) );
AO22x2_ASAP7_75t_L g850 ( .A1(n_293), .A2(n_851), .B1(n_904), .B2(n_905), .Y(n_850) );
INVxp67_ASAP7_75t_L g904 ( .A(n_293), .Y(n_904) );
INVx1_ASAP7_75t_L g687 ( .A(n_294), .Y(n_687) );
CKINVDCx5p33_ASAP7_75t_R g1419 ( .A(n_295), .Y(n_1419) );
INVx1_ASAP7_75t_L g1627 ( .A(n_296), .Y(n_1627) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_297), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_297), .B(n_354), .Y(n_511) );
AND2x2_ASAP7_75t_L g521 ( .A(n_297), .B(n_522), .Y(n_521) );
INVx1_ASAP7_75t_L g549 ( .A(n_297), .Y(n_549) );
CKINVDCx5p33_ASAP7_75t_R g1102 ( .A(n_298), .Y(n_1102) );
AOI21xp33_ASAP7_75t_L g742 ( .A1(n_299), .A2(n_743), .B(n_744), .Y(n_742) );
INVx1_ASAP7_75t_L g776 ( .A(n_299), .Y(n_776) );
AO22x2_ASAP7_75t_L g1464 ( .A1(n_300), .A2(n_1465), .B1(n_1466), .B2(n_1519), .Y(n_1464) );
INVxp67_ASAP7_75t_SL g1465 ( .A(n_300), .Y(n_1465) );
OR2x2_ASAP7_75t_L g417 ( .A(n_301), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g456 ( .A(n_301), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g1608 ( .A(n_303), .Y(n_1608) );
INVx1_ASAP7_75t_L g958 ( .A(n_305), .Y(n_958) );
OAI22xp33_ASAP7_75t_L g968 ( .A1(n_305), .A2(n_358), .B1(n_422), .B2(n_969), .Y(n_968) );
CKINVDCx5p33_ASAP7_75t_R g1646 ( .A(n_306), .Y(n_1646) );
INVx1_ASAP7_75t_L g1556 ( .A(n_307), .Y(n_1556) );
CKINVDCx5p33_ASAP7_75t_R g727 ( .A(n_308), .Y(n_727) );
CKINVDCx5p33_ASAP7_75t_R g669 ( .A(n_309), .Y(n_669) );
INVx1_ASAP7_75t_L g1548 ( .A(n_310), .Y(n_1548) );
INVx1_ASAP7_75t_L g941 ( .A(n_311), .Y(n_941) );
INVx1_ASAP7_75t_L g991 ( .A(n_312), .Y(n_991) );
OAI211xp5_ASAP7_75t_L g1008 ( .A1(n_312), .A2(n_517), .B(n_1009), .C(n_1014), .Y(n_1008) );
INVx1_ASAP7_75t_L g1675 ( .A(n_313), .Y(n_1675) );
INVx1_ASAP7_75t_L g420 ( .A(n_314), .Y(n_420) );
INVx1_ASAP7_75t_L g1312 ( .A(n_316), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g736 ( .A(n_317), .Y(n_736) );
INVx1_ASAP7_75t_L g1678 ( .A(n_318), .Y(n_1678) );
OAI22xp33_ASAP7_75t_L g1684 ( .A1(n_318), .A2(n_373), .B1(n_411), .B2(n_422), .Y(n_1684) );
INVxp67_ASAP7_75t_L g1949 ( .A(n_319), .Y(n_1949) );
OAI211xp5_ASAP7_75t_SL g1349 ( .A1(n_320), .A2(n_517), .B(n_1350), .C(n_1355), .Y(n_1349) );
INVx1_ASAP7_75t_L g1658 ( .A(n_322), .Y(n_1658) );
INVx1_ASAP7_75t_L g1036 ( .A(n_323), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1052 ( .A1(n_323), .A2(n_334), .B1(n_811), .B2(n_1053), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g680 ( .A(n_324), .Y(n_680) );
AOI22x1_ASAP7_75t_L g1071 ( .A1(n_326), .A2(n_1072), .B1(n_1073), .B2(n_1114), .Y(n_1071) );
INVxp67_ASAP7_75t_SL g1114 ( .A(n_326), .Y(n_1114) );
INVx1_ASAP7_75t_L g1032 ( .A(n_327), .Y(n_1032) );
AOI22xp5_ASAP7_75t_L g2007 ( .A1(n_328), .A2(n_356), .B1(n_1290), .B2(n_1499), .Y(n_2007) );
OAI22xp5_ASAP7_75t_L g2010 ( .A1(n_328), .A2(n_356), .B1(n_755), .B2(n_756), .Y(n_2010) );
INVx1_ASAP7_75t_L g1286 ( .A(n_331), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g1307 ( .A1(n_331), .A2(n_558), .B1(n_580), .B2(n_1308), .C(n_1309), .Y(n_1307) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_332), .A2(n_367), .B1(n_808), .B2(n_809), .Y(n_807) );
AOI22xp33_ASAP7_75t_L g824 ( .A1(n_332), .A2(n_367), .B1(n_649), .B2(n_825), .Y(n_824) );
CKINVDCx5p33_ASAP7_75t_R g458 ( .A(n_333), .Y(n_458) );
INVx1_ASAP7_75t_L g1035 ( .A(n_334), .Y(n_1035) );
CKINVDCx5p33_ASAP7_75t_R g981 ( .A(n_335), .Y(n_981) );
INVx1_ASAP7_75t_L g879 ( .A(n_336), .Y(n_879) );
INVx1_ASAP7_75t_L g2020 ( .A(n_337), .Y(n_2020) );
INVx1_ASAP7_75t_L g1012 ( .A(n_339), .Y(n_1012) );
INVx1_ASAP7_75t_L g577 ( .A(n_340), .Y(n_577) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_341), .Y(n_982) );
INVx1_ASAP7_75t_L g771 ( .A(n_342), .Y(n_771) );
HB1xp67_ASAP7_75t_L g384 ( .A(n_344), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g1701 ( .A(n_344), .B(n_382), .Y(n_1701) );
AND3x2_ASAP7_75t_L g1709 ( .A(n_344), .B(n_382), .C(n_1698), .Y(n_1709) );
CKINVDCx5p33_ASAP7_75t_R g1664 ( .A(n_345), .Y(n_1664) );
INVx2_ASAP7_75t_L g395 ( .A(n_346), .Y(n_395) );
CKINVDCx5p33_ASAP7_75t_R g921 ( .A(n_347), .Y(n_921) );
INVx1_ASAP7_75t_L g984 ( .A(n_348), .Y(n_984) );
AOI21xp33_ASAP7_75t_L g1006 ( .A1(n_348), .A2(n_694), .B(n_1007), .Y(n_1006) );
OAI221xp5_ASAP7_75t_L g1546 ( .A1(n_349), .A2(n_558), .B1(n_952), .B2(n_1547), .C(n_1552), .Y(n_1546) );
INVx1_ASAP7_75t_L g1098 ( .A(n_350), .Y(n_1098) );
INVx1_ASAP7_75t_L g964 ( .A(n_351), .Y(n_964) );
INVx1_ASAP7_75t_L g501 ( .A(n_352), .Y(n_501) );
INVx1_ASAP7_75t_L g1266 ( .A(n_353), .Y(n_1266) );
INVx1_ASAP7_75t_L g397 ( .A(n_354), .Y(n_397) );
INVx2_ASAP7_75t_L g522 ( .A(n_354), .Y(n_522) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_357), .Y(n_604) );
INVx1_ASAP7_75t_L g750 ( .A(n_359), .Y(n_750) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_359), .Y(n_774) );
OAI211xp5_ASAP7_75t_L g646 ( .A1(n_360), .A2(n_647), .B(n_651), .C(n_659), .Y(n_646) );
INVx1_ASAP7_75t_L g716 ( .A(n_360), .Y(n_716) );
INVx1_ASAP7_75t_L g1681 ( .A(n_362), .Y(n_1681) );
OAI211xp5_ASAP7_75t_SL g516 ( .A1(n_363), .A2(n_517), .B(n_527), .C(n_550), .Y(n_516) );
INVx1_ASAP7_75t_L g1478 ( .A(n_365), .Y(n_1478) );
CKINVDCx5p33_ASAP7_75t_R g1545 ( .A(n_368), .Y(n_1545) );
INVx1_ASAP7_75t_L g1254 ( .A(n_369), .Y(n_1254) );
INVx1_ASAP7_75t_L g2001 ( .A(n_370), .Y(n_2001) );
INVxp33_ASAP7_75t_SL g2015 ( .A(n_371), .Y(n_2015) );
INVx1_ASAP7_75t_L g1093 ( .A(n_372), .Y(n_1093) );
INVx1_ASAP7_75t_L g1205 ( .A(n_374), .Y(n_1205) );
AOI21xp5_ASAP7_75t_L g375 ( .A1(n_376), .A2(n_398), .B(n_1687), .Y(n_375) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx3_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_385), .Y(n_379) );
AND2x4_ASAP7_75t_L g1986 ( .A(n_380), .B(n_386), .Y(n_1986) );
NOR2xp33_ASAP7_75t_SL g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVx1_ASAP7_75t_SL g1991 ( .A(n_381), .Y(n_1991) );
NAND2xp5_ASAP7_75t_L g2030 ( .A(n_381), .B(n_383), .Y(n_2030) );
HB1xp67_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g1990 ( .A(n_383), .B(n_1991), .Y(n_1990) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_387), .B(n_391), .Y(n_386) );
INVxp67_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g601 ( .A(n_388), .B(n_493), .Y(n_601) );
OR2x6_ASAP7_75t_L g783 ( .A(n_388), .B(n_493), .Y(n_783) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g573 ( .A(n_389), .B(n_397), .Y(n_573) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
OR2x2_ASAP7_75t_L g694 ( .A(n_390), .B(n_609), .Y(n_694) );
INVx8_ASAP7_75t_L g603 ( .A(n_391), .Y(n_603) );
OR2x6_ASAP7_75t_L g391 ( .A(n_392), .B(n_396), .Y(n_391) );
BUFx6f_ASAP7_75t_L g569 ( .A(n_392), .Y(n_569) );
OR2x6_ASAP7_75t_L g794 ( .A(n_392), .B(n_608), .Y(n_794) );
INVx1_ASAP7_75t_L g950 ( .A(n_392), .Y(n_950) );
INVx2_ASAP7_75t_SL g1403 ( .A(n_392), .Y(n_1403) );
OR2x2_ASAP7_75t_L g1423 ( .A(n_392), .B(n_1394), .Y(n_1423) );
INVx2_ASAP7_75t_SL g1945 ( .A(n_392), .Y(n_1945) );
BUFx6f_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
AND2x2_ASAP7_75t_L g514 ( .A(n_394), .B(n_395), .Y(n_514) );
INVx1_ASAP7_75t_L g525 ( .A(n_394), .Y(n_525) );
INVx2_ASAP7_75t_L g532 ( .A(n_394), .Y(n_532) );
AND2x4_ASAP7_75t_L g538 ( .A(n_394), .B(n_526), .Y(n_538) );
INVx1_ASAP7_75t_L g565 ( .A(n_394), .Y(n_565) );
INVx2_ASAP7_75t_L g526 ( .A(n_395), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_395), .B(n_532), .Y(n_531) );
INVx1_ASAP7_75t_L g553 ( .A(n_395), .Y(n_553) );
INVx1_ASAP7_75t_L g564 ( .A(n_395), .Y(n_564) );
INVx1_ASAP7_75t_L g587 ( .A(n_395), .Y(n_587) );
AND2x4_ASAP7_75t_L g623 ( .A(n_396), .B(n_553), .Y(n_623) );
INVx2_ASAP7_75t_SL g396 ( .A(n_397), .Y(n_396) );
OR2x2_ASAP7_75t_L g1513 ( .A(n_397), .B(n_626), .Y(n_1513) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_399), .A2(n_400), .B1(n_1162), .B2(n_1163), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
XNOR2xp5_ASAP7_75t_L g400 ( .A(n_401), .B(n_593), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NAND3xp33_ASAP7_75t_L g405 ( .A(n_406), .B(n_500), .C(n_515), .Y(n_405) );
NOR2xp33_ASAP7_75t_L g406 ( .A(n_407), .B(n_443), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_408), .B(n_428), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B1(n_420), .B2(n_421), .Y(n_408) );
OAI221xp5_ASAP7_75t_L g527 ( .A1(n_409), .A2(n_438), .B1(n_528), .B2(n_533), .C(n_539), .Y(n_527) );
AOI22xp5_ASAP7_75t_L g777 ( .A1(n_410), .A2(n_421), .B1(n_738), .B2(n_740), .Y(n_777) );
AOI222xp33_ASAP7_75t_L g1110 ( .A1(n_410), .A2(n_430), .B1(n_503), .B2(n_1102), .C1(n_1105), .C2(n_1111), .Y(n_1110) );
AOI22xp5_ASAP7_75t_L g1150 ( .A1(n_410), .A2(n_421), .B1(n_1151), .B2(n_1152), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1340 ( .A1(n_410), .A2(n_421), .B1(n_1341), .B2(n_1342), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1572 ( .A1(n_410), .A2(n_421), .B1(n_1536), .B2(n_1542), .Y(n_1572) );
CKINVDCx6p67_ASAP7_75t_R g410 ( .A(n_411), .Y(n_410) );
OR2x6_ASAP7_75t_L g411 ( .A(n_412), .B(n_416), .Y(n_411) );
OR2x2_ASAP7_75t_L g969 ( .A(n_412), .B(n_416), .Y(n_969) );
INVx2_ASAP7_75t_L g1145 ( .A(n_412), .Y(n_1145) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx2_ASAP7_75t_L g477 ( .A(n_413), .Y(n_477) );
BUFx6f_ASAP7_75t_L g635 ( .A(n_413), .Y(n_635) );
INVx1_ASAP7_75t_L g768 ( .A(n_413), .Y(n_768) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_413), .Y(n_895) );
AND2x4_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g436 ( .A(n_414), .Y(n_436) );
AND2x2_ASAP7_75t_L g483 ( .A(n_414), .B(n_435), .Y(n_483) );
INVx1_ASAP7_75t_L g425 ( .A(n_415), .Y(n_425) );
OR2x6_ASAP7_75t_L g422 ( .A(n_416), .B(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g437 ( .A(n_416), .Y(n_437) );
OR2x2_ASAP7_75t_L g971 ( .A(n_416), .B(n_972), .Y(n_971) );
OR2x2_ASAP7_75t_L g973 ( .A(n_416), .B(n_974), .Y(n_973) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVx2_ASAP7_75t_L g1429 ( .A(n_417), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1459 ( .A(n_417), .B(n_641), .Y(n_1459) );
OR2x2_ASAP7_75t_L g1461 ( .A(n_417), .B(n_477), .Y(n_1461) );
INVx1_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
INVx1_ASAP7_75t_L g457 ( .A(n_419), .Y(n_457) );
AND2x4_ASAP7_75t_L g1380 ( .A(n_419), .B(n_521), .Y(n_1380) );
AOI22xp5_ASAP7_75t_L g1112 ( .A1(n_421), .A2(n_439), .B1(n_1103), .B2(n_1113), .Y(n_1112) );
CKINVDCx6p67_ASAP7_75t_R g421 ( .A(n_422), .Y(n_421) );
BUFx3_ASAP7_75t_L g684 ( .A(n_423), .Y(n_684) );
OAI221xp5_ASAP7_75t_L g1280 ( .A1(n_423), .A2(n_1173), .B1(n_1281), .B2(n_1282), .C(n_1283), .Y(n_1280) );
OAI22xp33_ASAP7_75t_L g1653 ( .A1(n_423), .A2(n_1174), .B1(n_1654), .B2(n_1655), .Y(n_1653) );
INVx2_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g682 ( .A(n_424), .Y(n_682) );
BUFx2_ASAP7_75t_L g925 ( .A(n_424), .Y(n_925) );
BUFx4f_ASAP7_75t_L g930 ( .A(n_424), .Y(n_930) );
INVx1_ASAP7_75t_L g1030 ( .A(n_424), .Y(n_1030) );
INVx1_ASAP7_75t_L g1971 ( .A(n_424), .Y(n_1971) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_426), .Y(n_424) );
OR2x2_ASAP7_75t_L g641 ( .A(n_425), .B(n_426), .Y(n_641) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
AND2x4_ASAP7_75t_L g442 ( .A(n_427), .B(n_435), .Y(n_442) );
AOI22xp33_ASAP7_75t_L g428 ( .A1(n_429), .A2(n_430), .B1(n_438), .B2(n_439), .Y(n_428) );
AOI222xp33_ASAP7_75t_L g775 ( .A1(n_430), .A2(n_439), .B1(n_503), .B2(n_736), .C1(n_746), .C2(n_776), .Y(n_775) );
AOI22xp5_ASAP7_75t_L g1153 ( .A1(n_430), .A2(n_439), .B1(n_1154), .B2(n_1155), .Y(n_1153) );
AOI22xp33_ASAP7_75t_L g1343 ( .A1(n_430), .A2(n_439), .B1(n_1344), .B2(n_1345), .Y(n_1343) );
AOI22xp33_ASAP7_75t_L g1573 ( .A1(n_430), .A2(n_439), .B1(n_1537), .B2(n_1541), .Y(n_1573) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_437), .Y(n_430) );
BUFx2_ASAP7_75t_L g1503 ( .A(n_431), .Y(n_1503) );
INVx2_ASAP7_75t_SL g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g1333 ( .A(n_432), .Y(n_1333) );
INVx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx2_ASAP7_75t_L g479 ( .A(n_433), .Y(n_479) );
INVx6_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
AND2x2_ASAP7_75t_L g504 ( .A(n_433), .B(n_453), .Y(n_504) );
AND2x4_ASAP7_75t_L g643 ( .A(n_433), .B(n_644), .Y(n_643) );
AND2x4_ASAP7_75t_L g433 ( .A(n_434), .B(n_436), .Y(n_433) );
INVx1_ASAP7_75t_L g463 ( .A(n_434), .Y(n_463) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g450 ( .A(n_436), .Y(n_450) );
AND2x2_ASAP7_75t_L g439 ( .A(n_437), .B(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
OAI22xp5_ASAP7_75t_L g686 ( .A1(n_441), .A2(n_687), .B1(n_688), .B2(n_689), .Y(n_686) );
INVx1_ASAP7_75t_L g1077 ( .A(n_441), .Y(n_1077) );
INVx2_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
BUFx2_ASAP7_75t_L g473 ( .A(n_442), .Y(n_473) );
BUFx6f_ASAP7_75t_L g490 ( .A(n_442), .Y(n_490) );
BUFx6f_ASAP7_75t_L g652 ( .A(n_442), .Y(n_652) );
BUFx6f_ASAP7_75t_L g767 ( .A(n_442), .Y(n_767) );
BUFx2_ASAP7_75t_L g822 ( .A(n_442), .Y(n_822) );
AND2x6_ASAP7_75t_L g845 ( .A(n_442), .B(n_639), .Y(n_845) );
BUFx3_ASAP7_75t_L g918 ( .A(n_442), .Y(n_918) );
BUFx6f_ASAP7_75t_L g1189 ( .A(n_442), .Y(n_1189) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_444), .B(n_464), .C(n_495), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_446), .B1(n_458), .B2(n_459), .Y(n_444) );
AOI22xp33_ASAP7_75t_L g550 ( .A1(n_445), .A2(n_458), .B1(n_551), .B2(n_554), .Y(n_550) );
INVx1_ASAP7_75t_L g1278 ( .A(n_446), .Y(n_1278) );
AOI22xp33_ASAP7_75t_L g1324 ( .A1(n_446), .A2(n_459), .B1(n_1325), .B2(n_1326), .Y(n_1324) );
INVx1_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g1086 ( .A(n_447), .Y(n_1086) );
HB1xp67_ASAP7_75t_L g1191 ( .A(n_447), .Y(n_1191) );
INVx1_ASAP7_75t_L g1562 ( .A(n_447), .Y(n_1562) );
NAND2x1p5_ASAP7_75t_L g447 ( .A(n_448), .B(n_451), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g1433 ( .A(n_449), .Y(n_1433) );
INVx1_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx1_ASAP7_75t_L g657 ( .A(n_450), .Y(n_657) );
INVx2_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
OR2x6_ASAP7_75t_L g460 ( .A(n_452), .B(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g499 ( .A(n_452), .Y(n_499) );
OR2x2_ASAP7_75t_L g1246 ( .A(n_452), .B(n_461), .Y(n_1246) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_453), .B(n_457), .Y(n_452) );
AND2x4_ASAP7_75t_L g1432 ( .A(n_453), .B(n_1433), .Y(n_1432) );
INVx1_ASAP7_75t_L g1435 ( .A(n_453), .Y(n_1435) );
AND2x2_ASAP7_75t_L g1594 ( .A(n_453), .B(n_462), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1965 ( .A(n_453), .B(n_462), .Y(n_1965) );
AND2x4_ASAP7_75t_L g453 ( .A(n_454), .B(n_455), .Y(n_453) );
AND2x4_ASAP7_75t_L g494 ( .A(n_455), .B(n_469), .Y(n_494) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AND2x2_ASAP7_75t_L g468 ( .A(n_456), .B(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g634 ( .A(n_456), .Y(n_634) );
INVx1_ASAP7_75t_L g640 ( .A(n_456), .Y(n_640) );
HB1xp67_ASAP7_75t_L g645 ( .A(n_456), .Y(n_645) );
OR2x6_ASAP7_75t_L g719 ( .A(n_457), .B(n_547), .Y(n_719) );
AOI221xp5_ASAP7_75t_L g1085 ( .A1(n_459), .A2(n_912), .B1(n_1086), .B2(n_1087), .C(n_1088), .Y(n_1085) );
AOI221xp5_ASAP7_75t_L g1156 ( .A1(n_459), .A2(n_912), .B1(n_1086), .B2(n_1157), .C(n_1158), .Y(n_1156) );
AOI22xp5_ASAP7_75t_L g1561 ( .A1(n_459), .A2(n_1544), .B1(n_1545), .B2(n_1562), .Y(n_1561) );
INVx2_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
OR2x2_ASAP7_75t_L g1434 ( .A(n_461), .B(n_1435), .Y(n_1434) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x6_ASAP7_75t_L g658 ( .A(n_463), .B(n_640), .Y(n_658) );
AOI33xp33_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_472), .A3(n_478), .B1(n_484), .B2(n_488), .B3(n_492), .Y(n_464) );
AOI221xp5_ASAP7_75t_L g759 ( .A1(n_465), .A2(n_691), .B1(n_760), .B2(n_769), .C(n_773), .Y(n_759) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_SL g1171 ( .A1(n_466), .A2(n_690), .B1(n_1172), .B2(n_1183), .Y(n_1171) );
OAI22xp5_ASAP7_75t_SL g1279 ( .A1(n_466), .A2(n_1238), .B1(n_1280), .B2(n_1285), .Y(n_1279) );
CKINVDCx5p33_ASAP7_75t_R g1328 ( .A(n_466), .Y(n_1328) );
CKINVDCx5p33_ASAP7_75t_R g1564 ( .A(n_466), .Y(n_1564) );
OAI22xp5_ASAP7_75t_SL g1999 ( .A1(n_466), .A2(n_1238), .B1(n_2000), .B2(n_2004), .Y(n_1999) );
OR2x6_ASAP7_75t_L g466 ( .A(n_467), .B(n_470), .Y(n_466) );
OR2x2_ASAP7_75t_L g667 ( .A(n_467), .B(n_470), .Y(n_667) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g899 ( .A(n_468), .Y(n_899) );
INVx2_ASAP7_75t_SL g1451 ( .A(n_468), .Y(n_1451) );
BUFx3_ASAP7_75t_L g1979 ( .A(n_468), .Y(n_1979) );
INVx1_ASAP7_75t_L g663 ( .A(n_469), .Y(n_663) );
INVx2_ASAP7_75t_L g506 ( .A(n_470), .Y(n_506) );
BUFx2_ASAP7_75t_L g592 ( .A(n_470), .Y(n_592) );
AND2x4_ASAP7_75t_L g806 ( .A(n_470), .B(n_573), .Y(n_806) );
OR2x2_ASAP7_75t_L g898 ( .A(n_470), .B(n_899), .Y(n_898) );
AND2x4_ASAP7_75t_L g1486 ( .A(n_470), .B(n_573), .Y(n_1486) );
OAI31xp33_ASAP7_75t_L g1531 ( .A1(n_470), .A2(n_1532), .A3(n_1533), .B(n_1546), .Y(n_1531) );
INVx2_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
BUFx2_ASAP7_75t_L g664 ( .A(n_471), .Y(n_664) );
OR2x6_ASAP7_75t_L g693 ( .A(n_471), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g491 ( .A(n_475), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g770 ( .A1(n_475), .A2(n_672), .B1(n_771), .B2(n_772), .Y(n_770) );
INVx2_ASAP7_75t_SL g1566 ( .A(n_475), .Y(n_1566) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
BUFx2_ASAP7_75t_L g1589 ( .A(n_476), .Y(n_1589) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g675 ( .A(n_477), .Y(n_675) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g1334 ( .A(n_481), .Y(n_1334) );
INVx1_ASAP7_75t_L g1568 ( .A(n_481), .Y(n_1568) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_482), .Y(n_498) );
INVx1_ASAP7_75t_L g829 ( .A(n_482), .Y(n_829) );
BUFx4f_ASAP7_75t_L g1079 ( .A(n_482), .Y(n_1079) );
BUFx3_ASAP7_75t_L g1336 ( .A(n_482), .Y(n_1336) );
AND2x4_ASAP7_75t_L g1447 ( .A(n_482), .B(n_1429), .Y(n_1447) );
INVx1_ASAP7_75t_L g1450 ( .A(n_482), .Y(n_1450) );
BUFx6f_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx6f_ASAP7_75t_L g650 ( .A(n_483), .Y(n_650) );
INVx4_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g1584 ( .A(n_486), .Y(n_1584) );
BUFx6f_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_487), .Y(n_764) );
INVx2_ASAP7_75t_L g826 ( .A(n_487), .Y(n_826) );
INVx2_ASAP7_75t_L g843 ( .A(n_487), .Y(n_843) );
INVx1_ASAP7_75t_L g902 ( .A(n_487), .Y(n_902) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_487), .Y(n_1083) );
BUFx4f_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g974 ( .A(n_490), .Y(n_974) );
BUFx2_ASAP7_75t_L g1180 ( .A(n_490), .Y(n_1180) );
AOI33xp33_ASAP7_75t_L g819 ( .A1(n_492), .A2(n_820), .A3(n_821), .B1(n_824), .B2(n_827), .B3(n_830), .Y(n_819) );
NAND3xp33_ASAP7_75t_L g900 ( .A(n_492), .B(n_901), .C(n_903), .Y(n_900) );
INVx1_ASAP7_75t_L g938 ( .A(n_492), .Y(n_938) );
INVx1_ASAP7_75t_L g1068 ( .A(n_492), .Y(n_1068) );
AOI33xp33_ASAP7_75t_L g1075 ( .A1(n_492), .A2(n_820), .A3(n_1076), .B1(n_1078), .B2(n_1080), .B3(n_1084), .Y(n_1075) );
AOI33xp33_ASAP7_75t_L g1143 ( .A1(n_492), .A2(n_897), .A3(n_1144), .B1(n_1146), .B2(n_1148), .B3(n_1149), .Y(n_1143) );
AND2x4_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
AND2x4_ASAP7_75t_L g503 ( .A(n_493), .B(n_504), .Y(n_503) );
AND2x4_ASAP7_75t_L g691 ( .A(n_493), .B(n_494), .Y(n_691) );
INVx2_ASAP7_75t_L g1443 ( .A(n_494), .Y(n_1443) );
INVx2_ASAP7_75t_SL g1974 ( .A(n_494), .Y(n_1974) );
NAND3xp33_ASAP7_75t_SL g1560 ( .A(n_495), .B(n_1561), .C(n_1563), .Y(n_1560) );
INVx1_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
NAND3xp33_ASAP7_75t_SL g1323 ( .A(n_497), .B(n_1324), .C(n_1327), .Y(n_1323) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_498), .B(n_499), .Y(n_497) );
INVx1_ASAP7_75t_L g1507 ( .A(n_498), .Y(n_1507) );
AND2x2_ASAP7_75t_L g912 ( .A(n_499), .B(n_913), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_501), .B(n_502), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_502), .B(n_941), .Y(n_940) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_502), .B(n_997), .Y(n_996) );
INVx1_ASAP7_75t_L g1119 ( .A(n_502), .Y(n_1119) );
NAND2xp5_ASAP7_75t_L g1192 ( .A(n_502), .B(n_1193), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1228 ( .A(n_502), .B(n_1229), .Y(n_1228) );
NAND2xp5_ASAP7_75t_L g1292 ( .A(n_502), .B(n_1293), .Y(n_1292) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_502), .B(n_1347), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1557 ( .A(n_502), .B(n_1558), .Y(n_1557) );
NAND2xp5_ASAP7_75t_L g1663 ( .A(n_502), .B(n_1664), .Y(n_1663) );
NAND2xp5_ASAP7_75t_L g1996 ( .A(n_502), .B(n_1997), .Y(n_1996) );
OR2x6_ASAP7_75t_L g502 ( .A(n_503), .B(n_505), .Y(n_502) );
INVx2_ASAP7_75t_L g1424 ( .A(n_503), .Y(n_1424) );
NOR2xp67_ASAP7_75t_L g505 ( .A(n_506), .B(n_507), .Y(n_505) );
INVx2_ASAP7_75t_L g758 ( .A(n_506), .Y(n_758) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .Y(n_507) );
AND2x2_ASAP7_75t_L g551 ( .A(n_508), .B(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g963 ( .A(n_508), .B(n_552), .Y(n_963) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
OR2x6_ASAP7_75t_L g555 ( .A(n_509), .B(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g580 ( .A(n_509), .B(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g753 ( .A(n_509), .Y(n_753) );
OR2x6_ASAP7_75t_L g952 ( .A(n_509), .B(n_581), .Y(n_952) );
INVx1_ASAP7_75t_L g1131 ( .A(n_509), .Y(n_1131) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
BUFx2_ASAP7_75t_L g808 ( .A(n_512), .Y(n_808) );
INVx2_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g743 ( .A(n_513), .Y(n_743) );
INVx2_ASAP7_75t_SL g1257 ( .A(n_513), .Y(n_1257) );
INVx3_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_514), .Y(n_544) );
OAI31xp33_ASAP7_75t_L g515 ( .A1(n_516), .A2(n_557), .A3(n_582), .B(n_590), .Y(n_515) );
INVx8_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AOI221xp5_ASAP7_75t_SL g1121 ( .A1(n_518), .A2(n_1122), .B1(n_1125), .B2(n_1128), .C(n_1129), .Y(n_1121) );
AND2x4_ASAP7_75t_L g518 ( .A(n_519), .B(n_523), .Y(n_518) );
AND2x4_ASAP7_75t_L g589 ( .A(n_519), .B(n_536), .Y(n_589) );
INVx1_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
AND2x4_ASAP7_75t_L g559 ( .A(n_521), .B(n_544), .Y(n_559) );
AND2x2_ASAP7_75t_L g584 ( .A(n_521), .B(n_585), .Y(n_584) );
INVx1_ASAP7_75t_L g548 ( .A(n_522), .Y(n_548) );
INVx1_ASAP7_75t_L g609 ( .A(n_522), .Y(n_609) );
INVx1_ASAP7_75t_L g541 ( .A(n_523), .Y(n_541) );
BUFx3_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
AND2x4_ASAP7_75t_L g616 ( .A(n_524), .B(n_617), .Y(n_616) );
BUFx6f_ASAP7_75t_L g799 ( .A(n_524), .Y(n_799) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_524), .Y(n_818) );
BUFx2_ASAP7_75t_L g877 ( .A(n_524), .Y(n_877) );
BUFx3_ASAP7_75t_L g960 ( .A(n_524), .Y(n_960) );
AND2x4_ASAP7_75t_L g524 ( .A(n_525), .B(n_526), .Y(n_524) );
BUFx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g576 ( .A(n_530), .Y(n_576) );
INVx1_ASAP7_75t_L g955 ( .A(n_530), .Y(n_955) );
HB1xp67_ASAP7_75t_L g1670 ( .A(n_530), .Y(n_1670) );
INVx1_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
BUFx2_ASAP7_75t_L g610 ( .A(n_531), .Y(n_610) );
INVx1_ASAP7_75t_L g704 ( .A(n_531), .Y(n_704) );
INVx1_ASAP7_75t_L g556 ( .A(n_532), .Y(n_556) );
AND2x4_ASAP7_75t_L g585 ( .A(n_532), .B(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_535), .A2(n_669), .B1(n_673), .B2(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g1300 ( .A(n_535), .Y(n_1300) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g1139 ( .A(n_537), .Y(n_1139) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g579 ( .A(n_538), .Y(n_579) );
INVx3_ASAP7_75t_L g708 ( .A(n_538), .Y(n_708) );
BUFx6f_ASAP7_75t_L g947 ( .A(n_538), .Y(n_947) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g1127 ( .A(n_541), .Y(n_1127) );
A2O1A1Ixp33_ASAP7_75t_L g1104 ( .A1(n_542), .A2(n_753), .B(n_1105), .C(n_1106), .Y(n_1104) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx2_ASAP7_75t_L g620 ( .A(n_543), .Y(n_620) );
INVx2_ASAP7_75t_SL g1007 ( .A(n_543), .Y(n_1007) );
INVx3_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
BUFx6f_ASAP7_75t_L g747 ( .A(n_544), .Y(n_747) );
BUFx2_ASAP7_75t_L g1126 ( .A(n_544), .Y(n_1126) );
INVx1_ASAP7_75t_L g1538 ( .A(n_545), .Y(n_1538) );
INVx2_ASAP7_75t_SL g545 ( .A(n_546), .Y(n_545) );
INVx1_ASAP7_75t_L g1303 ( .A(n_546), .Y(n_1303) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
BUFx2_ASAP7_75t_L g744 ( .A(n_547), .Y(n_744) );
NAND2x1p5_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
INVx1_ASAP7_75t_L g618 ( .A(n_548), .Y(n_618) );
AOI22xp33_ASAP7_75t_L g1217 ( .A1(n_551), .A2(n_554), .B1(n_1218), .B2(n_1219), .Y(n_1217) );
AOI22xp33_ASAP7_75t_L g1264 ( .A1(n_551), .A2(n_554), .B1(n_1265), .B2(n_1266), .Y(n_1264) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_551), .A2(n_554), .B1(n_1544), .B2(n_1545), .Y(n_1543) );
AOI22xp33_ASAP7_75t_L g1680 ( .A1(n_551), .A2(n_554), .B1(n_1681), .B2(n_1682), .Y(n_1680) );
AOI22xp33_ASAP7_75t_L g2022 ( .A1(n_551), .A2(n_554), .B1(n_2023), .B2(n_2024), .Y(n_2022) );
HB1xp67_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AOI22xp5_ASAP7_75t_L g749 ( .A1(n_553), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_749) );
INVx1_ASAP7_75t_L g1109 ( .A(n_553), .Y(n_1109) );
AOI22xp33_ASAP7_75t_L g961 ( .A1(n_554), .A2(n_962), .B1(n_963), .B2(n_964), .Y(n_961) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_554), .A2(n_963), .B1(n_1015), .B2(n_1016), .Y(n_1014) );
AOI22xp33_ASAP7_75t_L g1304 ( .A1(n_554), .A2(n_963), .B1(n_1305), .B2(n_1306), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_554), .A2(n_963), .B1(n_1325), .B2(n_1326), .Y(n_1355) );
CKINVDCx11_ASAP7_75t_R g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_L g752 ( .A(n_556), .Y(n_752) );
CKINVDCx6p67_ASAP7_75t_R g558 ( .A(n_559), .Y(n_558) );
AOI22xp5_ASAP7_75t_L g1094 ( .A1(n_559), .A2(n_1095), .B1(n_1097), .B2(n_1098), .Y(n_1094) );
AOI221xp5_ASAP7_75t_L g1135 ( .A1(n_559), .A2(n_1136), .B1(n_1137), .B2(n_1138), .C(n_1140), .Y(n_1135) );
OAI221xp5_ASAP7_75t_L g560 ( .A1(n_561), .A2(n_566), .B1(n_567), .B2(n_570), .C(n_571), .Y(n_560) );
OAI221xp5_ASAP7_75t_L g1308 ( .A1(n_561), .A2(n_951), .B1(n_1207), .B2(n_1281), .C(n_1282), .Y(n_1308) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
INVx1_ASAP7_75t_L g2013 ( .A(n_562), .Y(n_2013) );
BUFx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g581 ( .A(n_563), .Y(n_581) );
INVx3_ASAP7_75t_L g733 ( .A(n_563), .Y(n_733) );
INVx2_ASAP7_75t_L g741 ( .A(n_563), .Y(n_741) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g715 ( .A(n_564), .B(n_565), .Y(n_715) );
INVx1_ASAP7_75t_L g626 ( .A(n_565), .Y(n_626) );
OAI221xp5_ASAP7_75t_L g1534 ( .A1(n_567), .A2(n_1535), .B1(n_1536), .B2(n_1537), .C(n_1538), .Y(n_1534) );
OAI221xp5_ASAP7_75t_L g2012 ( .A1(n_567), .A2(n_571), .B1(n_2001), .B2(n_2002), .C(n_2013), .Y(n_2012) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
OAI22xp33_ASAP7_75t_L g695 ( .A1(n_569), .A2(n_677), .B1(n_680), .B2(n_696), .Y(n_695) );
OAI22xp33_ASAP7_75t_L g710 ( .A1(n_569), .A2(n_711), .B1(n_712), .B2(n_716), .Y(n_710) );
BUFx2_ASAP7_75t_L g1207 ( .A(n_569), .Y(n_1207) );
INVx1_ASAP7_75t_L g1555 ( .A(n_569), .Y(n_1555) );
OAI221xp5_ASAP7_75t_L g1672 ( .A1(n_569), .A2(n_571), .B1(n_714), .B2(n_1650), .C(n_1652), .Y(n_1672) );
OAI221xp5_ASAP7_75t_L g1206 ( .A1(n_571), .A2(n_741), .B1(n_1176), .B2(n_1177), .C(n_1207), .Y(n_1206) );
OAI221xp5_ASAP7_75t_L g1552 ( .A1(n_571), .A2(n_696), .B1(n_1553), .B2(n_1554), .C(n_1556), .Y(n_1552) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx2_ASAP7_75t_SL g951 ( .A(n_573), .Y(n_951) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_576), .B1(n_577), .B2(n_578), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g726 ( .A1(n_576), .A2(n_727), .B1(n_728), .B2(n_730), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g735 ( .A1(n_576), .A2(n_736), .B1(n_737), .B2(n_738), .Y(n_735) );
OAI22xp5_ASAP7_75t_L g1101 ( .A1(n_576), .A2(n_737), .B1(n_1102), .B2(n_1103), .Y(n_1101) );
BUFx2_ASAP7_75t_L g1540 ( .A(n_576), .Y(n_1540) );
OAI22xp5_ASAP7_75t_L g2014 ( .A1(n_576), .A2(n_946), .B1(n_2015), .B2(n_2016), .Y(n_2014) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g613 ( .A(n_579), .Y(n_613) );
INVx1_ASAP7_75t_L g697 ( .A(n_581), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_581), .B(n_749), .Y(n_748) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx3_ASAP7_75t_L g755 ( .A(n_584), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g1091 ( .A1(n_584), .A2(n_589), .B1(n_1092), .B2(n_1093), .Y(n_1091) );
AOI22xp33_ASAP7_75t_L g1132 ( .A1(n_584), .A2(n_589), .B1(n_1133), .B2(n_1134), .Y(n_1132) );
AND2x4_ASAP7_75t_L g787 ( .A(n_585), .B(n_608), .Y(n_787) );
INVx1_ASAP7_75t_L g812 ( .A(n_585), .Y(n_812) );
BUFx2_ASAP7_75t_L g1057 ( .A(n_585), .Y(n_1057) );
BUFx6f_ASAP7_75t_L g1096 ( .A(n_585), .Y(n_1096) );
BUFx6f_ASAP7_75t_L g1123 ( .A(n_585), .Y(n_1123) );
BUFx6f_ASAP7_75t_L g1388 ( .A(n_585), .Y(n_1388) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g588 ( .A(n_589), .Y(n_588) );
INVx3_ASAP7_75t_L g756 ( .A(n_589), .Y(n_756) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
CKINVDCx8_ASAP7_75t_R g591 ( .A(n_592), .Y(n_591) );
OAI31xp33_ASAP7_75t_SL g1194 ( .A1(n_592), .A2(n_1195), .A3(n_1196), .B(n_1208), .Y(n_1194) );
OAI31xp33_ASAP7_75t_L g1294 ( .A1(n_592), .A2(n_1295), .A3(n_1307), .B(n_1316), .Y(n_1294) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
OAI21x1_ASAP7_75t_L g594 ( .A1(n_595), .A2(n_1115), .B(n_1160), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
OR2x2_ASAP7_75t_L g1160 ( .A(n_596), .B(n_1161), .Y(n_1160) );
XNOR2xp5_ASAP7_75t_L g596 ( .A(n_597), .B(n_907), .Y(n_596) );
XNOR2x1_ASAP7_75t_L g597 ( .A(n_598), .B(n_778), .Y(n_597) );
XNOR2x1_ASAP7_75t_L g598 ( .A(n_599), .B(n_722), .Y(n_598) );
INVx1_ASAP7_75t_L g720 ( .A(n_600), .Y(n_720) );
OAI211xp5_ASAP7_75t_L g600 ( .A1(n_601), .A2(n_602), .B(n_629), .C(n_665), .Y(n_600) );
AOI31xp33_ASAP7_75t_L g1509 ( .A1(n_601), .A2(n_1510), .A3(n_1514), .B(n_1517), .Y(n_1509) );
AOI211xp5_ASAP7_75t_L g602 ( .A1(n_603), .A2(n_604), .B(n_605), .C(n_614), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g790 ( .A1(n_603), .A2(n_791), .B1(n_792), .B2(n_793), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g878 ( .A1(n_603), .A2(n_793), .B1(n_858), .B2(n_879), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_603), .A2(n_1033), .B1(n_1046), .B2(n_1047), .Y(n_1045) );
AOI22xp33_ASAP7_75t_SL g1517 ( .A1(n_603), .A2(n_1047), .B1(n_1472), .B2(n_1518), .Y(n_1517) );
OAI22xp33_ASAP7_75t_L g683 ( .A1(n_604), .A2(n_678), .B1(n_684), .B2(n_685), .Y(n_683) );
OR2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_610), .Y(n_606) );
AOI322xp5_ASAP7_75t_L g619 ( .A1(n_607), .A2(n_620), .A3(n_621), .B1(n_622), .B2(n_623), .C1(n_624), .C2(n_628), .Y(n_619) );
INVx1_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
AND2x4_ASAP7_75t_L g612 ( .A(n_608), .B(n_613), .Y(n_612) );
AND2x4_ASAP7_75t_L g789 ( .A(n_608), .B(n_613), .Y(n_789) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g700 ( .A(n_610), .Y(n_700) );
BUFx2_ASAP7_75t_L g1410 ( .A(n_610), .Y(n_1410) );
INVx5_ASAP7_75t_SL g611 ( .A(n_612), .Y(n_611) );
NAND4xp25_ASAP7_75t_SL g784 ( .A(n_615), .B(n_785), .C(n_790), .D(n_795), .Y(n_784) );
NAND4xp25_ASAP7_75t_SL g867 ( .A(n_615), .B(n_868), .C(n_871), .D(n_878), .Y(n_867) );
NAND4xp25_ASAP7_75t_SL g1037 ( .A(n_615), .B(n_1038), .C(n_1041), .D(n_1045), .Y(n_1037) );
CKINVDCx11_ASAP7_75t_R g615 ( .A(n_616), .Y(n_615) );
AOI211xp5_ASAP7_75t_L g1510 ( .A1(n_616), .A2(n_1127), .B(n_1511), .C(n_1512), .Y(n_1510) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
INVxp67_ASAP7_75t_L g627 ( .A(n_618), .Y(n_627) );
AOI322xp5_ASAP7_75t_L g651 ( .A1(n_622), .A2(n_628), .A3(n_652), .B1(n_653), .B2(n_654), .C1(n_655), .C2(n_658), .Y(n_651) );
INVx2_ASAP7_75t_L g802 ( .A(n_623), .Y(n_802) );
AOI222xp33_ASAP7_75t_L g871 ( .A1(n_623), .A2(n_624), .B1(n_872), .B2(n_873), .C1(n_874), .C2(n_875), .Y(n_871) );
AOI222xp33_ASAP7_75t_L g795 ( .A1(n_624), .A2(n_796), .B1(n_797), .B2(n_800), .C1(n_801), .C2(n_803), .Y(n_795) );
AOI222xp33_ASAP7_75t_L g1041 ( .A1(n_624), .A2(n_797), .B1(n_801), .B2(n_1042), .C1(n_1043), .C2(n_1044), .Y(n_1041) );
AND2x4_ASAP7_75t_L g624 ( .A(n_625), .B(n_627), .Y(n_624) );
AOI22xp5_ASAP7_75t_L g1107 ( .A1(n_625), .A2(n_1087), .B1(n_1088), .B2(n_1108), .Y(n_1107) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
OAI31xp33_ASAP7_75t_SL g629 ( .A1(n_630), .A2(n_636), .A3(n_646), .B(n_662), .Y(n_629) );
INVx4_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_632), .A2(n_845), .B1(n_846), .B2(n_847), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_632), .A2(n_854), .B1(n_855), .B2(n_856), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1034 ( .A1(n_632), .A2(n_845), .B1(n_1035), .B2(n_1036), .Y(n_1034) );
AOI22xp33_ASAP7_75t_L g1471 ( .A1(n_632), .A2(n_643), .B1(n_1472), .B2(n_1473), .Y(n_1471) );
AND2x6_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
AND2x4_ASAP7_75t_L g842 ( .A(n_633), .B(n_843), .Y(n_842) );
AND2x4_ASAP7_75t_L g854 ( .A(n_633), .B(n_843), .Y(n_854) );
INVx1_ASAP7_75t_SL g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g837 ( .A(n_634), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g689 ( .A(n_635), .Y(n_689) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_635), .Y(n_823) );
BUFx6f_ASAP7_75t_L g831 ( .A(n_635), .Y(n_831) );
BUFx6f_ASAP7_75t_L g936 ( .A(n_635), .Y(n_936) );
INVx2_ASAP7_75t_L g1291 ( .A(n_635), .Y(n_1291) );
INVx1_ASAP7_75t_L g1501 ( .A(n_635), .Y(n_1501) );
OR2x2_ASAP7_75t_L g637 ( .A(n_638), .B(n_641), .Y(n_637) );
INVx1_ASAP7_75t_L g653 ( .A(n_638), .Y(n_653) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g648 ( .A(n_639), .B(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g661 ( .A(n_639), .Y(n_661) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g679 ( .A(n_641), .Y(n_679) );
INVx1_ASAP7_75t_L g1175 ( .A(n_641), .Y(n_1175) );
BUFx2_ASAP7_75t_L g1233 ( .A(n_641), .Y(n_1233) );
INVx4_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_643), .A2(n_792), .B1(n_841), .B2(n_842), .Y(n_840) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_643), .A2(n_845), .B1(n_858), .B2(n_859), .C(n_860), .Y(n_857) );
AOI22xp33_ASAP7_75t_L g1031 ( .A1(n_643), .A2(n_854), .B1(n_1032), .B2(n_1033), .Y(n_1031) );
AND2x2_ASAP7_75t_SL g655 ( .A(n_644), .B(n_656), .Y(n_655) );
AND2x4_ASAP7_75t_L g1477 ( .A(n_644), .B(n_656), .Y(n_1477) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
AOI211xp5_ASAP7_75t_L g833 ( .A1(n_648), .A2(n_660), .B(n_834), .C(n_835), .Y(n_833) );
HB1xp67_ASAP7_75t_L g1504 ( .A(n_649), .Y(n_1504) );
BUFx6f_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x4_ASAP7_75t_L g660 ( .A(n_650), .B(n_661), .Y(n_660) );
INVx2_ASAP7_75t_L g762 ( .A(n_650), .Y(n_762) );
BUFx6f_ASAP7_75t_L g864 ( .A(n_650), .Y(n_864) );
INVx1_ASAP7_75t_L g914 ( .A(n_650), .Y(n_914) );
INVx2_ASAP7_75t_L g672 ( .A(n_652), .Y(n_672) );
INVx1_ASAP7_75t_L g933 ( .A(n_652), .Y(n_933) );
INVx2_ASAP7_75t_SL g980 ( .A(n_652), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g701 ( .A1(n_654), .A2(n_702), .B1(n_705), .B2(n_709), .Y(n_701) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g838 ( .A(n_657), .Y(n_838) );
INVx3_ASAP7_75t_L g839 ( .A(n_658), .Y(n_839) );
AOI222xp33_ASAP7_75t_L g1474 ( .A1(n_658), .A2(n_1336), .B1(n_1475), .B2(n_1476), .C1(n_1477), .C2(n_1478), .Y(n_1474) );
CKINVDCx8_ASAP7_75t_R g659 ( .A(n_660), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g1026 ( .A(n_660), .B(n_1027), .Y(n_1026) );
INVx5_ASAP7_75t_L g1479 ( .A(n_660), .Y(n_1479) );
OAI21xp33_ASAP7_75t_L g862 ( .A1(n_661), .A2(n_863), .B(n_864), .Y(n_862) );
INVx1_ASAP7_75t_SL g848 ( .A(n_662), .Y(n_848) );
AND2x4_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
AND2x4_ASAP7_75t_L g866 ( .A(n_663), .B(n_664), .Y(n_866) );
INVx2_ASAP7_75t_L g966 ( .A(n_664), .Y(n_966) );
BUFx2_ASAP7_75t_L g1463 ( .A(n_664), .Y(n_1463) );
NOR2xp33_ASAP7_75t_L g665 ( .A(n_666), .B(n_692), .Y(n_665) );
OAI33xp33_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_668), .A3(n_676), .B1(n_683), .B2(n_686), .B3(n_690), .Y(n_666) );
INVx1_ASAP7_75t_SL g820 ( .A(n_667), .Y(n_820) );
OAI33xp33_ASAP7_75t_L g915 ( .A1(n_667), .A2(n_916), .A3(n_922), .B1(n_927), .B2(n_932), .B3(n_938), .Y(n_915) );
OAI33xp33_ASAP7_75t_L g978 ( .A1(n_667), .A2(n_938), .A3(n_979), .B1(n_983), .B2(n_986), .B3(n_992), .Y(n_978) );
OAI22xp5_ASAP7_75t_L g1231 ( .A1(n_667), .A2(n_1232), .B1(n_1238), .B2(n_1240), .Y(n_1231) );
OAI33xp33_ASAP7_75t_L g1644 ( .A1(n_667), .A2(n_690), .A3(n_1645), .B1(n_1649), .B2(n_1653), .B3(n_1656), .Y(n_1644) );
OAI22xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_670), .B1(n_673), .B2(n_674), .Y(n_668) );
INVx1_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
OAI22xp33_ASAP7_75t_SL g676 ( .A1(n_677), .A2(n_678), .B1(n_680), .B2(n_681), .Y(n_676) );
OAI22xp33_ASAP7_75t_L g922 ( .A1(n_678), .A2(n_923), .B1(n_924), .B2(n_926), .Y(n_922) );
OAI22xp33_ASAP7_75t_L g927 ( .A1(n_678), .A2(n_928), .B1(n_929), .B2(n_931), .Y(n_927) );
OAI22xp33_ASAP7_75t_L g983 ( .A1(n_678), .A2(n_924), .B1(n_984), .B2(n_985), .Y(n_983) );
INVx2_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g972 ( .A(n_679), .Y(n_972) );
INVx2_ASAP7_75t_L g987 ( .A(n_679), .Y(n_987) );
INVx2_ASAP7_75t_L g1972 ( .A(n_679), .Y(n_1972) );
OAI221xp5_ASAP7_75t_L g1240 ( .A1(n_681), .A2(n_1233), .B1(n_1241), .B2(n_1242), .C(n_1243), .Y(n_1240) );
BUFx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g990 ( .A(n_682), .Y(n_990) );
INVx4_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
BUFx4f_ASAP7_75t_L g1239 ( .A(n_691), .Y(n_1239) );
BUFx4f_ASAP7_75t_L g1338 ( .A(n_691), .Y(n_1338) );
AOI33xp33_ASAP7_75t_L g1497 ( .A1(n_691), .A2(n_1328), .A3(n_1498), .B1(n_1502), .B2(n_1505), .B3(n_1508), .Y(n_1497) );
OAI33xp33_ASAP7_75t_L g692 ( .A1(n_693), .A2(n_695), .A3(n_698), .B1(n_701), .B2(n_710), .B3(n_717), .Y(n_692) );
OAI33xp33_ASAP7_75t_L g1399 ( .A1(n_693), .A2(n_717), .A3(n_1400), .B1(n_1408), .B2(n_1412), .B3(n_1416), .Y(n_1399) );
INVx1_ASAP7_75t_L g1625 ( .A(n_693), .Y(n_1625) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g1001 ( .A1(n_699), .A2(n_981), .B1(n_982), .B2(n_1002), .Y(n_1001) );
OAI221xp5_ASAP7_75t_L g1674 ( .A1(n_699), .A2(n_1675), .B1(n_1676), .B2(n_1678), .C(n_1679), .Y(n_1674) );
INVx2_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
OAI22xp5_ASAP7_75t_L g945 ( .A1(n_702), .A2(n_919), .B1(n_921), .B2(n_946), .Y(n_945) );
INVx2_ASAP7_75t_SL g702 ( .A(n_703), .Y(n_702) );
INVx2_ASAP7_75t_L g1251 ( .A(n_703), .Y(n_1251) );
INVx2_ASAP7_75t_L g1260 ( .A(n_703), .Y(n_1260) );
INVx2_ASAP7_75t_L g1364 ( .A(n_703), .Y(n_1364) );
BUFx3_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g1200 ( .A(n_704), .Y(n_1200) );
INVx1_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
INVx2_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g889 ( .A(n_707), .Y(n_889) );
INVx2_ASAP7_75t_L g1490 ( .A(n_707), .Y(n_1490) );
INVx2_ASAP7_75t_L g1550 ( .A(n_707), .Y(n_1550) );
INVx2_ASAP7_75t_L g1677 ( .A(n_707), .Y(n_1677) );
INVx3_ASAP7_75t_L g1951 ( .A(n_707), .Y(n_1951) );
BUFx6f_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx3_ASAP7_75t_L g729 ( .A(n_708), .Y(n_729) );
INVx3_ASAP7_75t_L g1003 ( .A(n_708), .Y(n_1003) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g1535 ( .A(n_713), .Y(n_1535) );
INVx1_ASAP7_75t_L g1628 ( .A(n_713), .Y(n_1628) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_714), .A2(n_923), .B1(n_926), .B2(n_949), .C(n_951), .Y(n_948) );
BUFx3_ASAP7_75t_L g1005 ( .A(n_714), .Y(n_1005) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_714), .B(n_1107), .Y(n_1106) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
AOI33xp33_ASAP7_75t_L g805 ( .A1(n_718), .A2(n_806), .A3(n_807), .B1(n_810), .B2(n_814), .B3(n_816), .Y(n_805) );
INVx6_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx5_ASAP7_75t_L g891 ( .A(n_719), .Y(n_891) );
NAND4xp25_ASAP7_75t_L g723 ( .A(n_724), .B(n_759), .C(n_775), .D(n_777), .Y(n_723) );
OAI31xp33_ASAP7_75t_L g724 ( .A1(n_725), .A2(n_754), .A3(n_757), .B(n_758), .Y(n_724) );
OAI221xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_731), .B1(n_735), .B2(n_739), .C(n_745), .Y(n_725) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_727), .A2(n_730), .B1(n_766), .B2(n_768), .Y(n_765) );
INVx2_ASAP7_75t_L g815 ( .A(n_728), .Y(n_815) );
INVx2_ASAP7_75t_SL g883 ( .A(n_728), .Y(n_883) );
INVx2_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
INVx2_ASAP7_75t_L g737 ( .A(n_729), .Y(n_737) );
INVx2_ASAP7_75t_L g1054 ( .A(n_729), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1124 ( .A(n_729), .Y(n_1124) );
INVx1_ASAP7_75t_L g1204 ( .A(n_729), .Y(n_1204) );
OAI21xp5_ASAP7_75t_L g731 ( .A1(n_732), .A2(n_733), .B(n_734), .Y(n_731) );
BUFx2_ASAP7_75t_L g1358 ( .A(n_733), .Y(n_1358) );
INVx1_ASAP7_75t_L g1406 ( .A(n_733), .Y(n_1406) );
INVx1_ASAP7_75t_L g813 ( .A(n_737), .Y(n_813) );
OAI21xp33_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B(n_742), .Y(n_739) );
A2O1A1Ixp33_ASAP7_75t_L g745 ( .A1(n_746), .A2(n_747), .B(n_748), .C(n_753), .Y(n_745) );
NAND2x1p5_ASAP7_75t_L g1396 ( .A(n_752), .B(n_1393), .Y(n_1396) );
INVx1_ASAP7_75t_L g1141 ( .A(n_758), .Y(n_1141) );
OAI31xp33_ASAP7_75t_L g1665 ( .A1(n_758), .A2(n_1666), .A3(n_1667), .B(n_1673), .Y(n_1665) );
OAI31xp33_ASAP7_75t_L g2009 ( .A1(n_758), .A2(n_2010), .A3(n_2011), .B(n_2017), .Y(n_2009) );
INVx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g1147 ( .A(n_762), .Y(n_1147) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g1330 ( .A(n_766), .Y(n_1330) );
INVx1_ASAP7_75t_L g1587 ( .A(n_766), .Y(n_1587) );
INVx2_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
AND2x4_ASAP7_75t_L g1428 ( .A(n_767), .B(n_1429), .Y(n_1428) );
BUFx3_ASAP7_75t_L g1437 ( .A(n_767), .Y(n_1437) );
OAI22xp33_ASAP7_75t_L g979 ( .A1(n_768), .A2(n_980), .B1(n_981), .B2(n_982), .Y(n_979) );
INVx1_ASAP7_75t_L g1284 ( .A(n_768), .Y(n_1284) );
INVx1_ASAP7_75t_L g1660 ( .A(n_768), .Y(n_1660) );
INVx1_ASAP7_75t_L g1969 ( .A(n_768), .Y(n_1969) );
OA22x2_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_849), .B1(n_850), .B2(n_906), .Y(n_778) );
INVx1_ASAP7_75t_L g906 ( .A(n_779), .Y(n_906) );
XNOR2xp5_ASAP7_75t_L g779 ( .A(n_780), .B(n_781), .Y(n_779) );
AOI211xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_784), .B(n_804), .C(n_832), .Y(n_781) );
AOI221x1_ASAP7_75t_L g851 ( .A1(n_782), .A2(n_852), .B1(n_865), .B2(n_867), .C(n_880), .Y(n_851) );
AOI221x1_ASAP7_75t_L g1024 ( .A1(n_782), .A2(n_865), .B1(n_1025), .B2(n_1037), .C(n_1048), .Y(n_1024) );
CKINVDCx16_ASAP7_75t_R g782 ( .A(n_783), .Y(n_782) );
AOI22xp5_ASAP7_75t_L g785 ( .A1(n_786), .A2(n_787), .B1(n_788), .B2(n_789), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_787), .A2(n_789), .B1(n_869), .B2(n_870), .Y(n_868) );
AOI22xp33_ASAP7_75t_L g1038 ( .A1(n_787), .A2(n_789), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
AOI22xp33_ASAP7_75t_SL g1514 ( .A1(n_787), .A2(n_789), .B1(n_1515), .B2(n_1516), .Y(n_1514) );
INVx4_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx5_ASAP7_75t_L g1047 ( .A(n_794), .Y(n_1047) );
INVx2_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx2_ASAP7_75t_SL g1496 ( .A(n_798), .Y(n_1496) );
INVx2_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
BUFx6f_ASAP7_75t_L g809 ( .A(n_799), .Y(n_809) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
NAND2xp5_ASAP7_75t_SL g804 ( .A(n_805), .B(n_819), .Y(n_804) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_806), .B(n_882), .C(n_884), .Y(n_881) );
NAND3xp33_ASAP7_75t_L g1055 ( .A(n_806), .B(n_1056), .C(n_1060), .Y(n_1055) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
BUFx2_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
INVx2_ASAP7_75t_SL g886 ( .A(n_818), .Y(n_886) );
HB1xp67_ASAP7_75t_L g1051 ( .A(n_818), .Y(n_1051) );
BUFx6f_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx1_ASAP7_75t_L g1454 ( .A(n_826), .Y(n_1454) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
AOI31xp33_ASAP7_75t_SL g832 ( .A1(n_833), .A2(n_840), .A3(n_844), .B(n_848), .Y(n_832) );
INVx2_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g861 ( .A(n_837), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g1468 ( .A1(n_842), .A2(n_845), .B1(n_1469), .B2(n_1470), .Y(n_1468) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
INVx1_ASAP7_75t_L g905 ( .A(n_851), .Y(n_905) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_857), .Y(n_852) );
AND2x4_ASAP7_75t_L g1455 ( .A(n_864), .B(n_1456), .Y(n_1455) );
INVx1_ASAP7_75t_L g1599 ( .A(n_864), .Y(n_1599) );
BUFx6f_ASAP7_75t_L g1977 ( .A(n_864), .Y(n_1977) );
BUFx6f_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx1_ASAP7_75t_L g1481 ( .A(n_866), .Y(n_1481) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND4xp25_ASAP7_75t_L g880 ( .A(n_881), .B(n_887), .C(n_892), .D(n_900), .Y(n_880) );
INVx2_ASAP7_75t_L g885 ( .A(n_886), .Y(n_885) );
NAND3xp33_ASAP7_75t_L g887 ( .A(n_888), .B(n_890), .C(n_891), .Y(n_887) );
INVx1_ASAP7_75t_L g1253 ( .A(n_889), .Y(n_1253) );
NAND3xp33_ASAP7_75t_L g1049 ( .A(n_891), .B(n_1050), .C(n_1052), .Y(n_1049) );
AOI33xp33_ASAP7_75t_L g1483 ( .A1(n_891), .A2(n_1484), .A3(n_1487), .B1(n_1491), .B2(n_1493), .B3(n_1495), .Y(n_1483) );
CKINVDCx8_ASAP7_75t_R g1637 ( .A(n_891), .Y(n_1637) );
NAND3xp33_ASAP7_75t_L g892 ( .A(n_893), .B(n_896), .C(n_897), .Y(n_892) );
BUFx6f_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g920 ( .A(n_895), .Y(n_920) );
INVx1_ASAP7_75t_L g1182 ( .A(n_895), .Y(n_1182) );
INVx1_ASAP7_75t_L g1439 ( .A(n_895), .Y(n_1439) );
BUFx3_ASAP7_75t_L g1603 ( .A(n_895), .Y(n_1603) );
NAND3xp33_ASAP7_75t_L g1061 ( .A(n_897), .B(n_1062), .C(n_1063), .Y(n_1061) );
INVx3_ASAP7_75t_L g897 ( .A(n_898), .Y(n_897) );
XNOR2xp5_ASAP7_75t_L g907 ( .A(n_908), .B(n_1020), .Y(n_907) );
XOR2xp5_ASAP7_75t_L g908 ( .A(n_909), .B(n_975), .Y(n_908) );
AND4x1_ASAP7_75t_L g910 ( .A(n_911), .B(n_940), .C(n_942), .D(n_967), .Y(n_910) );
NOR3xp33_ASAP7_75t_L g911 ( .A(n_912), .B(n_915), .C(n_939), .Y(n_911) );
NOR3xp33_ASAP7_75t_L g977 ( .A(n_912), .B(n_978), .C(n_995), .Y(n_977) );
BUFx2_ASAP7_75t_L g1170 ( .A(n_912), .Y(n_1170) );
NOR3xp33_ASAP7_75t_SL g1230 ( .A(n_912), .B(n_1231), .C(n_1244), .Y(n_1230) );
HB1xp67_ASAP7_75t_L g1643 ( .A(n_912), .Y(n_1643) );
INVx1_ASAP7_75t_L g913 ( .A(n_914), .Y(n_913) );
INVx1_ASAP7_75t_L g1583 ( .A(n_914), .Y(n_1583) );
OAI22xp33_ASAP7_75t_L g916 ( .A1(n_917), .A2(n_919), .B1(n_920), .B2(n_921), .Y(n_916) );
OAI22xp33_ASAP7_75t_L g1645 ( .A1(n_917), .A2(n_1646), .B1(n_1647), .B2(n_1648), .Y(n_1645) );
INVx2_ASAP7_75t_SL g917 ( .A(n_918), .Y(n_917) );
BUFx3_ASAP7_75t_L g1499 ( .A(n_918), .Y(n_1499) );
OAI22xp5_ASAP7_75t_L g992 ( .A1(n_920), .A2(n_933), .B1(n_993), .B2(n_994), .Y(n_992) );
INVx2_ASAP7_75t_SL g924 ( .A(n_925), .Y(n_924) );
BUFx2_ASAP7_75t_L g1178 ( .A(n_929), .Y(n_1178) );
INVx1_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g1235 ( .A(n_930), .Y(n_1235) );
INVx1_ASAP7_75t_L g1441 ( .A(n_930), .Y(n_1441) );
OAI22xp5_ASAP7_75t_L g932 ( .A1(n_933), .A2(n_934), .B1(n_935), .B2(n_937), .Y(n_932) );
INVx2_ASAP7_75t_SL g935 ( .A(n_936), .Y(n_935) );
OAI31xp33_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_944), .A3(n_953), .B(n_965), .Y(n_942) );
OAI221xp5_ASAP7_75t_L g1259 ( .A1(n_946), .A2(n_1260), .B1(n_1261), .B2(n_1262), .C(n_1263), .Y(n_1259) );
OAI22xp5_ASAP7_75t_L g1635 ( .A1(n_946), .A2(n_1590), .B1(n_1608), .B2(n_1631), .Y(n_1635) );
INVx4_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
INVx2_ASAP7_75t_SL g957 ( .A(n_947), .Y(n_957) );
INVx2_ASAP7_75t_SL g1011 ( .A(n_947), .Y(n_1011) );
BUFx3_ASAP7_75t_L g1367 ( .A(n_947), .Y(n_1367) );
INVx2_ASAP7_75t_SL g1414 ( .A(n_947), .Y(n_1414) );
OAI22xp33_ASAP7_75t_L g1626 ( .A1(n_949), .A2(n_1627), .B1(n_1628), .B2(n_1629), .Y(n_1626) );
INVx2_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx1_ASAP7_75t_L g1360 ( .A(n_950), .Y(n_1360) );
OAI221xp5_ASAP7_75t_L g1357 ( .A1(n_951), .A2(n_1358), .B1(n_1359), .B2(n_1360), .C(n_1361), .Y(n_1357) );
INVx2_ASAP7_75t_L g1140 ( .A(n_952), .Y(n_1140) );
OAI221xp5_ASAP7_75t_L g954 ( .A1(n_955), .A2(n_956), .B1(n_957), .B2(n_958), .C(n_959), .Y(n_954) );
OAI221xp5_ASAP7_75t_L g1009 ( .A1(n_955), .A2(n_1010), .B1(n_1011), .B2(n_1012), .C(n_1013), .Y(n_1009) );
INVx1_ASAP7_75t_L g1311 ( .A(n_955), .Y(n_1311) );
OAI22xp5_ASAP7_75t_L g1408 ( .A1(n_957), .A2(n_1409), .B1(n_1410), .B2(n_1411), .Y(n_1408) );
OAI22xp5_ASAP7_75t_L g1539 ( .A1(n_957), .A2(n_1540), .B1(n_1541), .B2(n_1542), .Y(n_1539) );
OAI22xp5_ASAP7_75t_L g1630 ( .A1(n_957), .A2(n_1631), .B1(n_1633), .B2(n_1634), .Y(n_1630) );
AND2x6_ASAP7_75t_L g1382 ( .A(n_960), .B(n_1380), .Y(n_1382) );
NAND2x1p5_ASAP7_75t_L g1398 ( .A(n_960), .B(n_1393), .Y(n_1398) );
OAI31xp33_ASAP7_75t_L g998 ( .A1(n_965), .A2(n_999), .A3(n_1000), .B(n_1008), .Y(n_998) );
OAI21xp5_ASAP7_75t_L g1089 ( .A1(n_965), .A2(n_1090), .B(n_1099), .Y(n_1089) );
OAI31xp33_ASAP7_75t_L g1247 ( .A1(n_965), .A2(n_1248), .A3(n_1249), .B(n_1258), .Y(n_1247) );
OAI31xp33_ASAP7_75t_L g1348 ( .A1(n_965), .A2(n_1349), .A3(n_1356), .B(n_1368), .Y(n_1348) );
BUFx8_ASAP7_75t_SL g965 ( .A(n_966), .Y(n_965) );
INVx2_ASAP7_75t_L g1579 ( .A(n_966), .Y(n_1579) );
NOR2xp33_ASAP7_75t_L g967 ( .A(n_968), .B(n_970), .Y(n_967) );
AND4x1_ASAP7_75t_L g976 ( .A(n_977), .B(n_996), .C(n_998), .D(n_1017), .Y(n_976) );
OAI21xp33_ASAP7_75t_SL g1004 ( .A1(n_985), .A2(n_1005), .B(n_1006), .Y(n_1004) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_988), .B1(n_989), .B2(n_991), .Y(n_986) );
OAI221xp5_ASAP7_75t_L g1183 ( .A1(n_987), .A2(n_989), .B1(n_1184), .B2(n_1185), .C(n_1186), .Y(n_1183) );
OAI221xp5_ASAP7_75t_L g1285 ( .A1(n_987), .A2(n_1178), .B1(n_1286), .B2(n_1287), .C(n_1288), .Y(n_1285) );
OAI221xp5_ASAP7_75t_L g2004 ( .A1(n_987), .A2(n_1235), .B1(n_2005), .B2(n_2006), .C(n_2007), .Y(n_2004) );
INVx2_ASAP7_75t_L g989 ( .A(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
INVx2_ASAP7_75t_L g1059 ( .A(n_1003), .Y(n_1059) );
BUFx3_ASAP7_75t_L g1314 ( .A(n_1003), .Y(n_1314) );
AND2x4_ASAP7_75t_L g1379 ( .A(n_1003), .B(n_1380), .Y(n_1379) );
OAI21xp33_ASAP7_75t_L g1255 ( .A1(n_1005), .A2(n_1236), .B(n_1256), .Y(n_1255) );
OAI22xp33_ASAP7_75t_L g1636 ( .A1(n_1005), .A2(n_1401), .B1(n_1605), .B2(n_1607), .Y(n_1636) );
OAI22xp33_ASAP7_75t_L g1942 ( .A1(n_1005), .A2(n_1943), .B1(n_1944), .B2(n_1946), .Y(n_1942) );
OAI22xp33_ASAP7_75t_L g1956 ( .A1(n_1005), .A2(n_1944), .B1(n_1957), .B2(n_1958), .Y(n_1956) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_1018), .B(n_1019), .Y(n_1017) );
OAI22x1_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1022), .B1(n_1070), .B2(n_1071), .Y(n_1020) );
INVx1_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
INVx1_ASAP7_75t_L g1069 ( .A(n_1024), .Y(n_1069) );
NAND3xp33_ASAP7_75t_L g1025 ( .A(n_1026), .B(n_1031), .C(n_1034), .Y(n_1025) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1029), .Y(n_1028) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
HB1xp67_ASAP7_75t_L g1651 ( .A(n_1030), .Y(n_1651) );
NAND4xp25_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1055), .C(n_1061), .D(n_1064), .Y(n_1048) );
INVx1_ASAP7_75t_L g1671 ( .A(n_1053), .Y(n_1671) );
INVx2_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1058 ( .A(n_1059), .Y(n_1058) );
NAND3xp33_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1066), .C(n_1067), .Y(n_1064) );
AOI33xp33_ASAP7_75t_L g1563 ( .A1(n_1067), .A2(n_1564), .A3(n_1565), .B1(n_1567), .B2(n_1569), .B3(n_1570), .Y(n_1563) );
INVx1_ASAP7_75t_L g1067 ( .A(n_1068), .Y(n_1067) );
INVx2_ASAP7_75t_SL g1070 ( .A(n_1071), .Y(n_1070) );
INVx2_ASAP7_75t_L g1072 ( .A(n_1073), .Y(n_1072) );
NAND4xp75_ASAP7_75t_L g1073 ( .A(n_1074), .B(n_1089), .C(n_1110), .D(n_1112), .Y(n_1073) );
AND2x2_ASAP7_75t_L g1074 ( .A(n_1075), .B(n_1085), .Y(n_1074) );
INVx2_ASAP7_75t_L g1081 ( .A(n_1082), .Y(n_1081) );
INVx1_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
INVx2_ASAP7_75t_L g1245 ( .A(n_1086), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1090 ( .A(n_1091), .B(n_1094), .Y(n_1090) );
BUFx3_ASAP7_75t_L g1488 ( .A(n_1096), .Y(n_1488) );
NAND2x1p5_ASAP7_75t_L g1130 ( .A(n_1108), .B(n_1131), .Y(n_1130) );
NAND2x1_ASAP7_75t_SL g1392 ( .A(n_1108), .B(n_1393), .Y(n_1392) );
INVx2_ASAP7_75t_L g1108 ( .A(n_1109), .Y(n_1108) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
INVx2_ASAP7_75t_L g1161 ( .A(n_1116), .Y(n_1161) );
XOR2x2_ASAP7_75t_L g1116 ( .A(n_1117), .B(n_1159), .Y(n_1116) );
NOR3xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1120), .C(n_1142), .Y(n_1117) );
AOI31xp33_ASAP7_75t_L g1120 ( .A1(n_1121), .A2(n_1132), .A3(n_1135), .B(n_1141), .Y(n_1120) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1139), .Y(n_1214) );
NAND4xp25_ASAP7_75t_L g1142 ( .A(n_1143), .B(n_1150), .C(n_1153), .D(n_1156), .Y(n_1142) );
INVx1_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
XNOR2xp5_ASAP7_75t_L g1163 ( .A(n_1164), .B(n_1223), .Y(n_1163) );
CKINVDCx14_ASAP7_75t_R g1164 ( .A(n_1165), .Y(n_1164) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1166), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_1167), .Y(n_1166) );
AND4x1_ASAP7_75t_L g1168 ( .A(n_1169), .B(n_1192), .C(n_1194), .D(n_1220), .Y(n_1168) );
NOR3xp33_ASAP7_75t_SL g1169 ( .A(n_1170), .B(n_1171), .C(n_1190), .Y(n_1169) );
NOR3xp33_ASAP7_75t_SL g1276 ( .A(n_1170), .B(n_1277), .C(n_1279), .Y(n_1276) );
NOR3xp33_ASAP7_75t_SL g1998 ( .A(n_1170), .B(n_1999), .C(n_2008), .Y(n_1998) );
OAI221xp5_ASAP7_75t_L g1172 ( .A1(n_1173), .A2(n_1176), .B1(n_1177), .B2(n_1178), .C(n_1179), .Y(n_1172) );
OAI221xp5_ASAP7_75t_L g2000 ( .A1(n_1173), .A2(n_1178), .B1(n_2001), .B2(n_2002), .C(n_2003), .Y(n_2000) );
BUFx2_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
INVx2_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g1181 ( .A(n_1182), .Y(n_1181) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
BUFx3_ASAP7_75t_L g1289 ( .A(n_1189), .Y(n_1289) );
BUFx2_ASAP7_75t_L g1597 ( .A(n_1189), .Y(n_1597) );
INVx1_ASAP7_75t_L g1657 ( .A(n_1189), .Y(n_1657) );
INVx2_ASAP7_75t_L g1968 ( .A(n_1189), .Y(n_1968) );
OAI22xp5_ASAP7_75t_L g1197 ( .A1(n_1198), .A2(n_1201), .B1(n_1202), .B2(n_1205), .Y(n_1197) );
OAI22xp5_ASAP7_75t_L g1947 ( .A1(n_1198), .A2(n_1948), .B1(n_1949), .B2(n_1950), .Y(n_1947) );
INVx2_ASAP7_75t_L g1198 ( .A(n_1199), .Y(n_1198) );
INVx2_ASAP7_75t_L g1210 ( .A(n_1199), .Y(n_1210) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1199), .Y(n_1297) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
BUFx2_ASAP7_75t_L g1351 ( .A(n_1200), .Y(n_1351) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1203), .Y(n_1202) );
INVx1_ASAP7_75t_L g1203 ( .A(n_1204), .Y(n_1203) );
OAI221xp5_ASAP7_75t_L g1209 ( .A1(n_1210), .A2(n_1211), .B1(n_1212), .B2(n_1215), .C(n_1216), .Y(n_1209) );
OAI221xp5_ASAP7_75t_L g2018 ( .A1(n_1210), .A2(n_1299), .B1(n_2019), .B2(n_2020), .C(n_2021), .Y(n_2018) );
OAI221xp5_ASAP7_75t_L g1350 ( .A1(n_1212), .A2(n_1341), .B1(n_1345), .B2(n_1351), .C(n_1352), .Y(n_1350) );
INVx1_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
NOR2xp33_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1222), .Y(n_1220) );
XNOR2xp5_ASAP7_75t_L g1223 ( .A(n_1224), .B(n_1270), .Y(n_1223) );
INVx1_ASAP7_75t_L g1224 ( .A(n_1225), .Y(n_1224) );
HB1xp67_ASAP7_75t_L g1225 ( .A(n_1226), .Y(n_1225) );
AND4x1_ASAP7_75t_L g1227 ( .A(n_1228), .B(n_1230), .C(n_1247), .D(n_1267), .Y(n_1227) );
OAI221xp5_ASAP7_75t_L g1232 ( .A1(n_1233), .A2(n_1234), .B1(n_1235), .B2(n_1236), .C(n_1237), .Y(n_1232) );
OAI221xp5_ASAP7_75t_L g1440 ( .A1(n_1233), .A2(n_1381), .B1(n_1384), .B2(n_1441), .C(n_1442), .Y(n_1440) );
OAI22xp33_ASAP7_75t_L g1649 ( .A1(n_1233), .A2(n_1650), .B1(n_1651), .B2(n_1652), .Y(n_1649) );
CKINVDCx5p33_ASAP7_75t_R g1238 ( .A(n_1239), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g1250 ( .A1(n_1251), .A2(n_1252), .B1(n_1253), .B2(n_1254), .Y(n_1250) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1257), .Y(n_1354) );
AND2x4_ASAP7_75t_L g1385 ( .A(n_1257), .B(n_1380), .Y(n_1385) );
BUFx3_ASAP7_75t_L g1492 ( .A(n_1257), .Y(n_1492) );
INVx2_ASAP7_75t_L g1632 ( .A(n_1260), .Y(n_1632) );
NOR2xp33_ASAP7_75t_L g1267 ( .A(n_1268), .B(n_1269), .Y(n_1267) );
AO22x2_ASAP7_75t_L g1270 ( .A1(n_1271), .A2(n_1524), .B1(n_1525), .B2(n_1686), .Y(n_1270) );
INVx2_ASAP7_75t_SL g1686 ( .A(n_1271), .Y(n_1686) );
AO22x2_ASAP7_75t_L g1271 ( .A1(n_1272), .A2(n_1273), .B1(n_1371), .B2(n_1523), .Y(n_1271) );
INVx1_ASAP7_75t_L g1272 ( .A(n_1273), .Y(n_1272) );
AO22x1_ASAP7_75t_L g1273 ( .A1(n_1274), .A2(n_1320), .B1(n_1369), .B2(n_1370), .Y(n_1273) );
INVx1_ASAP7_75t_L g1370 ( .A(n_1274), .Y(n_1370) );
AND4x1_ASAP7_75t_L g1275 ( .A(n_1276), .B(n_1292), .C(n_1294), .D(n_1317), .Y(n_1275) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1291), .Y(n_1290) );
INVx1_ASAP7_75t_L g1331 ( .A(n_1291), .Y(n_1331) );
OAI221xp5_ASAP7_75t_L g1296 ( .A1(n_1297), .A2(n_1298), .B1(n_1299), .B2(n_1301), .C(n_1302), .Y(n_1296) );
INVx1_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
OAI22xp5_ASAP7_75t_L g1309 ( .A1(n_1310), .A2(n_1312), .B1(n_1313), .B2(n_1315), .Y(n_1309) );
OAI22xp5_ASAP7_75t_L g1952 ( .A1(n_1310), .A2(n_1953), .B1(n_1954), .B2(n_1955), .Y(n_1952) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
CKINVDCx5p33_ASAP7_75t_R g1313 ( .A(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1955 ( .A(n_1314), .Y(n_1955) );
NOR2xp33_ASAP7_75t_L g1317 ( .A(n_1318), .B(n_1319), .Y(n_1317) );
INVx1_ASAP7_75t_L g1369 ( .A(n_1320), .Y(n_1369) );
AND3x1_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1346), .C(n_1348), .Y(n_1321) );
NOR2xp33_ASAP7_75t_L g1322 ( .A(n_1323), .B(n_1339), .Y(n_1322) );
AOI33xp33_ASAP7_75t_L g1327 ( .A1(n_1328), .A2(n_1329), .A3(n_1332), .B1(n_1335), .B2(n_1337), .B3(n_1338), .Y(n_1327) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1343), .Y(n_1339) );
OAI22xp5_ASAP7_75t_L g1547 ( .A1(n_1351), .A2(n_1548), .B1(n_1549), .B2(n_1551), .Y(n_1547) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1354), .Y(n_1353) );
OAI22xp5_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1364), .B1(n_1365), .B2(n_1366), .Y(n_1362) );
INVx1_ASAP7_75t_L g1366 ( .A(n_1367), .Y(n_1366) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1371), .Y(n_1523) );
AOI22x1_ASAP7_75t_L g1371 ( .A1(n_1372), .A2(n_1464), .B1(n_1520), .B2(n_1521), .Y(n_1371) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1420), .Y(n_1373) );
NOR3xp33_ASAP7_75t_L g1374 ( .A(n_1375), .B(n_1389), .C(n_1399), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1376), .B(n_1383), .Y(n_1375) );
AOI22xp33_ASAP7_75t_L g1376 ( .A1(n_1377), .A2(n_1378), .B1(n_1381), .B2(n_1382), .Y(n_1376) );
BUFx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
BUFx2_ASAP7_75t_L g1615 ( .A(n_1379), .Y(n_1615) );
BUFx2_ASAP7_75t_L g1934 ( .A(n_1379), .Y(n_1934) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1380), .B(n_1388), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1620 ( .A(n_1380), .B(n_1388), .Y(n_1620) );
AOI22xp33_ASAP7_75t_L g1613 ( .A1(n_1382), .A2(n_1614), .B1(n_1615), .B2(n_1616), .Y(n_1613) );
AOI22xp33_ASAP7_75t_L g1932 ( .A1(n_1382), .A2(n_1933), .B1(n_1934), .B2(n_1935), .Y(n_1932) );
AOI22xp33_ASAP7_75t_L g1383 ( .A1(n_1384), .A2(n_1385), .B1(n_1386), .B2(n_1387), .Y(n_1383) );
AOI22xp33_ASAP7_75t_L g1617 ( .A1(n_1385), .A2(n_1618), .B1(n_1619), .B2(n_1620), .Y(n_1617) );
AOI22xp33_ASAP7_75t_L g1936 ( .A1(n_1385), .A2(n_1387), .B1(n_1937), .B2(n_1938), .Y(n_1936) );
INVx2_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
INVx2_ASAP7_75t_SL g1622 ( .A(n_1391), .Y(n_1622) );
INVx2_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx3_ASAP7_75t_L g1393 ( .A(n_1394), .Y(n_1393) );
BUFx4f_ASAP7_75t_L g1395 ( .A(n_1396), .Y(n_1395) );
BUFx2_ASAP7_75t_L g1397 ( .A(n_1398), .Y(n_1397) );
BUFx3_ASAP7_75t_L g1940 ( .A(n_1398), .Y(n_1940) );
OAI22xp33_ASAP7_75t_L g1400 ( .A1(n_1401), .A2(n_1404), .B1(n_1405), .B2(n_1407), .Y(n_1400) );
OAI22xp33_ASAP7_75t_L g1416 ( .A1(n_1401), .A2(n_1417), .B1(n_1418), .B2(n_1419), .Y(n_1416) );
BUFx2_ASAP7_75t_L g1401 ( .A(n_1402), .Y(n_1401) );
INVx2_ASAP7_75t_L g1402 ( .A(n_1403), .Y(n_1402) );
INVx1_ASAP7_75t_L g1405 ( .A(n_1406), .Y(n_1405) );
INVx1_ASAP7_75t_L g1418 ( .A(n_1406), .Y(n_1418) );
OAI22xp5_ASAP7_75t_L g1412 ( .A1(n_1410), .A2(n_1413), .B1(n_1414), .B2(n_1415), .Y(n_1412) );
AOI211xp5_ASAP7_75t_L g1427 ( .A1(n_1413), .A2(n_1428), .B(n_1430), .C(n_1436), .Y(n_1427) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1414), .Y(n_1494) );
AOI22xp33_ASAP7_75t_L g1457 ( .A1(n_1415), .A2(n_1417), .B1(n_1458), .B2(n_1460), .Y(n_1457) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_1419), .A2(n_1445), .B1(n_1448), .B2(n_1452), .C(n_1455), .Y(n_1444) );
AOI21xp5_ASAP7_75t_L g1420 ( .A1(n_1421), .A2(n_1425), .B(n_1426), .Y(n_1420) );
INVx1_ASAP7_75t_L g1421 ( .A(n_1422), .Y(n_1421) );
INVx5_ASAP7_75t_L g1610 ( .A(n_1422), .Y(n_1610) );
AND2x4_ASAP7_75t_L g1422 ( .A(n_1423), .B(n_1424), .Y(n_1422) );
AOI31xp33_ASAP7_75t_L g1426 ( .A1(n_1427), .A2(n_1444), .A3(n_1457), .B(n_1462), .Y(n_1426) );
AOI221xp5_ASAP7_75t_L g1581 ( .A1(n_1428), .A2(n_1582), .B1(n_1586), .B2(n_1590), .C(n_1591), .Y(n_1581) );
AOI22xp33_ASAP7_75t_L g1981 ( .A1(n_1428), .A2(n_1458), .B1(n_1953), .B2(n_1957), .Y(n_1981) );
INVx2_ASAP7_75t_SL g1431 ( .A(n_1432), .Y(n_1431) );
INVx2_ASAP7_75t_L g1592 ( .A(n_1432), .Y(n_1592) );
INVx1_ASAP7_75t_L g1963 ( .A(n_1432), .Y(n_1963) );
INVx1_ASAP7_75t_SL g1456 ( .A(n_1435), .Y(n_1456) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1442 ( .A(n_1443), .Y(n_1442) );
BUFx2_ASAP7_75t_L g1585 ( .A(n_1443), .Y(n_1585) );
INVx1_ASAP7_75t_L g1445 ( .A(n_1446), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
BUFx6f_ASAP7_75t_L g1604 ( .A(n_1447), .Y(n_1604) );
INVx1_ASAP7_75t_L g1449 ( .A(n_1450), .Y(n_1449) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1451), .Y(n_1601) );
INVx2_ASAP7_75t_L g1453 ( .A(n_1454), .Y(n_1453) );
AOI221xp5_ASAP7_75t_L g1595 ( .A1(n_1455), .A2(n_1596), .B1(n_1602), .B2(n_1604), .C(n_1605), .Y(n_1595) );
AOI221xp5_ASAP7_75t_L g1975 ( .A1(n_1455), .A2(n_1604), .B1(n_1958), .B2(n_1976), .C(n_1980), .Y(n_1975) );
AOI22xp33_ASAP7_75t_L g1606 ( .A1(n_1458), .A2(n_1460), .B1(n_1607), .B2(n_1608), .Y(n_1606) );
INVx6_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
AOI211xp5_ASAP7_75t_L g1961 ( .A1(n_1460), .A2(n_1954), .B(n_1962), .C(n_1966), .Y(n_1961) );
INVx4_ASAP7_75t_L g1460 ( .A(n_1461), .Y(n_1460) );
INVx2_ASAP7_75t_L g1462 ( .A(n_1463), .Y(n_1462) );
AOI22xp5_ASAP7_75t_L g1959 ( .A1(n_1463), .A2(n_1610), .B1(n_1960), .B2(n_1982), .Y(n_1959) );
INVx2_ASAP7_75t_L g1520 ( .A(n_1464), .Y(n_1520) );
INVx1_ASAP7_75t_L g1519 ( .A(n_1466), .Y(n_1519) );
AOI211x1_ASAP7_75t_L g1466 ( .A1(n_1467), .A2(n_1480), .B(n_1482), .C(n_1509), .Y(n_1466) );
NAND4xp25_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1471), .C(n_1474), .D(n_1479), .Y(n_1467) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1483), .B(n_1497), .Y(n_1482) );
INVx2_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx2_ASAP7_75t_L g1485 ( .A(n_1486), .Y(n_1485) );
HB1xp67_ASAP7_75t_L g1489 ( .A(n_1490), .Y(n_1489) );
INVx1_ASAP7_75t_L g1500 ( .A(n_1501), .Y(n_1500) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
INVx3_ASAP7_75t_SL g1521 ( .A(n_1522), .Y(n_1521) );
INVx1_ASAP7_75t_L g1524 ( .A(n_1525), .Y(n_1524) );
XOR2xp5_ASAP7_75t_L g1525 ( .A(n_1526), .B(n_1638), .Y(n_1525) );
INVx1_ASAP7_75t_L g1526 ( .A(n_1527), .Y(n_1526) );
AOI22x1_ASAP7_75t_L g1527 ( .A1(n_1528), .A2(n_1529), .B1(n_1574), .B2(n_1575), .Y(n_1527) );
INVx2_ASAP7_75t_L g1528 ( .A(n_1529), .Y(n_1528) );
NAND3xp33_ASAP7_75t_L g1530 ( .A(n_1531), .B(n_1557), .C(n_1559), .Y(n_1530) );
INVx1_ASAP7_75t_L g1549 ( .A(n_1550), .Y(n_1549) );
INVx1_ASAP7_75t_L g1554 ( .A(n_1555), .Y(n_1554) );
NOR2xp33_ASAP7_75t_SL g1559 ( .A(n_1560), .B(n_1571), .Y(n_1559) );
INVx1_ASAP7_75t_L g1647 ( .A(n_1566), .Y(n_1647) );
NAND2xp5_ASAP7_75t_L g1571 ( .A(n_1572), .B(n_1573), .Y(n_1571) );
INVx2_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
XNOR2x1_ASAP7_75t_L g1575 ( .A(n_1576), .B(n_1577), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1577 ( .A(n_1578), .B(n_1611), .Y(n_1577) );
AOI22xp33_ASAP7_75t_L g1578 ( .A1(n_1579), .A2(n_1580), .B1(n_1609), .B2(n_1610), .Y(n_1578) );
NAND3xp33_ASAP7_75t_L g1580 ( .A(n_1581), .B(n_1595), .C(n_1606), .Y(n_1580) );
HB1xp67_ASAP7_75t_L g1588 ( .A(n_1589), .Y(n_1588) );
INVx2_ASAP7_75t_SL g1593 ( .A(n_1594), .Y(n_1593) );
INVx1_ASAP7_75t_L g1598 ( .A(n_1599), .Y(n_1598) );
INVx1_ASAP7_75t_L g1600 ( .A(n_1601), .Y(n_1600) );
NOR3xp33_ASAP7_75t_SL g1611 ( .A(n_1612), .B(n_1621), .C(n_1623), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1612 ( .A(n_1613), .B(n_1617), .Y(n_1612) );
OAI33xp33_ASAP7_75t_L g1623 ( .A1(n_1624), .A2(n_1626), .A3(n_1630), .B1(n_1635), .B2(n_1636), .B3(n_1637), .Y(n_1623) );
OAI33xp33_ASAP7_75t_L g1941 ( .A1(n_1624), .A2(n_1637), .A3(n_1942), .B1(n_1947), .B2(n_1952), .B3(n_1956), .Y(n_1941) );
INVx1_ASAP7_75t_L g1624 ( .A(n_1625), .Y(n_1624) );
INVx2_ASAP7_75t_L g1631 ( .A(n_1632), .Y(n_1631) );
HB1xp67_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1639 ( .A(n_1640), .Y(n_1639) );
AND4x1_ASAP7_75t_L g1641 ( .A(n_1642), .B(n_1663), .C(n_1665), .D(n_1683), .Y(n_1641) );
NOR3xp33_ASAP7_75t_L g1642 ( .A(n_1643), .B(n_1644), .C(n_1662), .Y(n_1642) );
OAI22xp5_ASAP7_75t_L g1668 ( .A1(n_1646), .A2(n_1648), .B1(n_1669), .B2(n_1671), .Y(n_1668) );
OAI22xp5_ASAP7_75t_L g1656 ( .A1(n_1657), .A2(n_1658), .B1(n_1659), .B2(n_1661), .Y(n_1656) );
INVx1_ASAP7_75t_L g1659 ( .A(n_1660), .Y(n_1659) );
INVx1_ASAP7_75t_L g1669 ( .A(n_1670), .Y(n_1669) );
INVx1_ASAP7_75t_L g1676 ( .A(n_1677), .Y(n_1676) );
NOR2xp33_ASAP7_75t_L g1683 ( .A(n_1684), .B(n_1685), .Y(n_1683) );
OAI221xp5_ASAP7_75t_L g1687 ( .A1(n_1688), .A2(n_1924), .B1(n_1926), .B2(n_1983), .C(n_1987), .Y(n_1687) );
NOR2x1_ASAP7_75t_L g1688 ( .A(n_1689), .B(n_1859), .Y(n_1688) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_1690), .B(n_1782), .Y(n_1689) );
A2O1A1Ixp33_ASAP7_75t_SL g1690 ( .A1(n_1691), .A2(n_1723), .B(n_1743), .C(n_1774), .Y(n_1690) );
AND2x2_ASAP7_75t_L g1809 ( .A(n_1691), .B(n_1772), .Y(n_1809) );
NAND2xp5_ASAP7_75t_L g1838 ( .A(n_1691), .B(n_1839), .Y(n_1838) );
INVx1_ASAP7_75t_L g1863 ( .A(n_1691), .Y(n_1863) );
AND2x2_ASAP7_75t_L g1691 ( .A(n_1692), .B(n_1711), .Y(n_1691) );
INVx2_ASAP7_75t_L g1759 ( .A(n_1692), .Y(n_1759) );
BUFx3_ASAP7_75t_L g1799 ( .A(n_1692), .Y(n_1799) );
OR2x2_ASAP7_75t_L g1847 ( .A(n_1692), .B(n_1795), .Y(n_1847) );
AND2x2_ASAP7_75t_L g1857 ( .A(n_1692), .B(n_1851), .Y(n_1857) );
AND2x2_ASAP7_75t_L g1886 ( .A(n_1692), .B(n_1815), .Y(n_1886) );
AND2x2_ASAP7_75t_L g1889 ( .A(n_1692), .B(n_1777), .Y(n_1889) );
AND2x2_ASAP7_75t_L g1692 ( .A(n_1693), .B(n_1705), .Y(n_1692) );
AND2x4_ASAP7_75t_L g1694 ( .A(n_1695), .B(n_1700), .Y(n_1694) );
OAI21xp33_ASAP7_75t_SL g2029 ( .A1(n_1695), .A2(n_1991), .B(n_2030), .Y(n_2029) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
OR2x2_ASAP7_75t_L g1716 ( .A(n_1696), .B(n_1701), .Y(n_1716) );
NAND2xp5_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1699), .Y(n_1696) );
INVx1_ASAP7_75t_L g1697 ( .A(n_1698), .Y(n_1697) );
INVx1_ASAP7_75t_L g1708 ( .A(n_1699), .Y(n_1708) );
AND2x4_ASAP7_75t_L g1702 ( .A(n_1700), .B(n_1703), .Y(n_1702) );
INVx1_ASAP7_75t_L g1700 ( .A(n_1701), .Y(n_1700) );
OR2x2_ASAP7_75t_L g1718 ( .A(n_1701), .B(n_1704), .Y(n_1718) );
INVx1_ASAP7_75t_L g1703 ( .A(n_1704), .Y(n_1703) );
INVx1_ASAP7_75t_L g1727 ( .A(n_1706), .Y(n_1727) );
AND2x4_ASAP7_75t_L g1706 ( .A(n_1707), .B(n_1709), .Y(n_1706) );
AND2x2_ASAP7_75t_L g1751 ( .A(n_1707), .B(n_1709), .Y(n_1751) );
INVx1_ASAP7_75t_L g1707 ( .A(n_1708), .Y(n_1707) );
AND2x4_ASAP7_75t_L g1710 ( .A(n_1708), .B(n_1709), .Y(n_1710) );
INVx2_ASAP7_75t_L g1729 ( .A(n_1710), .Y(n_1729) );
AND2x2_ASAP7_75t_L g1773 ( .A(n_1711), .B(n_1759), .Y(n_1773) );
AND2x2_ASAP7_75t_L g1803 ( .A(n_1711), .B(n_1804), .Y(n_1803) );
NAND2xp5_ASAP7_75t_L g1823 ( .A(n_1711), .B(n_1824), .Y(n_1823) );
INVx1_ASAP7_75t_L g1904 ( .A(n_1711), .Y(n_1904) );
AND2x2_ASAP7_75t_L g1711 ( .A(n_1712), .B(n_1719), .Y(n_1711) );
AND2x2_ASAP7_75t_L g1765 ( .A(n_1712), .B(n_1766), .Y(n_1765) );
INVx2_ASAP7_75t_L g1778 ( .A(n_1712), .Y(n_1778) );
OAI22xp5_ASAP7_75t_L g1713 ( .A1(n_1714), .A2(n_1715), .B1(n_1717), .B2(n_1718), .Y(n_1713) );
OAI22xp33_ASAP7_75t_L g1720 ( .A1(n_1715), .A2(n_1718), .B1(n_1721), .B2(n_1722), .Y(n_1720) );
BUFx3_ASAP7_75t_L g1732 ( .A(n_1715), .Y(n_1732) );
OAI22xp33_ASAP7_75t_L g1739 ( .A1(n_1715), .A2(n_1740), .B1(n_1741), .B2(n_1742), .Y(n_1739) );
BUFx6f_ASAP7_75t_L g1715 ( .A(n_1716), .Y(n_1715) );
INVx1_ASAP7_75t_L g1735 ( .A(n_1718), .Y(n_1735) );
HB1xp67_ASAP7_75t_L g1742 ( .A(n_1718), .Y(n_1742) );
INVx1_ASAP7_75t_L g1766 ( .A(n_1719), .Y(n_1766) );
AND2x2_ASAP7_75t_L g1777 ( .A(n_1719), .B(n_1778), .Y(n_1777) );
INVx1_ASAP7_75t_L g1851 ( .A(n_1719), .Y(n_1851) );
INVx1_ASAP7_75t_L g1723 ( .A(n_1724), .Y(n_1723) );
AOI211xp5_ASAP7_75t_SL g1849 ( .A1(n_1724), .A2(n_1772), .B(n_1850), .C(n_1852), .Y(n_1849) );
NAND2xp5_ASAP7_75t_L g1724 ( .A(n_1725), .B(n_1736), .Y(n_1724) );
INVx1_ASAP7_75t_L g1825 ( .A(n_1725), .Y(n_1825) );
AND2x2_ASAP7_75t_L g1842 ( .A(n_1725), .B(n_1737), .Y(n_1842) );
NOR2xp33_ASAP7_75t_L g1848 ( .A(n_1725), .B(n_1736), .Y(n_1848) );
BUFx3_ASAP7_75t_L g1866 ( .A(n_1725), .Y(n_1866) );
INVx1_ASAP7_75t_L g1726 ( .A(n_1727), .Y(n_1726) );
INVx2_ASAP7_75t_L g1728 ( .A(n_1729), .Y(n_1728) );
OAI22xp33_ASAP7_75t_L g1730 ( .A1(n_1731), .A2(n_1732), .B1(n_1733), .B2(n_1734), .Y(n_1730) );
INVx1_ASAP7_75t_L g1925 ( .A(n_1732), .Y(n_1925) );
INVx1_ASAP7_75t_L g1734 ( .A(n_1735), .Y(n_1734) );
OAI211xp5_ASAP7_75t_L g1854 ( .A1(n_1736), .A2(n_1855), .B(n_1857), .C(n_1858), .Y(n_1854) );
OAI31xp33_ASAP7_75t_L g1901 ( .A1(n_1736), .A2(n_1806), .A3(n_1902), .B(n_1903), .Y(n_1901) );
NOR3xp33_ASAP7_75t_L g1920 ( .A(n_1736), .B(n_1852), .C(n_1862), .Y(n_1920) );
INVx2_ASAP7_75t_L g1736 ( .A(n_1737), .Y(n_1736) );
AND2x2_ASAP7_75t_L g1824 ( .A(n_1737), .B(n_1779), .Y(n_1824) );
INVx2_ASAP7_75t_L g1839 ( .A(n_1737), .Y(n_1839) );
INVx2_ASAP7_75t_L g1737 ( .A(n_1738), .Y(n_1737) );
INVx2_ASAP7_75t_SL g1788 ( .A(n_1738), .Y(n_1788) );
AND2x2_ASAP7_75t_L g1896 ( .A(n_1738), .B(n_1781), .Y(n_1896) );
OR2x2_ASAP7_75t_L g1900 ( .A(n_1738), .B(n_1755), .Y(n_1900) );
AOI22xp5_ASAP7_75t_L g1743 ( .A1(n_1744), .A2(n_1753), .B1(n_1767), .B2(n_1768), .Y(n_1743) );
NAND2xp5_ASAP7_75t_L g1796 ( .A(n_1744), .B(n_1793), .Y(n_1796) );
O2A1O1Ixp33_ASAP7_75t_L g1836 ( .A1(n_1744), .A2(n_1793), .B(n_1837), .C(n_1840), .Y(n_1836) );
AND2x2_ASAP7_75t_L g1744 ( .A(n_1745), .B(n_1749), .Y(n_1744) );
INVx1_ASAP7_75t_SL g1745 ( .A(n_1746), .Y(n_1745) );
CKINVDCx5p33_ASAP7_75t_R g1756 ( .A(n_1746), .Y(n_1756) );
AND2x2_ASAP7_75t_L g1779 ( .A(n_1746), .B(n_1749), .Y(n_1779) );
AND2x2_ASAP7_75t_L g1780 ( .A(n_1746), .B(n_1781), .Y(n_1780) );
INVx1_ASAP7_75t_L g1789 ( .A(n_1746), .Y(n_1789) );
AND2x2_ASAP7_75t_L g1801 ( .A(n_1746), .B(n_1793), .Y(n_1801) );
INVx1_ASAP7_75t_L g1853 ( .A(n_1746), .Y(n_1853) );
OR2x2_ASAP7_75t_L g1862 ( .A(n_1746), .B(n_1762), .Y(n_1862) );
INVx1_ASAP7_75t_L g1871 ( .A(n_1746), .Y(n_1871) );
NAND2xp5_ASAP7_75t_L g1887 ( .A(n_1746), .B(n_1791), .Y(n_1887) );
AND2x2_ASAP7_75t_L g1746 ( .A(n_1747), .B(n_1748), .Y(n_1746) );
CKINVDCx5p33_ASAP7_75t_R g1767 ( .A(n_1749), .Y(n_1767) );
CKINVDCx6p67_ASAP7_75t_R g1781 ( .A(n_1749), .Y(n_1781) );
AND2x2_ASAP7_75t_L g1787 ( .A(n_1749), .B(n_1788), .Y(n_1787) );
OAI32xp33_ASAP7_75t_L g1890 ( .A1(n_1749), .A2(n_1828), .A3(n_1866), .B1(n_1891), .B2(n_1892), .Y(n_1890) );
NAND2xp5_ASAP7_75t_L g1892 ( .A(n_1749), .B(n_1825), .Y(n_1892) );
OR2x6_ASAP7_75t_L g1749 ( .A(n_1750), .B(n_1752), .Y(n_1749) );
INVx1_ASAP7_75t_L g1753 ( .A(n_1754), .Y(n_1753) );
NOR2xp33_ASAP7_75t_L g1754 ( .A(n_1755), .B(n_1757), .Y(n_1754) );
NAND2xp5_ASAP7_75t_L g1822 ( .A(n_1755), .B(n_1788), .Y(n_1822) );
NAND3xp33_ASAP7_75t_L g1835 ( .A(n_1755), .B(n_1803), .C(n_1812), .Y(n_1835) );
INVx3_ASAP7_75t_L g1755 ( .A(n_1756), .Y(n_1755) );
AND2x2_ASAP7_75t_L g1769 ( .A(n_1756), .B(n_1770), .Y(n_1769) );
AND2x2_ASAP7_75t_L g1807 ( .A(n_1756), .B(n_1781), .Y(n_1807) );
NAND2xp5_ASAP7_75t_L g1817 ( .A(n_1756), .B(n_1812), .Y(n_1817) );
NOR2xp33_ASAP7_75t_L g1867 ( .A(n_1756), .B(n_1868), .Y(n_1867) );
OAI211xp5_ASAP7_75t_L g1861 ( .A1(n_1757), .A2(n_1862), .B(n_1863), .C(n_1864), .Y(n_1861) );
INVx1_ASAP7_75t_L g1757 ( .A(n_1758), .Y(n_1757) );
AND2x2_ASAP7_75t_L g1758 ( .A(n_1759), .B(n_1760), .Y(n_1758) );
OR2x2_ASAP7_75t_L g1775 ( .A(n_1759), .B(n_1776), .Y(n_1775) );
AND2x2_ASAP7_75t_L g1792 ( .A(n_1759), .B(n_1793), .Y(n_1792) );
NAND2xp5_ASAP7_75t_L g1850 ( .A(n_1759), .B(n_1851), .Y(n_1850) );
NAND2xp5_ASAP7_75t_L g1876 ( .A(n_1759), .B(n_1815), .Y(n_1876) );
INVx1_ASAP7_75t_L g1760 ( .A(n_1761), .Y(n_1760) );
NAND2xp5_ASAP7_75t_L g1761 ( .A(n_1762), .B(n_1765), .Y(n_1761) );
INVx3_ASAP7_75t_L g1772 ( .A(n_1762), .Y(n_1772) );
NAND2xp5_ASAP7_75t_L g1784 ( .A(n_1762), .B(n_1777), .Y(n_1784) );
INVx4_ASAP7_75t_L g1793 ( .A(n_1762), .Y(n_1793) );
AND2x2_ASAP7_75t_L g1804 ( .A(n_1762), .B(n_1799), .Y(n_1804) );
NAND2xp5_ASAP7_75t_L g1814 ( .A(n_1762), .B(n_1815), .Y(n_1814) );
NAND3xp33_ASAP7_75t_L g1841 ( .A(n_1762), .B(n_1780), .C(n_1842), .Y(n_1841) );
NOR2xp67_ASAP7_75t_SL g1915 ( .A(n_1762), .B(n_1798), .Y(n_1915) );
AND2x4_ASAP7_75t_L g1762 ( .A(n_1763), .B(n_1764), .Y(n_1762) );
AND2x2_ASAP7_75t_L g1791 ( .A(n_1765), .B(n_1792), .Y(n_1791) );
INVx1_ASAP7_75t_L g1795 ( .A(n_1765), .Y(n_1795) );
AND2x2_ASAP7_75t_L g1880 ( .A(n_1765), .B(n_1793), .Y(n_1880) );
NAND2xp5_ASAP7_75t_L g1909 ( .A(n_1765), .B(n_1804), .Y(n_1909) );
AND2x2_ASAP7_75t_L g1815 ( .A(n_1766), .B(n_1778), .Y(n_1815) );
INVx1_ASAP7_75t_L g1768 ( .A(n_1769), .Y(n_1768) );
OAI21xp5_ASAP7_75t_SL g1881 ( .A1(n_1769), .A2(n_1882), .B(n_1893), .Y(n_1881) );
O2A1O1Ixp33_ASAP7_75t_L g1894 ( .A1(n_1770), .A2(n_1895), .B(n_1896), .C(n_1897), .Y(n_1894) );
AND2x2_ASAP7_75t_L g1770 ( .A(n_1771), .B(n_1773), .Y(n_1770) );
OR2x2_ASAP7_75t_L g1870 ( .A(n_1771), .B(n_1856), .Y(n_1870) );
INVx2_ASAP7_75t_L g1771 ( .A(n_1772), .Y(n_1771) );
NAND2xp5_ASAP7_75t_L g1776 ( .A(n_1772), .B(n_1777), .Y(n_1776) );
NOR2xp33_ASAP7_75t_L g1818 ( .A(n_1772), .B(n_1819), .Y(n_1818) );
OR2x2_ASAP7_75t_L g1875 ( .A(n_1772), .B(n_1876), .Y(n_1875) );
AOI21xp5_ASAP7_75t_L g1774 ( .A1(n_1775), .A2(n_1779), .B(n_1780), .Y(n_1774) );
INVx1_ASAP7_75t_L g1811 ( .A(n_1775), .Y(n_1811) );
INVx1_ASAP7_75t_L g1891 ( .A(n_1776), .Y(n_1891) );
INVx1_ASAP7_75t_L g1830 ( .A(n_1777), .Y(n_1830) );
NAND2xp5_ASAP7_75t_L g1798 ( .A(n_1778), .B(n_1799), .Y(n_1798) );
INVx2_ASAP7_75t_L g1820 ( .A(n_1778), .Y(n_1820) );
NOR2xp33_ASAP7_75t_L g1833 ( .A(n_1778), .B(n_1799), .Y(n_1833) );
NAND2xp5_ASAP7_75t_L g1888 ( .A(n_1779), .B(n_1889), .Y(n_1888) );
AOI211xp5_ASAP7_75t_L g1790 ( .A1(n_1780), .A2(n_1791), .B(n_1794), .C(n_1797), .Y(n_1790) );
NAND2xp5_ASAP7_75t_L g1802 ( .A(n_1780), .B(n_1803), .Y(n_1802) );
NAND2xp5_ASAP7_75t_L g1883 ( .A(n_1780), .B(n_1884), .Y(n_1883) );
AND2x4_ASAP7_75t_SL g1812 ( .A(n_1781), .B(n_1788), .Y(n_1812) );
NOR2xp33_ASAP7_75t_L g1864 ( .A(n_1781), .B(n_1865), .Y(n_1864) );
NAND2xp5_ASAP7_75t_L g1873 ( .A(n_1781), .B(n_1866), .Y(n_1873) );
OR2x2_ASAP7_75t_L g1911 ( .A(n_1781), .B(n_1788), .Y(n_1911) );
O2A1O1Ixp33_ASAP7_75t_L g1782 ( .A1(n_1783), .A2(n_1805), .B(n_1825), .C(n_1826), .Y(n_1782) );
OAI211xp5_ASAP7_75t_SL g1783 ( .A1(n_1784), .A2(n_1785), .B(n_1790), .C(n_1802), .Y(n_1783) );
OR2x2_ASAP7_75t_L g1868 ( .A(n_1784), .B(n_1799), .Y(n_1868) );
AOI21xp5_ASAP7_75t_L g1921 ( .A1(n_1784), .A2(n_1822), .B(n_1922), .Y(n_1921) );
INVx1_ASAP7_75t_L g1785 ( .A(n_1786), .Y(n_1785) );
AND2x2_ASAP7_75t_L g1786 ( .A(n_1787), .B(n_1789), .Y(n_1786) );
INVx2_ASAP7_75t_L g1843 ( .A(n_1787), .Y(n_1843) );
OAI221xp5_ASAP7_75t_L g1898 ( .A1(n_1791), .A2(n_1822), .B1(n_1899), .B2(n_1900), .C(n_1901), .Y(n_1898) );
NAND2xp5_ASAP7_75t_L g1844 ( .A(n_1792), .B(n_1815), .Y(n_1844) );
INVx1_ASAP7_75t_L g1832 ( .A(n_1793), .Y(n_1832) );
NOR2xp33_ASAP7_75t_L g1794 ( .A(n_1795), .B(n_1796), .Y(n_1794) );
INVx1_ASAP7_75t_L g1858 ( .A(n_1796), .Y(n_1858) );
NOR2xp33_ASAP7_75t_L g1797 ( .A(n_1798), .B(n_1800), .Y(n_1797) );
NAND2xp5_ASAP7_75t_L g1819 ( .A(n_1799), .B(n_1820), .Y(n_1819) );
OR2x2_ASAP7_75t_L g1829 ( .A(n_1799), .B(n_1830), .Y(n_1829) );
OR2x2_ASAP7_75t_L g1856 ( .A(n_1799), .B(n_1851), .Y(n_1856) );
AND2x2_ASAP7_75t_L g1923 ( .A(n_1799), .B(n_1880), .Y(n_1923) );
INVx1_ASAP7_75t_L g1800 ( .A(n_1801), .Y(n_1800) );
INVx1_ASAP7_75t_L g1902 ( .A(n_1804), .Y(n_1902) );
OAI211xp5_ASAP7_75t_L g1805 ( .A1(n_1806), .A2(n_1808), .B(n_1810), .C(n_1823), .Y(n_1805) );
INVx1_ASAP7_75t_L g1806 ( .A(n_1807), .Y(n_1806) );
OAI21xp5_ASAP7_75t_L g1878 ( .A1(n_1807), .A2(n_1879), .B(n_1880), .Y(n_1878) );
INVx1_ASAP7_75t_L g1808 ( .A(n_1809), .Y(n_1808) );
AOI222xp33_ASAP7_75t_L g1810 ( .A1(n_1811), .A2(n_1812), .B1(n_1813), .B2(n_1816), .C1(n_1818), .C2(n_1821), .Y(n_1810) );
INVx1_ASAP7_75t_L g1918 ( .A(n_1812), .Y(n_1918) );
A2O1A1Ixp33_ASAP7_75t_L g1905 ( .A1(n_1813), .A2(n_1866), .B(n_1906), .C(n_1910), .Y(n_1905) );
INVx1_ASAP7_75t_L g1813 ( .A(n_1814), .Y(n_1813) );
INVx1_ASAP7_75t_L g1852 ( .A(n_1815), .Y(n_1852) );
INVx1_ASAP7_75t_L g1816 ( .A(n_1817), .Y(n_1816) );
OAI22xp33_ASAP7_75t_L g1840 ( .A1(n_1820), .A2(n_1841), .B1(n_1843), .B2(n_1844), .Y(n_1840) );
INVx1_ASAP7_75t_L g1821 ( .A(n_1822), .Y(n_1821) );
O2A1O1Ixp33_ASAP7_75t_SL g1827 ( .A1(n_1824), .A2(n_1828), .B(n_1831), .C(n_1834), .Y(n_1827) );
NAND4xp25_ASAP7_75t_L g1826 ( .A(n_1827), .B(n_1836), .C(n_1845), .D(n_1854), .Y(n_1826) );
INVx1_ASAP7_75t_L g1828 ( .A(n_1829), .Y(n_1828) );
AND2x2_ASAP7_75t_L g1831 ( .A(n_1832), .B(n_1833), .Y(n_1831) );
INVxp67_ASAP7_75t_SL g1834 ( .A(n_1835), .Y(n_1834) );
INVx1_ASAP7_75t_L g1837 ( .A(n_1838), .Y(n_1837) );
OAI211xp5_ASAP7_75t_L g1913 ( .A1(n_1843), .A2(n_1914), .B(n_1916), .C(n_1919), .Y(n_1913) );
INVx1_ASAP7_75t_L g1899 ( .A(n_1844), .Y(n_1899) );
A2O1A1Ixp33_ASAP7_75t_L g1845 ( .A1(n_1846), .A2(n_1848), .B(n_1849), .C(n_1853), .Y(n_1845) );
INVx1_ASAP7_75t_L g1846 ( .A(n_1847), .Y(n_1846) );
NAND2xp5_ASAP7_75t_L g1884 ( .A(n_1847), .B(n_1885), .Y(n_1884) );
INVxp67_ASAP7_75t_L g1893 ( .A(n_1848), .Y(n_1893) );
NAND2xp5_ASAP7_75t_L g1903 ( .A(n_1852), .B(n_1904), .Y(n_1903) );
INVx1_ASAP7_75t_L g1907 ( .A(n_1853), .Y(n_1907) );
INVx1_ASAP7_75t_L g1855 ( .A(n_1856), .Y(n_1855) );
OAI211xp5_ASAP7_75t_L g1859 ( .A1(n_1860), .A2(n_1881), .B(n_1894), .C(n_1912), .Y(n_1859) );
O2A1O1Ixp33_ASAP7_75t_SL g1860 ( .A1(n_1861), .A2(n_1867), .B(n_1869), .C(n_1874), .Y(n_1860) );
INVx2_ASAP7_75t_L g1865 ( .A(n_1866), .Y(n_1865) );
OAI21xp5_ASAP7_75t_L g1912 ( .A1(n_1866), .A2(n_1913), .B(n_1921), .Y(n_1912) );
OAI21xp33_ASAP7_75t_L g1869 ( .A1(n_1870), .A2(n_1871), .B(n_1872), .Y(n_1869) );
NOR2xp33_ASAP7_75t_L g1917 ( .A(n_1870), .B(n_1918), .Y(n_1917) );
INVx1_ASAP7_75t_L g1877 ( .A(n_1871), .Y(n_1877) );
INVxp33_ASAP7_75t_L g1872 ( .A(n_1873), .Y(n_1872) );
OAI21xp5_ASAP7_75t_L g1874 ( .A1(n_1875), .A2(n_1877), .B(n_1878), .Y(n_1874) );
INVx1_ASAP7_75t_L g1879 ( .A(n_1876), .Y(n_1879) );
NAND4xp25_ASAP7_75t_L g1882 ( .A(n_1883), .B(n_1887), .C(n_1888), .D(n_1890), .Y(n_1882) );
INVx1_ASAP7_75t_L g1885 ( .A(n_1886), .Y(n_1885) );
INVx1_ASAP7_75t_L g1895 ( .A(n_1887), .Y(n_1895) );
NAND2xp5_ASAP7_75t_L g1897 ( .A(n_1898), .B(n_1905), .Y(n_1897) );
AND2x2_ASAP7_75t_L g1906 ( .A(n_1907), .B(n_1908), .Y(n_1906) );
INVx1_ASAP7_75t_L g1908 ( .A(n_1909), .Y(n_1908) );
INVx1_ASAP7_75t_L g1910 ( .A(n_1911), .Y(n_1910) );
INVx1_ASAP7_75t_L g1914 ( .A(n_1915), .Y(n_1914) );
INVxp67_ASAP7_75t_SL g1916 ( .A(n_1917), .Y(n_1916) );
INVxp67_ASAP7_75t_SL g1919 ( .A(n_1920), .Y(n_1919) );
INVx1_ASAP7_75t_L g1922 ( .A(n_1923), .Y(n_1922) );
CKINVDCx16_ASAP7_75t_R g1924 ( .A(n_1925), .Y(n_1924) );
INVx1_ASAP7_75t_L g1926 ( .A(n_1927), .Y(n_1926) );
XNOR2x1_ASAP7_75t_SL g1927 ( .A(n_1928), .B(n_1929), .Y(n_1927) );
AND2x2_ASAP7_75t_L g1929 ( .A(n_1930), .B(n_1959), .Y(n_1929) );
NOR3xp33_ASAP7_75t_SL g1930 ( .A(n_1931), .B(n_1939), .C(n_1941), .Y(n_1930) );
NAND2xp5_ASAP7_75t_L g1931 ( .A(n_1932), .B(n_1936), .Y(n_1931) );
OAI221xp5_ASAP7_75t_L g1970 ( .A1(n_1935), .A2(n_1937), .B1(n_1971), .B2(n_1972), .C(n_1973), .Y(n_1970) );
INVx3_ASAP7_75t_L g1944 ( .A(n_1945), .Y(n_1944) );
INVx1_ASAP7_75t_L g1950 ( .A(n_1951), .Y(n_1950) );
NAND3xp33_ASAP7_75t_L g1960 ( .A(n_1961), .B(n_1975), .C(n_1981), .Y(n_1960) );
INVx3_ASAP7_75t_L g1964 ( .A(n_1965), .Y(n_1964) );
INVx1_ASAP7_75t_L g1967 ( .A(n_1968), .Y(n_1967) );
INVx1_ASAP7_75t_L g1973 ( .A(n_1974), .Y(n_1973) );
INVx1_ASAP7_75t_L g1978 ( .A(n_1979), .Y(n_1978) );
INVx4_ASAP7_75t_SL g1983 ( .A(n_1984), .Y(n_1983) );
BUFx3_ASAP7_75t_L g1984 ( .A(n_1985), .Y(n_1984) );
BUFx2_ASAP7_75t_L g1985 ( .A(n_1986), .Y(n_1985) );
INVx2_ASAP7_75t_L g1988 ( .A(n_1989), .Y(n_1988) );
CKINVDCx5p33_ASAP7_75t_R g1989 ( .A(n_1990), .Y(n_1989) );
INVxp33_ASAP7_75t_L g1992 ( .A(n_1993), .Y(n_1992) );
HB1xp67_ASAP7_75t_L g1994 ( .A(n_1995), .Y(n_1994) );
AND4x1_ASAP7_75t_L g1995 ( .A(n_1996), .B(n_1998), .C(n_2009), .D(n_2025), .Y(n_1995) );
NOR2xp33_ASAP7_75t_L g2025 ( .A(n_2026), .B(n_2027), .Y(n_2025) );
HB1xp67_ASAP7_75t_L g2028 ( .A(n_2029), .Y(n_2028) );
endmodule