module fake_netlist_1_1372_n_636 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_636);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_636;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_446;
wire n_342;
wire n_423;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_261;
wire n_110;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_60), .Y(n_73) );
BUFx3_ASAP7_75t_L g74 ( .A(n_49), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_19), .Y(n_75) );
CKINVDCx5p33_ASAP7_75t_R g76 ( .A(n_57), .Y(n_76) );
INVx2_ASAP7_75t_L g77 ( .A(n_62), .Y(n_77) );
INVxp67_ASAP7_75t_SL g78 ( .A(n_56), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_43), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_28), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_47), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_46), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_55), .Y(n_83) );
INVxp67_ASAP7_75t_L g84 ( .A(n_22), .Y(n_84) );
INVxp67_ASAP7_75t_SL g85 ( .A(n_29), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_14), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_13), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_59), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_6), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_34), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_20), .Y(n_91) );
INVxp33_ASAP7_75t_SL g92 ( .A(n_1), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_36), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_61), .Y(n_94) );
INVx2_ASAP7_75t_SL g95 ( .A(n_45), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_53), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_13), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_21), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_58), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_69), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_41), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_10), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_48), .Y(n_103) );
CKINVDCx16_ASAP7_75t_R g104 ( .A(n_31), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_65), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_6), .Y(n_106) );
INVxp67_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_5), .Y(n_108) );
CKINVDCx20_ASAP7_75t_R g109 ( .A(n_24), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_35), .Y(n_110) );
BUFx3_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_4), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_11), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_7), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_3), .Y(n_115) );
INVxp33_ASAP7_75t_L g116 ( .A(n_70), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_14), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_2), .Y(n_118) );
BUFx6f_ASAP7_75t_L g119 ( .A(n_74), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_79), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_79), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_104), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_109), .Y(n_123) );
BUFx6f_ASAP7_75t_L g124 ( .A(n_74), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_80), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_109), .Y(n_126) );
INVx3_ASAP7_75t_L g127 ( .A(n_111), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_80), .Y(n_128) );
BUFx3_ASAP7_75t_L g129 ( .A(n_95), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_76), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_76), .Y(n_131) );
NOR2xp33_ASAP7_75t_R g132 ( .A(n_81), .B(n_33), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g133 ( .A(n_81), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_82), .Y(n_134) );
AND2x2_ASAP7_75t_L g135 ( .A(n_113), .B(n_0), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
BUFx2_ASAP7_75t_L g137 ( .A(n_113), .Y(n_137) );
INVx2_ASAP7_75t_L g138 ( .A(n_77), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g139 ( .A(n_111), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_83), .Y(n_140) );
HB1xp67_ASAP7_75t_L g141 ( .A(n_86), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_83), .Y(n_142) );
BUFx2_ASAP7_75t_L g143 ( .A(n_86), .Y(n_143) );
INVx3_ASAP7_75t_L g144 ( .A(n_88), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_88), .Y(n_145) );
OR2x2_ASAP7_75t_L g146 ( .A(n_87), .B(n_0), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_95), .B(n_1), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_77), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_73), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_92), .Y(n_150) );
AND2x2_ASAP7_75t_L g151 ( .A(n_116), .B(n_3), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_100), .Y(n_152) );
BUFx6f_ASAP7_75t_L g153 ( .A(n_100), .Y(n_153) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_75), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g155 ( .A(n_87), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_89), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_92), .Y(n_157) );
BUFx6f_ASAP7_75t_L g158 ( .A(n_90), .Y(n_158) );
INVx2_ASAP7_75t_L g159 ( .A(n_91), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_153), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_156), .Y(n_161) );
AND2x4_ASAP7_75t_L g162 ( .A(n_143), .B(n_118), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_137), .B(n_107), .Y(n_163) );
AND2x2_ASAP7_75t_L g164 ( .A(n_137), .B(n_118), .Y(n_164) );
AND2x2_ASAP7_75t_L g165 ( .A(n_143), .B(n_117), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_153), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_156), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_156), .Y(n_169) );
INVx2_ASAP7_75t_SL g170 ( .A(n_129), .Y(n_170) );
BUFx3_ASAP7_75t_L g171 ( .A(n_129), .Y(n_171) );
NAND3x1_ASAP7_75t_L g172 ( .A(n_135), .B(n_117), .C(n_115), .Y(n_172) );
HB1xp67_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_153), .Y(n_175) );
BUFx3_ASAP7_75t_L g176 ( .A(n_129), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_153), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_144), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_131), .B(n_84), .Y(n_179) );
HB1xp67_ASAP7_75t_L g180 ( .A(n_133), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_119), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_144), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_144), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_149), .B(n_101), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_119), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_135), .B(n_115), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_141), .B(n_89), .Y(n_188) );
INVx1_ASAP7_75t_L g189 ( .A(n_154), .Y(n_189) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_119), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_154), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_154), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_120), .B(n_114), .Y(n_193) );
AND2x4_ASAP7_75t_L g194 ( .A(n_120), .B(n_112), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_149), .B(n_98), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_154), .Y(n_196) );
AND2x4_ASAP7_75t_L g197 ( .A(n_121), .B(n_102), .Y(n_197) );
BUFx2_ASAP7_75t_L g198 ( .A(n_139), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_151), .B(n_97), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_119), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_121), .B(n_99), .Y(n_201) );
NOR2x1p5_ASAP7_75t_L g202 ( .A(n_122), .B(n_106), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_119), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_124), .Y(n_204) );
INVx2_ASAP7_75t_L g205 ( .A(n_124), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_124), .Y(n_206) );
INVx2_ASAP7_75t_L g207 ( .A(n_124), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_124), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_154), .Y(n_209) );
INVx1_ASAP7_75t_L g210 ( .A(n_158), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_158), .Y(n_211) );
AO22x2_ASAP7_75t_L g212 ( .A1(n_146), .A2(n_108), .B1(n_96), .B2(n_105), .Y(n_212) );
OR2x2_ASAP7_75t_L g213 ( .A(n_146), .B(n_4), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_158), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_158), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_158), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_162), .B(n_151), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_162), .B(n_134), .Y(n_218) );
AND2x2_ASAP7_75t_SL g219 ( .A(n_213), .B(n_134), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_162), .B(n_159), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_213), .Y(n_221) );
OAI21xp5_ASAP7_75t_L g222 ( .A1(n_178), .A2(n_145), .B(n_128), .Y(n_222) );
NOR2xp33_ASAP7_75t_R g223 ( .A(n_173), .B(n_123), .Y(n_223) );
HB1xp67_ASAP7_75t_L g224 ( .A(n_162), .Y(n_224) );
INVx3_ASAP7_75t_L g225 ( .A(n_171), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_187), .B(n_159), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_198), .Y(n_227) );
CKINVDCx5p33_ASAP7_75t_R g228 ( .A(n_198), .Y(n_228) );
BUFx2_ASAP7_75t_L g229 ( .A(n_180), .Y(n_229) );
BUFx2_ASAP7_75t_L g230 ( .A(n_212), .Y(n_230) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_202), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_161), .Y(n_232) );
INVx5_ASAP7_75t_L g233 ( .A(n_214), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_164), .B(n_157), .Y(n_234) );
NOR3xp33_ASAP7_75t_SL g235 ( .A(n_163), .B(n_126), .C(n_150), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_161), .Y(n_236) );
AND2x2_ASAP7_75t_L g237 ( .A(n_164), .B(n_155), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_168), .Y(n_238) );
HB1xp67_ASAP7_75t_L g239 ( .A(n_188), .Y(n_239) );
INVx1_ASAP7_75t_SL g240 ( .A(n_188), .Y(n_240) );
OR2x6_ASAP7_75t_L g241 ( .A(n_172), .B(n_147), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_168), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_169), .Y(n_243) );
NAND2xp33_ASAP7_75t_L g244 ( .A(n_172), .B(n_132), .Y(n_244) );
CKINVDCx6p67_ASAP7_75t_R g245 ( .A(n_187), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_187), .B(n_125), .Y(n_246) );
NAND2xp33_ASAP7_75t_SL g247 ( .A(n_202), .B(n_136), .Y(n_247) );
INVx5_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_171), .Y(n_249) );
AND2x6_ASAP7_75t_L g250 ( .A(n_187), .B(n_125), .Y(n_250) );
INVxp67_ASAP7_75t_L g251 ( .A(n_165), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_169), .Y(n_252) );
CKINVDCx5p33_ASAP7_75t_R g253 ( .A(n_179), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_165), .Y(n_254) );
AOI22xp5_ASAP7_75t_L g255 ( .A1(n_212), .A2(n_128), .B1(n_145), .B2(n_142), .Y(n_255) );
INVx2_ASAP7_75t_L g256 ( .A(n_174), .Y(n_256) );
BUFx6f_ASAP7_75t_L g257 ( .A(n_181), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_212), .Y(n_258) );
BUFx2_ASAP7_75t_SL g259 ( .A(n_212), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_199), .B(n_197), .Y(n_260) );
BUFx8_ASAP7_75t_L g261 ( .A(n_199), .Y(n_261) );
HB1xp67_ASAP7_75t_L g262 ( .A(n_197), .Y(n_262) );
BUFx12f_ASAP7_75t_L g263 ( .A(n_193), .Y(n_263) );
NOR2xp33_ASAP7_75t_R g264 ( .A(n_170), .B(n_127), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_193), .B(n_136), .Y(n_265) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_197), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_193), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_174), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_193), .B(n_142), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_194), .B(n_140), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_178), .Y(n_271) );
BUFx2_ASAP7_75t_L g272 ( .A(n_176), .Y(n_272) );
HB1xp67_ASAP7_75t_L g273 ( .A(n_194), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_182), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_176), .Y(n_275) );
INVx3_ASAP7_75t_L g276 ( .A(n_170), .Y(n_276) );
NAND2xp5_ASAP7_75t_SL g277 ( .A(n_182), .B(n_183), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_262), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_273), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_250), .Y(n_280) );
NOR2x1_ASAP7_75t_SL g281 ( .A(n_263), .B(n_201), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_224), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_263), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_240), .B(n_194), .Y(n_284) );
NOR2xp67_ASAP7_75t_L g285 ( .A(n_231), .B(n_195), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_260), .Y(n_286) );
INVx5_ASAP7_75t_L g287 ( .A(n_250), .Y(n_287) );
INVx2_ASAP7_75t_SL g288 ( .A(n_250), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_217), .B(n_194), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_226), .Y(n_290) );
NAND2xp5_ASAP7_75t_SL g291 ( .A(n_255), .B(n_183), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_236), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_250), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_217), .B(n_185), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_226), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_217), .B(n_184), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_267), .B(n_184), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_219), .A2(n_140), .B1(n_127), .B2(n_138), .Y(n_298) );
INVx2_ASAP7_75t_L g299 ( .A(n_236), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_252), .Y(n_300) );
BUFx2_ASAP7_75t_L g301 ( .A(n_261), .Y(n_301) );
BUFx3_ASAP7_75t_L g302 ( .A(n_250), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g303 ( .A1(n_259), .A2(n_127), .B1(n_148), .B2(n_138), .Y(n_303) );
INVx2_ASAP7_75t_L g304 ( .A(n_252), .Y(n_304) );
INVxp67_ASAP7_75t_SL g305 ( .A(n_261), .Y(n_305) );
A2O1A1Ixp33_ASAP7_75t_L g306 ( .A1(n_222), .A2(n_152), .B(n_148), .C(n_127), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_226), .Y(n_307) );
INVx3_ASAP7_75t_L g308 ( .A(n_225), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_270), .Y(n_309) );
AOI21xp5_ASAP7_75t_L g310 ( .A1(n_277), .A2(n_196), .B(n_215), .Y(n_310) );
BUFx6f_ASAP7_75t_L g311 ( .A(n_257), .Y(n_311) );
CKINVDCx8_ASAP7_75t_R g312 ( .A(n_229), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_230), .B(n_258), .Y(n_313) );
BUFx12f_ASAP7_75t_L g314 ( .A(n_261), .Y(n_314) );
INVx5_ASAP7_75t_L g315 ( .A(n_225), .Y(n_315) );
CKINVDCx20_ASAP7_75t_R g316 ( .A(n_223), .Y(n_316) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_266), .A2(n_78), .B1(n_110), .B2(n_85), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_219), .A2(n_152), .B1(n_94), .B2(n_103), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_220), .Y(n_319) );
AND2x4_ASAP7_75t_L g320 ( .A(n_220), .B(n_93), .Y(n_320) );
INVx2_ASAP7_75t_SL g321 ( .A(n_245), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_256), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_220), .B(n_5), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_246), .Y(n_324) );
NOR2xp33_ASAP7_75t_L g325 ( .A(n_312), .B(n_254), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_280), .B(n_221), .Y(n_326) );
BUFx10_ASAP7_75t_L g327 ( .A(n_321), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_292), .Y(n_328) );
AOI22xp33_ASAP7_75t_L g329 ( .A1(n_286), .A2(n_254), .B1(n_234), .B2(n_237), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_284), .B(n_239), .Y(n_330) );
INVx3_ASAP7_75t_L g331 ( .A(n_280), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_324), .B(n_251), .Y(n_332) );
O2A1O1Ixp33_ASAP7_75t_L g333 ( .A1(n_318), .A2(n_244), .B(n_218), .C(n_241), .Y(n_333) );
CKINVDCx20_ASAP7_75t_R g334 ( .A(n_312), .Y(n_334) );
INVx4_ASAP7_75t_L g335 ( .A(n_280), .Y(n_335) );
BUFx3_ASAP7_75t_L g336 ( .A(n_280), .Y(n_336) );
NAND2xp33_ASAP7_75t_SL g337 ( .A(n_288), .B(n_223), .Y(n_337) );
AOI221xp5_ASAP7_75t_L g338 ( .A1(n_309), .A2(n_247), .B1(n_227), .B2(n_228), .C(n_253), .Y(n_338) );
AOI22xp33_ASAP7_75t_L g339 ( .A1(n_313), .A2(n_241), .B1(n_247), .B2(n_244), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_313), .B(n_265), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_292), .Y(n_341) );
AOI22xp33_ASAP7_75t_L g342 ( .A1(n_313), .A2(n_241), .B1(n_253), .B2(n_228), .Y(n_342) );
AND2x4_ASAP7_75t_L g343 ( .A(n_287), .B(n_269), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_313), .A2(n_227), .B1(n_272), .B2(n_243), .Y(n_344) );
CKINVDCx6p67_ASAP7_75t_R g345 ( .A(n_314), .Y(n_345) );
AOI22xp33_ASAP7_75t_L g346 ( .A1(n_282), .A2(n_238), .B1(n_232), .B2(n_242), .Y(n_346) );
INVx4_ASAP7_75t_SL g347 ( .A(n_293), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_299), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_299), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_298), .A2(n_275), .B1(n_268), .B2(n_274), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_300), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_294), .B(n_275), .Y(n_352) );
AOI21xp5_ASAP7_75t_L g353 ( .A1(n_291), .A2(n_277), .B(n_274), .Y(n_353) );
BUFx8_ASAP7_75t_L g354 ( .A(n_314), .Y(n_354) );
OAI21xp33_ASAP7_75t_L g355 ( .A1(n_329), .A2(n_235), .B(n_297), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_332), .B(n_290), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_341), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_325), .A2(n_316), .B1(n_301), .B2(n_320), .Y(n_358) );
AOI221xp5_ASAP7_75t_L g359 ( .A1(n_332), .A2(n_289), .B1(n_278), .B2(n_295), .C(n_307), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_330), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_334), .A2(n_316), .B1(n_305), .B2(n_287), .Y(n_361) );
BUFx3_ASAP7_75t_L g362 ( .A(n_354), .Y(n_362) );
INVx1_ASAP7_75t_SL g363 ( .A(n_345), .Y(n_363) );
OAI22xp5_ASAP7_75t_L g364 ( .A1(n_350), .A2(n_303), .B1(n_302), .B2(n_293), .Y(n_364) );
OAI221xp5_ASAP7_75t_L g365 ( .A1(n_338), .A2(n_317), .B1(n_285), .B2(n_297), .C(n_321), .Y(n_365) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_340), .A2(n_320), .B1(n_323), .B2(n_279), .Y(n_366) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_333), .A2(n_303), .B(n_320), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_283), .B1(n_319), .B2(n_296), .C(n_306), .Y(n_368) );
BUFx12f_ASAP7_75t_L g369 ( .A(n_354), .Y(n_369) );
AOI22xp33_ASAP7_75t_SL g370 ( .A1(n_354), .A2(n_281), .B1(n_302), .B2(n_283), .Y(n_370) );
AOI221xp5_ASAP7_75t_L g371 ( .A1(n_330), .A2(n_306), .B1(n_291), .B2(n_300), .C(n_304), .Y(n_371) );
BUFx2_ASAP7_75t_L g372 ( .A(n_354), .Y(n_372) );
OAI211xp5_ASAP7_75t_SL g373 ( .A1(n_344), .A2(n_308), .B(n_189), .C(n_211), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_340), .B(n_304), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g375 ( .A1(n_339), .A2(n_287), .B1(n_288), .B2(n_308), .Y(n_375) );
OAI221xp5_ASAP7_75t_L g376 ( .A1(n_352), .A2(n_308), .B1(n_322), .B2(n_287), .C(n_276), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_346), .B(n_322), .Y(n_377) );
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_326), .A2(n_225), .B1(n_249), .B2(n_315), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_350), .A2(n_315), .B1(n_249), .B2(n_276), .Y(n_379) );
BUFx5_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
OAI22xp5_ASAP7_75t_L g381 ( .A1(n_328), .A2(n_315), .B1(n_249), .B2(n_276), .Y(n_381) );
HB1xp67_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_357), .Y(n_383) );
AND2x2_ASAP7_75t_L g384 ( .A(n_374), .B(n_328), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_377), .Y(n_385) );
NAND3xp33_ASAP7_75t_L g386 ( .A(n_355), .B(n_337), .C(n_349), .Y(n_386) );
INVx2_ASAP7_75t_L g387 ( .A(n_380), .Y(n_387) );
AOI22xp33_ASAP7_75t_L g388 ( .A1(n_365), .A2(n_326), .B1(n_343), .B2(n_345), .Y(n_388) );
AO21x2_ASAP7_75t_L g389 ( .A1(n_367), .A2(n_353), .B(n_349), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_360), .Y(n_390) );
OAI221xp5_ASAP7_75t_SL g391 ( .A1(n_358), .A2(n_351), .B1(n_348), .B2(n_341), .C(n_310), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_356), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_380), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_380), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_380), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_366), .B(n_348), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_380), .Y(n_397) );
INVx3_ASAP7_75t_SL g398 ( .A(n_362), .Y(n_398) );
INVx3_ASAP7_75t_L g399 ( .A(n_380), .Y(n_399) );
AND2x2_ASAP7_75t_L g400 ( .A(n_371), .B(n_351), .Y(n_400) );
AOI31xp33_ASAP7_75t_L g401 ( .A1(n_370), .A2(n_326), .A3(n_343), .B(n_327), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_379), .Y(n_402) );
OAI31xp33_ASAP7_75t_L g403 ( .A1(n_373), .A2(n_326), .A3(n_343), .B(n_336), .Y(n_403) );
OR2x2_ASAP7_75t_L g404 ( .A(n_372), .B(n_343), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_368), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_381), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_364), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_359), .B(n_331), .Y(n_408) );
NOR4xp25_ASAP7_75t_L g409 ( .A(n_373), .B(n_203), .C(n_200), .D(n_186), .Y(n_409) );
AOI22xp33_ASAP7_75t_SL g410 ( .A1(n_369), .A2(n_336), .B1(n_335), .B2(n_331), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_370), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_378), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_361), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g415 ( .A1(n_363), .A2(n_331), .B1(n_335), .B2(n_315), .C(n_271), .Y(n_415) );
AND2x2_ASAP7_75t_SL g416 ( .A(n_412), .B(n_335), .Y(n_416) );
INVx2_ASAP7_75t_L g417 ( .A(n_383), .Y(n_417) );
INVx3_ASAP7_75t_L g418 ( .A(n_399), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_385), .B(n_375), .Y(n_419) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_398), .B(n_327), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_385), .B(n_331), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_383), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_384), .B(n_7), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_393), .Y(n_425) );
INVx2_ASAP7_75t_SL g426 ( .A(n_399), .Y(n_426) );
INVx1_ASAP7_75t_SL g427 ( .A(n_382), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_394), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_392), .B(n_327), .Y(n_429) );
NAND2xp33_ASAP7_75t_L g430 ( .A(n_398), .B(n_264), .Y(n_430) );
HB1xp67_ASAP7_75t_L g431 ( .A(n_384), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_394), .Y(n_432) );
HB1xp67_ASAP7_75t_L g433 ( .A(n_404), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_397), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_407), .B(n_8), .Y(n_435) );
OR2x2_ASAP7_75t_L g436 ( .A(n_407), .B(n_8), .Y(n_436) );
NAND2xp5_ASAP7_75t_SL g437 ( .A(n_412), .B(n_327), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_412), .B(n_9), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_397), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_387), .Y(n_440) );
INVx2_ASAP7_75t_SL g441 ( .A(n_399), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_387), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_390), .B(n_9), .Y(n_443) );
NAND3xp33_ASAP7_75t_SL g444 ( .A(n_388), .B(n_264), .C(n_335), .Y(n_444) );
AND2x4_ASAP7_75t_L g445 ( .A(n_412), .B(n_347), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_392), .B(n_10), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_395), .Y(n_447) );
OAI21x1_ASAP7_75t_L g448 ( .A1(n_399), .A2(n_204), .B(n_186), .Y(n_448) );
INVx2_ASAP7_75t_L g449 ( .A(n_395), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_390), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_400), .B(n_11), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_396), .B(n_12), .Y(n_452) );
OAI21xp5_ASAP7_75t_L g453 ( .A1(n_405), .A2(n_192), .B(n_196), .Y(n_453) );
BUFx3_ASAP7_75t_L g454 ( .A(n_404), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_400), .B(n_12), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_402), .B(n_204), .Y(n_456) );
AND2x4_ASAP7_75t_L g457 ( .A(n_402), .B(n_347), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_405), .B(n_347), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_406), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_408), .B(n_347), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_408), .B(n_205), .Y(n_461) );
OR2x2_ASAP7_75t_L g462 ( .A(n_396), .B(n_190), .Y(n_462) );
CKINVDCx16_ASAP7_75t_R g463 ( .A(n_398), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_450), .B(n_414), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_431), .B(n_413), .Y(n_465) );
BUFx2_ASAP7_75t_L g466 ( .A(n_463), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_454), .B(n_414), .Y(n_467) );
OR2x2_ASAP7_75t_L g468 ( .A(n_427), .B(n_413), .Y(n_468) );
OAI22xp5_ASAP7_75t_L g469 ( .A1(n_438), .A2(n_401), .B1(n_391), .B2(n_386), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_417), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_417), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_454), .B(n_389), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_450), .Y(n_473) );
NAND3xp33_ASAP7_75t_L g474 ( .A(n_438), .B(n_386), .C(n_403), .Y(n_474) );
OR2x2_ASAP7_75t_L g475 ( .A(n_427), .B(n_389), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g476 ( .A(n_463), .B(n_410), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_428), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_420), .Y(n_478) );
AOI22xp33_ASAP7_75t_L g479 ( .A1(n_451), .A2(n_411), .B1(n_389), .B2(n_415), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_428), .Y(n_480) );
INVx1_ASAP7_75t_SL g481 ( .A(n_424), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_433), .B(n_409), .Y(n_482) );
AND2x2_ASAP7_75t_L g483 ( .A(n_424), .B(n_411), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g484 ( .A(n_446), .B(n_15), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_416), .B(n_347), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_422), .B(n_190), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_430), .A2(n_315), .B1(n_271), .B2(n_256), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_452), .B(n_208), .Y(n_488) );
INVx1_ASAP7_75t_L g489 ( .A(n_432), .Y(n_489) );
NOR2x1_ASAP7_75t_L g490 ( .A(n_435), .B(n_203), .Y(n_490) );
NAND4xp25_ASAP7_75t_SL g491 ( .A(n_452), .B(n_16), .C(n_17), .D(n_18), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_422), .B(n_208), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_422), .B(n_190), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_432), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_423), .Y(n_495) );
AOI211xp5_ASAP7_75t_L g496 ( .A1(n_451), .A2(n_189), .B(n_191), .C(n_215), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_455), .B(n_25), .Y(n_497) );
NAND2x1_ASAP7_75t_L g498 ( .A(n_445), .B(n_181), .Y(n_498) );
AND2x2_ASAP7_75t_L g499 ( .A(n_443), .B(n_207), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_436), .B(n_190), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_455), .B(n_190), .Y(n_501) );
INVx1_ASAP7_75t_SL g502 ( .A(n_443), .Y(n_502) );
NOR2xp33_ASAP7_75t_L g503 ( .A(n_436), .B(n_181), .Y(n_503) );
AND2x4_ASAP7_75t_L g504 ( .A(n_445), .B(n_26), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_423), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_425), .B(n_181), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_425), .B(n_181), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_461), .B(n_206), .Y(n_508) );
INVx2_ASAP7_75t_SL g509 ( .A(n_429), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_425), .Y(n_510) );
HB1xp67_ASAP7_75t_L g511 ( .A(n_440), .Y(n_511) );
OR2x2_ASAP7_75t_L g512 ( .A(n_434), .B(n_205), .Y(n_512) );
BUFx2_ASAP7_75t_L g513 ( .A(n_445), .Y(n_513) );
INVx1_ASAP7_75t_SL g514 ( .A(n_416), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_481), .B(n_419), .Y(n_515) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_482), .A2(n_437), .B(n_458), .Y(n_516) );
AOI211x1_ASAP7_75t_L g517 ( .A1(n_469), .A2(n_491), .B(n_474), .C(n_485), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_465), .B(n_419), .Y(n_518) );
INVx2_ASAP7_75t_L g519 ( .A(n_511), .Y(n_519) );
OAI31xp33_ASAP7_75t_L g520 ( .A1(n_466), .A2(n_445), .A3(n_460), .B(n_457), .Y(n_520) );
AOI22xp5_ASAP7_75t_L g521 ( .A1(n_476), .A2(n_416), .B1(n_457), .B2(n_444), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_502), .B(n_439), .Y(n_522) );
NAND3xp33_ASAP7_75t_L g523 ( .A(n_475), .B(n_434), .C(n_439), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_473), .Y(n_524) );
OAI211xp5_ASAP7_75t_SL g525 ( .A1(n_478), .A2(n_421), .B(n_439), .C(n_434), .Y(n_525) );
AND2x2_ASAP7_75t_L g526 ( .A(n_467), .B(n_457), .Y(n_526) );
AND2x2_ASAP7_75t_SL g527 ( .A(n_504), .B(n_513), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_468), .B(n_421), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_477), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_480), .Y(n_530) );
AOI32xp33_ASAP7_75t_L g531 ( .A1(n_469), .A2(n_459), .A3(n_441), .B1(n_426), .B2(n_418), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_489), .Y(n_532) );
HB1xp67_ASAP7_75t_L g533 ( .A(n_511), .Y(n_533) );
OAI222xp33_ASAP7_75t_L g534 ( .A1(n_514), .A2(n_441), .B1(n_426), .B2(n_459), .C1(n_418), .C2(n_442), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_494), .Y(n_535) );
AOI31xp33_ASAP7_75t_L g536 ( .A1(n_479), .A2(n_447), .A3(n_440), .B(n_442), .Y(n_536) );
AND2x2_ASAP7_75t_SL g537 ( .A(n_504), .B(n_418), .Y(n_537) );
OAI22xp5_ASAP7_75t_L g538 ( .A1(n_490), .A2(n_440), .B1(n_442), .B2(n_449), .Y(n_538) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_497), .A2(n_491), .B1(n_483), .B2(n_509), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_464), .Y(n_540) );
AOI221xp5_ASAP7_75t_L g541 ( .A1(n_464), .A2(n_456), .B1(n_453), .B2(n_447), .C(n_449), .Y(n_541) );
AOI22xp5_ASAP7_75t_L g542 ( .A1(n_484), .A2(n_456), .B1(n_418), .B2(n_449), .Y(n_542) );
OAI22xp33_ASAP7_75t_SL g543 ( .A1(n_498), .A2(n_447), .B1(n_462), .B2(n_453), .Y(n_543) );
AOI21xp33_ASAP7_75t_SL g544 ( .A1(n_487), .A2(n_462), .B(n_30), .Y(n_544) );
NOR2xp33_ASAP7_75t_L g545 ( .A(n_488), .B(n_27), .Y(n_545) );
OAI31xp33_ASAP7_75t_L g546 ( .A1(n_479), .A2(n_200), .A3(n_175), .B(n_191), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_470), .B(n_448), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_505), .Y(n_548) );
INVxp67_ASAP7_75t_SL g549 ( .A(n_471), .Y(n_549) );
OAI221xp5_ASAP7_75t_L g550 ( .A1(n_496), .A2(n_210), .B1(n_192), .B2(n_211), .C(n_175), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_510), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_499), .B(n_32), .Y(n_552) );
NOR2xp33_ASAP7_75t_L g553 ( .A(n_501), .B(n_37), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_500), .A2(n_448), .B1(n_311), .B2(n_210), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_495), .B(n_177), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_486), .Y(n_556) );
OAI221xp5_ASAP7_75t_L g557 ( .A1(n_500), .A2(n_209), .B1(n_166), .B2(n_167), .C(n_177), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
OAI21xp5_ASAP7_75t_L g559 ( .A1(n_503), .A2(n_167), .B(n_166), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_472), .B(n_160), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_540), .B(n_508), .Y(n_561) );
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_539), .A2(n_507), .B1(n_506), .B2(n_493), .Y(n_562) );
BUFx3_ASAP7_75t_L g563 ( .A(n_522), .Y(n_563) );
INVxp67_ASAP7_75t_L g564 ( .A(n_533), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_518), .B(n_507), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_515), .B(n_512), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g567 ( .A(n_516), .B(n_493), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_524), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_529), .Y(n_569) );
OAI211xp5_ASAP7_75t_L g570 ( .A1(n_517), .A2(n_486), .B(n_492), .C(n_160), .Y(n_570) );
INVxp67_ASAP7_75t_SL g571 ( .A(n_549), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_530), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_526), .B(n_527), .Y(n_573) );
XOR2x2_ASAP7_75t_L g574 ( .A(n_537), .B(n_38), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_532), .Y(n_575) );
CKINVDCx16_ASAP7_75t_R g576 ( .A(n_521), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_535), .Y(n_577) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_543), .A2(n_311), .B(n_257), .Y(n_578) );
NAND4xp25_ASAP7_75t_L g579 ( .A(n_531), .B(n_209), .C(n_40), .D(n_42), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_528), .B(n_216), .Y(n_580) );
XNOR2x2_ASAP7_75t_L g581 ( .A(n_538), .B(n_39), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_558), .B(n_44), .Y(n_582) );
NOR2x1_ASAP7_75t_L g583 ( .A(n_525), .B(n_311), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_519), .B(n_216), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g585 ( .A1(n_542), .A2(n_216), .B1(n_214), .B2(n_257), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_548), .Y(n_586) );
NOR3xp33_ASAP7_75t_SL g587 ( .A(n_534), .B(n_50), .C(n_51), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_551), .B(n_216), .Y(n_588) );
AND2x2_ASAP7_75t_L g589 ( .A(n_520), .B(n_52), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g590 ( .A1(n_544), .A2(n_214), .B1(n_311), .B2(n_248), .Y(n_590) );
OR2x2_ASAP7_75t_L g591 ( .A(n_571), .B(n_523), .Y(n_591) );
O2A1O1Ixp33_ASAP7_75t_L g592 ( .A1(n_579), .A2(n_536), .B(n_538), .C(n_546), .Y(n_592) );
AOI222xp33_ASAP7_75t_L g593 ( .A1(n_564), .A2(n_541), .B1(n_556), .B2(n_560), .C1(n_545), .C2(n_553), .Y(n_593) );
NOR2x1_ASAP7_75t_L g594 ( .A(n_583), .B(n_570), .Y(n_594) );
NOR2xp33_ASAP7_75t_L g595 ( .A(n_576), .B(n_536), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_578), .A2(n_554), .B(n_559), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_571), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_586), .Y(n_598) );
INVx1_ASAP7_75t_SL g599 ( .A(n_563), .Y(n_599) );
AOI21xp33_ASAP7_75t_L g600 ( .A1(n_570), .A2(n_552), .B(n_547), .Y(n_600) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_578), .B(n_554), .Y(n_601) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_562), .A2(n_559), .B1(n_555), .B2(n_550), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_567), .B(n_214), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_567), .B(n_557), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_564), .B(n_54), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_568), .Y(n_606) );
OAI21xp33_ASAP7_75t_SL g607 ( .A1(n_573), .A2(n_63), .B(n_64), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_569), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_597), .Y(n_609) );
AND2x4_ASAP7_75t_L g610 ( .A(n_599), .B(n_577), .Y(n_610) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_594), .B(n_589), .Y(n_611) );
AOI221xp5_ASAP7_75t_L g612 ( .A1(n_595), .A2(n_602), .B1(n_604), .B2(n_606), .C(n_598), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_607), .A2(n_587), .B(n_574), .Y(n_613) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_591), .Y(n_614) );
OAI221xp5_ASAP7_75t_L g615 ( .A1(n_601), .A2(n_587), .B1(n_565), .B2(n_561), .C(n_572), .Y(n_615) );
OA22x2_ASAP7_75t_L g616 ( .A1(n_608), .A2(n_575), .B1(n_581), .B2(n_590), .Y(n_616) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_593), .A2(n_566), .B1(n_582), .B2(n_580), .Y(n_617) );
INVx1_ASAP7_75t_SL g618 ( .A(n_605), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g619 ( .A(n_603), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g620 ( .A1(n_592), .A2(n_585), .B1(n_588), .B2(n_584), .Y(n_620) );
AOI311xp33_ASAP7_75t_L g621 ( .A1(n_600), .A2(n_66), .A3(n_67), .B(n_68), .C(n_71), .Y(n_621) );
OAI22xp5_ASAP7_75t_L g622 ( .A1(n_592), .A2(n_233), .B1(n_248), .B2(n_72), .Y(n_622) );
AOI211xp5_ASAP7_75t_L g623 ( .A1(n_596), .A2(n_233), .B(n_248), .C(n_607), .Y(n_623) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_596), .B(n_517), .C(n_595), .D(n_593), .Y(n_624) );
INVx1_ASAP7_75t_SL g625 ( .A(n_610), .Y(n_625) );
NOR2x1_ASAP7_75t_L g626 ( .A(n_624), .B(n_611), .Y(n_626) );
CKINVDCx5p33_ASAP7_75t_R g627 ( .A(n_610), .Y(n_627) );
NOR2xp33_ASAP7_75t_L g628 ( .A(n_614), .B(n_612), .Y(n_628) );
OAI22xp5_ASAP7_75t_L g629 ( .A1(n_626), .A2(n_616), .B1(n_617), .B2(n_615), .Y(n_629) );
NOR3xp33_ASAP7_75t_L g630 ( .A(n_628), .B(n_622), .C(n_613), .Y(n_630) );
NAND3xp33_ASAP7_75t_L g631 ( .A(n_627), .B(n_621), .C(n_623), .Y(n_631) );
NOR2xp33_ASAP7_75t_R g632 ( .A(n_631), .B(n_625), .Y(n_632) );
BUFx2_ASAP7_75t_L g633 ( .A(n_629), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_632), .Y(n_634) );
AOI22xp5_ASAP7_75t_SL g635 ( .A1(n_634), .A2(n_633), .B1(n_616), .B2(n_630), .Y(n_635) );
AOI221xp5_ASAP7_75t_L g636 ( .A1(n_635), .A2(n_620), .B1(n_609), .B2(n_618), .C(n_619), .Y(n_636) );
endmodule