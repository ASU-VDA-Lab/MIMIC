module fake_netlist_5_2468_n_878 (n_137, n_168, n_164, n_191, n_91, n_82, n_122, n_194, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_188, n_190, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_878);

input n_137;
input n_168;
input n_164;
input n_191;
input n_91;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_188;
input n_190;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_878;

wire n_676;
wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_653;
wire n_611;
wire n_444;
wire n_642;
wire n_469;
wire n_615;
wire n_851;
wire n_316;
wire n_785;
wire n_389;
wire n_843;
wire n_855;
wire n_549;
wire n_684;
wire n_850;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_523;
wire n_451;
wire n_532;
wire n_705;
wire n_619;
wire n_408;
wire n_865;
wire n_678;
wire n_664;
wire n_376;
wire n_697;
wire n_503;
wire n_235;
wire n_226;
wire n_605;
wire n_776;
wire n_667;
wire n_515;
wire n_790;
wire n_353;
wire n_351;
wire n_367;
wire n_620;
wire n_643;
wire n_452;
wire n_397;
wire n_493;
wire n_525;
wire n_703;
wire n_698;
wire n_483;
wire n_544;
wire n_683;
wire n_780;
wire n_649;
wire n_552;
wire n_547;
wire n_721;
wire n_841;
wire n_467;
wire n_564;
wire n_802;
wire n_423;
wire n_840;
wire n_284;
wire n_501;
wire n_245;
wire n_823;
wire n_725;
wire n_280;
wire n_744;
wire n_590;
wire n_629;
wire n_672;
wire n_873;
wire n_378;
wire n_551;
wire n_762;
wire n_581;
wire n_688;
wire n_382;
wire n_554;
wire n_800;
wire n_254;
wire n_690;
wire n_583;
wire n_671;
wire n_718;
wire n_819;
wire n_302;
wire n_265;
wire n_526;
wire n_719;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_677;
wire n_859;
wire n_864;
wire n_821;
wire n_198;
wire n_714;
wire n_447;
wire n_314;
wire n_368;
wire n_247;
wire n_433;
wire n_604;
wire n_321;
wire n_292;
wire n_625;
wire n_854;
wire n_621;
wire n_753;
wire n_455;
wire n_674;
wire n_417;
wire n_612;
wire n_212;
wire n_385;
wire n_498;
wire n_516;
wire n_788;
wire n_507;
wire n_497;
wire n_689;
wire n_738;
wire n_606;
wire n_559;
wire n_275;
wire n_640;
wire n_252;
wire n_624;
wire n_825;
wire n_295;
wire n_330;
wire n_877;
wire n_508;
wire n_739;
wire n_506;
wire n_737;
wire n_610;
wire n_692;
wire n_755;
wire n_509;
wire n_568;
wire n_373;
wire n_820;
wire n_757;
wire n_307;
wire n_633;
wire n_439;
wire n_530;
wire n_556;
wire n_209;
wire n_259;
wire n_448;
wire n_758;
wire n_668;
wire n_733;
wire n_375;
wire n_301;
wire n_828;
wire n_779;
wire n_576;
wire n_804;
wire n_867;
wire n_537;
wire n_587;
wire n_659;
wire n_492;
wire n_792;
wire n_563;
wire n_756;
wire n_524;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_579;
wire n_741;
wire n_548;
wire n_543;
wire n_260;
wire n_812;
wire n_842;
wire n_298;
wire n_650;
wire n_320;
wire n_694;
wire n_518;
wire n_505;
wire n_286;
wire n_282;
wire n_752;
wire n_331;
wire n_406;
wire n_519;
wire n_470;
wire n_782;
wire n_325;
wire n_449;
wire n_862;
wire n_724;
wire n_856;
wire n_546;
wire n_760;
wire n_658;
wire n_281;
wire n_240;
wire n_381;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_731;
wire n_456;
wire n_371;
wire n_481;
wire n_535;
wire n_709;
wire n_540;
wire n_317;
wire n_618;
wire n_323;
wire n_569;
wire n_769;
wire n_356;
wire n_227;
wire n_592;
wire n_271;
wire n_831;
wire n_826;
wire n_335;
wire n_654;
wire n_370;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_514;
wire n_457;
wire n_570;
wire n_833;
wire n_297;
wire n_853;
wire n_603;
wire n_225;
wire n_377;
wire n_751;
wire n_484;
wire n_775;
wire n_219;
wire n_442;
wire n_814;
wire n_636;
wire n_786;
wire n_600;
wire n_660;
wire n_223;
wire n_392;
wire n_655;
wire n_704;
wire n_787;
wire n_264;
wire n_669;
wire n_472;
wire n_742;
wire n_750;
wire n_454;
wire n_387;
wire n_771;
wire n_374;
wire n_276;
wire n_339;
wire n_243;
wire n_398;
wire n_396;
wire n_635;
wire n_347;
wire n_763;
wire n_550;
wire n_522;
wire n_255;
wire n_696;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_662;
wire n_459;
wire n_646;
wire n_211;
wire n_218;
wire n_400;
wire n_436;
wire n_290;
wire n_580;
wire n_221;
wire n_622;
wire n_723;
wire n_386;
wire n_578;
wire n_287;
wire n_344;
wire n_848;
wire n_555;
wire n_783;
wire n_473;
wire n_422;
wire n_475;
wire n_777;
wire n_661;
wire n_682;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_849;
wire n_486;
wire n_670;
wire n_816;
wire n_336;
wire n_584;
wire n_681;
wire n_591;
wire n_521;
wire n_614;
wire n_663;
wire n_845;
wire n_430;
wire n_337;
wire n_313;
wire n_631;
wire n_673;
wire n_837;
wire n_479;
wire n_528;
wire n_510;
wire n_216;
wire n_680;
wire n_432;
wire n_395;
wire n_553;
wire n_727;
wire n_839;
wire n_311;
wire n_813;
wire n_830;
wire n_773;
wire n_208;
wire n_743;
wire n_214;
wire n_328;
wire n_801;
wire n_299;
wire n_303;
wire n_369;
wire n_675;
wire n_296;
wire n_613;
wire n_871;
wire n_241;
wire n_637;
wire n_357;
wire n_875;
wire n_598;
wire n_685;
wire n_608;
wire n_446;
wire n_445;
wire n_749;
wire n_829;
wire n_858;
wire n_772;
wire n_691;
wire n_717;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_517;
wire n_588;
wire n_361;
wire n_464;
wire n_789;
wire n_363;
wire n_413;
wire n_402;
wire n_734;
wire n_638;
wire n_700;
wire n_197;
wire n_796;
wire n_573;
wire n_866;
wire n_236;
wire n_388;
wire n_761;
wire n_249;
wire n_740;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_577;
wire n_384;
wire n_582;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_571;
wire n_461;
wire n_333;
wire n_693;
wire n_309;
wire n_512;
wire n_836;
wire n_462;
wire n_322;
wire n_567;
wire n_258;
wire n_652;
wire n_778;
wire n_306;
wire n_722;
wire n_458;
wire n_288;
wire n_770;
wire n_844;
wire n_201;
wire n_263;
wire n_471;
wire n_609;
wire n_852;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_711;
wire n_781;
wire n_834;
wire n_474;
wire n_765;
wire n_542;
wire n_488;
wire n_463;
wire n_595;
wire n_736;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_630;
wire n_489;
wire n_632;
wire n_699;
wire n_617;
wire n_310;
wire n_593;
wire n_504;
wire n_511;
wire n_748;
wire n_586;
wire n_846;
wire n_874;
wire n_465;
wire n_838;
wire n_358;
wire n_362;
wire n_876;
wire n_332;
wire n_273;
wire n_585;
wire n_349;
wire n_270;
wire n_616;
wire n_230;
wire n_601;
wire n_279;
wire n_253;
wire n_261;
wire n_289;
wire n_745;
wire n_627;
wire n_767;
wire n_206;
wire n_217;
wire n_440;
wire n_726;
wire n_478;
wire n_793;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_648;
wire n_312;
wire n_476;
wire n_818;
wire n_429;
wire n_861;
wire n_534;
wire n_345;
wire n_210;
wire n_494;
wire n_641;
wire n_628;
wire n_365;
wire n_774;
wire n_730;
wire n_729;
wire n_557;
wire n_354;
wire n_575;
wire n_647;
wire n_480;
wire n_607;
wire n_237;
wire n_425;
wire n_513;
wire n_407;
wire n_527;
wire n_707;
wire n_679;
wire n_710;
wire n_832;
wire n_695;
wire n_795;
wire n_857;
wire n_560;
wire n_656;
wire n_340;
wire n_207;
wire n_561;
wire n_346;
wire n_393;
wire n_229;
wire n_495;
wire n_487;
wire n_602;
wire n_665;
wire n_574;
wire n_437;
wire n_453;
wire n_403;
wire n_421;
wire n_720;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_863;
wire n_490;
wire n_805;
wire n_326;
wire n_794;
wire n_768;
wire n_233;
wire n_404;
wire n_686;
wire n_205;
wire n_366;
wire n_572;
wire n_712;
wire n_754;
wire n_847;
wire n_815;
wire n_246;
wire n_596;
wire n_410;
wire n_558;
wire n_708;
wire n_269;
wire n_529;
wire n_735;
wire n_702;
wire n_285;
wire n_822;
wire n_412;
wire n_232;
wire n_327;
wire n_657;
wire n_644;
wire n_728;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_791;
wire n_732;
wire n_251;
wire n_352;
wire n_566;
wire n_426;
wire n_520;
wire n_565;
wire n_808;
wire n_409;
wire n_797;
wire n_589;
wire n_716;
wire n_597;
wire n_500;
wire n_562;
wire n_300;
wire n_651;
wire n_435;
wire n_809;
wire n_870;
wire n_334;
wire n_599;
wire n_766;
wire n_811;
wire n_541;
wire n_807;
wire n_391;
wire n_701;
wire n_434;
wire n_645;
wire n_539;
wire n_835;
wire n_538;
wire n_666;
wire n_262;
wire n_803;
wire n_868;
wire n_238;
wire n_639;
wire n_799;
wire n_687;
wire n_715;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_536;
wire n_531;
wire n_242;
wire n_817;
wire n_872;
wire n_360;
wire n_594;
wire n_764;
wire n_200;
wire n_759;
wire n_222;
wire n_438;
wire n_806;
wire n_713;
wire n_869;
wire n_324;
wire n_810;
wire n_634;
wire n_416;
wire n_199;
wire n_827;
wire n_401;
wire n_348;
wire n_626;
wire n_424;
wire n_706;
wire n_746;
wire n_256;
wire n_305;
wire n_533;
wire n_747;
wire n_278;
wire n_784;

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_72),
.Y(n_196)
);

BUFx2_ASAP7_75t_L g197 ( 
.A(n_139),
.Y(n_197)
);

BUFx10_ASAP7_75t_L g198 ( 
.A(n_24),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_155),
.Y(n_200)
);

BUFx2_ASAP7_75t_L g201 ( 
.A(n_164),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_173),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_170),
.Y(n_203)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_193),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_120),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_118),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g208 ( 
.A(n_152),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_147),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_162),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_17),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_53),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_23),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_158),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_106),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_179),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_144),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_54),
.Y(n_219)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_180),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_189),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_77),
.Y(n_222)
);

INVx1_ASAP7_75t_SL g223 ( 
.A(n_112),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_117),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_43),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_135),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_125),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_55),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_100),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_130),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_12),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_11),
.Y(n_233)
);

INVx2_ASAP7_75t_L g234 ( 
.A(n_98),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_160),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_32),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_97),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_6),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_63),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_192),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_40),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_129),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_4),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_4),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_92),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_107),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_148),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_163),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_12),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_19),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_116),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_153),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_122),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_16),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_86),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_85),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_172),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_11),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_103),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_62),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_68),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g263 ( 
.A(n_99),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_10),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_41),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_177),
.Y(n_266)
);

INVx1_ASAP7_75t_SL g267 ( 
.A(n_67),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_29),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_31),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_90),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_69),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_114),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_109),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_142),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_131),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_39),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_102),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_0),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_20),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_105),
.Y(n_280)
);

INVxp33_ASAP7_75t_R g281 ( 
.A(n_42),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_136),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g283 ( 
.A(n_211),
.B(n_0),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_196),
.Y(n_284)
);

INVxp67_ASAP7_75t_SL g285 ( 
.A(n_197),
.Y(n_285)
);

BUFx6f_ASAP7_75t_SL g286 ( 
.A(n_198),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_232),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_233),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_208),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_201),
.B(n_1),
.Y(n_290)
);

INVxp33_ASAP7_75t_SL g291 ( 
.A(n_238),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_244),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_259),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_251),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_199),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_206),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_207),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_212),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_203),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_216),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_219),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_224),
.Y(n_303)
);

BUFx2_ASAP7_75t_SL g304 ( 
.A(n_198),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_225),
.Y(n_305)
);

CKINVDCx16_ASAP7_75t_R g306 ( 
.A(n_198),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_205),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_209),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_226),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_210),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_229),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_200),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_250),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_231),
.Y(n_314)
);

INVxp67_ASAP7_75t_SL g315 ( 
.A(n_228),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVxp67_ASAP7_75t_SL g317 ( 
.A(n_237),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_239),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_214),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_215),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_243),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_242),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_254),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_256),
.Y(n_324)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_204),
.Y(n_325)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_264),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_223),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_260),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_265),
.Y(n_329)
);

INVxp33_ASAP7_75t_SL g330 ( 
.A(n_278),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g331 ( 
.A(n_271),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_255),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_272),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_243),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_312),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_312),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_312),
.B(n_282),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g338 ( 
.A(n_285),
.B(n_267),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_312),
.Y(n_339)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_321),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_287),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_295),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_321),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_288),
.Y(n_344)
);

INVx6_ASAP7_75t_L g345 ( 
.A(n_306),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_296),
.Y(n_346)
);

OAI21x1_ASAP7_75t_L g347 ( 
.A1(n_297),
.A2(n_202),
.B(n_200),
.Y(n_347)
);

CKINVDCx8_ASAP7_75t_R g348 ( 
.A(n_304),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_293),
.Y(n_349)
);

AND2x6_ASAP7_75t_L g350 ( 
.A(n_283),
.B(n_202),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_299),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_301),
.Y(n_353)
);

AND2x2_ASAP7_75t_L g354 ( 
.A(n_315),
.B(n_282),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_284),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_302),
.Y(n_356)
);

BUFx6f_ASAP7_75t_L g357 ( 
.A(n_303),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_305),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_309),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_311),
.Y(n_360)
);

INVx3_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_316),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_318),
.Y(n_363)
);

NAND2xp33_ASAP7_75t_SL g364 ( 
.A(n_332),
.B(n_220),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_322),
.Y(n_365)
);

BUFx6f_ASAP7_75t_L g366 ( 
.A(n_323),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g367 ( 
.A1(n_325),
.A2(n_269),
.B1(n_217),
.B2(n_252),
.Y(n_367)
);

HB1xp67_ASAP7_75t_L g368 ( 
.A(n_334),
.Y(n_368)
);

AND2x2_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_324),
.Y(n_370)
);

BUFx6f_ASAP7_75t_L g371 ( 
.A(n_328),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

HB1xp67_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_317),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_289),
.B(n_220),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_331),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_290),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_290),
.Y(n_378)
);

INVx3_ASAP7_75t_L g379 ( 
.A(n_300),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_307),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_332),
.A2(n_234),
.B1(n_281),
.B2(n_279),
.Y(n_381)
);

AND2x6_ASAP7_75t_L g382 ( 
.A(n_286),
.B(n_234),
.Y(n_382)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_310),
.Y(n_383)
);

BUFx2_ASAP7_75t_L g384 ( 
.A(n_292),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_320),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_286),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_291),
.B(n_263),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_348),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_336),
.B(n_263),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_342),
.Y(n_390)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_375),
.B(n_274),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_339),
.B(n_263),
.Y(n_392)
);

INVx4_ASAP7_75t_L g393 ( 
.A(n_383),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_335),
.Y(n_394)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_357),
.Y(n_395)
);

AND2x6_ASAP7_75t_L g396 ( 
.A(n_380),
.B(n_383),
.Y(n_396)
);

BUFx10_ASAP7_75t_L g397 ( 
.A(n_345),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

BUFx2_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_352),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_353),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_351),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_374),
.B(n_326),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_368),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_356),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_383),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_358),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_345),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_338),
.B(n_308),
.Y(n_409)
);

BUFx3_ASAP7_75t_L g410 ( 
.A(n_383),
.Y(n_410)
);

BUFx3_ASAP7_75t_L g411 ( 
.A(n_385),
.Y(n_411)
);

AND3x2_ASAP7_75t_L g412 ( 
.A(n_340),
.B(n_280),
.C(n_294),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_360),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_377),
.B(n_330),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_350),
.B(n_263),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_376),
.B(n_319),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g417 ( 
.A(n_387),
.B(n_292),
.Y(n_417)
);

INVx4_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

AND2x4_ASAP7_75t_L g419 ( 
.A(n_373),
.B(n_221),
.Y(n_419)
);

HB1xp67_ASAP7_75t_L g420 ( 
.A(n_368),
.Y(n_420)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_357),
.Y(n_421)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_363),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_387),
.B(n_313),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_350),
.B(n_263),
.Y(n_424)
);

OR2x6_ASAP7_75t_L g425 ( 
.A(n_345),
.B(n_385),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_362),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_350),
.B(n_263),
.Y(n_428)
);

AOI22xp33_ASAP7_75t_L g429 ( 
.A1(n_377),
.A2(n_313),
.B1(n_277),
.B2(n_276),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_357),
.Y(n_430)
);

AND2x4_ASAP7_75t_L g431 ( 
.A(n_373),
.B(n_222),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_350),
.B(n_227),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_340),
.Y(n_434)
);

AOI22xp33_ASAP7_75t_L g435 ( 
.A1(n_377),
.A2(n_275),
.B1(n_273),
.B2(n_270),
.Y(n_435)
);

AND2x4_ASAP7_75t_L g436 ( 
.A(n_337),
.B(n_230),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_377),
.B(n_235),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_337),
.B(n_240),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_355),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_378),
.B(n_241),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_378),
.B(n_268),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_370),
.Y(n_442)
);

INVx6_ASAP7_75t_L g443 ( 
.A(n_355),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_359),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_359),
.Y(n_445)
);

BUFx6f_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_384),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_343),
.B(n_245),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_350),
.B(n_246),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_359),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g451 ( 
.A(n_343),
.B(n_247),
.Y(n_451)
);

BUFx4f_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g453 ( 
.A(n_372),
.B(n_378),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_390),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_388),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_400),
.Y(n_456)
);

AND2x4_ASAP7_75t_L g457 ( 
.A(n_410),
.B(n_379),
.Y(n_457)
);

AOI22xp5_ASAP7_75t_L g458 ( 
.A1(n_417),
.A2(n_354),
.B1(n_379),
.B2(n_364),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_405),
.Y(n_460)
);

AND2x4_ASAP7_75t_L g461 ( 
.A(n_411),
.B(n_341),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_434),
.Y(n_462)
);

AO22x2_ASAP7_75t_L g463 ( 
.A1(n_409),
.A2(n_404),
.B1(n_451),
.B2(n_414),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_407),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_413),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_437),
.B(n_367),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_426),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_403),
.B(n_381),
.Y(n_468)
);

INVx1_ASAP7_75t_SL g469 ( 
.A(n_420),
.Y(n_469)
);

AO22x2_ASAP7_75t_L g470 ( 
.A1(n_404),
.A2(n_386),
.B1(n_364),
.B2(n_3),
.Y(n_470)
);

INVxp67_ASAP7_75t_L g471 ( 
.A(n_448),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_402),
.Y(n_472)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_416),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_406),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_419),
.Y(n_475)
);

AO22x2_ASAP7_75t_L g476 ( 
.A1(n_419),
.A2(n_431),
.B1(n_453),
.B2(n_440),
.Y(n_476)
);

INVx2_ASAP7_75t_SL g477 ( 
.A(n_397),
.Y(n_477)
);

OR2x2_ASAP7_75t_L g478 ( 
.A(n_453),
.B(n_344),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_431),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_423),
.A2(n_382),
.B1(n_266),
.B2(n_262),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_432),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_399),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g483 ( 
.A1(n_441),
.A2(n_382),
.B1(n_248),
.B2(n_261),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g484 ( 
.A(n_443),
.B(n_366),
.Y(n_484)
);

AO22x2_ASAP7_75t_L g485 ( 
.A1(n_391),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_443),
.B(n_344),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_442),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_422),
.Y(n_488)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_427),
.B(n_361),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_452),
.B(n_436),
.Y(n_490)
);

AOI22xp33_ASAP7_75t_L g491 ( 
.A1(n_436),
.A2(n_361),
.B1(n_371),
.B2(n_366),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_389),
.Y(n_492)
);

BUFx8_ASAP7_75t_L g493 ( 
.A(n_396),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_452),
.B(n_366),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_389),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_392),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_425),
.B(n_349),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_392),
.Y(n_498)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_438),
.Y(n_499)
);

INVx2_ASAP7_75t_SL g500 ( 
.A(n_397),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_394),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_393),
.B(n_346),
.Y(n_502)
);

NAND2x1p5_ASAP7_75t_L g503 ( 
.A(n_393),
.B(n_346),
.Y(n_503)
);

AO22x2_ASAP7_75t_L g504 ( 
.A1(n_438),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_430),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_444),
.Y(n_506)
);

AND2x4_ASAP7_75t_L g507 ( 
.A(n_418),
.B(n_382),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_L g508 ( 
.A(n_395),
.B(n_366),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_450),
.Y(n_509)
);

AO22x2_ASAP7_75t_L g510 ( 
.A1(n_412),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_510)
);

NAND2x1p5_ASAP7_75t_L g511 ( 
.A(n_418),
.B(n_371),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_425),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_408),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_415),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_439),
.B(n_371),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_424),
.Y(n_517)
);

OAI221xp5_ASAP7_75t_L g518 ( 
.A1(n_435),
.A2(n_371),
.B1(n_258),
.B2(n_257),
.C(n_253),
.Y(n_518)
);

AO22x2_ASAP7_75t_L g519 ( 
.A1(n_412),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_395),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_429),
.B(n_249),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_408),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_466),
.B(n_446),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_473),
.B(n_446),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_SL g525 ( 
.A(n_458),
.B(n_446),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_478),
.B(n_396),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_457),
.B(n_433),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_SL g528 ( 
.A(n_499),
.B(n_433),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_492),
.B(n_396),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_457),
.B(n_449),
.Y(n_530)
);

NAND2xp33_ASAP7_75t_SL g531 ( 
.A(n_477),
.B(n_449),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_471),
.B(n_447),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_495),
.B(n_396),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_490),
.B(n_445),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_468),
.B(n_486),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_502),
.B(n_445),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_502),
.B(n_398),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_491),
.B(n_398),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_496),
.B(n_498),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g540 ( 
.A(n_514),
.B(n_421),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_500),
.B(n_424),
.Y(n_541)
);

AND2x4_ASAP7_75t_L g542 ( 
.A(n_454),
.B(n_425),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_SL g543 ( 
.A(n_522),
.B(n_513),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_SL g544 ( 
.A(n_475),
.B(n_421),
.Y(n_544)
);

NAND2xp33_ASAP7_75t_SL g545 ( 
.A(n_474),
.B(n_428),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_479),
.B(n_428),
.Y(n_546)
);

NAND2xp33_ASAP7_75t_SL g547 ( 
.A(n_455),
.B(n_382),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g548 ( 
.A(n_489),
.B(n_347),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_469),
.B(n_382),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_515),
.B(n_9),
.Y(n_550)
);

NAND2xp33_ASAP7_75t_SL g551 ( 
.A(n_497),
.B(n_10),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_461),
.B(n_21),
.Y(n_552)
);

NAND2xp33_ASAP7_75t_SL g553 ( 
.A(n_521),
.B(n_13),
.Y(n_553)
);

NAND2xp33_ASAP7_75t_SL g554 ( 
.A(n_516),
.B(n_13),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g555 ( 
.A(n_461),
.B(n_22),
.Y(n_555)
);

NAND2xp33_ASAP7_75t_SL g556 ( 
.A(n_507),
.B(n_14),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_507),
.B(n_14),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_SL g558 ( 
.A(n_462),
.B(n_456),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_459),
.B(n_25),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_460),
.B(n_26),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_464),
.B(n_27),
.Y(n_561)
);

NAND2xp33_ASAP7_75t_SL g562 ( 
.A(n_465),
.B(n_15),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_467),
.B(n_28),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_481),
.B(n_30),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_487),
.B(n_482),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_480),
.B(n_484),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_SL g567 ( 
.A(n_517),
.B(n_494),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_476),
.B(n_472),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_488),
.B(n_33),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_SL g570 ( 
.A(n_483),
.B(n_34),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_503),
.B(n_35),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_493),
.B(n_15),
.Y(n_572)
);

OR2x2_ASAP7_75t_L g573 ( 
.A(n_512),
.B(n_16),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_511),
.B(n_36),
.Y(n_574)
);

AND2x2_ASAP7_75t_SL g575 ( 
.A(n_485),
.B(n_37),
.Y(n_575)
);

AND2x2_ASAP7_75t_L g576 ( 
.A(n_463),
.B(n_476),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_508),
.B(n_520),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_SL g578 ( 
.A(n_501),
.B(n_38),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_505),
.B(n_17),
.Y(n_579)
);

NAND3xp33_ASAP7_75t_L g580 ( 
.A(n_535),
.B(n_518),
.C(n_506),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_539),
.A2(n_509),
.B(n_463),
.Y(n_581)
);

A2O1A1Ixp33_ASAP7_75t_L g582 ( 
.A1(n_550),
.A2(n_553),
.B(n_554),
.C(n_545),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_567),
.B(n_470),
.Y(n_583)
);

INVx1_ASAP7_75t_SL g584 ( 
.A(n_576),
.Y(n_584)
);

BUFx2_ASAP7_75t_L g585 ( 
.A(n_542),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_546),
.B(n_540),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_527),
.A2(n_530),
.B(n_536),
.Y(n_587)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_549),
.B(n_470),
.Y(n_588)
);

OAI22xp5_ASAP7_75t_L g589 ( 
.A1(n_575),
.A2(n_485),
.B1(n_504),
.B2(n_510),
.Y(n_589)
);

OA21x2_ASAP7_75t_L g590 ( 
.A1(n_568),
.A2(n_504),
.B(n_519),
.Y(n_590)
);

NAND2x1p5_ASAP7_75t_L g591 ( 
.A(n_542),
.B(n_44),
.Y(n_591)
);

AOI21x1_ASAP7_75t_L g592 ( 
.A1(n_523),
.A2(n_566),
.B(n_526),
.Y(n_592)
);

AOI21xp5_ASAP7_75t_L g593 ( 
.A1(n_529),
.A2(n_533),
.B(n_548),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_577),
.A2(n_121),
.B(n_46),
.Y(n_594)
);

BUFx3_ASAP7_75t_L g595 ( 
.A(n_573),
.Y(n_595)
);

OA21x2_ASAP7_75t_L g596 ( 
.A1(n_525),
.A2(n_519),
.B(n_510),
.Y(n_596)
);

INVx2_ASAP7_75t_SL g597 ( 
.A(n_565),
.Y(n_597)
);

AO31x2_ASAP7_75t_L g598 ( 
.A1(n_528),
.A2(n_18),
.A3(n_47),
.B(n_48),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_534),
.A2(n_123),
.B(n_49),
.Y(n_599)
);

OAI21x1_ASAP7_75t_L g600 ( 
.A1(n_538),
.A2(n_124),
.B(n_50),
.Y(n_600)
);

AND2x2_ASAP7_75t_L g601 ( 
.A(n_542),
.B(n_18),
.Y(n_601)
);

CKINVDCx16_ASAP7_75t_R g602 ( 
.A(n_547),
.Y(n_602)
);

AOI21xp5_ASAP7_75t_L g603 ( 
.A1(n_537),
.A2(n_51),
.B(n_52),
.Y(n_603)
);

BUFx12f_ASAP7_75t_L g604 ( 
.A(n_575),
.Y(n_604)
);

OAI22xp5_ASAP7_75t_L g605 ( 
.A1(n_524),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_544),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_L g607 ( 
.A(n_552),
.B(n_59),
.Y(n_607)
);

AO21x2_ASAP7_75t_L g608 ( 
.A1(n_570),
.A2(n_60),
.B(n_61),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_571),
.A2(n_64),
.B(n_65),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_532),
.B(n_66),
.Y(n_610)
);

AOI21xp5_ASAP7_75t_SL g611 ( 
.A1(n_574),
.A2(n_70),
.B(n_71),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_543),
.Y(n_612)
);

CKINVDCx20_ASAP7_75t_R g613 ( 
.A(n_558),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_555),
.B(n_73),
.Y(n_614)
);

AO32x2_ASAP7_75t_L g615 ( 
.A1(n_551),
.A2(n_195),
.A3(n_75),
.B1(n_76),
.B2(n_78),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_531),
.Y(n_616)
);

OAI21xp5_ASAP7_75t_L g617 ( 
.A1(n_559),
.A2(n_194),
.B(n_79),
.Y(n_617)
);

OAI21x1_ASAP7_75t_L g618 ( 
.A1(n_578),
.A2(n_561),
.B(n_564),
.Y(n_618)
);

BUFx2_ASAP7_75t_L g619 ( 
.A(n_556),
.Y(n_619)
);

BUFx10_ASAP7_75t_L g620 ( 
.A(n_562),
.Y(n_620)
);

OAI22xp5_ASAP7_75t_L g621 ( 
.A1(n_560),
.A2(n_74),
.B1(n_80),
.B2(n_81),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_557),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_579),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_541),
.Y(n_624)
);

BUFx2_ASAP7_75t_L g625 ( 
.A(n_585),
.Y(n_625)
);

OAI21x1_ASAP7_75t_L g626 ( 
.A1(n_593),
.A2(n_592),
.B(n_600),
.Y(n_626)
);

CKINVDCx20_ASAP7_75t_R g627 ( 
.A(n_613),
.Y(n_627)
);

AND2x4_ASAP7_75t_L g628 ( 
.A(n_597),
.B(n_563),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_606),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_587),
.A2(n_569),
.B(n_83),
.Y(n_630)
);

AOI22xp33_ASAP7_75t_L g631 ( 
.A1(n_589),
.A2(n_572),
.B1(n_84),
.B2(n_87),
.Y(n_631)
);

OAI21x1_ASAP7_75t_SL g632 ( 
.A1(n_617),
.A2(n_82),
.B(n_88),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_623),
.Y(n_633)
);

CKINVDCx8_ASAP7_75t_R g634 ( 
.A(n_612),
.Y(n_634)
);

OA21x2_ASAP7_75t_L g635 ( 
.A1(n_581),
.A2(n_89),
.B(n_91),
.Y(n_635)
);

OA21x2_ASAP7_75t_L g636 ( 
.A1(n_580),
.A2(n_93),
.B(n_94),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_586),
.B(n_95),
.Y(n_637)
);

AOI21x1_ASAP7_75t_L g638 ( 
.A1(n_580),
.A2(n_96),
.B(n_101),
.Y(n_638)
);

OAI21x1_ASAP7_75t_L g639 ( 
.A1(n_599),
.A2(n_108),
.B(n_110),
.Y(n_639)
);

OR2x2_ASAP7_75t_L g640 ( 
.A(n_584),
.B(n_111),
.Y(n_640)
);

OAI21x1_ASAP7_75t_L g641 ( 
.A1(n_594),
.A2(n_113),
.B(n_115),
.Y(n_641)
);

AOI22xp33_ASAP7_75t_L g642 ( 
.A1(n_589),
.A2(n_119),
.B1(n_126),
.B2(n_127),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_591),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_622),
.Y(n_644)
);

OAI21x1_ASAP7_75t_L g645 ( 
.A1(n_618),
.A2(n_128),
.B(n_132),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_624),
.B(n_133),
.Y(n_646)
);

AOI21xp5_ASAP7_75t_L g647 ( 
.A1(n_582),
.A2(n_134),
.B(n_137),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_584),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_588),
.B(n_138),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_583),
.Y(n_650)
);

AOI22xp33_ASAP7_75t_L g651 ( 
.A1(n_604),
.A2(n_140),
.B1(n_141),
.B2(n_143),
.Y(n_651)
);

INVx4_ASAP7_75t_L g652 ( 
.A(n_591),
.Y(n_652)
);

NOR2xp67_ASAP7_75t_SL g653 ( 
.A(n_611),
.B(n_145),
.Y(n_653)
);

AND2x4_ASAP7_75t_L g654 ( 
.A(n_619),
.B(n_146),
.Y(n_654)
);

OAI21x1_ASAP7_75t_L g655 ( 
.A1(n_624),
.A2(n_149),
.B(n_150),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_617),
.A2(n_151),
.B(n_154),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_595),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_601),
.Y(n_658)
);

CKINVDCx16_ASAP7_75t_R g659 ( 
.A(n_602),
.Y(n_659)
);

CKINVDCx11_ASAP7_75t_R g660 ( 
.A(n_620),
.Y(n_660)
);

HB1xp67_ASAP7_75t_L g661 ( 
.A(n_596),
.Y(n_661)
);

INVxp67_ASAP7_75t_L g662 ( 
.A(n_590),
.Y(n_662)
);

OAI222xp33_ASAP7_75t_L g663 ( 
.A1(n_621),
.A2(n_156),
.B1(n_157),
.B2(n_159),
.C1(n_161),
.C2(n_165),
.Y(n_663)
);

AOI22xp33_ASAP7_75t_L g664 ( 
.A1(n_596),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_620),
.B(n_171),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_608),
.Y(n_666)
);

OAI21x1_ASAP7_75t_L g667 ( 
.A1(n_603),
.A2(n_174),
.B(n_175),
.Y(n_667)
);

AO31x2_ASAP7_75t_L g668 ( 
.A1(n_666),
.A2(n_647),
.A3(n_637),
.B(n_650),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_644),
.Y(n_669)
);

AOI21x1_ASAP7_75t_L g670 ( 
.A1(n_638),
.A2(n_614),
.B(n_607),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_R g671 ( 
.A(n_627),
.B(n_634),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_626),
.A2(n_621),
.B(n_605),
.Y(n_672)
);

OR2x6_ASAP7_75t_L g673 ( 
.A(n_647),
.B(n_590),
.Y(n_673)
);

AO21x2_ASAP7_75t_L g674 ( 
.A1(n_632),
.A2(n_608),
.B(n_609),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_629),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_633),
.Y(n_676)
);

INVx1_ASAP7_75t_L g677 ( 
.A(n_648),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_635),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_649),
.B(n_615),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_661),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_661),
.Y(n_681)
);

INVx3_ASAP7_75t_SL g682 ( 
.A(n_659),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_662),
.Y(n_683)
);

BUFx2_ASAP7_75t_L g684 ( 
.A(n_662),
.Y(n_684)
);

AOI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_654),
.A2(n_610),
.B1(n_616),
.B2(n_609),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_645),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_641),
.Y(n_687)
);

AO31x2_ASAP7_75t_L g688 ( 
.A1(n_637),
.A2(n_615),
.A3(n_598),
.B(n_181),
.Y(n_688)
);

INVx3_ASAP7_75t_L g689 ( 
.A(n_667),
.Y(n_689)
);

CKINVDCx5p33_ASAP7_75t_R g690 ( 
.A(n_660),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_657),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_649),
.B(n_615),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_658),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_639),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_625),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_640),
.Y(n_696)
);

INVx3_ASAP7_75t_L g697 ( 
.A(n_643),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_636),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_654),
.B(n_176),
.Y(n_699)
);

INVx2_ASAP7_75t_L g700 ( 
.A(n_636),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_643),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_628),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_628),
.Y(n_703)
);

INVx1_ASAP7_75t_SL g704 ( 
.A(n_643),
.Y(n_704)
);

INVx2_ASAP7_75t_SL g705 ( 
.A(n_652),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_665),
.Y(n_706)
);

OR2x2_ASAP7_75t_L g707 ( 
.A(n_652),
.B(n_598),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_630),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_665),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_656),
.Y(n_710)
);

AND2x2_ASAP7_75t_L g711 ( 
.A(n_642),
.B(n_598),
.Y(n_711)
);

INVxp33_ASAP7_75t_L g712 ( 
.A(n_631),
.Y(n_712)
);

BUFx3_ASAP7_75t_L g713 ( 
.A(n_646),
.Y(n_713)
);

NAND2xp33_ASAP7_75t_R g714 ( 
.A(n_671),
.B(n_655),
.Y(n_714)
);

XNOR2xp5_ASAP7_75t_L g715 ( 
.A(n_690),
.B(n_651),
.Y(n_715)
);

CKINVDCx8_ASAP7_75t_R g716 ( 
.A(n_690),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_684),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_R g718 ( 
.A(n_701),
.B(n_646),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_713),
.B(n_646),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_R g720 ( 
.A(n_701),
.B(n_646),
.Y(n_720)
);

BUFx3_ASAP7_75t_L g721 ( 
.A(n_691),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_R g722 ( 
.A(n_706),
.B(n_646),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_684),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_R g724 ( 
.A(n_699),
.B(n_178),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_696),
.B(n_631),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_680),
.Y(n_726)
);

OR2x4_ASAP7_75t_L g727 ( 
.A(n_702),
.B(n_703),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_709),
.B(n_642),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_R g729 ( 
.A(n_706),
.B(n_651),
.Y(n_729)
);

OR2x6_ASAP7_75t_L g730 ( 
.A(n_713),
.B(n_663),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_R g731 ( 
.A(n_691),
.B(n_664),
.Y(n_731)
);

CKINVDCx6p67_ASAP7_75t_R g732 ( 
.A(n_682),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_677),
.B(n_664),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_681),
.Y(n_734)
);

INVxp67_ASAP7_75t_L g735 ( 
.A(n_695),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_682),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_R g737 ( 
.A(n_697),
.B(n_182),
.Y(n_737)
);

XOR2xp5_ASAP7_75t_L g738 ( 
.A(n_685),
.B(n_183),
.Y(n_738)
);

INVxp67_ASAP7_75t_L g739 ( 
.A(n_693),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_697),
.B(n_184),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_SL g741 ( 
.A(n_712),
.B(n_653),
.Y(n_741)
);

OR2x6_ASAP7_75t_L g742 ( 
.A(n_705),
.B(n_663),
.Y(n_742)
);

CKINVDCx11_ASAP7_75t_R g743 ( 
.A(n_704),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_R g744 ( 
.A(n_697),
.B(n_186),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_R g745 ( 
.A(n_705),
.B(n_676),
.Y(n_745)
);

NOR2xp33_ASAP7_75t_R g746 ( 
.A(n_707),
.B(n_670),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_675),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_669),
.B(n_188),
.Y(n_748)
);

XNOR2xp5_ASAP7_75t_L g749 ( 
.A(n_675),
.B(n_190),
.Y(n_749)
);

NAND2xp33_ASAP7_75t_R g750 ( 
.A(n_673),
.B(n_707),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_735),
.B(n_739),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_743),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_734),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_747),
.B(n_683),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_725),
.B(n_683),
.Y(n_755)
);

AND2x2_ASAP7_75t_L g756 ( 
.A(n_717),
.B(n_711),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_726),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_723),
.B(n_711),
.Y(n_758)
);

BUFx2_ASAP7_75t_L g759 ( 
.A(n_746),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_730),
.B(n_679),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_727),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_728),
.B(n_669),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_730),
.B(n_692),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_733),
.Y(n_764)
);

OAI21xp5_ASAP7_75t_SL g765 ( 
.A1(n_715),
.A2(n_738),
.B(n_749),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_745),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_721),
.Y(n_767)
);

AND2x2_ASAP7_75t_L g768 ( 
.A(n_742),
.B(n_692),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_742),
.Y(n_769)
);

HB1xp67_ASAP7_75t_L g770 ( 
.A(n_750),
.Y(n_770)
);

AND2x4_ASAP7_75t_L g771 ( 
.A(n_719),
.B(n_681),
.Y(n_771)
);

AOI222xp33_ASAP7_75t_L g772 ( 
.A1(n_741),
.A2(n_679),
.B1(n_710),
.B2(n_672),
.C1(n_698),
.C2(n_700),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_748),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_732),
.B(n_668),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_719),
.B(n_688),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_736),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_722),
.B(n_688),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_731),
.B(n_688),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_718),
.Y(n_779)
);

BUFx2_ASAP7_75t_L g780 ( 
.A(n_769),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_761),
.A2(n_729),
.B1(n_673),
.B2(n_720),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_760),
.B(n_698),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_760),
.B(n_700),
.Y(n_783)
);

BUFx3_ASAP7_75t_L g784 ( 
.A(n_766),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_764),
.B(n_668),
.Y(n_785)
);

OAI31xp33_ASAP7_75t_SL g786 ( 
.A1(n_778),
.A2(n_724),
.A3(n_714),
.B(n_672),
.Y(n_786)
);

OR2x2_ASAP7_75t_L g787 ( 
.A(n_756),
.B(n_668),
.Y(n_787)
);

AND2x2_ASAP7_75t_L g788 ( 
.A(n_763),
.B(n_688),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_775),
.B(n_673),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_753),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_763),
.B(n_688),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_768),
.B(n_673),
.Y(n_792)
);

OAI22xp5_ASAP7_75t_L g793 ( 
.A1(n_765),
.A2(n_716),
.B1(n_710),
.B2(n_708),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_768),
.B(n_668),
.Y(n_794)
);

AND2x4_ASAP7_75t_L g795 ( 
.A(n_775),
.B(n_708),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_753),
.Y(n_796)
);

AND2x2_ASAP7_75t_L g797 ( 
.A(n_756),
.B(n_668),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_758),
.B(n_678),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_790),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_790),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_780),
.B(n_770),
.Y(n_801)
);

AND3x2_ASAP7_75t_L g802 ( 
.A(n_786),
.B(n_759),
.C(n_776),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_796),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_780),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_792),
.B(n_758),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_785),
.B(n_764),
.Y(n_806)
);

AND2x2_ASAP7_75t_L g807 ( 
.A(n_792),
.B(n_777),
.Y(n_807)
);

AND2x2_ASAP7_75t_L g808 ( 
.A(n_782),
.B(n_777),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_798),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_809),
.Y(n_810)
);

NAND2xp33_ASAP7_75t_SL g811 ( 
.A(n_801),
.B(n_759),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_806),
.B(n_791),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_806),
.B(n_794),
.Y(n_813)
);

OR2x2_ASAP7_75t_L g814 ( 
.A(n_812),
.B(n_805),
.Y(n_814)
);

INVx1_ASAP7_75t_SL g815 ( 
.A(n_811),
.Y(n_815)
);

OR2x2_ASAP7_75t_L g816 ( 
.A(n_813),
.B(n_787),
.Y(n_816)
);

INVx1_ASAP7_75t_SL g817 ( 
.A(n_810),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_810),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_815),
.A2(n_793),
.B(n_752),
.C(n_778),
.Y(n_819)
);

AND2x2_ASAP7_75t_L g820 ( 
.A(n_817),
.B(n_807),
.Y(n_820)
);

AOI21xp33_ASAP7_75t_L g821 ( 
.A1(n_818),
.A2(n_774),
.B(n_779),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_814),
.Y(n_822)
);

AOI21xp33_ASAP7_75t_L g823 ( 
.A1(n_822),
.A2(n_774),
.B(n_776),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_820),
.Y(n_824)
);

OR2x2_ASAP7_75t_L g825 ( 
.A(n_819),
.B(n_816),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_824),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_825),
.B(n_821),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_823),
.Y(n_828)
);

INVx1_ASAP7_75t_SL g829 ( 
.A(n_824),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_826),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_829),
.B(n_827),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_828),
.Y(n_832)
);

NOR3xp33_ASAP7_75t_L g833 ( 
.A(n_827),
.B(n_751),
.C(n_767),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_SL g834 ( 
.A(n_827),
.B(n_737),
.C(n_740),
.Y(n_834)
);

AOI21xp33_ASAP7_75t_L g835 ( 
.A1(n_827),
.A2(n_784),
.B(n_754),
.Y(n_835)
);

NAND3xp33_ASAP7_75t_L g836 ( 
.A(n_827),
.B(n_802),
.C(n_784),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_831),
.A2(n_804),
.B(n_803),
.Y(n_837)
);

AOI21xp33_ASAP7_75t_R g838 ( 
.A1(n_832),
.A2(n_800),
.B(n_799),
.Y(n_838)
);

AOI211xp5_ASAP7_75t_L g839 ( 
.A1(n_836),
.A2(n_744),
.B(n_802),
.C(n_791),
.Y(n_839)
);

NAND4xp25_ASAP7_75t_L g840 ( 
.A(n_833),
.B(n_781),
.C(n_762),
.D(n_772),
.Y(n_840)
);

INVxp33_ASAP7_75t_L g841 ( 
.A(n_834),
.Y(n_841)
);

O2A1O1Ixp5_ASAP7_75t_L g842 ( 
.A1(n_830),
.A2(n_799),
.B(n_757),
.C(n_788),
.Y(n_842)
);

OAI21xp33_ASAP7_75t_L g843 ( 
.A1(n_835),
.A2(n_788),
.B(n_794),
.Y(n_843)
);

NAND4xp25_ASAP7_75t_L g844 ( 
.A(n_831),
.B(n_755),
.C(n_773),
.D(n_789),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_837),
.Y(n_845)
);

INVx2_ASAP7_75t_SL g846 ( 
.A(n_838),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_844),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_840),
.B(n_808),
.Y(n_848)
);

NOR3xp33_ASAP7_75t_L g849 ( 
.A(n_839),
.B(n_670),
.C(n_783),
.Y(n_849)
);

NAND4xp75_ASAP7_75t_L g850 ( 
.A(n_842),
.B(n_797),
.C(n_783),
.D(n_782),
.Y(n_850)
);

INVx2_ASAP7_75t_L g851 ( 
.A(n_841),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_843),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_845),
.B(n_771),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_851),
.B(n_797),
.Y(n_854)
);

NOR2xp33_ASAP7_75t_R g855 ( 
.A(n_846),
.B(n_847),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_852),
.B(n_795),
.Y(n_856)
);

XNOR2xp5_ASAP7_75t_L g857 ( 
.A(n_848),
.B(n_771),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_SL g858 ( 
.A(n_849),
.B(n_771),
.Y(n_858)
);

XNOR2xp5_ASAP7_75t_L g859 ( 
.A(n_850),
.B(n_789),
.Y(n_859)
);

HB1xp67_ASAP7_75t_L g860 ( 
.A(n_855),
.Y(n_860)
);

INVxp67_ASAP7_75t_L g861 ( 
.A(n_853),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_857),
.Y(n_862)
);

HB1xp67_ASAP7_75t_L g863 ( 
.A(n_856),
.Y(n_863)
);

NAND3xp33_ASAP7_75t_SL g864 ( 
.A(n_854),
.B(n_787),
.C(n_798),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_859),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_858),
.Y(n_866)
);

INVx2_ASAP7_75t_L g867 ( 
.A(n_860),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_865),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_863),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_861),
.Y(n_870)
);

AO22x1_ASAP7_75t_L g871 ( 
.A1(n_869),
.A2(n_862),
.B1(n_866),
.B2(n_864),
.Y(n_871)
);

BUFx2_ASAP7_75t_L g872 ( 
.A(n_867),
.Y(n_872)
);

AOI31xp33_ASAP7_75t_L g873 ( 
.A1(n_872),
.A2(n_870),
.A3(n_868),
.B(n_789),
.Y(n_873)
);

OAI322xp33_ASAP7_75t_L g874 ( 
.A1(n_873),
.A2(n_871),
.A3(n_686),
.B1(n_687),
.B2(n_694),
.C1(n_689),
.C2(n_191),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_874),
.A2(n_694),
.B(n_687),
.Y(n_875)
);

INVxp67_ASAP7_75t_SL g876 ( 
.A(n_875),
.Y(n_876)
);

AOI22xp33_ASAP7_75t_L g877 ( 
.A1(n_876),
.A2(n_795),
.B1(n_674),
.B2(n_689),
.Y(n_877)
);

AOI211xp5_ASAP7_75t_L g878 ( 
.A1(n_877),
.A2(n_795),
.B(n_686),
.C(n_678),
.Y(n_878)
);


endmodule