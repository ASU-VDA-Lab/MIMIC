module fake_jpeg_31646_n_441 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_441);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_441;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_12),
.B(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx13_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx1_ASAP7_75t_SL g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_2),
.B(n_12),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_15),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_46),
.Y(n_98)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

BUFx2_ASAP7_75t_SL g109 ( 
.A(n_47),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_19),
.B(n_15),
.Y(n_48)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_59),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_22),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_49),
.B(n_50),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_22),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_51),
.Y(n_121)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_53),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_54),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_55),
.Y(n_118)
);

INVx8_ASAP7_75t_SL g56 ( 
.A(n_23),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_56),
.Y(n_93)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_57),
.Y(n_101)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_29),
.Y(n_61)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_61),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_62),
.Y(n_123)
);

BUFx8_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_64),
.B(n_79),
.Y(n_112)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_23),
.Y(n_65)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_25),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_66),
.Y(n_127)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_67),
.Y(n_138)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_68),
.Y(n_131)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_70),
.Y(n_110)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_20),
.Y(n_71)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_71),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx6_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_73),
.Y(n_117)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_29),
.Y(n_74)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_74),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_75),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g76 ( 
.A(n_18),
.Y(n_76)
);

NAND2xp33_ASAP7_75t_SL g119 ( 
.A(n_76),
.B(n_36),
.Y(n_119)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_29),
.Y(n_77)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_18),
.Y(n_78)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_14),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_20),
.Y(n_80)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_81),
.Y(n_94)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_18),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_83),
.B(n_84),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_13),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_85),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_39),
.Y(n_86)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_86),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_39),
.Y(n_87)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_87),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_41),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_88),
.B(n_90),
.Y(n_124)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_39),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_44),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_91),
.B(n_42),
.Y(n_128)
);

OA22x2_ASAP7_75t_L g100 ( 
.A1(n_46),
.A2(n_32),
.B1(n_17),
.B2(n_34),
.Y(n_100)
);

OAI32xp33_ASAP7_75t_L g183 ( 
.A1(n_100),
.A2(n_125),
.A3(n_90),
.B1(n_21),
.B2(n_63),
.Y(n_183)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_81),
.A2(n_32),
.B1(n_21),
.B2(n_33),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_111),
.A2(n_67),
.B1(n_86),
.B2(n_89),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_47),
.A2(n_43),
.B1(n_44),
.B2(n_42),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

OR2x4_ASAP7_75t_L g165 ( 
.A(n_119),
.B(n_109),
.Y(n_165)
);

OA22x2_ASAP7_75t_L g125 ( 
.A1(n_68),
.A2(n_17),
.B1(n_36),
.B2(n_34),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_128),
.B(n_10),
.Y(n_174)
);

OAI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_82),
.A2(n_37),
.B1(n_35),
.B2(n_31),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_134),
.B1(n_135),
.B2(n_136),
.Y(n_160)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_61),
.Y(n_133)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_133),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_53),
.A2(n_31),
.B1(n_35),
.B2(n_37),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_54),
.A2(n_37),
.B1(n_35),
.B2(n_31),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g136 ( 
.A1(n_73),
.A2(n_39),
.B1(n_37),
.B2(n_35),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_55),
.A2(n_31),
.B1(n_28),
.B2(n_45),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_142),
.A2(n_143),
.B1(n_75),
.B2(n_69),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_62),
.A2(n_28),
.B1(n_45),
.B2(n_27),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_66),
.A2(n_33),
.B1(n_21),
.B2(n_17),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_144),
.A2(n_90),
.B1(n_33),
.B2(n_21),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_74),
.A2(n_45),
.B1(n_27),
.B2(n_11),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_105),
.Y(n_146)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_146),
.Y(n_229)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_147),
.Y(n_225)
);

INVx11_ASAP7_75t_L g148 ( 
.A(n_92),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g203 ( 
.A(n_148),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_114),
.B(n_27),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_151),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_96),
.B(n_76),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_150),
.B(n_172),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_72),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_152),
.B(n_156),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_110),
.A2(n_77),
.B1(n_78),
.B2(n_60),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_153),
.A2(n_181),
.B1(n_191),
.B2(n_97),
.Y(n_206)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_140),
.Y(n_154)
);

INVx4_ASAP7_75t_L g212 ( 
.A(n_154),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g155 ( 
.A(n_106),
.Y(n_155)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_155),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_112),
.B(n_11),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_137),
.B(n_87),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_157),
.B(n_161),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g158 ( 
.A(n_121),
.Y(n_158)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

INVx3_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_159),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g161 ( 
.A(n_96),
.B(n_11),
.Y(n_161)
);

INVx6_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_124),
.B(n_51),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_164),
.B(n_170),
.Y(n_218)
);

OAI21xp33_ASAP7_75t_L g214 ( 
.A1(n_165),
.A2(n_102),
.B(n_131),
.Y(n_214)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_171),
.Y(n_198)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_104),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_168),
.Y(n_230)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_169),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_125),
.B(n_65),
.Y(n_170)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_138),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_113),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_173),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_174),
.B(n_176),
.Y(n_220)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_101),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_175),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_125),
.B(n_65),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_93),
.B(n_85),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_103),
.B(n_63),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_178),
.B(n_185),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_93),
.B(n_33),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_179),
.B(n_184),
.Y(n_226)
);

OA22x2_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_183),
.B1(n_144),
.B2(n_136),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_129),
.A2(n_52),
.B1(n_33),
.B2(n_21),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_117),
.Y(n_182)
);

CKINVDCx14_ASAP7_75t_R g231 ( 
.A(n_182),
.Y(n_231)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_122),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_100),
.B(n_0),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_100),
.B(n_0),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_186),
.B(n_5),
.Y(n_227)
);

OAI22xp33_ASAP7_75t_SL g187 ( 
.A1(n_117),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_187)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_187),
.A2(n_97),
.B1(n_127),
.B2(n_115),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_111),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_188),
.B(n_190),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g189 ( 
.A(n_92),
.Y(n_189)
);

BUFx24_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_94),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_94),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_130),
.A2(n_1),
.B1(n_3),
.B2(n_5),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_192),
.A2(n_127),
.B1(n_123),
.B2(n_118),
.Y(n_208)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_95),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_132),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_194),
.Y(n_211)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_95),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_195),
.Y(n_232)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_99),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_196),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_204),
.A2(n_207),
.B1(n_208),
.B2(n_216),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_206),
.A2(n_189),
.B1(n_172),
.B2(n_163),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_149),
.B(n_108),
.C(n_126),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_213),
.B(n_221),
.C(n_235),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_214),
.B(n_227),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_98),
.B1(n_131),
.B2(n_115),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_162),
.B(n_98),
.C(n_123),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_162),
.B(n_3),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_224),
.B(n_148),
.Y(n_268)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_197),
.A2(n_5),
.B(n_7),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_233),
.A2(n_165),
.B(n_8),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_186),
.B(n_118),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_151),
.B(n_9),
.C(n_7),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_236),
.B(n_233),
.C(n_202),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_160),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_239),
.A2(n_180),
.B1(n_192),
.B2(n_155),
.Y(n_248)
);

AO22x1_ASAP7_75t_SL g240 ( 
.A1(n_183),
.A2(n_8),
.B1(n_170),
.B2(n_176),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_240),
.B(n_197),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_241),
.Y(n_286)
);

INVx5_ASAP7_75t_L g242 ( 
.A(n_203),
.Y(n_242)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_242),
.Y(n_283)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_243),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_245),
.B(n_252),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_246),
.B(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_200),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_248),
.A2(n_257),
.B1(n_264),
.B2(n_271),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_199),
.B(n_157),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_249),
.B(n_266),
.Y(n_298)
);

OAI21xp5_ASAP7_75t_L g309 ( 
.A1(n_251),
.A2(n_261),
.B(n_225),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_205),
.B(n_146),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_226),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_253),
.B(n_254),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_201),
.B(n_224),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_237),
.Y(n_255)
);

CKINVDCx14_ASAP7_75t_R g311 ( 
.A(n_255),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_205),
.B(n_166),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_256),
.B(n_258),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_198),
.A2(n_160),
.B1(n_167),
.B2(n_182),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_235),
.B(n_147),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_154),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_259),
.B(n_263),
.Y(n_294)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_260),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_218),
.A2(n_196),
.B(n_194),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_229),
.Y(n_262)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_262),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_228),
.B(n_169),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_198),
.A2(n_173),
.B1(n_159),
.B2(n_184),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_229),
.Y(n_265)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_265),
.Y(n_302)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_200),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_267),
.B(n_270),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g281 ( 
.A(n_268),
.B(n_232),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_8),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g304 ( 
.A(n_269),
.B(n_273),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_213),
.B(n_220),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_198),
.A2(n_239),
.B1(n_216),
.B2(n_204),
.Y(n_271)
);

INVx5_ASAP7_75t_L g272 ( 
.A(n_203),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_SL g308 ( 
.A1(n_272),
.A2(n_209),
.B1(n_200),
.B2(n_217),
.Y(n_308)
);

OR2x2_ASAP7_75t_L g273 ( 
.A(n_221),
.B(n_202),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_236),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_275),
.B(n_276),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_240),
.B(n_208),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_234),
.C(n_215),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_232),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_278),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_280),
.Y(n_317)
);

CKINVDCx14_ASAP7_75t_R g327 ( 
.A(n_281),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_271),
.A2(n_204),
.B1(n_223),
.B2(n_209),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_284),
.A2(n_310),
.B1(n_253),
.B2(n_248),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_262),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_288),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_265),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_291),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_268),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_296),
.B(n_243),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_251),
.A2(n_204),
.B(n_200),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_297),
.A2(n_305),
.B(n_273),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_277),
.A2(n_211),
.B1(n_231),
.B2(n_222),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_301),
.A2(n_303),
.B1(n_264),
.B2(n_261),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_244),
.A2(n_211),
.B1(n_223),
.B2(n_234),
.Y(n_303)
);

AOI21xp33_ASAP7_75t_L g305 ( 
.A1(n_275),
.A2(n_230),
.B(n_215),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g318 ( 
.A(n_306),
.B(n_274),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_256),
.B(n_225),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_307),
.B(n_309),
.Y(n_315)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_308),
.A2(n_267),
.B1(n_272),
.B2(n_242),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_257),
.A2(n_212),
.B1(n_225),
.B2(n_244),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_285),
.Y(n_312)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_312),
.Y(n_341)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_285),
.Y(n_313)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_313),
.Y(n_351)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_314),
.B(n_320),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_316),
.A2(n_324),
.B1(n_332),
.B2(n_301),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_SL g360 ( 
.A(n_318),
.B(n_323),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_289),
.B(n_246),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_319),
.B(n_329),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_281),
.B(n_252),
.Y(n_320)
);

NAND3xp33_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_270),
.C(n_263),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_321),
.B(n_326),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g322 ( 
.A(n_299),
.B(n_274),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_322),
.B(n_334),
.C(n_337),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_284),
.A2(n_250),
.B1(n_245),
.B2(n_273),
.Y(n_324)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_283),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_299),
.B(n_250),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_328),
.B(n_304),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_276),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_330),
.A2(n_336),
.B1(n_286),
.B2(n_310),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_331),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_303),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_296),
.B(n_266),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_333),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_212),
.C(n_247),
.Y(n_334)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_304),
.B(n_267),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_298),
.B(n_307),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_338),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_311),
.B(n_298),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_339),
.B(n_320),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_340),
.A2(n_357),
.B1(n_361),
.B2(n_332),
.Y(n_371)
);

OAI21xp5_ASAP7_75t_L g343 ( 
.A1(n_315),
.A2(n_297),
.B(n_309),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_343),
.A2(n_323),
.B(n_330),
.Y(n_366)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_327),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_344),
.B(n_356),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_345),
.B(n_349),
.C(n_354),
.Y(n_374)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_318),
.B(n_295),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_317),
.B(n_300),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g368 ( 
.A(n_353),
.Y(n_368)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_322),
.B(n_306),
.C(n_294),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_355),
.A2(n_315),
.B1(n_333),
.B2(n_335),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_317),
.B(n_300),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_316),
.A2(n_292),
.B1(n_297),
.B2(n_282),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_359),
.B(n_279),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_324),
.A2(n_292),
.B1(n_282),
.B2(n_305),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_328),
.B(n_294),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_362),
.B(n_363),
.C(n_354),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_293),
.C(n_280),
.Y(n_363)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_364),
.A2(n_382),
.B(n_361),
.Y(n_397)
);

AOI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_366),
.A2(n_379),
.B(n_372),
.Y(n_392)
);

CKINVDCx16_ASAP7_75t_R g367 ( 
.A(n_347),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_370),
.Y(n_394)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_347),
.Y(n_369)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_369),
.Y(n_395)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_341),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_L g390 ( 
.A1(n_371),
.A2(n_375),
.B1(n_381),
.B2(n_363),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_346),
.B(n_335),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_372),
.B(n_373),
.Y(n_391)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_341),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_325),
.B1(n_338),
.B2(n_279),
.Y(n_375)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_376),
.B(n_380),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g398 ( 
.A(n_377),
.B(n_379),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_342),
.B(n_334),
.C(n_293),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_378),
.B(n_345),
.C(n_362),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_358),
.B(n_325),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_SL g380 ( 
.A(n_352),
.B(n_313),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_357),
.A2(n_314),
.B1(n_312),
.B2(n_288),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_351),
.B(n_291),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_351),
.B(n_287),
.Y(n_383)
);

OAI21xp33_ASAP7_75t_L g396 ( 
.A1(n_383),
.A2(n_290),
.B(n_302),
.Y(n_396)
);

AOI32xp33_ASAP7_75t_L g385 ( 
.A1(n_368),
.A2(n_348),
.A3(n_343),
.B1(n_360),
.B2(n_355),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_385),
.B(n_396),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_342),
.C(n_349),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_386),
.B(n_389),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_366),
.B(n_360),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_SL g410 ( 
.A(n_387),
.B(n_383),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_370),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_388),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_393),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_392),
.B(n_375),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_376),
.B(n_374),
.C(n_378),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g408 ( 
.A(n_397),
.B(n_382),
.Y(n_408)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g409 ( 
.A1(n_399),
.A2(n_326),
.B1(n_290),
.B2(n_302),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_393),
.B(n_371),
.C(n_364),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_402),
.Y(n_415)
);

A2O1A1Ixp33_ASAP7_75t_SL g403 ( 
.A1(n_392),
.A2(n_367),
.B(n_381),
.C(n_340),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g420 ( 
.A(n_403),
.Y(n_420)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_395),
.A2(n_373),
.B1(n_380),
.B2(n_377),
.Y(n_406)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_406),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_408),
.Y(n_414)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_409),
.Y(n_417)
);

XNOR2x1_ASAP7_75t_SL g421 ( 
.A(n_410),
.B(n_387),
.Y(n_421)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_384),
.Y(n_411)
);

BUFx24_ASAP7_75t_SL g412 ( 
.A(n_411),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_384),
.C(n_389),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_419),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_391),
.B(n_394),
.Y(n_418)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_418),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_365),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_421),
.B(n_410),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g431 ( 
.A(n_422),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_SL g423 ( 
.A(n_420),
.B(n_405),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_423),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g425 ( 
.A1(n_414),
.A2(n_398),
.B(n_365),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_426),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_415),
.B(n_399),
.C(n_403),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_420),
.B(n_388),
.Y(n_427)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_427),
.Y(n_430)
);

O2A1O1Ixp33_ASAP7_75t_SL g433 ( 
.A1(n_432),
.A2(n_427),
.B(n_428),
.C(n_403),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_433),
.B(n_434),
.Y(n_436)
);

CKINVDCx14_ASAP7_75t_R g434 ( 
.A(n_429),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_430),
.B(n_424),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_435),
.B(n_431),
.Y(n_437)
);

OAI21xp5_ASAP7_75t_L g438 ( 
.A1(n_437),
.A2(n_413),
.B(n_412),
.Y(n_438)
);

AO21x2_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_436),
.B(n_396),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g440 ( 
.A1(n_439),
.A2(n_283),
.B1(n_417),
.B2(n_327),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_440),
.Y(n_441)
);


endmodule