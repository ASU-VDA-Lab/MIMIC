module fake_jpeg_3758_n_288 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_288);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_288;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_223;
wire n_57;
wire n_21;
wire n_187;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_270;
wire n_260;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

BUFx4f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx5_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_32),
.Y(n_44)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx12f_ASAP7_75t_SL g32 ( 
.A(n_17),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_18),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_37),
.B(n_38),
.Y(n_62)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_20),
.Y(n_56)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_49),
.B(n_52),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_19),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_50),
.B(n_44),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_38),
.A2(n_37),
.B1(n_36),
.B2(n_15),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_51),
.B(n_65),
.C(n_20),
.Y(n_80)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_38),
.A2(n_35),
.B1(n_29),
.B2(n_15),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_54),
.A2(n_42),
.B1(n_39),
.B2(n_52),
.Y(n_71)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_58),
.Y(n_75)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_56),
.Y(n_68)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_59),
.B(n_61),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_45),
.Y(n_63)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_63),
.Y(n_76)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_45),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_15),
.B1(n_29),
.B2(n_35),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g83 ( 
.A1(n_66),
.A2(n_39),
.B1(n_46),
.B2(n_43),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_67),
.A2(n_73),
.B(n_78),
.Y(n_91)
);

AOI32xp33_ASAP7_75t_L g69 ( 
.A1(n_62),
.A2(n_48),
.A3(n_19),
.B1(n_33),
.B2(n_42),
.Y(n_69)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_69),
.B(n_80),
.CI(n_14),
.CON(n_104),
.SN(n_104)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_50),
.A2(n_42),
.B1(n_46),
.B2(n_41),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_70),
.A2(n_81),
.B1(n_63),
.B2(n_61),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_71),
.A2(n_84),
.B1(n_66),
.B2(n_64),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_49),
.B(n_41),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_56),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_SL g73 ( 
.A(n_50),
.B(n_14),
.C(n_18),
.Y(n_73)
);

FAx1_ASAP7_75t_SL g77 ( 
.A(n_54),
.B(n_48),
.CI(n_43),
.CON(n_77),
.SN(n_77)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_77),
.B(n_43),
.Y(n_90)
);

FAx1_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_14),
.CI(n_46),
.CON(n_78),
.SN(n_78)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_46),
.B1(n_39),
.B2(n_13),
.Y(n_81)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_39),
.B1(n_13),
.B2(n_30),
.Y(n_84)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_86),
.B(n_96),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_68),
.B(n_58),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g117 ( 
.A(n_90),
.B(n_98),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_68),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_92),
.B(n_99),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_93),
.A2(n_81),
.B1(n_78),
.B2(n_71),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_94),
.A2(n_82),
.B1(n_77),
.B2(n_31),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_80),
.B(n_84),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_95),
.B(n_97),
.C(n_73),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_72),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_33),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_53),
.Y(n_100)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_100),
.Y(n_107)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_76),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_79),
.B(n_59),
.Y(n_102)
);

INVxp33_ASAP7_75t_L g106 ( 
.A(n_102),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_57),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_103),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g108 ( 
.A1(n_104),
.A2(n_69),
.B(n_78),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_97),
.B(n_78),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_105),
.B(n_108),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_109),
.A2(n_122),
.B1(n_88),
.B2(n_101),
.Y(n_129)
);

MAJx2_ASAP7_75t_L g112 ( 
.A(n_91),
.B(n_67),
.C(n_77),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g126 ( 
.A(n_112),
.B(n_104),
.Y(n_126)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_114),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_116),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_87),
.B(n_82),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_85),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_125),
.C(n_95),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_20),
.B(n_76),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_120),
.A2(n_89),
.B(n_99),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_90),
.A2(n_13),
.B(n_21),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_121),
.A2(n_115),
.B(n_107),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_93),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_94),
.A2(n_22),
.B1(n_24),
.B2(n_27),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_88),
.B1(n_98),
.B2(n_102),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_85),
.B1(n_34),
.B2(n_27),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_86),
.B1(n_85),
.B2(n_103),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_95),
.B(n_34),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_126),
.B(n_119),
.Y(n_156)
);

XNOR2x1_ASAP7_75t_SL g127 ( 
.A(n_112),
.B(n_104),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_127),
.B(n_25),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_117),
.A2(n_108),
.B(n_112),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g162 ( 
.A1(n_128),
.A2(n_132),
.B(n_134),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_129),
.A2(n_141),
.B1(n_134),
.B2(n_123),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_111),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_140),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_96),
.B(n_92),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_145),
.C(n_125),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g164 ( 
.A(n_135),
.Y(n_164)
);

OA21x2_ASAP7_75t_L g136 ( 
.A1(n_111),
.A2(n_100),
.B(n_97),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_136),
.A2(n_138),
.B(n_122),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_118),
.B(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_146),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_121),
.B(n_104),
.Y(n_140)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_142),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_114),
.Y(n_143)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_143),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_125),
.B(n_34),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_106),
.B(n_86),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_147),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_109),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_148),
.A2(n_120),
.B1(n_110),
.B2(n_107),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_150),
.A2(n_164),
.B1(n_149),
.B2(n_157),
.Y(n_183)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_151),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_144),
.A2(n_119),
.B1(n_105),
.B2(n_120),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_147),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_153),
.B(n_131),
.Y(n_177)
);

OAI21xp33_ASAP7_75t_L g155 ( 
.A1(n_127),
.A2(n_113),
.B(n_105),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_155),
.B(n_156),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_159),
.C(n_166),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_113),
.C(n_110),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_163),
.A2(n_167),
.B(n_138),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g165 ( 
.A(n_136),
.Y(n_165)
);

CKINVDCx16_ASAP7_75t_R g174 ( 
.A(n_165),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_25),
.C(n_26),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g167 ( 
.A1(n_128),
.A2(n_25),
.B(n_26),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_129),
.A2(n_23),
.B1(n_25),
.B2(n_26),
.Y(n_168)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_146),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_169),
.B(n_137),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_170),
.B(n_136),
.Y(n_178)
);

INVxp67_ASAP7_75t_SL g171 ( 
.A(n_136),
.Y(n_171)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_171),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_126),
.B(n_26),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_172),
.B(n_148),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_131),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_173),
.Y(n_176)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_179),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_152),
.B(n_126),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g201 ( 
.A1(n_180),
.A2(n_189),
.B(n_162),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_158),
.B(n_145),
.C(n_139),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_195),
.C(n_166),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_183),
.A2(n_149),
.B1(n_167),
.B2(n_172),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_169),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_184),
.Y(n_212)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_186),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_161),
.B(n_132),
.Y(n_188)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_188),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_140),
.B(n_144),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_135),
.Y(n_190)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_190),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_194),
.B(n_160),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_23),
.C(n_1),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_174),
.A2(n_181),
.B(n_180),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_211),
.Y(n_217)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_199),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_200),
.B(n_195),
.C(n_178),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_201),
.B(n_204),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_175),
.B(n_154),
.C(n_170),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_202),
.B(n_213),
.C(n_215),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_176),
.A2(n_163),
.B1(n_157),
.B2(n_150),
.Y(n_203)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_203),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g205 ( 
.A(n_183),
.Y(n_205)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_205),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_206),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_191),
.A2(n_23),
.B1(n_1),
.B2(n_2),
.Y(n_207)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_207),
.Y(n_229)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_0),
.C(n_2),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_185),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_214),
.A2(n_190),
.B1(n_192),
.B2(n_12),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_182),
.B(n_0),
.C(n_3),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_196),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_209),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_179),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_219),
.B(n_221),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_193),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_230),
.C(n_231),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_197),
.B(n_189),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_223),
.A2(n_214),
.B(n_4),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_206),
.B(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_224),
.B(n_215),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_204),
.B(n_187),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_210),
.B(n_185),
.C(n_188),
.Y(n_231)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_232),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_223),
.A2(n_205),
.B1(n_208),
.B2(n_212),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_233),
.A2(n_237),
.B1(n_238),
.B2(n_235),
.Y(n_259)
);

AOI21xp33_ASAP7_75t_L g234 ( 
.A1(n_217),
.A2(n_201),
.B(n_198),
.Y(n_234)
);

INVxp33_ASAP7_75t_L g257 ( 
.A(n_234),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_216),
.B(n_208),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_236),
.B(n_242),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_220),
.B1(n_228),
.B2(n_231),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_230),
.B(n_210),
.C(n_197),
.Y(n_238)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_238),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_240),
.B(n_241),
.Y(n_253)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_226),
.Y(n_241)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_226),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_247),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_225),
.B(n_213),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_245),
.B(n_4),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_246),
.A2(n_12),
.B(n_11),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_225),
.B(n_218),
.C(n_229),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_249),
.B(n_252),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_3),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_259),
.Y(n_266)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_247),
.B(n_12),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_4),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_255),
.B(n_256),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_5),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_258),
.B(n_5),
.Y(n_264)
);

AOI211xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_235),
.B(n_244),
.C(n_7),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_261),
.A2(n_263),
.B(n_265),
.Y(n_275)
);

NOR2xp67_ASAP7_75t_L g263 ( 
.A(n_257),
.B(n_244),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_264),
.B(n_10),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g265 ( 
.A(n_252),
.B(n_5),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_253),
.B(n_5),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_267),
.B(n_251),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_6),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.C(n_262),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_248),
.B(n_6),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_271),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_6),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_272),
.B(n_10),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_266),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_273),
.A2(n_275),
.B(n_9),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_8),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_276),
.C(n_8),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_260),
.B(n_8),
.Y(n_276)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_277),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_273),
.C(n_9),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_282),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_8),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_285),
.B(n_280),
.C(n_281),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_287),
.B(n_10),
.C(n_280),
.Y(n_288)
);


endmodule