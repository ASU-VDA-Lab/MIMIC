module fake_ariane_2358_n_1839 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1839);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1839;

wire n_913;
wire n_1681;
wire n_1507;
wire n_1486;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_645;
wire n_242;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_238;
wire n_365;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_851;
wire n_444;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_348;
wire n_552;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_604;
wire n_677;
wire n_439;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_727;
wire n_590;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_221;
wire n_321;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1429;
wire n_1324;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_166;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_978;
wire n_1011;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_485;
wire n_401;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_548;
wire n_289;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_484;
wire n_411;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_796;
wire n_573;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_131),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_99),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_45),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_18),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_50),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_76),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_116),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_75),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_61),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_12),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_86),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_118),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_156),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_17),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_110),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_45),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_111),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_80),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_112),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

BUFx3_ASAP7_75t_L g190 ( 
.A(n_84),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_81),
.Y(n_191)
);

INVx2_ASAP7_75t_SL g192 ( 
.A(n_44),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_6),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_141),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_49),
.Y(n_196)
);

BUFx10_ASAP7_75t_L g197 ( 
.A(n_25),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_128),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_51),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_104),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_66),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g202 ( 
.A(n_135),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_82),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_12),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_2),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_163),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_44),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_145),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_137),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_126),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_10),
.Y(n_212)
);

BUFx4f_ASAP7_75t_SL g213 ( 
.A(n_49),
.Y(n_213)
);

BUFx8_ASAP7_75t_SL g214 ( 
.A(n_40),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_122),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_40),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g217 ( 
.A(n_64),
.Y(n_217)
);

BUFx3_ASAP7_75t_L g218 ( 
.A(n_66),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_93),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_106),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_62),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_46),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_42),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_72),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_42),
.Y(n_225)
);

INVxp33_ASAP7_75t_R g226 ( 
.A(n_16),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_31),
.Y(n_227)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_120),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_102),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_150),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_27),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_89),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_32),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_132),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_31),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_20),
.Y(n_236)
);

BUFx2_ASAP7_75t_L g237 ( 
.A(n_125),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_164),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_71),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_18),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_70),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_90),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_20),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_56),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_3),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_114),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_6),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_157),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_119),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_136),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_24),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_139),
.Y(n_252)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_50),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_79),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_27),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_32),
.Y(n_256)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_96),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_103),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_59),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_62),
.Y(n_260)
);

BUFx3_ASAP7_75t_L g261 ( 
.A(n_24),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_108),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_107),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_23),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_11),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_23),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_9),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_127),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_92),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_59),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_100),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_61),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_41),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_52),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_140),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_48),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_39),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_95),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_67),
.Y(n_282)
);

INVx2_ASAP7_75t_SL g283 ( 
.A(n_57),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_17),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_134),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_28),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_109),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_25),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_53),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_85),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_51),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_159),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_83),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_133),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g295 ( 
.A(n_35),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_161),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_60),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_147),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_69),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_98),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_8),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_58),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_60),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_46),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_38),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_123),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_8),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_77),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_1),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_88),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_22),
.Y(n_311)
);

INVx2_ASAP7_75t_SL g312 ( 
.A(n_94),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_63),
.Y(n_313)
);

INVx2_ASAP7_75t_SL g314 ( 
.A(n_21),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_9),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_35),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_39),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_97),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_130),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_36),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_48),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_43),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_52),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_146),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_55),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_138),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_28),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_36),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_38),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_30),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_47),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_16),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_168),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_172),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_214),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_251),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_237),
.B(n_0),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_237),
.B(n_0),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_175),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_189),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_195),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_219),
.Y(n_342)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_172),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_168),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_271),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_300),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_179),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_179),
.Y(n_348)
);

INVxp67_ASAP7_75t_SL g349 ( 
.A(n_322),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_182),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_182),
.Y(n_351)
);

CKINVDCx16_ASAP7_75t_R g352 ( 
.A(n_251),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_318),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_188),
.Y(n_354)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_205),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_170),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g357 ( 
.A(n_199),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_199),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_192),
.B(n_2),
.Y(n_359)
);

INVx1_ASAP7_75t_SL g360 ( 
.A(n_253),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_235),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_171),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_273),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_188),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_275),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_198),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_198),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_203),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_176),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_203),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_177),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_183),
.Y(n_372)
);

NAND2xp33_ASAP7_75t_R g373 ( 
.A(n_167),
.B(n_142),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_209),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_209),
.Y(n_375)
);

INVx2_ASAP7_75t_L g376 ( 
.A(n_217),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_185),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_193),
.Y(n_378)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_231),
.B(n_4),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_196),
.Y(n_380)
);

INVxp67_ASAP7_75t_SL g381 ( 
.A(n_322),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_215),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_201),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_218),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_166),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_322),
.Y(n_386)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_212),
.Y(n_387)
);

INVxp67_ASAP7_75t_SL g388 ( 
.A(n_218),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_206),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_208),
.Y(n_390)
);

INVx2_ASAP7_75t_L g391 ( 
.A(n_217),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_215),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_229),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_216),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g395 ( 
.A(n_190),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_223),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_229),
.B(n_4),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_234),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_234),
.Y(n_399)
);

CKINVDCx16_ASAP7_75t_R g400 ( 
.A(n_178),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_190),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_225),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_190),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g404 ( 
.A(n_212),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_227),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_217),
.Y(n_406)
);

INVxp67_ASAP7_75t_SL g407 ( 
.A(n_261),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_239),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_239),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_249),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_202),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_233),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_236),
.Y(n_413)
);

NOR2xp67_ASAP7_75t_L g414 ( 
.A(n_192),
.B(n_5),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_202),
.Y(n_415)
);

OA21x2_ASAP7_75t_L g416 ( 
.A1(n_376),
.A2(n_274),
.B(n_249),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_333),
.Y(n_417)
);

AND2x4_ASAP7_75t_L g418 ( 
.A(n_333),
.B(n_261),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_344),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_347),
.B(n_274),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_376),
.Y(n_422)
);

BUFx2_ASAP7_75t_L g423 ( 
.A(n_360),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_347),
.B(n_281),
.Y(n_424)
);

INVx3_ASAP7_75t_L g425 ( 
.A(n_376),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_348),
.B(n_281),
.Y(n_426)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_391),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_391),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_348),
.B(n_350),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_350),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

AND2x4_ASAP7_75t_L g432 ( 
.A(n_351),
.B(n_283),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_354),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_354),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_391),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_406),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_336),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_364),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_406),
.Y(n_439)
);

OAI21x1_ASAP7_75t_L g440 ( 
.A1(n_397),
.A2(n_296),
.B(n_293),
.Y(n_440)
);

OAI21x1_ASAP7_75t_L g441 ( 
.A1(n_397),
.A2(n_296),
.B(n_293),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_364),
.B(n_326),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_341),
.Y(n_443)
);

AND2x4_ASAP7_75t_L g444 ( 
.A(n_366),
.B(n_283),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_366),
.Y(n_445)
);

INVx2_ASAP7_75t_L g446 ( 
.A(n_406),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_367),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_367),
.Y(n_448)
);

BUFx2_ASAP7_75t_L g449 ( 
.A(n_360),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_352),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_368),
.B(n_326),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_352),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_368),
.B(n_314),
.Y(n_453)
);

INVx2_ASAP7_75t_L g454 ( 
.A(n_370),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_370),
.B(n_282),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_374),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_374),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_375),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_375),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_382),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_382),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_392),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_392),
.Y(n_463)
);

NAND2xp33_ASAP7_75t_L g464 ( 
.A(n_337),
.B(n_217),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_393),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_345),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_393),
.B(n_282),
.Y(n_467)
);

INVx4_ASAP7_75t_L g468 ( 
.A(n_398),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_400),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_398),
.Y(n_470)
);

INVx3_ASAP7_75t_L g471 ( 
.A(n_399),
.Y(n_471)
);

INVx4_ASAP7_75t_L g472 ( 
.A(n_399),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_379),
.Y(n_473)
);

NAND2xp33_ASAP7_75t_L g474 ( 
.A(n_337),
.B(n_217),
.Y(n_474)
);

AND2x4_ASAP7_75t_L g475 ( 
.A(n_408),
.B(n_314),
.Y(n_475)
);

INVx3_ASAP7_75t_L g476 ( 
.A(n_408),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_353),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_409),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_409),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_349),
.B(n_312),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_410),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_410),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_379),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_400),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_381),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_386),
.B(n_312),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_388),
.Y(n_487)
);

INVx6_ASAP7_75t_L g488 ( 
.A(n_373),
.Y(n_488)
);

INVxp33_ASAP7_75t_SL g489 ( 
.A(n_335),
.Y(n_489)
);

BUFx8_ASAP7_75t_L g490 ( 
.A(n_385),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_338),
.Y(n_491)
);

INVx3_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

INVx4_ASAP7_75t_L g493 ( 
.A(n_488),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_470),
.Y(n_494)
);

INVxp33_ASAP7_75t_SL g495 ( 
.A(n_443),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_425),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_356),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_480),
.B(n_362),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_425),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_369),
.Y(n_500)
);

INVx8_ASAP7_75t_L g501 ( 
.A(n_491),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_473),
.B(n_486),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_425),
.Y(n_503)
);

INVx4_ASAP7_75t_SL g504 ( 
.A(n_470),
.Y(n_504)
);

NAND3xp33_ASAP7_75t_L g505 ( 
.A(n_491),
.B(n_372),
.C(n_371),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_443),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_484),
.B(n_377),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_425),
.Y(n_508)
);

OAI22xp5_ASAP7_75t_L g509 ( 
.A1(n_473),
.A2(n_359),
.B1(n_414),
.B2(n_327),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_423),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_L g511 ( 
.A(n_485),
.B(n_378),
.Y(n_511)
);

INVx4_ASAP7_75t_L g512 ( 
.A(n_488),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_487),
.B(n_380),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_473),
.B(n_383),
.Y(n_514)
);

AOI22xp33_ASAP7_75t_L g515 ( 
.A1(n_488),
.A2(n_359),
.B1(n_414),
.B2(n_401),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_425),
.Y(n_516)
);

BUFx3_ASAP7_75t_L g517 ( 
.A(n_488),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_427),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_487),
.B(n_389),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_470),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_470),
.Y(n_521)
);

INVx4_ASAP7_75t_L g522 ( 
.A(n_488),
.Y(n_522)
);

INVx4_ASAP7_75t_SL g523 ( 
.A(n_470),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_473),
.B(n_390),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_427),
.Y(n_525)
);

OR2x6_ASAP7_75t_L g526 ( 
.A(n_473),
.B(n_334),
.Y(n_526)
);

BUFx3_ASAP7_75t_L g527 ( 
.A(n_488),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_470),
.Y(n_528)
);

AO21x2_ASAP7_75t_L g529 ( 
.A1(n_440),
.A2(n_250),
.B(n_181),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_427),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_473),
.B(n_394),
.Y(n_531)
);

XOR2xp5_ASAP7_75t_L g532 ( 
.A(n_469),
.B(n_339),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_477),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_491),
.B(n_396),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_470),
.Y(n_535)
);

NAND3xp33_ASAP7_75t_L g536 ( 
.A(n_491),
.B(n_405),
.C(n_402),
.Y(n_536)
);

AOI22xp5_ASAP7_75t_L g537 ( 
.A1(n_491),
.A2(n_295),
.B1(n_297),
.B2(n_240),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_432),
.B(n_407),
.Y(n_538)
);

AOI22xp33_ASAP7_75t_L g539 ( 
.A1(n_491),
.A2(n_444),
.B1(n_453),
.B2(n_432),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_471),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_471),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_427),
.Y(n_542)
);

BUFx3_ASAP7_75t_L g543 ( 
.A(n_471),
.Y(n_543)
);

INVx2_ASAP7_75t_SL g544 ( 
.A(n_423),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_428),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_486),
.B(n_412),
.Y(n_546)
);

AND2x2_ASAP7_75t_L g547 ( 
.A(n_423),
.B(n_384),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_468),
.B(n_413),
.Y(n_548)
);

NAND3xp33_ASAP7_75t_L g549 ( 
.A(n_491),
.B(n_357),
.C(n_343),
.Y(n_549)
);

INVx2_ASAP7_75t_SL g550 ( 
.A(n_449),
.Y(n_550)
);

BUFx6f_ASAP7_75t_L g551 ( 
.A(n_422),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_471),
.Y(n_552)
);

INVx4_ASAP7_75t_L g553 ( 
.A(n_471),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_476),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_449),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_491),
.A2(n_415),
.B1(n_411),
.B2(n_403),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_476),
.Y(n_557)
);

AOI22xp33_ASAP7_75t_L g558 ( 
.A1(n_432),
.A2(n_395),
.B1(n_279),
.B2(n_256),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g559 ( 
.A(n_449),
.B(n_358),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_468),
.B(n_387),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_476),
.Y(n_561)
);

INVx2_ASAP7_75t_SL g562 ( 
.A(n_484),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_484),
.B(n_197),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_450),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_484),
.B(n_404),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_484),
.B(n_468),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_476),
.Y(n_567)
);

INVx4_ASAP7_75t_SL g568 ( 
.A(n_422),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_476),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_481),
.Y(n_570)
);

INVx5_ASAP7_75t_L g571 ( 
.A(n_422),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_477),
.Y(n_572)
);

BUFx6f_ASAP7_75t_L g573 ( 
.A(n_422),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_481),
.Y(n_574)
);

INVx2_ASAP7_75t_L g575 ( 
.A(n_428),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g576 ( 
.A1(n_483),
.A2(n_267),
.B1(n_265),
.B2(n_284),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_428),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_468),
.B(n_340),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_481),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_481),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_481),
.Y(n_581)
);

INVx3_ASAP7_75t_L g582 ( 
.A(n_468),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_428),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_466),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_472),
.B(n_342),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_454),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_454),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_436),
.Y(n_588)
);

BUFx4f_ASAP7_75t_L g589 ( 
.A(n_416),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_436),
.Y(n_590)
);

INVx6_ASAP7_75t_L g591 ( 
.A(n_472),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_429),
.B(n_197),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_472),
.B(n_346),
.Y(n_593)
);

INVxp67_ASAP7_75t_SL g594 ( 
.A(n_429),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_472),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_436),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_436),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_469),
.B(n_221),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g599 ( 
.A(n_472),
.B(n_238),
.Y(n_599)
);

AND2x6_ASAP7_75t_L g600 ( 
.A(n_454),
.B(n_202),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_417),
.B(n_169),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_446),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_446),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_454),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_417),
.B(n_419),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_457),
.Y(n_606)
);

AOI22xp33_ASAP7_75t_L g607 ( 
.A1(n_432),
.A2(n_279),
.B1(n_231),
.B2(n_256),
.Y(n_607)
);

AOI22xp33_ASAP7_75t_L g608 ( 
.A1(n_432),
.A2(n_268),
.B1(n_332),
.B2(n_331),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_SL g609 ( 
.A(n_483),
.B(n_197),
.Y(n_609)
);

INVx1_ASAP7_75t_SL g610 ( 
.A(n_450),
.Y(n_610)
);

INVx3_ASAP7_75t_L g611 ( 
.A(n_457),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_444),
.B(n_197),
.Y(n_612)
);

NOR3xp33_ASAP7_75t_L g613 ( 
.A(n_452),
.B(n_222),
.C(n_221),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_444),
.A2(n_269),
.B1(n_332),
.B2(n_331),
.Y(n_614)
);

INVxp33_ASAP7_75t_L g615 ( 
.A(n_437),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_446),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_SL g617 ( 
.A1(n_421),
.A2(n_288),
.B1(n_291),
.B2(n_329),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_457),
.Y(n_618)
);

NOR2xp33_ASAP7_75t_L g619 ( 
.A(n_419),
.B(n_420),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_446),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_457),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_461),
.Y(n_622)
);

INVx3_ASAP7_75t_L g623 ( 
.A(n_461),
.Y(n_623)
);

AOI22xp5_ASAP7_75t_L g624 ( 
.A1(n_464),
.A2(n_259),
.B1(n_255),
.B2(n_301),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_461),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_461),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_462),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_420),
.B(n_173),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_464),
.A2(n_245),
.B1(n_260),
.B2(n_328),
.Y(n_629)
);

OR2x6_ASAP7_75t_L g630 ( 
.A(n_444),
.B(n_222),
.Y(n_630)
);

INVx2_ASAP7_75t_SL g631 ( 
.A(n_452),
.Y(n_631)
);

OAI22xp33_ASAP7_75t_L g632 ( 
.A1(n_437),
.A2(n_302),
.B1(n_313),
.B2(n_303),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_462),
.Y(n_633)
);

BUFx3_ASAP7_75t_L g634 ( 
.A(n_430),
.Y(n_634)
);

NOR2xp33_ASAP7_75t_L g635 ( 
.A(n_430),
.B(n_431),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_431),
.B(n_174),
.Y(n_636)
);

INVx3_ASAP7_75t_L g637 ( 
.A(n_462),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_462),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_465),
.Y(n_639)
);

BUFx4f_ASAP7_75t_L g640 ( 
.A(n_416),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_465),
.Y(n_641)
);

OAI22x1_ASAP7_75t_L g642 ( 
.A1(n_444),
.A2(n_226),
.B1(n_307),
.B2(n_304),
.Y(n_642)
);

AOI22xp5_ASAP7_75t_L g643 ( 
.A1(n_474),
.A2(n_311),
.B1(n_325),
.B2(n_213),
.Y(n_643)
);

INVx2_ASAP7_75t_SL g644 ( 
.A(n_453),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_594),
.B(n_433),
.Y(n_645)
);

AND2x2_ASAP7_75t_L g646 ( 
.A(n_544),
.B(n_453),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_544),
.B(n_418),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_565),
.B(n_433),
.Y(n_648)
);

AND2x6_ASAP7_75t_L g649 ( 
.A(n_517),
.B(n_453),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_634),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_546),
.B(n_434),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_502),
.B(n_592),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_592),
.B(n_434),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_634),
.Y(n_654)
);

INVx2_ASAP7_75t_SL g655 ( 
.A(n_550),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_534),
.B(n_438),
.Y(n_656)
);

INVx8_ASAP7_75t_L g657 ( 
.A(n_526),
.Y(n_657)
);

NOR3xp33_ASAP7_75t_L g658 ( 
.A(n_506),
.B(n_572),
.C(n_533),
.Y(n_658)
);

INVx2_ASAP7_75t_SL g659 ( 
.A(n_550),
.Y(n_659)
);

NAND3xp33_ASAP7_75t_L g660 ( 
.A(n_500),
.B(n_474),
.C(n_467),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_L g661 ( 
.A(n_644),
.B(n_438),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_644),
.B(n_445),
.Y(n_662)
);

AND2x4_ASAP7_75t_L g663 ( 
.A(n_555),
.B(n_418),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_540),
.Y(n_664)
);

AND2x4_ASAP7_75t_L g665 ( 
.A(n_538),
.B(n_418),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_611),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_511),
.B(n_445),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_559),
.B(n_453),
.Y(n_668)
);

INVxp67_ASAP7_75t_L g669 ( 
.A(n_564),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_SL g670 ( 
.A(n_584),
.B(n_489),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_611),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_540),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_541),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_611),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_497),
.B(n_447),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_513),
.B(n_447),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_519),
.B(n_448),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_493),
.B(n_448),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_498),
.B(n_456),
.Y(n_679)
);

INVx2_ASAP7_75t_SL g680 ( 
.A(n_631),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_623),
.Y(n_681)
);

NOR2x1p5_ASAP7_75t_L g682 ( 
.A(n_584),
.B(n_506),
.Y(n_682)
);

HB1xp67_ASAP7_75t_L g683 ( 
.A(n_610),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_493),
.B(n_456),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_493),
.B(n_458),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_562),
.B(n_458),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_623),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_514),
.B(n_459),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_533),
.Y(n_689)
);

INVx8_ASAP7_75t_L g690 ( 
.A(n_526),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_562),
.B(n_538),
.Y(n_691)
);

NOR2xp67_ASAP7_75t_SL g692 ( 
.A(n_512),
.B(n_243),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_543),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_538),
.B(n_459),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_554),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_623),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_512),
.B(n_522),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_589),
.A2(n_416),
.B1(n_475),
.B2(n_440),
.Y(n_698)
);

NAND2x1p5_ASAP7_75t_L g699 ( 
.A(n_512),
.B(n_460),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_566),
.B(n_460),
.Y(n_700)
);

BUFx6f_ASAP7_75t_SL g701 ( 
.A(n_631),
.Y(n_701)
);

INVx3_ASAP7_75t_L g702 ( 
.A(n_553),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_554),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_SL g704 ( 
.A(n_522),
.B(n_463),
.Y(n_704)
);

INVx8_ASAP7_75t_L g705 ( 
.A(n_526),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_522),
.B(n_463),
.Y(n_706)
);

BUFx2_ASAP7_75t_L g707 ( 
.A(n_510),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_557),
.Y(n_708)
);

AOI21xp5_ASAP7_75t_L g709 ( 
.A1(n_501),
.A2(n_467),
.B(n_455),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_539),
.B(n_560),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_557),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_537),
.A2(n_475),
.B1(n_455),
.B2(n_418),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_619),
.B(n_478),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_637),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_635),
.B(n_478),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_561),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_524),
.B(n_475),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_537),
.A2(n_440),
.B(n_441),
.C(n_482),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_589),
.A2(n_416),
.B1(n_475),
.B2(n_441),
.Y(n_719)
);

NOR2xp67_ASAP7_75t_L g720 ( 
.A(n_572),
.B(n_421),
.Y(n_720)
);

INVxp67_ASAP7_75t_L g721 ( 
.A(n_564),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_637),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_589),
.A2(n_416),
.B1(n_475),
.B2(n_441),
.Y(n_723)
);

NAND2xp33_ASAP7_75t_L g724 ( 
.A(n_501),
.B(n_465),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_547),
.B(n_615),
.Y(n_725)
);

O2A1O1Ixp33_ASAP7_75t_L g726 ( 
.A1(n_605),
.A2(n_465),
.B(n_479),
.C(n_482),
.Y(n_726)
);

NOR3xp33_ASAP7_75t_L g727 ( 
.A(n_578),
.B(n_244),
.C(n_243),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_640),
.A2(n_416),
.B1(n_479),
.B2(n_482),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_561),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_517),
.B(n_479),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_531),
.B(n_418),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_567),
.Y(n_732)
);

BUFx3_ASAP7_75t_L g733 ( 
.A(n_543),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_552),
.B(n_479),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_552),
.B(n_482),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_567),
.Y(n_736)
);

NOR2xp33_ASAP7_75t_R g737 ( 
.A(n_510),
.B(n_490),
.Y(n_737)
);

OR2x6_ASAP7_75t_L g738 ( 
.A(n_526),
.B(n_490),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_547),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_527),
.B(n_585),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_637),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_509),
.A2(n_424),
.B1(n_451),
.B2(n_442),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_621),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_621),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_527),
.B(n_553),
.Y(n_745)
);

INVxp67_ASAP7_75t_L g746 ( 
.A(n_532),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_552),
.B(n_424),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_L g748 ( 
.A(n_548),
.B(n_426),
.Y(n_748)
);

AOI22xp33_ASAP7_75t_L g749 ( 
.A1(n_640),
.A2(n_426),
.B1(n_442),
.B2(n_451),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_630),
.B(n_244),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_R g751 ( 
.A(n_593),
.B(n_490),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_574),
.B(n_247),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_626),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_574),
.B(n_247),
.Y(n_754)
);

NOR3xp33_ASAP7_75t_L g755 ( 
.A(n_632),
.B(n_276),
.C(n_289),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_SL g756 ( 
.A(n_553),
.B(n_489),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_626),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_574),
.B(n_262),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_582),
.B(n_262),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_507),
.B(n_263),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_569),
.Y(n_761)
);

AOI22xp5_ASAP7_75t_L g762 ( 
.A1(n_630),
.A2(n_211),
.B1(n_210),
.B2(n_324),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_640),
.A2(n_305),
.B1(n_263),
.B2(n_268),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_SL g764 ( 
.A(n_569),
.B(n_181),
.Y(n_764)
);

O2A1O1Ixp5_ASAP7_75t_L g765 ( 
.A1(n_599),
.A2(n_276),
.B(n_289),
.C(n_286),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_551),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_630),
.A2(n_204),
.B1(n_186),
.B2(n_184),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_582),
.B(n_269),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_582),
.B(n_270),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_591),
.Y(n_770)
);

NOR2xp67_ASAP7_75t_L g771 ( 
.A(n_505),
.B(n_180),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_641),
.Y(n_772)
);

INVxp67_ASAP7_75t_L g773 ( 
.A(n_598),
.Y(n_773)
);

NOR2xp33_ASAP7_75t_L g774 ( 
.A(n_612),
.B(n_270),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_SL g775 ( 
.A(n_570),
.B(n_250),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_570),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_595),
.B(n_277),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_SL g778 ( 
.A(n_515),
.B(n_490),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_608),
.A2(n_614),
.B1(n_558),
.B2(n_607),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_579),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_595),
.B(n_277),
.Y(n_781)
);

BUFx4_ASAP7_75t_L g782 ( 
.A(n_495),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_SL g783 ( 
.A(n_495),
.B(n_490),
.Y(n_783)
);

OAI22xp5_ASAP7_75t_L g784 ( 
.A1(n_549),
.A2(n_315),
.B1(n_316),
.B2(n_280),
.Y(n_784)
);

NAND2xp33_ASAP7_75t_L g785 ( 
.A(n_501),
.B(n_217),
.Y(n_785)
);

AO21x2_ASAP7_75t_L g786 ( 
.A1(n_529),
.A2(n_315),
.B(n_280),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_579),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_536),
.B(n_187),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_L g789 ( 
.A(n_595),
.B(n_286),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_630),
.A2(n_191),
.B1(n_194),
.B2(n_200),
.Y(n_790)
);

OAI22xp33_ASAP7_75t_L g791 ( 
.A1(n_629),
.A2(n_317),
.B1(n_305),
.B2(n_309),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_580),
.B(n_309),
.Y(n_792)
);

OR2x2_ASAP7_75t_L g793 ( 
.A(n_598),
.B(n_355),
.Y(n_793)
);

NOR3xp33_ASAP7_75t_L g794 ( 
.A(n_617),
.B(n_316),
.C(n_317),
.Y(n_794)
);

NOR2x1p5_ASAP7_75t_L g795 ( 
.A(n_601),
.B(n_320),
.Y(n_795)
);

BUFx5_ASAP7_75t_L g796 ( 
.A(n_580),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_581),
.B(n_628),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_556),
.B(n_361),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_609),
.B(n_563),
.Y(n_799)
);

AOI22xp33_ASAP7_75t_SL g800 ( 
.A1(n_642),
.A2(n_363),
.B1(n_365),
.B2(n_600),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_581),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_586),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_591),
.B(n_320),
.Y(n_803)
);

NAND2xp33_ASAP7_75t_L g804 ( 
.A(n_501),
.B(n_323),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_L g805 ( 
.A(n_636),
.B(n_321),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_551),
.B(n_257),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_586),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_591),
.B(n_321),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_587),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_591),
.B(n_587),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_604),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_604),
.A2(n_330),
.B1(n_230),
.B2(n_178),
.Y(n_812)
);

AOI21x1_ASAP7_75t_L g813 ( 
.A1(n_730),
.A2(n_618),
.B(n_606),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_675),
.B(n_629),
.Y(n_814)
);

OAI22xp5_ASAP7_75t_L g815 ( 
.A1(n_667),
.A2(n_576),
.B1(n_622),
.B2(n_639),
.Y(n_815)
);

O2A1O1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_652),
.A2(n_618),
.B(n_606),
.C(n_622),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_676),
.A2(n_633),
.B1(n_625),
.B2(n_639),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_656),
.A2(n_521),
.B(n_494),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_702),
.B(n_551),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_700),
.A2(n_521),
.B(n_494),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_702),
.B(n_551),
.Y(n_821)
);

OAI21xp5_ASAP7_75t_L g822 ( 
.A1(n_698),
.A2(n_627),
.B(n_625),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_675),
.B(n_613),
.Y(n_823)
);

AOI21xp5_ASAP7_75t_L g824 ( 
.A1(n_745),
.A2(n_535),
.B(n_528),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_745),
.A2(n_535),
.B(n_528),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_651),
.B(n_627),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_651),
.B(n_633),
.Y(n_827)
);

O2A1O1Ixp33_ASAP7_75t_L g828 ( 
.A1(n_677),
.A2(n_638),
.B(n_641),
.C(n_503),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_748),
.B(n_638),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_748),
.B(n_624),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_664),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_653),
.A2(n_496),
.B(n_516),
.C(n_499),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_725),
.B(n_642),
.Y(n_833)
);

BUFx6f_ASAP7_75t_L g834 ( 
.A(n_766),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_SL g835 ( 
.A(n_796),
.B(n_551),
.Y(n_835)
);

AOI21x1_ASAP7_75t_L g836 ( 
.A1(n_730),
.A2(n_575),
.B(n_620),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_678),
.A2(n_492),
.B(n_520),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_679),
.B(n_643),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_665),
.B(n_504),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_678),
.A2(n_492),
.B(n_520),
.Y(n_840)
);

AOI22xp5_ASAP7_75t_L g841 ( 
.A1(n_727),
.A2(n_492),
.B1(n_520),
.B2(n_600),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_684),
.A2(n_573),
.B(n_499),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_646),
.B(n_496),
.Y(n_843)
);

OAI21xp33_ASAP7_75t_SL g844 ( 
.A1(n_688),
.A2(n_503),
.B(n_508),
.Y(n_844)
);

INVxp67_ASAP7_75t_L g845 ( 
.A(n_683),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_739),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_668),
.B(n_508),
.Y(n_847)
);

INVxp67_ASAP7_75t_L g848 ( 
.A(n_707),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_688),
.B(n_516),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_694),
.B(n_518),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_689),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_655),
.B(n_518),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_648),
.A2(n_330),
.B1(n_573),
.B2(n_603),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_749),
.B(n_525),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_684),
.A2(n_573),
.B(n_529),
.Y(n_855)
);

NOR2xp33_ASAP7_75t_SL g856 ( 
.A(n_670),
.B(n_178),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_685),
.A2(n_573),
.B(n_529),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_749),
.B(n_665),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_720),
.B(n_620),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_663),
.B(n_525),
.Y(n_860)
);

AOI22xp33_ASAP7_75t_L g861 ( 
.A1(n_763),
.A2(n_600),
.B1(n_616),
.B2(n_602),
.Y(n_861)
);

OAI21xp5_ASAP7_75t_L g862 ( 
.A1(n_698),
.A2(n_616),
.B(n_603),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_796),
.B(n_573),
.Y(n_863)
);

AOI21x1_ASAP7_75t_L g864 ( 
.A1(n_692),
.A2(n_602),
.B(n_530),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_663),
.B(n_530),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_666),
.Y(n_866)
);

INVx2_ASAP7_75t_SL g867 ( 
.A(n_782),
.Y(n_867)
);

AOI21x1_ASAP7_75t_L g868 ( 
.A1(n_685),
.A2(n_706),
.B(n_704),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_704),
.A2(n_571),
.B(n_597),
.Y(n_869)
);

OAI21xp33_ASAP7_75t_L g870 ( 
.A1(n_717),
.A2(n_323),
.B(n_597),
.Y(n_870)
);

OR2x2_ASAP7_75t_L g871 ( 
.A(n_793),
.B(n_542),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_706),
.A2(n_571),
.B(n_596),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_672),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_666),
.Y(n_874)
);

AOI22x1_ASAP7_75t_L g875 ( 
.A1(n_709),
.A2(n_577),
.B1(n_596),
.B2(n_590),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_671),
.Y(n_876)
);

AND2x2_ASAP7_75t_L g877 ( 
.A(n_773),
.B(n_542),
.Y(n_877)
);

BUFx3_ASAP7_75t_L g878 ( 
.A(n_680),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_659),
.B(n_545),
.Y(n_879)
);

CKINVDCx20_ASAP7_75t_R g880 ( 
.A(n_737),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_797),
.A2(n_571),
.B(n_590),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_691),
.B(n_545),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_671),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_669),
.B(n_575),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_721),
.B(n_746),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_658),
.B(n_798),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_750),
.B(n_577),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_803),
.B(n_583),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_803),
.B(n_583),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_697),
.A2(n_571),
.B(n_588),
.Y(n_890)
);

AOI21xp5_ASAP7_75t_L g891 ( 
.A1(n_747),
.A2(n_571),
.B(n_588),
.Y(n_891)
);

NAND2x1p5_ASAP7_75t_L g892 ( 
.A(n_693),
.B(n_571),
.Y(n_892)
);

OAI21xp5_ASAP7_75t_L g893 ( 
.A1(n_719),
.A2(n_600),
.B(n_504),
.Y(n_893)
);

INVx2_ASAP7_75t_L g894 ( 
.A(n_674),
.Y(n_894)
);

INVx1_ASAP7_75t_SL g895 ( 
.A(n_737),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_713),
.B(n_600),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_715),
.B(n_600),
.Y(n_897)
);

NOR2xp33_ASAP7_75t_L g898 ( 
.A(n_647),
.B(n_5),
.Y(n_898)
);

AOI22xp5_ASAP7_75t_L g899 ( 
.A1(n_657),
.A2(n_600),
.B1(n_504),
.B2(n_523),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_799),
.B(n_7),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_742),
.B(n_504),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_673),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_766),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_760),
.A2(n_228),
.B(n_323),
.C(n_422),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_695),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_719),
.A2(n_523),
.B(n_272),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_645),
.B(n_523),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_724),
.A2(n_266),
.B(n_224),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_SL g909 ( 
.A(n_783),
.B(n_178),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_731),
.B(n_523),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_810),
.A2(n_278),
.B(n_220),
.Y(n_911)
);

AND2x2_ASAP7_75t_L g912 ( 
.A(n_750),
.B(n_230),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_734),
.A2(n_287),
.B(n_232),
.Y(n_913)
);

BUFx4f_ASAP7_75t_L g914 ( 
.A(n_738),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_731),
.B(n_568),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_681),
.Y(n_916)
);

OAI22xp5_ASAP7_75t_L g917 ( 
.A1(n_661),
.A2(n_323),
.B1(n_228),
.B2(n_207),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_796),
.B(n_568),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_779),
.B(n_568),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_735),
.A2(n_290),
.B(n_246),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_686),
.A2(n_292),
.B(n_248),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_657),
.A2(n_294),
.B1(n_241),
.B2(n_242),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_681),
.Y(n_923)
);

NOR3xp33_ASAP7_75t_L g924 ( 
.A(n_755),
.B(n_228),
.C(n_252),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_690),
.A2(n_306),
.B1(n_254),
.B2(n_258),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_779),
.B(n_568),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_796),
.B(n_435),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_662),
.A2(n_308),
.B(n_264),
.Y(n_928)
);

BUFx6f_ASAP7_75t_L g929 ( 
.A(n_766),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_687),
.Y(n_930)
);

AOI21xp5_ASAP7_75t_L g931 ( 
.A1(n_687),
.A2(n_310),
.B(n_285),
.Y(n_931)
);

AND2x4_ASAP7_75t_L g932 ( 
.A(n_738),
.B(n_435),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_791),
.A2(n_756),
.B(n_777),
.C(n_781),
.Y(n_933)
);

O2A1O1Ixp33_ASAP7_75t_L g934 ( 
.A1(n_756),
.A2(n_7),
.B(n_10),
.C(n_13),
.Y(n_934)
);

A2O1A1Ixp33_ASAP7_75t_L g935 ( 
.A1(n_760),
.A2(n_323),
.B(n_435),
.C(n_422),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_759),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_696),
.A2(n_319),
.B(n_298),
.Y(n_937)
);

AOI21xp33_ASAP7_75t_L g938 ( 
.A1(n_763),
.A2(n_299),
.B(n_435),
.Y(n_938)
);

AND2x6_ASAP7_75t_SL g939 ( 
.A(n_738),
.B(n_14),
.Y(n_939)
);

NOR2xp33_ASAP7_75t_L g940 ( 
.A(n_799),
.B(n_15),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_690),
.Y(n_941)
);

INVx2_ASAP7_75t_L g942 ( 
.A(n_696),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_712),
.B(n_323),
.Y(n_943)
);

NOR3xp33_ASAP7_75t_L g944 ( 
.A(n_794),
.B(n_805),
.C(n_765),
.Y(n_944)
);

OAI22xp5_ASAP7_75t_L g945 ( 
.A1(n_710),
.A2(n_439),
.B1(n_435),
.B2(n_422),
.Y(n_945)
);

NOR2xp33_ASAP7_75t_L g946 ( 
.A(n_650),
.B(n_19),
.Y(n_946)
);

AOI21xp5_ASAP7_75t_L g947 ( 
.A1(n_714),
.A2(n_439),
.B(n_435),
.Y(n_947)
);

BUFx6f_ASAP7_75t_L g948 ( 
.A(n_766),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_751),
.B(n_230),
.Y(n_949)
);

OAI21xp5_ASAP7_75t_L g950 ( 
.A1(n_723),
.A2(n_439),
.B(n_435),
.Y(n_950)
);

HB1xp67_ASAP7_75t_L g951 ( 
.A(n_690),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_703),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_796),
.B(n_699),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_714),
.A2(n_439),
.B(n_435),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_654),
.B(n_774),
.Y(n_955)
);

NOR2xp33_ASAP7_75t_L g956 ( 
.A(n_705),
.B(n_778),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_722),
.A2(n_439),
.B(n_422),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_722),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_774),
.B(n_230),
.Y(n_959)
);

AOI21xp5_ASAP7_75t_L g960 ( 
.A1(n_741),
.A2(n_785),
.B(n_804),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_741),
.A2(n_439),
.B(n_257),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_705),
.B(n_19),
.Y(n_962)
);

O2A1O1Ixp33_ASAP7_75t_L g963 ( 
.A1(n_768),
.A2(n_21),
.B(n_22),
.C(n_26),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_705),
.B(n_26),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_649),
.B(n_29),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_708),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_693),
.Y(n_967)
);

BUFx2_ASAP7_75t_L g968 ( 
.A(n_751),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_711),
.A2(n_439),
.B(n_257),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_716),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_729),
.A2(n_439),
.B(n_257),
.Y(n_971)
);

AOI21xp5_ASAP7_75t_L g972 ( 
.A1(n_732),
.A2(n_257),
.B(n_87),
.Y(n_972)
);

INVx3_ASAP7_75t_L g973 ( 
.A(n_733),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_736),
.A2(n_257),
.B(n_78),
.Y(n_974)
);

BUFx6f_ASAP7_75t_L g975 ( 
.A(n_733),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_649),
.Y(n_976)
);

INVx2_ASAP7_75t_SL g977 ( 
.A(n_682),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_649),
.B(n_29),
.Y(n_978)
);

A2O1A1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_660),
.A2(n_30),
.B(n_33),
.C(n_34),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_761),
.Y(n_980)
);

AOI21xp5_ASAP7_75t_L g981 ( 
.A1(n_776),
.A2(n_91),
.B(n_162),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_649),
.B(n_33),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_780),
.Y(n_983)
);

O2A1O1Ixp33_ASAP7_75t_L g984 ( 
.A1(n_769),
.A2(n_34),
.B(n_37),
.C(n_41),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_649),
.B(n_812),
.Y(n_985)
);

AOI21xp5_ASAP7_75t_L g986 ( 
.A1(n_787),
.A2(n_105),
.B(n_160),
.Y(n_986)
);

OAI21xp5_ASAP7_75t_L g987 ( 
.A1(n_723),
.A2(n_101),
.B(n_154),
.Y(n_987)
);

INVx2_ASAP7_75t_SL g988 ( 
.A(n_795),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_812),
.B(n_37),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_770),
.Y(n_990)
);

BUFx2_ASAP7_75t_L g991 ( 
.A(n_808),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_770),
.Y(n_992)
);

AND2x2_ASAP7_75t_SL g993 ( 
.A(n_728),
.B(n_43),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_801),
.A2(n_789),
.B(n_809),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_752),
.B(n_47),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_802),
.A2(n_113),
.B(n_153),
.Y(n_996)
);

NAND2xp5_ASAP7_75t_L g997 ( 
.A(n_754),
.B(n_53),
.Y(n_997)
);

OAI21xp5_ASAP7_75t_L g998 ( 
.A1(n_718),
.A2(n_117),
.B(n_152),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_807),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_758),
.B(n_54),
.Y(n_1000)
);

INVxp67_ASAP7_75t_L g1001 ( 
.A(n_701),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_823),
.B(n_800),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_814),
.B(n_762),
.Y(n_1003)
);

BUFx2_ASAP7_75t_L g1004 ( 
.A(n_845),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_830),
.A2(n_767),
.B1(n_790),
.B2(n_699),
.Y(n_1005)
);

O2A1O1Ixp33_ASAP7_75t_L g1006 ( 
.A1(n_900),
.A2(n_792),
.B(n_726),
.C(n_764),
.Y(n_1006)
);

INVx2_ASAP7_75t_SL g1007 ( 
.A(n_851),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_829),
.A2(n_740),
.B(n_788),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_877),
.B(n_900),
.Y(n_1009)
);

BUFx6f_ASAP7_75t_L g1010 ( 
.A(n_941),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_831),
.Y(n_1011)
);

BUFx3_ASAP7_75t_L g1012 ( 
.A(n_867),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_846),
.B(n_784),
.Y(n_1013)
);

NOR2xp33_ASAP7_75t_L g1014 ( 
.A(n_885),
.B(n_701),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_940),
.B(n_811),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_940),
.B(n_884),
.Y(n_1016)
);

NOR2xp33_ASAP7_75t_L g1017 ( 
.A(n_848),
.B(n_856),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_848),
.B(n_772),
.Y(n_1018)
);

AO32x2_ASAP7_75t_L g1019 ( 
.A1(n_945),
.A2(n_786),
.A3(n_728),
.B1(n_764),
.B2(n_775),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_826),
.A2(n_775),
.B(n_744),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_976),
.B(n_796),
.Y(n_1021)
);

INVx2_ASAP7_75t_L g1022 ( 
.A(n_866),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_880),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_846),
.B(n_757),
.Y(n_1024)
);

INVx3_ASAP7_75t_L g1025 ( 
.A(n_976),
.Y(n_1025)
);

AOI22xp5_ASAP7_75t_L g1026 ( 
.A1(n_993),
.A2(n_771),
.B1(n_743),
.B2(n_772),
.Y(n_1026)
);

BUFx2_ASAP7_75t_SL g1027 ( 
.A(n_977),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_L g1028 ( 
.A(n_884),
.B(n_757),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_878),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_874),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_876),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_967),
.Y(n_1032)
);

A2O1A1Ixp33_ASAP7_75t_L g1033 ( 
.A1(n_987),
.A2(n_753),
.B(n_744),
.C(n_743),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_895),
.B(n_753),
.Y(n_1034)
);

BUFx12f_ASAP7_75t_L g1035 ( 
.A(n_939),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_967),
.Y(n_1036)
);

A2O1A1Ixp33_ASAP7_75t_L g1037 ( 
.A1(n_933),
.A2(n_806),
.B(n_786),
.C(n_56),
.Y(n_1037)
);

O2A1O1Ixp33_ASAP7_75t_L g1038 ( 
.A1(n_979),
.A2(n_806),
.B(n_55),
.C(n_57),
.Y(n_1038)
);

CKINVDCx20_ASAP7_75t_R g1039 ( 
.A(n_1001),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_838),
.A2(n_54),
.B(n_58),
.C(n_63),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_898),
.B(n_64),
.Y(n_1041)
);

OAI22xp5_ASAP7_75t_L g1042 ( 
.A1(n_993),
.A2(n_65),
.B1(n_68),
.B2(n_73),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_827),
.A2(n_65),
.B(n_129),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_898),
.B(n_991),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_873),
.Y(n_1045)
);

AOI22x1_ASAP7_75t_L g1046 ( 
.A1(n_994),
.A2(n_143),
.B1(n_148),
.B2(n_149),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_883),
.Y(n_1047)
);

INVx2_ASAP7_75t_L g1048 ( 
.A(n_894),
.Y(n_1048)
);

AND2x6_ASAP7_75t_L g1049 ( 
.A(n_976),
.B(n_151),
.Y(n_1049)
);

AOI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_849),
.A2(n_165),
.B(n_998),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_886),
.B(n_912),
.Y(n_1051)
);

O2A1O1Ixp33_ASAP7_75t_L g1052 ( 
.A1(n_815),
.A2(n_944),
.B(n_989),
.C(n_858),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_924),
.A2(n_946),
.B(n_959),
.C(n_955),
.Y(n_1053)
);

BUFx2_ASAP7_75t_L g1054 ( 
.A(n_962),
.Y(n_1054)
);

O2A1O1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_944),
.A2(n_936),
.B(n_984),
.C(n_963),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_L g1056 ( 
.A(n_871),
.B(n_968),
.Y(n_1056)
);

AND2x4_ASAP7_75t_L g1057 ( 
.A(n_951),
.B(n_839),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_949),
.B(n_887),
.Y(n_1058)
);

BUFx4f_ASAP7_75t_L g1059 ( 
.A(n_976),
.Y(n_1059)
);

NAND3xp33_ASAP7_75t_SL g1060 ( 
.A(n_924),
.B(n_909),
.C(n_934),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_999),
.A2(n_980),
.B1(n_970),
.B2(n_902),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_833),
.B(n_988),
.Y(n_1062)
);

AOI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_822),
.A2(n_855),
.B(n_857),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_1001),
.B(n_964),
.Y(n_1064)
);

BUFx4f_ASAP7_75t_L g1065 ( 
.A(n_839),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_967),
.B(n_975),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_905),
.B(n_952),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_946),
.A2(n_879),
.B(n_901),
.C(n_816),
.Y(n_1068)
);

A2O1A1Ixp33_ASAP7_75t_SL g1069 ( 
.A1(n_913),
.A2(n_920),
.B(n_921),
.C(n_928),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_916),
.Y(n_1070)
);

AOI22xp33_ASAP7_75t_L g1071 ( 
.A1(n_914),
.A2(n_985),
.B1(n_966),
.B2(n_983),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_923),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_950),
.A2(n_927),
.B(n_953),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_875),
.A2(n_836),
.B(n_813),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_L g1075 ( 
.A(n_951),
.B(n_879),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_847),
.A2(n_817),
.B1(n_843),
.B2(n_973),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_973),
.B(n_956),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_930),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_927),
.A2(n_953),
.B(n_835),
.Y(n_1079)
);

BUFx2_ASAP7_75t_SL g1080 ( 
.A(n_967),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_956),
.B(n_850),
.Y(n_1081)
);

INVx3_ASAP7_75t_L g1082 ( 
.A(n_975),
.Y(n_1082)
);

INVx3_ASAP7_75t_L g1083 ( 
.A(n_975),
.Y(n_1083)
);

NAND2x1p5_ASAP7_75t_L g1084 ( 
.A(n_975),
.B(n_932),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_922),
.B(n_925),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_SL g1086 ( 
.A(n_965),
.B(n_978),
.Y(n_1086)
);

AOI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_835),
.A2(n_863),
.B(n_820),
.Y(n_1087)
);

OAI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_982),
.A2(n_997),
.B1(n_995),
.B2(n_1000),
.Y(n_1088)
);

NAND2x1p5_ASAP7_75t_L g1089 ( 
.A(n_932),
.B(n_834),
.Y(n_1089)
);

AOI22xp5_ASAP7_75t_L g1090 ( 
.A1(n_852),
.A2(n_853),
.B1(n_860),
.B2(n_865),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_942),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_958),
.Y(n_1092)
);

AND2x2_ASAP7_75t_L g1093 ( 
.A(n_992),
.B(n_859),
.Y(n_1093)
);

OAI21x1_ASAP7_75t_L g1094 ( 
.A1(n_862),
.A2(n_825),
.B(n_824),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_896),
.A2(n_897),
.B1(n_861),
.B2(n_888),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_889),
.B(n_882),
.Y(n_1096)
);

NAND2x1p5_ASAP7_75t_L g1097 ( 
.A(n_834),
.B(n_903),
.Y(n_1097)
);

NAND3xp33_ASAP7_75t_SL g1098 ( 
.A(n_841),
.B(n_906),
.C(n_986),
.Y(n_1098)
);

BUFx3_ASAP7_75t_L g1099 ( 
.A(n_990),
.Y(n_1099)
);

A2O1A1Ixp33_ASAP7_75t_L g1100 ( 
.A1(n_844),
.A2(n_828),
.B(n_832),
.C(n_910),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_863),
.A2(n_881),
.B(n_818),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_992),
.B(n_990),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_854),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_SL g1104 ( 
.A(n_981),
.B(n_996),
.C(n_908),
.Y(n_1104)
);

INVx2_ASAP7_75t_L g1105 ( 
.A(n_990),
.Y(n_1105)
);

AOI21xp5_ASAP7_75t_L g1106 ( 
.A1(n_891),
.A2(n_915),
.B(n_960),
.Y(n_1106)
);

BUFx2_ASAP7_75t_L g1107 ( 
.A(n_834),
.Y(n_1107)
);

INVx3_ASAP7_75t_SL g1108 ( 
.A(n_834),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_903),
.B(n_948),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_990),
.B(n_903),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_SL g1111 ( 
.A(n_903),
.B(n_948),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_907),
.A2(n_943),
.B(n_893),
.C(n_904),
.Y(n_1112)
);

AOI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_861),
.A2(n_926),
.B1(n_919),
.B2(n_819),
.Y(n_1113)
);

O2A1O1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_904),
.A2(n_917),
.B(n_935),
.C(n_821),
.Y(n_1114)
);

A2O1A1Ixp33_ASAP7_75t_SL g1115 ( 
.A1(n_911),
.A2(n_837),
.B(n_840),
.C(n_931),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_819),
.A2(n_821),
.B(n_842),
.Y(n_1116)
);

O2A1O1Ixp33_ASAP7_75t_L g1117 ( 
.A1(n_935),
.A2(n_937),
.B(n_918),
.C(n_969),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_929),
.Y(n_1118)
);

OAI22xp5_ASAP7_75t_L g1119 ( 
.A1(n_929),
.A2(n_948),
.B1(n_892),
.B2(n_868),
.Y(n_1119)
);

INVx2_ASAP7_75t_L g1120 ( 
.A(n_929),
.Y(n_1120)
);

NOR3xp33_ASAP7_75t_L g1121 ( 
.A(n_918),
.B(n_864),
.C(n_938),
.Y(n_1121)
);

AO32x2_ASAP7_75t_L g1122 ( 
.A1(n_870),
.A2(n_971),
.A3(n_961),
.B1(n_957),
.B2(n_954),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_929),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_948),
.B(n_892),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_899),
.B(n_947),
.Y(n_1125)
);

HB1xp67_ASAP7_75t_L g1126 ( 
.A(n_869),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_872),
.A2(n_890),
.B(n_974),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_972),
.A2(n_829),
.B(n_656),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_866),
.Y(n_1129)
);

AOI22xp33_ASAP7_75t_L g1130 ( 
.A1(n_993),
.A2(n_798),
.B1(n_556),
.B2(n_800),
.Y(n_1130)
);

AOI21xp5_ASAP7_75t_L g1131 ( 
.A1(n_829),
.A2(n_656),
.B(n_826),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_823),
.B(n_814),
.Y(n_1132)
);

NAND2x1p5_ASAP7_75t_L g1133 ( 
.A(n_976),
.B(n_839),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_823),
.B(n_814),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_829),
.A2(n_656),
.B(n_826),
.Y(n_1135)
);

AOI21xp5_ASAP7_75t_L g1136 ( 
.A1(n_829),
.A2(n_656),
.B(n_826),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_831),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_829),
.A2(n_656),
.B(n_826),
.Y(n_1138)
);

BUFx10_ASAP7_75t_L g1139 ( 
.A(n_851),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_829),
.A2(n_656),
.B(n_826),
.Y(n_1140)
);

AND2x2_ASAP7_75t_L g1141 ( 
.A(n_846),
.B(n_544),
.Y(n_1141)
);

BUFx12f_ASAP7_75t_L g1142 ( 
.A(n_867),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_831),
.Y(n_1143)
);

NAND2xp5_ASAP7_75t_SL g1144 ( 
.A(n_856),
.B(n_680),
.Y(n_1144)
);

NOR3xp33_ASAP7_75t_SL g1145 ( 
.A(n_851),
.B(n_689),
.C(n_533),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_814),
.A2(n_940),
.B(n_900),
.C(n_830),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_SL g1147 ( 
.A(n_856),
.B(n_680),
.Y(n_1147)
);

INVx1_ASAP7_75t_L g1148 ( 
.A(n_831),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_829),
.A2(n_656),
.B(n_826),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_831),
.Y(n_1150)
);

INVx8_ASAP7_75t_L g1151 ( 
.A(n_839),
.Y(n_1151)
);

BUFx6f_ASAP7_75t_L g1152 ( 
.A(n_941),
.Y(n_1152)
);

AOI21x1_ASAP7_75t_L g1153 ( 
.A1(n_855),
.A2(n_857),
.B(n_945),
.Y(n_1153)
);

AOI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1011),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1131),
.A2(n_1136),
.B(n_1135),
.Y(n_1156)
);

AND2x2_ASAP7_75t_L g1157 ( 
.A(n_1141),
.B(n_1051),
.Y(n_1157)
);

AO21x2_ASAP7_75t_L g1158 ( 
.A1(n_1063),
.A2(n_1050),
.B(n_1153),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1045),
.Y(n_1159)
);

NOR4xp25_ASAP7_75t_L g1160 ( 
.A(n_1053),
.B(n_1016),
.C(n_1055),
.D(n_1040),
.Y(n_1160)
);

OAI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1132),
.A2(n_1134),
.B1(n_1041),
.B2(n_1015),
.Y(n_1161)
);

NAND3xp33_ASAP7_75t_L g1162 ( 
.A(n_1055),
.B(n_1042),
.C(n_1052),
.Y(n_1162)
);

AO31x2_ASAP7_75t_L g1163 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1163)
);

OAI21x1_ASAP7_75t_L g1164 ( 
.A1(n_1106),
.A2(n_1087),
.B(n_1101),
.Y(n_1164)
);

AO31x2_ASAP7_75t_L g1165 ( 
.A1(n_1033),
.A2(n_1101),
.A3(n_1100),
.B(n_1127),
.Y(n_1165)
);

OAI21x1_ASAP7_75t_L g1166 ( 
.A1(n_1127),
.A2(n_1094),
.B(n_1116),
.Y(n_1166)
);

OAI21x1_ASAP7_75t_L g1167 ( 
.A1(n_1116),
.A2(n_1079),
.B(n_1073),
.Y(n_1167)
);

HB1xp67_ASAP7_75t_L g1168 ( 
.A(n_1004),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_1030),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_SL g1170 ( 
.A1(n_1009),
.A2(n_1096),
.B(n_1068),
.Y(n_1170)
);

AOI221x1_ASAP7_75t_L g1171 ( 
.A1(n_1060),
.A2(n_1043),
.B1(n_1037),
.B2(n_1098),
.C(n_1005),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1136),
.A2(n_1140),
.B(n_1149),
.Y(n_1172)
);

A2O1A1Ixp33_ASAP7_75t_L g1173 ( 
.A1(n_1003),
.A2(n_1052),
.B(n_1002),
.C(n_1085),
.Y(n_1173)
);

AOI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1138),
.A2(n_1140),
.B(n_1149),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1031),
.Y(n_1175)
);

AO31x2_ASAP7_75t_L g1176 ( 
.A1(n_1073),
.A2(n_1128),
.A3(n_1138),
.B(n_1103),
.Y(n_1176)
);

AOI221x1_ASAP7_75t_L g1177 ( 
.A1(n_1060),
.A2(n_1043),
.B1(n_1098),
.B2(n_1008),
.C(n_1121),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1038),
.A2(n_1006),
.B(n_1130),
.C(n_1044),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1065),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1059),
.Y(n_1180)
);

INVx3_ASAP7_75t_L g1181 ( 
.A(n_1059),
.Y(n_1181)
);

BUFx8_ASAP7_75t_L g1182 ( 
.A(n_1035),
.Y(n_1182)
);

OAI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1128),
.A2(n_1008),
.B(n_1114),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_1137),
.Y(n_1184)
);

NAND2x1p5_ASAP7_75t_L g1185 ( 
.A(n_1065),
.B(n_1057),
.Y(n_1185)
);

OAI21x1_ASAP7_75t_L g1186 ( 
.A1(n_1079),
.A2(n_1125),
.B(n_1117),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1056),
.B(n_1013),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_1143),
.Y(n_1188)
);

INVxp67_ASAP7_75t_SL g1189 ( 
.A(n_1018),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1148),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1081),
.B(n_1028),
.Y(n_1191)
);

INVx1_ASAP7_75t_SL g1192 ( 
.A(n_1108),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1104),
.A2(n_1088),
.B(n_1076),
.Y(n_1193)
);

AOI221x1_ASAP7_75t_L g1194 ( 
.A1(n_1075),
.A2(n_1020),
.B1(n_1104),
.B2(n_1119),
.C(n_1058),
.Y(n_1194)
);

AND2x2_ASAP7_75t_L g1195 ( 
.A(n_1062),
.B(n_1057),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_1150),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1047),
.Y(n_1197)
);

OAI21x1_ASAP7_75t_L g1198 ( 
.A1(n_1117),
.A2(n_1020),
.B(n_1114),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1067),
.Y(n_1199)
);

INVx3_ASAP7_75t_L g1200 ( 
.A(n_1133),
.Y(n_1200)
);

OAI21xp5_ASAP7_75t_L g1201 ( 
.A1(n_1113),
.A2(n_1086),
.B(n_1026),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1115),
.A2(n_1069),
.B(n_1021),
.Y(n_1202)
);

NOR2x1_ASAP7_75t_SL g1203 ( 
.A(n_1080),
.B(n_1036),
.Y(n_1203)
);

OR2x2_ASAP7_75t_L g1204 ( 
.A(n_1014),
.B(n_1024),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1038),
.A2(n_1126),
.B(n_1061),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1078),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1092),
.Y(n_1207)
);

CKINVDCx20_ASAP7_75t_R g1208 ( 
.A(n_1023),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1109),
.A2(n_1111),
.B(n_1124),
.Y(n_1209)
);

INVx2_ASAP7_75t_L g1210 ( 
.A(n_1048),
.Y(n_1210)
);

OAI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_1093),
.A2(n_1090),
.B(n_1077),
.Y(n_1211)
);

AOI22xp5_ASAP7_75t_L g1212 ( 
.A1(n_1144),
.A2(n_1147),
.B1(n_1064),
.B2(n_1029),
.Y(n_1212)
);

AOI21xp5_ASAP7_75t_L g1213 ( 
.A1(n_1102),
.A2(n_1110),
.B(n_1097),
.Y(n_1213)
);

INVx6_ASAP7_75t_L g1214 ( 
.A(n_1139),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1054),
.B(n_1034),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1071),
.B(n_1070),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_1072),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1046),
.A2(n_1097),
.B(n_1066),
.Y(n_1218)
);

AO22x2_ASAP7_75t_L g1219 ( 
.A1(n_1091),
.A2(n_1129),
.B1(n_1012),
.B2(n_1105),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1010),
.B(n_1152),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_1120),
.A2(n_1123),
.B(n_1118),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1084),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1118),
.A2(n_1107),
.B(n_1089),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1025),
.B(n_1133),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1007),
.B(n_1039),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_SL g1226 ( 
.A(n_1036),
.B(n_1025),
.Y(n_1226)
);

INVx2_ASAP7_75t_L g1227 ( 
.A(n_1032),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_L g1228 ( 
.A1(n_1118),
.A2(n_1089),
.B(n_1082),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1139),
.Y(n_1229)
);

INVx5_ASAP7_75t_L g1230 ( 
.A(n_1151),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1083),
.A2(n_1099),
.B(n_1027),
.C(n_1019),
.Y(n_1231)
);

INVx2_ASAP7_75t_SL g1232 ( 
.A(n_1010),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1151),
.Y(n_1233)
);

AOI21xp5_ASAP7_75t_L g1234 ( 
.A1(n_1151),
.A2(n_1122),
.B(n_1019),
.Y(n_1234)
);

A2O1A1Ixp33_ASAP7_75t_L g1235 ( 
.A1(n_1010),
.A2(n_1152),
.B(n_1019),
.C(n_1049),
.Y(n_1235)
);

OAI21xp5_ASAP7_75t_L g1236 ( 
.A1(n_1049),
.A2(n_1122),
.B(n_1152),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1049),
.B(n_1142),
.Y(n_1237)
);

NOR2xp67_ASAP7_75t_L g1238 ( 
.A(n_1049),
.B(n_1122),
.Y(n_1238)
);

OAI21x1_ASAP7_75t_L g1239 ( 
.A1(n_1074),
.A2(n_1106),
.B(n_1087),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1141),
.B(n_544),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_L g1241 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1022),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1243)
);

HB1xp67_ASAP7_75t_L g1244 ( 
.A(n_1004),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1146),
.A2(n_1134),
.B(n_1132),
.Y(n_1245)
);

NAND3xp33_ASAP7_75t_L g1246 ( 
.A(n_1146),
.B(n_1016),
.C(n_940),
.Y(n_1246)
);

INVx2_ASAP7_75t_SL g1247 ( 
.A(n_1139),
.Y(n_1247)
);

AND2x2_ASAP7_75t_L g1248 ( 
.A(n_1141),
.B(n_544),
.Y(n_1248)
);

AOI21x1_ASAP7_75t_L g1249 ( 
.A1(n_1050),
.A2(n_1153),
.B(n_1063),
.Y(n_1249)
);

NAND2xp5_ASAP7_75t_L g1250 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1250)
);

BUFx10_ASAP7_75t_L g1251 ( 
.A(n_1017),
.Y(n_1251)
);

OA21x2_ASAP7_75t_L g1252 ( 
.A1(n_1106),
.A2(n_1063),
.B(n_1074),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1254)
);

BUFx4f_ASAP7_75t_L g1255 ( 
.A(n_1151),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1256)
);

INVx5_ASAP7_75t_L g1257 ( 
.A(n_1151),
.Y(n_1257)
);

INVxp67_ASAP7_75t_SL g1258 ( 
.A(n_1009),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1259)
);

OAI22x1_ASAP7_75t_L g1260 ( 
.A1(n_1051),
.A2(n_1002),
.B1(n_532),
.B2(n_533),
.Y(n_1260)
);

AO31x2_ASAP7_75t_L g1261 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1261)
);

AOI221xp5_ASAP7_75t_L g1262 ( 
.A1(n_1146),
.A2(n_823),
.B1(n_791),
.B2(n_727),
.C(n_814),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_1151),
.Y(n_1263)
);

AOI21xp5_ASAP7_75t_L g1264 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1264)
);

AOI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1050),
.A2(n_1153),
.B(n_1063),
.Y(n_1265)
);

AOI31xp67_ASAP7_75t_L g1266 ( 
.A1(n_1086),
.A2(n_1125),
.A3(n_1026),
.B(n_1113),
.Y(n_1266)
);

NOR2xp33_ASAP7_75t_SL g1267 ( 
.A(n_1042),
.B(n_993),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1145),
.Y(n_1268)
);

INVx2_ASAP7_75t_L g1269 ( 
.A(n_1022),
.Y(n_1269)
);

INVxp67_ASAP7_75t_L g1270 ( 
.A(n_1004),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1271)
);

A2O1A1Ixp33_ASAP7_75t_L g1272 ( 
.A1(n_1146),
.A2(n_814),
.B(n_1016),
.C(n_940),
.Y(n_1272)
);

AOI21xp5_ASAP7_75t_L g1273 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1074),
.A2(n_1106),
.B(n_1087),
.Y(n_1274)
);

O2A1O1Ixp33_ASAP7_75t_L g1275 ( 
.A1(n_1146),
.A2(n_823),
.B(n_1016),
.C(n_1053),
.Y(n_1275)
);

AO21x1_ASAP7_75t_L g1276 ( 
.A1(n_1088),
.A2(n_1016),
.B(n_1050),
.Y(n_1276)
);

OAI21xp5_ASAP7_75t_L g1277 ( 
.A1(n_1146),
.A2(n_1134),
.B(n_1132),
.Y(n_1277)
);

A2O1A1Ixp33_ASAP7_75t_L g1278 ( 
.A1(n_1146),
.A2(n_814),
.B(n_1016),
.C(n_940),
.Y(n_1278)
);

AOI21xp5_ASAP7_75t_L g1279 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1280)
);

INVxp67_ASAP7_75t_L g1281 ( 
.A(n_1004),
.Y(n_1281)
);

OAI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1146),
.A2(n_1134),
.B(n_1132),
.Y(n_1282)
);

INVxp67_ASAP7_75t_L g1283 ( 
.A(n_1004),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1146),
.A2(n_1135),
.B(n_1131),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1011),
.Y(n_1285)
);

OR2x2_ASAP7_75t_L g1286 ( 
.A(n_1002),
.B(n_544),
.Y(n_1286)
);

AO31x2_ASAP7_75t_L g1287 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1287)
);

AO31x2_ASAP7_75t_L g1288 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1288)
);

CKINVDCx12_ASAP7_75t_R g1289 ( 
.A(n_1062),
.Y(n_1289)
);

INVxp67_ASAP7_75t_SL g1290 ( 
.A(n_1009),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1132),
.B(n_1134),
.Y(n_1291)
);

BUFx8_ASAP7_75t_L g1292 ( 
.A(n_1004),
.Y(n_1292)
);

A2O1A1Ixp33_ASAP7_75t_L g1293 ( 
.A1(n_1146),
.A2(n_814),
.B(n_1016),
.C(n_940),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1023),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1022),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1141),
.B(n_544),
.Y(n_1296)
);

AO31x2_ASAP7_75t_L g1297 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1297)
);

AOI221xp5_ASAP7_75t_SL g1298 ( 
.A1(n_1146),
.A2(n_1041),
.B1(n_1016),
.B2(n_940),
.C(n_900),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1074),
.A2(n_1106),
.B(n_1087),
.Y(n_1299)
);

OAI21xp5_ASAP7_75t_L g1300 ( 
.A1(n_1146),
.A2(n_1134),
.B(n_1132),
.Y(n_1300)
);

O2A1O1Ixp33_ASAP7_75t_L g1301 ( 
.A1(n_1146),
.A2(n_823),
.B(n_1016),
.C(n_1053),
.Y(n_1301)
);

AO31x2_ASAP7_75t_L g1302 ( 
.A1(n_1063),
.A2(n_1050),
.A3(n_1112),
.B(n_1095),
.Y(n_1302)
);

AO21x1_ASAP7_75t_L g1303 ( 
.A1(n_1088),
.A2(n_1016),
.B(n_1050),
.Y(n_1303)
);

BUFx10_ASAP7_75t_L g1304 ( 
.A(n_1225),
.Y(n_1304)
);

BUFx12f_ASAP7_75t_L g1305 ( 
.A(n_1182),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_SL g1306 ( 
.A1(n_1272),
.A2(n_1293),
.B(n_1278),
.Y(n_1306)
);

BUFx2_ASAP7_75t_L g1307 ( 
.A(n_1292),
.Y(n_1307)
);

CKINVDCx6p67_ASAP7_75t_R g1308 ( 
.A(n_1208),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1220),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1246),
.A2(n_1162),
.B1(n_1262),
.B2(n_1161),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1159),
.Y(n_1311)
);

BUFx4f_ASAP7_75t_SL g1312 ( 
.A(n_1294),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1255),
.Y(n_1313)
);

INVx2_ASAP7_75t_SL g1314 ( 
.A(n_1214),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1267),
.A2(n_1260),
.B1(n_1246),
.B2(n_1161),
.Y(n_1315)
);

HB1xp67_ASAP7_75t_L g1316 ( 
.A(n_1167),
.Y(n_1316)
);

AOI22xp5_ASAP7_75t_L g1317 ( 
.A1(n_1267),
.A2(n_1189),
.B1(n_1157),
.B2(n_1173),
.Y(n_1317)
);

INVx3_ASAP7_75t_L g1318 ( 
.A(n_1255),
.Y(n_1318)
);

INVx6_ASAP7_75t_L g1319 ( 
.A(n_1230),
.Y(n_1319)
);

AOI22xp33_ASAP7_75t_L g1320 ( 
.A1(n_1245),
.A2(n_1282),
.B1(n_1300),
.B2(n_1277),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1184),
.Y(n_1321)
);

BUFx2_ASAP7_75t_L g1322 ( 
.A(n_1292),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1188),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_1229),
.Y(n_1324)
);

AOI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1245),
.A2(n_1282),
.B1(n_1300),
.B2(n_1277),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1162),
.A2(n_1250),
.B1(n_1254),
.B2(n_1241),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1190),
.Y(n_1327)
);

AOI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1204),
.A2(n_1187),
.B1(n_1243),
.B2(n_1250),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1196),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1243),
.A2(n_1254),
.B1(n_1280),
.B2(n_1291),
.Y(n_1330)
);

BUFx2_ASAP7_75t_L g1331 ( 
.A(n_1168),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1176),
.Y(n_1332)
);

AOI22xp5_ASAP7_75t_L g1333 ( 
.A1(n_1298),
.A2(n_1212),
.B1(n_1258),
.B2(n_1290),
.Y(n_1333)
);

OAI21xp5_ASAP7_75t_SL g1334 ( 
.A1(n_1275),
.A2(n_1301),
.B(n_1193),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1285),
.Y(n_1335)
);

INVx6_ASAP7_75t_L g1336 ( 
.A(n_1257),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1286),
.A2(n_1205),
.B1(n_1201),
.B2(n_1199),
.Y(n_1337)
);

INVx3_ASAP7_75t_SL g1338 ( 
.A(n_1268),
.Y(n_1338)
);

BUFx3_ASAP7_75t_L g1339 ( 
.A(n_1220),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1244),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1206),
.Y(n_1341)
);

OAI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1171),
.A2(n_1191),
.B1(n_1215),
.B2(n_1177),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1191),
.A2(n_1303),
.B1(n_1276),
.B2(n_1240),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1270),
.Y(n_1344)
);

BUFx2_ASAP7_75t_L g1345 ( 
.A(n_1281),
.Y(n_1345)
);

OAI22xp5_ASAP7_75t_L g1346 ( 
.A1(n_1178),
.A2(n_1283),
.B1(n_1248),
.B2(n_1296),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1257),
.B(n_1263),
.Y(n_1347)
);

AOI22xp33_ASAP7_75t_L g1348 ( 
.A1(n_1216),
.A2(n_1207),
.B1(n_1211),
.B2(n_1217),
.Y(n_1348)
);

BUFx12f_ASAP7_75t_L g1349 ( 
.A(n_1182),
.Y(n_1349)
);

INVx6_ASAP7_75t_L g1350 ( 
.A(n_1263),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1169),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1214),
.Y(n_1352)
);

OAI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1170),
.A2(n_1154),
.B1(n_1253),
.B2(n_1256),
.Y(n_1353)
);

NAND2x1p5_ASAP7_75t_L g1354 ( 
.A(n_1263),
.B(n_1179),
.Y(n_1354)
);

CKINVDCx14_ASAP7_75t_R g1355 ( 
.A(n_1195),
.Y(n_1355)
);

CKINVDCx14_ASAP7_75t_R g1356 ( 
.A(n_1251),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1192),
.B(n_1232),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1216),
.A2(n_1211),
.B1(n_1238),
.B2(n_1197),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1175),
.A2(n_1210),
.B1(n_1269),
.B2(n_1242),
.Y(n_1359)
);

AOI22xp33_ASAP7_75t_L g1360 ( 
.A1(n_1295),
.A2(n_1273),
.B1(n_1259),
.B2(n_1264),
.Y(n_1360)
);

INVx1_ASAP7_75t_SL g1361 ( 
.A(n_1192),
.Y(n_1361)
);

INVx6_ASAP7_75t_L g1362 ( 
.A(n_1179),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_1247),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1219),
.Y(n_1364)
);

CKINVDCx11_ASAP7_75t_R g1365 ( 
.A(n_1179),
.Y(n_1365)
);

BUFx8_ASAP7_75t_SL g1366 ( 
.A(n_1237),
.Y(n_1366)
);

BUFx10_ASAP7_75t_L g1367 ( 
.A(n_1233),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_SL g1368 ( 
.A1(n_1236),
.A2(n_1183),
.B1(n_1234),
.B2(n_1298),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1289),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1227),
.Y(n_1370)
);

AOI22xp33_ASAP7_75t_L g1371 ( 
.A1(n_1279),
.A2(n_1284),
.B1(n_1183),
.B2(n_1236),
.Y(n_1371)
);

CKINVDCx11_ASAP7_75t_R g1372 ( 
.A(n_1222),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1231),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1224),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1224),
.Y(n_1375)
);

NAND2xp5_ASAP7_75t_L g1376 ( 
.A(n_1160),
.B(n_1185),
.Y(n_1376)
);

AOI22xp33_ASAP7_75t_L g1377 ( 
.A1(n_1156),
.A2(n_1172),
.B1(n_1174),
.B2(n_1185),
.Y(n_1377)
);

CKINVDCx8_ASAP7_75t_R g1378 ( 
.A(n_1252),
.Y(n_1378)
);

BUFx3_ASAP7_75t_L g1379 ( 
.A(n_1180),
.Y(n_1379)
);

AND2x2_ASAP7_75t_L g1380 ( 
.A(n_1180),
.B(n_1181),
.Y(n_1380)
);

BUFx8_ASAP7_75t_L g1381 ( 
.A(n_1160),
.Y(n_1381)
);

AOI22xp5_ASAP7_75t_SL g1382 ( 
.A1(n_1181),
.A2(n_1200),
.B1(n_1223),
.B2(n_1213),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1266),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1198),
.Y(n_1384)
);

BUFx6f_ASAP7_75t_L g1385 ( 
.A(n_1200),
.Y(n_1385)
);

OAI22xp33_ASAP7_75t_L g1386 ( 
.A1(n_1194),
.A2(n_1228),
.B1(n_1209),
.B2(n_1226),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1218),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_SL g1388 ( 
.A1(n_1235),
.A2(n_1252),
.B1(n_1297),
.B2(n_1163),
.Y(n_1388)
);

INVx6_ASAP7_75t_L g1389 ( 
.A(n_1203),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1158),
.A2(n_1186),
.B1(n_1221),
.B2(n_1202),
.Y(n_1390)
);

OAI22xp5_ASAP7_75t_L g1391 ( 
.A1(n_1249),
.A2(n_1265),
.B1(n_1302),
.B2(n_1163),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1163),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1165),
.Y(n_1393)
);

CKINVDCx11_ASAP7_75t_R g1394 ( 
.A(n_1261),
.Y(n_1394)
);

BUFx12f_ASAP7_75t_L g1395 ( 
.A(n_1261),
.Y(n_1395)
);

AOI22xp33_ASAP7_75t_SL g1396 ( 
.A1(n_1158),
.A2(n_1271),
.B1(n_1297),
.B2(n_1288),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1261),
.A2(n_1271),
.B1(n_1297),
.B2(n_1288),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1164),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1165),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1165),
.Y(n_1400)
);

BUFx8_ASAP7_75t_L g1401 ( 
.A(n_1287),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1287),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_SL g1403 ( 
.A1(n_1287),
.A2(n_1302),
.B1(n_1288),
.B2(n_1166),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1302),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1239),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1274),
.Y(n_1406)
);

INVx6_ASAP7_75t_L g1407 ( 
.A(n_1299),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_SL g1408 ( 
.A1(n_1267),
.A2(n_993),
.B1(n_340),
.B2(n_342),
.Y(n_1408)
);

OAI22xp33_ASAP7_75t_L g1409 ( 
.A1(n_1267),
.A2(n_1016),
.B1(n_1246),
.B2(n_1002),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1155),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1220),
.Y(n_1411)
);

AOI22xp33_ASAP7_75t_L g1412 ( 
.A1(n_1267),
.A2(n_1130),
.B1(n_1002),
.B2(n_993),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1155),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1182),
.Y(n_1414)
);

INVx1_ASAP7_75t_SL g1415 ( 
.A(n_1208),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1208),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1220),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1155),
.Y(n_1418)
);

INVx6_ASAP7_75t_L g1419 ( 
.A(n_1230),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1229),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_L g1421 ( 
.A1(n_1267),
.A2(n_1130),
.B1(n_1002),
.B2(n_993),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1155),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1267),
.A2(n_993),
.B1(n_340),
.B2(n_342),
.Y(n_1423)
);

INVx3_ASAP7_75t_L g1424 ( 
.A(n_1255),
.Y(n_1424)
);

OAI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1246),
.A2(n_1016),
.B1(n_1146),
.B2(n_1272),
.Y(n_1425)
);

CKINVDCx11_ASAP7_75t_R g1426 ( 
.A(n_1208),
.Y(n_1426)
);

AOI22xp33_ASAP7_75t_SL g1427 ( 
.A1(n_1267),
.A2(n_993),
.B1(n_340),
.B2(n_342),
.Y(n_1427)
);

CKINVDCx6p67_ASAP7_75t_R g1428 ( 
.A(n_1208),
.Y(n_1428)
);

BUFx2_ASAP7_75t_SL g1429 ( 
.A(n_1208),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1157),
.B(n_1195),
.Y(n_1430)
);

BUFx6f_ASAP7_75t_L g1431 ( 
.A(n_1179),
.Y(n_1431)
);

CKINVDCx6p67_ASAP7_75t_R g1432 ( 
.A(n_1208),
.Y(n_1432)
);

AO21x2_ASAP7_75t_L g1433 ( 
.A1(n_1383),
.A2(n_1391),
.B(n_1332),
.Y(n_1433)
);

AOI22xp5_ASAP7_75t_L g1434 ( 
.A1(n_1408),
.A2(n_1423),
.B1(n_1427),
.B2(n_1421),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1374),
.Y(n_1435)
);

O2A1O1Ixp33_ASAP7_75t_L g1436 ( 
.A1(n_1310),
.A2(n_1409),
.B(n_1334),
.C(n_1425),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1375),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1393),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1399),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1353),
.A2(n_1390),
.B(n_1377),
.Y(n_1440)
);

OR2x2_ASAP7_75t_L g1441 ( 
.A(n_1392),
.B(n_1400),
.Y(n_1441)
);

AOI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1412),
.A2(n_1421),
.B1(n_1409),
.B2(n_1381),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1311),
.Y(n_1443)
);

BUFx2_ASAP7_75t_L g1444 ( 
.A(n_1401),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1390),
.A2(n_1377),
.B(n_1360),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1368),
.B(n_1394),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1321),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1323),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1327),
.Y(n_1449)
);

HB1xp67_ASAP7_75t_L g1450 ( 
.A(n_1331),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1329),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1335),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1410),
.Y(n_1453)
);

O2A1O1Ixp33_ASAP7_75t_L g1454 ( 
.A1(n_1315),
.A2(n_1346),
.B(n_1342),
.C(n_1325),
.Y(n_1454)
);

HB1xp67_ASAP7_75t_L g1455 ( 
.A(n_1340),
.Y(n_1455)
);

BUFx6f_ASAP7_75t_L g1456 ( 
.A(n_1395),
.Y(n_1456)
);

BUFx3_ASAP7_75t_L g1457 ( 
.A(n_1339),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1360),
.A2(n_1383),
.B(n_1384),
.Y(n_1458)
);

NOR2xp33_ASAP7_75t_L g1459 ( 
.A(n_1312),
.B(n_1416),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1413),
.Y(n_1460)
);

HB1xp67_ASAP7_75t_L g1461 ( 
.A(n_1418),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1422),
.Y(n_1462)
);

AND2x6_ASAP7_75t_L g1463 ( 
.A(n_1317),
.B(n_1364),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1341),
.Y(n_1464)
);

NAND2xp5_ASAP7_75t_L g1465 ( 
.A(n_1328),
.B(n_1330),
.Y(n_1465)
);

NOR2xp33_ASAP7_75t_L g1466 ( 
.A(n_1312),
.B(n_1415),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1402),
.Y(n_1467)
);

AOI21xp33_ASAP7_75t_L g1468 ( 
.A1(n_1315),
.A2(n_1342),
.B(n_1412),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1330),
.B(n_1326),
.Y(n_1469)
);

AND2x2_ASAP7_75t_L g1470 ( 
.A(n_1320),
.B(n_1325),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1320),
.B(n_1371),
.Y(n_1471)
);

HB1xp67_ASAP7_75t_L g1472 ( 
.A(n_1344),
.Y(n_1472)
);

INVxp67_ASAP7_75t_L g1473 ( 
.A(n_1430),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1371),
.A2(n_1404),
.B(n_1343),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1316),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1397),
.B(n_1396),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1316),
.Y(n_1477)
);

AOI221xp5_ASAP7_75t_L g1478 ( 
.A1(n_1306),
.A2(n_1337),
.B1(n_1343),
.B2(n_1333),
.C(n_1373),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1351),
.Y(n_1479)
);

AO21x1_ASAP7_75t_SL g1480 ( 
.A1(n_1376),
.A2(n_1358),
.B(n_1348),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1388),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1378),
.Y(n_1482)
);

AOI221xp5_ASAP7_75t_L g1483 ( 
.A1(n_1348),
.A2(n_1386),
.B1(n_1361),
.B2(n_1357),
.C(n_1403),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1387),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1387),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1398),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1406),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1345),
.B(n_1417),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1379),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1386),
.Y(n_1490)
);

INVx1_ASAP7_75t_SL g1491 ( 
.A(n_1429),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1406),
.Y(n_1492)
);

AND2x2_ASAP7_75t_L g1493 ( 
.A(n_1355),
.B(n_1405),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1411),
.B(n_1417),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1380),
.A2(n_1407),
.B(n_1382),
.Y(n_1495)
);

OA22x2_ASAP7_75t_L g1496 ( 
.A1(n_1370),
.A2(n_1322),
.B1(n_1307),
.B2(n_1338),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1347),
.A2(n_1354),
.B(n_1359),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1407),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1407),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1379),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1359),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1385),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1385),
.Y(n_1503)
);

AND2x4_ASAP7_75t_L g1504 ( 
.A(n_1411),
.B(n_1385),
.Y(n_1504)
);

OAI21x1_ASAP7_75t_L g1505 ( 
.A1(n_1347),
.A2(n_1354),
.B(n_1313),
.Y(n_1505)
);

AOI22xp5_ASAP7_75t_L g1506 ( 
.A1(n_1369),
.A2(n_1356),
.B1(n_1372),
.B2(n_1365),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1431),
.B(n_1424),
.Y(n_1507)
);

NOR2xp33_ASAP7_75t_L g1508 ( 
.A(n_1426),
.B(n_1432),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1367),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1367),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_SL g1511 ( 
.A(n_1305),
.B(n_1349),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1309),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1314),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1356),
.B(n_1352),
.Y(n_1514)
);

INVx2_ASAP7_75t_L g1515 ( 
.A(n_1389),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1304),
.B(n_1431),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1304),
.B(n_1431),
.Y(n_1517)
);

INVx3_ASAP7_75t_L g1518 ( 
.A(n_1319),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1493),
.B(n_1308),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1440),
.A2(n_1363),
.B(n_1420),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1493),
.B(n_1428),
.Y(n_1521)
);

A2O1A1Ixp33_ASAP7_75t_L g1522 ( 
.A1(n_1436),
.A2(n_1313),
.B(n_1318),
.C(n_1424),
.Y(n_1522)
);

BUFx10_ASAP7_75t_L g1523 ( 
.A(n_1459),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1461),
.B(n_1338),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1454),
.A2(n_1318),
.B(n_1324),
.C(n_1366),
.Y(n_1525)
);

AO22x2_ASAP7_75t_L g1526 ( 
.A1(n_1441),
.A2(n_1362),
.B1(n_1414),
.B2(n_1389),
.Y(n_1526)
);

AO21x2_ASAP7_75t_L g1527 ( 
.A1(n_1468),
.A2(n_1389),
.B(n_1419),
.Y(n_1527)
);

AND2x6_ASAP7_75t_L g1528 ( 
.A(n_1442),
.B(n_1336),
.Y(n_1528)
);

INVx4_ASAP7_75t_L g1529 ( 
.A(n_1507),
.Y(n_1529)
);

AOI22xp5_ASAP7_75t_L g1530 ( 
.A1(n_1434),
.A2(n_1350),
.B1(n_1419),
.B2(n_1470),
.Y(n_1530)
);

A2O1A1Ixp33_ASAP7_75t_L g1531 ( 
.A1(n_1434),
.A2(n_1478),
.B(n_1446),
.C(n_1483),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1473),
.B(n_1450),
.Y(n_1532)
);

INVx3_ASAP7_75t_L g1533 ( 
.A(n_1509),
.Y(n_1533)
);

BUFx3_ASAP7_75t_L g1534 ( 
.A(n_1514),
.Y(n_1534)
);

AOI21xp5_ASAP7_75t_L g1535 ( 
.A1(n_1471),
.A2(n_1469),
.B(n_1440),
.Y(n_1535)
);

OAI21xp5_ASAP7_75t_L g1536 ( 
.A1(n_1471),
.A2(n_1490),
.B(n_1465),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1455),
.B(n_1488),
.Y(n_1537)
);

NOR2x1_ASAP7_75t_SL g1538 ( 
.A(n_1480),
.B(n_1495),
.Y(n_1538)
);

O2A1O1Ixp33_ASAP7_75t_L g1539 ( 
.A1(n_1490),
.A2(n_1481),
.B(n_1472),
.C(n_1513),
.Y(n_1539)
);

OA21x2_ASAP7_75t_L g1540 ( 
.A1(n_1445),
.A2(n_1474),
.B(n_1458),
.Y(n_1540)
);

A2O1A1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1446),
.A2(n_1476),
.B(n_1474),
.C(n_1482),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1488),
.B(n_1500),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1491),
.B(n_1466),
.Y(n_1543)
);

A2O1A1Ixp33_ASAP7_75t_L g1544 ( 
.A1(n_1480),
.A2(n_1444),
.B(n_1445),
.C(n_1506),
.Y(n_1544)
);

NOR2x1_ASAP7_75t_SL g1545 ( 
.A(n_1495),
.B(n_1457),
.Y(n_1545)
);

O2A1O1Ixp33_ASAP7_75t_SL g1546 ( 
.A1(n_1508),
.A2(n_1506),
.B(n_1489),
.C(n_1510),
.Y(n_1546)
);

NAND3xp33_ASAP7_75t_L g1547 ( 
.A(n_1510),
.B(n_1475),
.C(n_1477),
.Y(n_1547)
);

AO21x1_ASAP7_75t_L g1548 ( 
.A1(n_1443),
.A2(n_1453),
.B(n_1464),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1496),
.A2(n_1448),
.B1(n_1462),
.B2(n_1460),
.Y(n_1549)
);

INVx3_ASAP7_75t_L g1550 ( 
.A(n_1509),
.Y(n_1550)
);

OAI21xp33_ASAP7_75t_L g1551 ( 
.A1(n_1496),
.A2(n_1475),
.B(n_1477),
.Y(n_1551)
);

NOR2xp33_ASAP7_75t_L g1552 ( 
.A(n_1496),
.B(n_1511),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1463),
.A2(n_1505),
.B(n_1458),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1516),
.B(n_1517),
.Y(n_1554)
);

NAND2xp33_ASAP7_75t_R g1555 ( 
.A(n_1444),
.B(n_1516),
.Y(n_1555)
);

OAI22xp5_ASAP7_75t_L g1556 ( 
.A1(n_1447),
.A2(n_1464),
.B1(n_1451),
.B2(n_1449),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1517),
.B(n_1494),
.Y(n_1557)
);

OAI22xp5_ASAP7_75t_L g1558 ( 
.A1(n_1449),
.A2(n_1460),
.B1(n_1462),
.B2(n_1453),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1494),
.B(n_1457),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1463),
.A2(n_1437),
.B1(n_1435),
.B2(n_1452),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1437),
.A2(n_1507),
.B1(n_1501),
.B2(n_1441),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1438),
.A2(n_1439),
.B1(n_1467),
.B2(n_1492),
.C(n_1485),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1479),
.B(n_1502),
.Y(n_1563)
);

AO32x2_ASAP7_75t_L g1564 ( 
.A1(n_1463),
.A2(n_1479),
.A3(n_1484),
.B1(n_1467),
.B2(n_1438),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1439),
.Y(n_1565)
);

AOI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1463),
.A2(n_1504),
.B1(n_1515),
.B2(n_1512),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1487),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1503),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1565),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1548),
.Y(n_1570)
);

INVx2_ASAP7_75t_L g1571 ( 
.A(n_1540),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1520),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1564),
.B(n_1498),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1558),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1567),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1558),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1547),
.Y(n_1577)
);

INVxp67_ASAP7_75t_L g1578 ( 
.A(n_1547),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1564),
.B(n_1498),
.Y(n_1579)
);

AND2x4_ASAP7_75t_L g1580 ( 
.A(n_1553),
.B(n_1498),
.Y(n_1580)
);

AOI22xp33_ASAP7_75t_SL g1581 ( 
.A1(n_1549),
.A2(n_1463),
.B1(n_1456),
.B2(n_1433),
.Y(n_1581)
);

INVx2_ASAP7_75t_L g1582 ( 
.A(n_1540),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1535),
.B(n_1433),
.Y(n_1583)
);

BUFx2_ASAP7_75t_L g1584 ( 
.A(n_1520),
.Y(n_1584)
);

NOR2xp33_ASAP7_75t_L g1585 ( 
.A(n_1546),
.B(n_1499),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1551),
.B(n_1433),
.Y(n_1586)
);

NOR2x1p5_ASAP7_75t_L g1587 ( 
.A(n_1524),
.B(n_1518),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1556),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1563),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1568),
.Y(n_1590)
);

INVx2_ASAP7_75t_L g1591 ( 
.A(n_1545),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1549),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1538),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1537),
.B(n_1557),
.Y(n_1594)
);

HB1xp67_ASAP7_75t_L g1595 ( 
.A(n_1533),
.Y(n_1595)
);

OAI21xp33_ASAP7_75t_SL g1596 ( 
.A1(n_1560),
.A2(n_1497),
.B(n_1486),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1550),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1561),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1592),
.B(n_1542),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1573),
.B(n_1554),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1569),
.Y(n_1601)
);

OR2x2_ASAP7_75t_L g1602 ( 
.A(n_1592),
.B(n_1532),
.Y(n_1602)
);

HB1xp67_ASAP7_75t_L g1603 ( 
.A(n_1577),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1577),
.B(n_1561),
.Y(n_1604)
);

INVx2_ASAP7_75t_SL g1605 ( 
.A(n_1593),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1571),
.Y(n_1607)
);

INVx2_ASAP7_75t_L g1608 ( 
.A(n_1571),
.Y(n_1608)
);

AND2x4_ASAP7_75t_L g1609 ( 
.A(n_1593),
.B(n_1529),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1593),
.Y(n_1610)
);

AOI222xp33_ASAP7_75t_L g1611 ( 
.A1(n_1578),
.A2(n_1531),
.B1(n_1536),
.B2(n_1552),
.C1(n_1541),
.C2(n_1528),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1579),
.B(n_1559),
.Y(n_1612)
);

AOI221xp5_ASAP7_75t_L g1613 ( 
.A1(n_1578),
.A2(n_1539),
.B1(n_1536),
.B2(n_1544),
.C(n_1525),
.Y(n_1613)
);

HB1xp67_ASAP7_75t_L g1614 ( 
.A(n_1574),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1574),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1571),
.Y(n_1616)
);

BUFx3_ASAP7_75t_L g1617 ( 
.A(n_1575),
.Y(n_1617)
);

OR2x6_ASAP7_75t_L g1618 ( 
.A(n_1580),
.B(n_1526),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1571),
.Y(n_1619)
);

AO21x2_ASAP7_75t_L g1620 ( 
.A1(n_1586),
.A2(n_1527),
.B(n_1530),
.Y(n_1620)
);

AND4x1_ASAP7_75t_L g1621 ( 
.A(n_1585),
.B(n_1522),
.C(n_1530),
.D(n_1543),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1576),
.B(n_1562),
.Y(n_1622)
);

NAND4xp25_ASAP7_75t_L g1623 ( 
.A(n_1576),
.B(n_1519),
.C(n_1521),
.D(n_1534),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1597),
.B(n_1594),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1594),
.B(n_1598),
.Y(n_1625)
);

AND2x4_ASAP7_75t_L g1626 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1614),
.B(n_1588),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1614),
.B(n_1588),
.Y(n_1628)
);

AND2x2_ASAP7_75t_SL g1629 ( 
.A(n_1604),
.B(n_1621),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1572),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1601),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1606),
.B(n_1572),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1606),
.B(n_1572),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1606),
.B(n_1584),
.Y(n_1634)
);

INVx1_ASAP7_75t_L g1635 ( 
.A(n_1601),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1600),
.B(n_1584),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1601),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1600),
.B(n_1612),
.Y(n_1638)
);

OR2x2_ASAP7_75t_L g1639 ( 
.A(n_1615),
.B(n_1590),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1600),
.B(n_1584),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1600),
.B(n_1594),
.Y(n_1642)
);

OAI22xp33_ASAP7_75t_L g1643 ( 
.A1(n_1613),
.A2(n_1570),
.B1(n_1566),
.B2(n_1598),
.Y(n_1643)
);

NAND2xp5_ASAP7_75t_L g1644 ( 
.A(n_1615),
.B(n_1570),
.Y(n_1644)
);

INVx4_ASAP7_75t_L g1645 ( 
.A(n_1603),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1603),
.B(n_1589),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1617),
.B(n_1591),
.Y(n_1647)
);

INVx2_ASAP7_75t_L g1648 ( 
.A(n_1619),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1619),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1622),
.B(n_1625),
.Y(n_1650)
);

INVx5_ASAP7_75t_L g1651 ( 
.A(n_1618),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1619),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1619),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1622),
.B(n_1589),
.Y(n_1654)
);

INVxp67_ASAP7_75t_SL g1655 ( 
.A(n_1604),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1612),
.B(n_1595),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1609),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1612),
.B(n_1624),
.Y(n_1658)
);

OR2x2_ASAP7_75t_L g1659 ( 
.A(n_1604),
.B(n_1590),
.Y(n_1659)
);

INVx2_ASAP7_75t_L g1660 ( 
.A(n_1658),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1629),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1650),
.B(n_1599),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1659),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1655),
.B(n_1625),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1658),
.Y(n_1666)
);

OAI222xp33_ASAP7_75t_L g1667 ( 
.A1(n_1643),
.A2(n_1581),
.B1(n_1651),
.B2(n_1650),
.C1(n_1630),
.C2(n_1633),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1627),
.B(n_1599),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1629),
.B(n_1625),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1638),
.B(n_1605),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1638),
.B(n_1642),
.Y(n_1671)
);

AOI22xp5_ASAP7_75t_L g1672 ( 
.A1(n_1629),
.A2(n_1611),
.B1(n_1613),
.B2(n_1581),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1642),
.B(n_1638),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1642),
.B(n_1624),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1629),
.B(n_1602),
.Y(n_1675)
);

INVx1_ASAP7_75t_L g1676 ( 
.A(n_1639),
.Y(n_1676)
);

INVx2_ASAP7_75t_L g1677 ( 
.A(n_1658),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1639),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1639),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1681)
);

INVx2_ASAP7_75t_L g1682 ( 
.A(n_1636),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1645),
.B(n_1605),
.Y(n_1683)
);

NOR2xp33_ASAP7_75t_L g1684 ( 
.A(n_1627),
.B(n_1623),
.Y(n_1684)
);

INVxp67_ASAP7_75t_L g1685 ( 
.A(n_1654),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1659),
.Y(n_1686)
);

NAND2x1p5_ASAP7_75t_L g1687 ( 
.A(n_1645),
.B(n_1621),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1659),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1654),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1646),
.Y(n_1690)
);

INVx2_ASAP7_75t_L g1691 ( 
.A(n_1636),
.Y(n_1691)
);

NOR2xp33_ASAP7_75t_SL g1692 ( 
.A(n_1651),
.B(n_1623),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1628),
.B(n_1599),
.Y(n_1693)
);

OR2x2_ASAP7_75t_L g1694 ( 
.A(n_1628),
.B(n_1602),
.Y(n_1694)
);

NAND2x1_ASAP7_75t_L g1695 ( 
.A(n_1645),
.B(n_1610),
.Y(n_1695)
);

INVxp33_ASAP7_75t_L g1696 ( 
.A(n_1644),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1630),
.B(n_1624),
.Y(n_1697)
);

AOI22x1_ASAP7_75t_L g1698 ( 
.A1(n_1645),
.A2(n_1611),
.B1(n_1619),
.B2(n_1587),
.Y(n_1698)
);

NAND2xp5_ASAP7_75t_L g1699 ( 
.A(n_1643),
.B(n_1602),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1644),
.B(n_1523),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1646),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1636),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1661),
.B(n_1630),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1685),
.B(n_1632),
.Y(n_1704)
);

INVx1_ASAP7_75t_SL g1705 ( 
.A(n_1675),
.Y(n_1705)
);

HB1xp67_ASAP7_75t_L g1706 ( 
.A(n_1664),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1687),
.B(n_1632),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1689),
.B(n_1632),
.Y(n_1708)
);

AND2x2_ASAP7_75t_SL g1709 ( 
.A(n_1672),
.B(n_1699),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1662),
.B(n_1633),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1664),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1687),
.B(n_1633),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1688),
.Y(n_1714)
);

NOR2x1_ASAP7_75t_L g1715 ( 
.A(n_1669),
.B(n_1657),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1684),
.B(n_1634),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1676),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1690),
.B(n_1634),
.Y(n_1718)
);

NAND2x1p5_ASAP7_75t_L g1719 ( 
.A(n_1698),
.B(n_1621),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1701),
.B(n_1634),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1680),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1687),
.B(n_1657),
.Y(n_1723)
);

NAND3x1_ASAP7_75t_L g1724 ( 
.A(n_1663),
.B(n_1640),
.C(n_1656),
.Y(n_1724)
);

NAND2x1p5_ASAP7_75t_L g1725 ( 
.A(n_1698),
.B(n_1651),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1671),
.B(n_1657),
.Y(n_1726)
);

OR2x2_ASAP7_75t_L g1727 ( 
.A(n_1662),
.B(n_1631),
.Y(n_1727)
);

OR2x2_ASAP7_75t_L g1728 ( 
.A(n_1694),
.B(n_1668),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1694),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1671),
.B(n_1673),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1660),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1692),
.A2(n_1651),
.B1(n_1620),
.B2(n_1583),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1660),
.Y(n_1733)
);

NAND2x1_ASAP7_75t_L g1734 ( 
.A(n_1670),
.B(n_1679),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1671),
.B(n_1640),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1668),
.Y(n_1736)
);

AND2x4_ASAP7_75t_L g1737 ( 
.A(n_1673),
.B(n_1651),
.Y(n_1737)
);

NAND3xp33_ASAP7_75t_L g1738 ( 
.A(n_1696),
.B(n_1619),
.C(n_1585),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1729),
.B(n_1696),
.Y(n_1739)
);

INVx1_ASAP7_75t_SL g1740 ( 
.A(n_1707),
.Y(n_1740)
);

OAI21xp5_ASAP7_75t_L g1741 ( 
.A1(n_1719),
.A2(n_1667),
.B(n_1665),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_SL g1742 ( 
.A(n_1719),
.B(n_1679),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1730),
.B(n_1700),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1706),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1711),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1729),
.B(n_1697),
.Y(n_1746)
);

A2O1A1Ixp33_ASAP7_75t_L g1747 ( 
.A1(n_1709),
.A2(n_1651),
.B(n_1596),
.C(n_1640),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1709),
.A2(n_1620),
.B1(n_1651),
.B2(n_1583),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1711),
.Y(n_1749)
);

NOR3xp33_ASAP7_75t_L g1750 ( 
.A(n_1705),
.B(n_1693),
.C(n_1695),
.Y(n_1750)
);

INVx1_ASAP7_75t_L g1751 ( 
.A(n_1717),
.Y(n_1751)
);

INVx3_ASAP7_75t_L g1752 ( 
.A(n_1725),
.Y(n_1752)
);

AOI32xp33_ASAP7_75t_L g1753 ( 
.A1(n_1707),
.A2(n_1702),
.A3(n_1682),
.B1(n_1691),
.B2(n_1697),
.Y(n_1753)
);

AOI22xp33_ASAP7_75t_L g1754 ( 
.A1(n_1719),
.A2(n_1651),
.B1(n_1620),
.B2(n_1582),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1730),
.B(n_1666),
.Y(n_1755)
);

AOI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1716),
.A2(n_1616),
.B1(n_1608),
.B2(n_1607),
.C(n_1586),
.Y(n_1756)
);

OAI22xp33_ASAP7_75t_L g1757 ( 
.A1(n_1725),
.A2(n_1651),
.B1(n_1618),
.B2(n_1693),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_L g1758 ( 
.A(n_1736),
.B(n_1682),
.Y(n_1758)
);

INVxp67_ASAP7_75t_L g1759 ( 
.A(n_1723),
.Y(n_1759)
);

AOI221x1_ASAP7_75t_SL g1760 ( 
.A1(n_1703),
.A2(n_1702),
.B1(n_1691),
.B2(n_1677),
.C(n_1666),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1717),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1721),
.Y(n_1762)
);

NOR2x1p5_ASAP7_75t_L g1763 ( 
.A(n_1734),
.B(n_1695),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1728),
.B(n_1523),
.Y(n_1764)
);

NAND2xp33_ASAP7_75t_SL g1765 ( 
.A(n_1742),
.B(n_1712),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1748),
.A2(n_1712),
.B1(n_1725),
.B2(n_1732),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1745),
.Y(n_1767)
);

AND2x4_ASAP7_75t_L g1768 ( 
.A(n_1759),
.B(n_1726),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1749),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1751),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1761),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1762),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1742),
.Y(n_1773)
);

OAI32xp33_ASAP7_75t_L g1774 ( 
.A1(n_1741),
.A2(n_1710),
.A3(n_1704),
.B1(n_1728),
.B2(n_1738),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1755),
.Y(n_1775)
);

AND2x2_ASAP7_75t_L g1776 ( 
.A(n_1740),
.B(n_1735),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1752),
.Y(n_1777)
);

INVx1_ASAP7_75t_SL g1778 ( 
.A(n_1739),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_SL g1779 ( 
.A1(n_1747),
.A2(n_1734),
.B(n_1710),
.C(n_1721),
.Y(n_1779)
);

OAI21xp33_ASAP7_75t_L g1780 ( 
.A1(n_1753),
.A2(n_1720),
.B(n_1718),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1760),
.B(n_1722),
.Y(n_1781)
);

INVx1_ASAP7_75t_L g1782 ( 
.A(n_1758),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1744),
.Y(n_1783)
);

A2O1A1Ixp33_ASAP7_75t_L g1784 ( 
.A1(n_1747),
.A2(n_1723),
.B(n_1715),
.C(n_1708),
.Y(n_1784)
);

OR2x2_ASAP7_75t_L g1785 ( 
.A(n_1775),
.B(n_1746),
.Y(n_1785)
);

AOI21xp5_ASAP7_75t_L g1786 ( 
.A1(n_1779),
.A2(n_1764),
.B(n_1750),
.Y(n_1786)
);

OAI21xp33_ASAP7_75t_L g1787 ( 
.A1(n_1780),
.A2(n_1764),
.B(n_1743),
.Y(n_1787)
);

INVx1_ASAP7_75t_SL g1788 ( 
.A(n_1778),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1774),
.A2(n_1754),
.B1(n_1756),
.B2(n_1757),
.C(n_1752),
.Y(n_1789)
);

OAI321xp33_ASAP7_75t_L g1790 ( 
.A1(n_1784),
.A2(n_1754),
.A3(n_1714),
.B1(n_1713),
.B2(n_1731),
.C(n_1733),
.Y(n_1790)
);

NOR2x1_ASAP7_75t_L g1791 ( 
.A(n_1777),
.B(n_1763),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_L g1792 ( 
.A(n_1775),
.B(n_1713),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1776),
.Y(n_1793)
);

AND2x2_ASAP7_75t_L g1794 ( 
.A(n_1768),
.B(n_1773),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1767),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1769),
.Y(n_1796)
);

NAND3xp33_ASAP7_75t_L g1797 ( 
.A(n_1794),
.B(n_1765),
.C(n_1784),
.Y(n_1797)
);

AOI33xp33_ASAP7_75t_L g1798 ( 
.A1(n_1788),
.A2(n_1779),
.A3(n_1768),
.B1(n_1783),
.B2(n_1782),
.B3(n_1770),
.Y(n_1798)
);

OAI21xp5_ASAP7_75t_SL g1799 ( 
.A1(n_1786),
.A2(n_1781),
.B(n_1777),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1788),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1793),
.B(n_1735),
.Y(n_1801)
);

NAND3xp33_ASAP7_75t_L g1802 ( 
.A(n_1789),
.B(n_1765),
.C(n_1771),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1785),
.Y(n_1803)
);

AND3x1_ASAP7_75t_L g1804 ( 
.A(n_1787),
.B(n_1772),
.C(n_1752),
.Y(n_1804)
);

AOI322xp5_ASAP7_75t_L g1805 ( 
.A1(n_1795),
.A2(n_1766),
.A3(n_1714),
.B1(n_1733),
.B2(n_1731),
.C1(n_1724),
.C2(n_1737),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_SL g1806 ( 
.A(n_1796),
.B(n_1726),
.C(n_1727),
.Y(n_1806)
);

OAI21xp33_ASAP7_75t_SL g1807 ( 
.A1(n_1791),
.A2(n_1724),
.B(n_1727),
.Y(n_1807)
);

OAI22xp5_ASAP7_75t_L g1808 ( 
.A1(n_1797),
.A2(n_1737),
.B1(n_1792),
.B2(n_1677),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1802),
.A2(n_1737),
.B1(n_1790),
.B2(n_1616),
.Y(n_1809)
);

NAND2xp67_ASAP7_75t_SL g1810 ( 
.A(n_1801),
.B(n_1674),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1799),
.A2(n_1607),
.B1(n_1608),
.B2(n_1616),
.C(n_1619),
.Y(n_1811)
);

A2O1A1Ixp33_ASAP7_75t_L g1812 ( 
.A1(n_1807),
.A2(n_1683),
.B(n_1681),
.C(n_1679),
.Y(n_1812)
);

OAI211xp5_ASAP7_75t_L g1813 ( 
.A1(n_1809),
.A2(n_1805),
.B(n_1800),
.C(n_1803),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1808),
.Y(n_1814)
);

AOI221x1_ASAP7_75t_L g1815 ( 
.A1(n_1812),
.A2(n_1806),
.B1(n_1798),
.B2(n_1804),
.C(n_1683),
.Y(n_1815)
);

OAI22xp5_ASAP7_75t_SL g1816 ( 
.A1(n_1810),
.A2(n_1806),
.B1(n_1670),
.B2(n_1683),
.Y(n_1816)
);

AOI211x1_ASAP7_75t_L g1817 ( 
.A1(n_1811),
.A2(n_1674),
.B(n_1635),
.C(n_1637),
.Y(n_1817)
);

AOI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1811),
.A2(n_1620),
.B1(n_1582),
.B2(n_1619),
.Y(n_1818)
);

AND2x4_ASAP7_75t_L g1819 ( 
.A(n_1814),
.B(n_1670),
.Y(n_1819)
);

NOR2xp33_ASAP7_75t_L g1820 ( 
.A(n_1813),
.B(n_1681),
.Y(n_1820)
);

XOR2xp5_ASAP7_75t_L g1821 ( 
.A(n_1816),
.B(n_1526),
.Y(n_1821)
);

AOI22xp5_ASAP7_75t_L g1822 ( 
.A1(n_1818),
.A2(n_1681),
.B1(n_1607),
.B2(n_1608),
.Y(n_1822)
);

OAI211xp5_ASAP7_75t_L g1823 ( 
.A1(n_1815),
.A2(n_1653),
.B(n_1652),
.C(n_1648),
.Y(n_1823)
);

OAI211xp5_ASAP7_75t_L g1824 ( 
.A1(n_1820),
.A2(n_1817),
.B(n_1652),
.C(n_1653),
.Y(n_1824)
);

NOR2xp67_ASAP7_75t_L g1825 ( 
.A(n_1819),
.B(n_1648),
.Y(n_1825)
);

NOR2xp67_ASAP7_75t_L g1826 ( 
.A(n_1823),
.B(n_1648),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1825),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1827),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1828),
.Y(n_1829)
);

OA21x2_ASAP7_75t_L g1830 ( 
.A1(n_1828),
.A2(n_1824),
.B(n_1826),
.Y(n_1830)
);

OR2x2_ASAP7_75t_L g1831 ( 
.A(n_1829),
.B(n_1821),
.Y(n_1831)
);

OAI22x1_ASAP7_75t_L g1832 ( 
.A1(n_1830),
.A2(n_1822),
.B1(n_1648),
.B2(n_1649),
.Y(n_1832)
);

INVxp67_ASAP7_75t_L g1833 ( 
.A(n_1831),
.Y(n_1833)
);

AOI22xp5_ASAP7_75t_L g1834 ( 
.A1(n_1832),
.A2(n_1830),
.B1(n_1626),
.B2(n_1641),
.Y(n_1834)
);

AOI21xp5_ASAP7_75t_L g1835 ( 
.A1(n_1833),
.A2(n_1649),
.B(n_1652),
.Y(n_1835)
);

AOI22xp5_ASAP7_75t_L g1836 ( 
.A1(n_1835),
.A2(n_1834),
.B1(n_1652),
.B2(n_1653),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1836),
.Y(n_1837)
);

OAI221xp5_ASAP7_75t_R g1838 ( 
.A1(n_1837),
.A2(n_1555),
.B1(n_1641),
.B2(n_1626),
.C(n_1647),
.Y(n_1838)
);

AOI211xp5_ASAP7_75t_L g1839 ( 
.A1(n_1838),
.A2(n_1653),
.B(n_1649),
.C(n_1641),
.Y(n_1839)
);


endmodule