module fake_jpeg_21370_n_229 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_229);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_11;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx3_ASAP7_75t_L g12 ( 
.A(n_10),
.Y(n_12)
);

INVx8_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

INVx8_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_25),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_23),
.B(n_0),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_27),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_SL g32 ( 
.A(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_21),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_13),
.B1(n_19),
.B2(n_20),
.Y(n_34)
);

O2A1O1Ixp33_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_39),
.B(n_30),
.C(n_27),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_24),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_26),
.A2(n_13),
.B1(n_19),
.B2(n_22),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_36),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_42),
.B(n_43),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_35),
.B(n_24),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_36),
.Y(n_45)
);

AO21x1_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_56),
.B(n_57),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_36),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_46),
.B(n_49),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_35),
.A2(n_25),
.B(n_18),
.C(n_15),
.Y(n_47)
);

A2O1A1Ixp33_ASAP7_75t_L g64 ( 
.A1(n_47),
.A2(n_40),
.B(n_41),
.C(n_19),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_48),
.A2(n_33),
.B1(n_41),
.B2(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_25),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_37),
.B(n_22),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_50),
.B(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_34),
.B(n_15),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_18),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_53),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_39),
.B(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_18),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_41),
.A2(n_19),
.B1(n_13),
.B2(n_30),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_58),
.A2(n_33),
.B1(n_32),
.B2(n_31),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_54),
.A2(n_41),
.B1(n_40),
.B2(n_27),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_63),
.A2(n_69),
.B1(n_74),
.B2(n_48),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_55),
.Y(n_65)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_56),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_67),
.B(n_43),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_33),
.Y(n_69)
);

AOI32xp33_ASAP7_75t_L g70 ( 
.A1(n_49),
.A2(n_38),
.A3(n_40),
.B1(n_13),
.B2(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_72),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_45),
.B(n_38),
.C(n_28),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_71),
.B(n_50),
.Y(n_87)
);

OAI22xp33_ASAP7_75t_SL g74 ( 
.A1(n_42),
.A2(n_38),
.B1(n_33),
.B2(n_32),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_75),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_61),
.A2(n_46),
.B1(n_51),
.B2(n_52),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_80),
.B1(n_90),
.B2(n_69),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_77),
.B(n_81),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_78),
.B(n_79),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_66),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_61),
.A2(n_48),
.B1(n_44),
.B2(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_66),
.Y(n_83)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_83),
.Y(n_94)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_63),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_85),
.A2(n_73),
.B(n_62),
.Y(n_99)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_47),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_59),
.Y(n_88)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_88),
.B(n_59),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_21),
.Y(n_89)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_89),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_95),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_85),
.B(n_60),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_109),
.Y(n_128)
);

INVxp33_ASAP7_75t_L g97 ( 
.A(n_77),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_97),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_104),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_100),
.A2(n_108),
.B1(n_33),
.B2(n_31),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_82),
.A2(n_72),
.B(n_64),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_102),
.A2(n_75),
.B(n_90),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_71),
.C(n_73),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g105 ( 
.A(n_80),
.B(n_72),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_107),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_82),
.A2(n_68),
.B(n_70),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_101),
.B(n_108),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_83),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_76),
.A2(n_75),
.B1(n_68),
.B2(n_58),
.Y(n_108)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_79),
.Y(n_114)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_111),
.Y(n_116)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_114),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_115),
.A2(n_121),
.B(n_123),
.Y(n_148)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_47),
.C(n_86),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_21),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_29),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_102),
.Y(n_124)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_124),
.Y(n_146)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_126),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_101),
.A2(n_31),
.B1(n_28),
.B2(n_29),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_129),
.A2(n_136),
.B1(n_0),
.B2(n_1),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_101),
.A2(n_21),
.B(n_14),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_130),
.B(n_131),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_95),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_96),
.B(n_103),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_132),
.B(n_134),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g133 ( 
.A(n_97),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_133),
.Y(n_154)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_100),
.Y(n_134)
);

OA21x2_ASAP7_75t_SL g135 ( 
.A1(n_109),
.A2(n_21),
.B(n_14),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_135),
.B(n_8),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_0),
.B(n_1),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_120),
.B(n_104),
.C(n_106),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_139),
.B(n_150),
.C(n_152),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_140),
.A2(n_151),
.B1(n_112),
.B2(n_122),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_143),
.B(n_144),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_118),
.B(n_8),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_147),
.B(n_136),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_127),
.A2(n_17),
.B1(n_16),
.B2(n_14),
.Y(n_149)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_12),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_119),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_113),
.B(n_17),
.C(n_16),
.Y(n_152)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_155),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_128),
.B(n_12),
.Y(n_157)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_157),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_156),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_160),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_122),
.B1(n_124),
.B2(n_138),
.Y(n_160)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_137),
.Y(n_163)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_163),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_164),
.A2(n_172),
.B1(n_173),
.B2(n_130),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_146),
.A2(n_112),
.B1(n_121),
.B2(n_133),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_165),
.B(n_169),
.Y(n_176)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_141),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_167),
.Y(n_182)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_170),
.B(n_171),
.Y(n_179)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_148),
.A2(n_129),
.B1(n_115),
.B2(n_128),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_154),
.A2(n_147),
.B1(n_123),
.B2(n_148),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_174),
.B(n_178),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_139),
.C(n_150),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_177),
.B(n_183),
.C(n_159),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_160),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_161),
.B(n_152),
.Y(n_181)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_181),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_168),
.B(n_157),
.C(n_143),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_142),
.B(n_123),
.Y(n_184)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_185),
.B(n_186),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_165),
.A2(n_116),
.B(n_151),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_172),
.C(n_166),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_188),
.B(n_190),
.Y(n_203)
);

A2O1A1Ixp33_ASAP7_75t_SL g189 ( 
.A1(n_185),
.A2(n_140),
.B(n_166),
.C(n_125),
.Y(n_189)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_16),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_180),
.B(n_170),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_183),
.B(n_162),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_192),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_8),
.B1(n_9),
.B2(n_7),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_182),
.Y(n_197)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_197),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_196),
.B1(n_187),
.B2(n_194),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_192),
.B(n_179),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_189),
.A2(n_175),
.B(n_176),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_202),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_186),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_201),
.B(n_12),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_16),
.C(n_17),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_205),
.B(n_2),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_203),
.B(n_17),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_206),
.B(n_212),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g214 ( 
.A(n_208),
.B(n_213),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_210),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_204),
.B(n_5),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_201),
.B(n_5),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_209),
.B(n_202),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_2),
.Y(n_222)
);

NOR2xp67_ASAP7_75t_SL g216 ( 
.A(n_211),
.B(n_205),
.Y(n_216)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_216),
.Y(n_221)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_210),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_218),
.A2(n_207),
.B1(n_5),
.B2(n_4),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_220),
.A2(n_222),
.B(n_3),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_214),
.B(n_3),
.C(n_4),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_223),
.A2(n_217),
.B(n_219),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_224),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_225),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_223),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_221),
.Y(n_229)
);


endmodule