module real_jpeg_21390_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_307, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_307;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_292;
wire n_221;
wire n_249;
wire n_288;
wire n_300;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_301;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_299;
wire n_173;
wire n_115;
wire n_255;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_293;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_178;
wire n_76;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_305;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_304;
wire n_112;
wire n_42;
wire n_268;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_302;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_298;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_296;
wire n_134;
wire n_270;
wire n_223;
wire n_72;
wire n_159;
wire n_303;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_195;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_297;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_128;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_295;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

AOI22xp33_ASAP7_75t_L g148 ( 
.A1(n_0),
.A2(n_30),
.B1(n_31),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_0),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g161 ( 
.A1(n_0),
.A2(n_57),
.B1(n_58),
.B2(n_149),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_0),
.A2(n_49),
.B1(n_50),
.B2(n_149),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_0),
.A2(n_38),
.B1(n_39),
.B2(n_149),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_1),
.A2(n_57),
.B1(n_58),
.B2(n_89),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_1),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_1),
.A2(n_38),
.B1(n_39),
.B2(n_89),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_1),
.A2(n_30),
.B1(n_31),
.B2(n_89),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_1),
.A2(n_49),
.B1(n_50),
.B2(n_89),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_2),
.A2(n_57),
.B1(n_58),
.B2(n_65),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_2),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_2),
.A2(n_30),
.B1(n_31),
.B2(n_65),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_2),
.A2(n_38),
.B1(n_39),
.B2(n_65),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_65),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_3),
.A2(n_38),
.B1(n_39),
.B2(n_52),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_3),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_3),
.A2(n_49),
.B1(n_50),
.B2(n_52),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_3),
.A2(n_30),
.B1(n_31),
.B2(n_52),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_5),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_5),
.B(n_63),
.Y(n_181)
);

AOI21xp33_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_16),
.B(n_49),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_5),
.A2(n_38),
.B1(n_39),
.B2(n_153),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_5),
.A2(n_79),
.B1(n_80),
.B2(n_210),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_5),
.B(n_42),
.Y(n_222)
);

AOI21xp33_ASAP7_75t_L g239 ( 
.A1(n_5),
.A2(n_30),
.B(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_6),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g122 ( 
.A1(n_6),
.A2(n_30),
.B1(n_31),
.B2(n_56),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_6),
.A2(n_38),
.B1(n_39),
.B2(n_56),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_6),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_7),
.A2(n_30),
.B1(n_31),
.B2(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_7),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_7),
.A2(n_38),
.B1(n_39),
.B2(n_41),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_7),
.A2(n_41),
.B1(n_49),
.B2(n_50),
.Y(n_116)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_8),
.Y(n_80)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_8),
.Y(n_117)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_9),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_10),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_10),
.A2(n_30),
.B1(n_31),
.B2(n_126),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g197 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_126),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_10),
.A2(n_38),
.B1(n_39),
.B2(n_126),
.Y(n_243)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_12),
.A2(n_57),
.B1(n_58),
.B2(n_155),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_12),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_12),
.A2(n_30),
.B1(n_31),
.B2(n_155),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_12),
.A2(n_38),
.B1(n_39),
.B2(n_155),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_155),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g29 ( 
.A1(n_13),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_13),
.A2(n_32),
.B1(n_38),
.B2(n_39),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_13),
.A2(n_32),
.B1(n_57),
.B2(n_58),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_13),
.A2(n_32),
.B1(n_49),
.B2(n_50),
.Y(n_139)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_14),
.A2(n_35),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_14),
.A2(n_30),
.A3(n_39),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_15),
.A2(n_30),
.B1(n_31),
.B2(n_61),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_16),
.A2(n_38),
.B1(n_39),
.B2(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_16),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_16),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

BUFx3_ASAP7_75t_SL g39 ( 
.A(n_17),
.Y(n_39)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_104),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_90),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_22),
.B(n_90),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_69),
.C(n_75),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_23),
.A2(n_24),
.B1(n_69),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_25),
.A2(n_53),
.B1(n_67),
.B2(n_68),
.Y(n_24)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_25),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_43),
.B2(n_44),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_27),
.B(n_43),
.C(n_53),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_33),
.B1(n_40),
.B2(n_42),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_29),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_29),
.A2(n_34),
.B1(n_37),
.B2(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_30),
.B(n_61),
.Y(n_167)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

A2O1A1Ixp33_ASAP7_75t_L g34 ( 
.A1(n_31),
.A2(n_35),
.B(n_36),
.C(n_37),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_35),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_31),
.A2(n_62),
.B1(n_152),
.B2(n_167),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_31),
.B(n_153),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_33),
.A2(n_40),
.B1(n_42),
.B2(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_33),
.A2(n_42),
.B1(n_72),
.B2(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_33),
.A2(n_42),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_34),
.A2(n_37),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_34),
.A2(n_37),
.B1(n_150),
.B2(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_34),
.A2(n_37),
.B1(n_179),
.B2(n_239),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_34),
.A2(n_37),
.B1(n_122),
.B2(n_163),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_35),
.B(n_38),
.Y(n_235)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

A2O1A1Ixp33_ASAP7_75t_L g200 ( 
.A1(n_39),
.A2(n_47),
.B(n_153),
.C(n_201),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_43),
.A2(n_44),
.B1(n_98),
.B2(n_99),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_45),
.A2(n_48),
.B(n_51),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_45),
.A2(n_48),
.B1(n_51),
.B2(n_74),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_45),
.A2(n_48),
.B1(n_74),
.B2(n_85),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_45),
.A2(n_48),
.B1(n_85),
.B2(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_45),
.A2(n_48),
.B1(n_119),
.B2(n_141),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_45),
.A2(n_48),
.B1(n_141),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_45),
.A2(n_48),
.B1(n_204),
.B2(n_205),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_45),
.A2(n_48),
.B1(n_205),
.B2(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_45),
.A2(n_48),
.B1(n_225),
.B2(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_45),
.A2(n_48),
.B1(n_145),
.B2(n_243),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_48),
.B(n_153),
.Y(n_208)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_49),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_50),
.B(n_213),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_53),
.A2(n_68),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_59),
.B1(n_64),
.B2(n_66),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_55),
.A2(n_60),
.B1(n_63),
.B2(n_87),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_57),
.Y(n_58)
);

O2A1O1Ixp33_ASAP7_75t_L g60 ( 
.A1(n_57),
.A2(n_61),
.B(n_62),
.C(n_63),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_61),
.Y(n_62)
);

HAxp5_ASAP7_75t_SL g152 ( 
.A(n_57),
.B(n_153),
.CON(n_152),
.SN(n_152)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_59),
.A2(n_64),
.B1(n_66),
.B2(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_59),
.A2(n_66),
.B1(n_88),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_59),
.A2(n_66),
.B1(n_160),
.B2(n_161),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_59),
.A2(n_66),
.B1(n_125),
.B2(n_161),
.Y(n_281)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_60),
.A2(n_63),
.B1(n_152),
.B2(n_154),
.Y(n_151)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_69),
.A2(n_70),
.B(n_73),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g130 ( 
.A(n_69),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_73),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_72),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_75),
.A2(n_76),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_86),
.B2(n_307),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_84),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_78),
.A2(n_86),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_78),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_78),
.A2(n_84),
.B1(n_110),
.B2(n_296),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_81),
.B(n_83),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_79),
.A2(n_83),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_79),
.A2(n_116),
.B1(n_117),
.B2(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_79),
.A2(n_117),
.B1(n_139),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_79),
.A2(n_80),
.B1(n_169),
.B2(n_184),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_79),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_79),
.A2(n_80),
.B1(n_195),
.B2(n_210),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_79),
.A2(n_81),
.B1(n_197),
.B2(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_79),
.A2(n_80),
.B1(n_184),
.B2(n_227),
.Y(n_233)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_82),
.A2(n_193),
.B1(n_194),
.B2(n_196),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_84),
.Y(n_296)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_102),
.Y(n_90)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_97),
.B2(n_101),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_94),
.Y(n_101)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_131),
.B(n_305),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_127),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_106),
.B(n_127),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_111),
.C(n_112),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_107),
.B(n_111),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g301 ( 
.A1(n_112),
.A2(n_113),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_114),
.B(n_120),
.C(n_123),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_114),
.B(n_292),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_115),
.B(n_118),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_117),
.B(n_153),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_120),
.A2(n_123),
.B1(n_124),
.B2(n_293),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_120),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_299),
.B(n_304),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_133),
.A2(n_286),
.B(n_298),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_134),
.A2(n_185),
.B(n_268),
.C(n_285),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_170),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_135),
.B(n_170),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_156),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_137),
.B(n_142),
.C(n_156),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_138),
.B(n_140),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_146),
.C(n_151),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_148),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_157),
.B(n_165),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_158),
.A2(n_159),
.B1(n_162),
.B2(n_164),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_158),
.B(n_164),
.C(n_165),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_162),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_168),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_166),
.B(n_168),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_173),
.C(n_175),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_171),
.B(n_265),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_176),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_181),
.C(n_182),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_177),
.B(n_253),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_181),
.A2(n_182),
.B1(n_183),
.B2(n_254),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_181),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_183),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_186),
.B(n_267),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_262),
.B(n_266),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_248),
.B(n_261),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_229),
.B(n_247),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_190),
.A2(n_217),
.B(n_228),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_206),
.B(n_216),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_198),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_198),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_199),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_200),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_202),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_211),
.B(n_215),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_208),
.B(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_219),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_226),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_224),
.C(n_226),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_230),
.B(n_231),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_237),
.B1(n_245),
.B2(n_246),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_232),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_234),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_236),
.Y(n_240)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_237),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_241),
.B1(n_242),
.B2(n_244),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_238),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_244),
.C(n_245),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_249),
.B(n_250),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_255),
.B2(n_256),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_251),
.B(n_258),
.C(n_259),
.Y(n_263)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_257),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_258),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_263),
.B(n_264),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_269),
.B(n_270),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_271),
.A2(n_272),
.B1(n_273),
.B2(n_284),
.Y(n_270)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_271),
.Y(n_284)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_276),
.B2(n_277),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_274),
.B(n_277),
.C(n_284),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_280),
.C(n_283),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_281),
.B1(n_282),
.B2(n_283),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_281),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_282),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_287),
.B(n_288),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_297),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_294),
.B2(n_295),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_290),
.B(n_295),
.C(n_297),
.Y(n_300)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_300),
.B(n_301),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);


endmodule