module real_jpeg_29173_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_201;
wire n_49;
wire n_114;
wire n_252;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_194;
wire n_104;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_184;
wire n_56;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_155;
wire n_120;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_203;
wire n_192;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_195;
wire n_61;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_217;
wire n_210;
wire n_53;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_101;
wire n_182;
wire n_253;
wire n_96;
wire n_89;

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_0),
.A2(n_63),
.B1(n_64),
.B2(n_80),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_0),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_0),
.A2(n_57),
.B1(n_58),
.B2(n_80),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_0),
.A2(n_40),
.B1(n_41),
.B2(n_80),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_80),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_1),
.A2(n_32),
.B1(n_40),
.B2(n_41),
.Y(n_86)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

HB1xp67_ASAP7_75t_L g216 ( 
.A(n_2),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_SL g96 ( 
.A1(n_3),
.A2(n_58),
.B(n_62),
.C(n_97),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_3),
.Y(n_98)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_98),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_60),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_40),
.Y(n_181)
);

A2O1A1O1Ixp25_ASAP7_75t_L g183 ( 
.A1(n_3),
.A2(n_40),
.B(n_44),
.C(n_181),
.D(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_3),
.B(n_72),
.Y(n_188)
);

OAI21xp33_ASAP7_75t_L g212 ( 
.A1(n_3),
.A2(n_25),
.B(n_194),
.Y(n_212)
);

A2O1A1O1Ixp25_ASAP7_75t_L g224 ( 
.A1(n_3),
.A2(n_64),
.B(n_76),
.C(n_110),
.D(n_225),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_3),
.B(n_64),
.Y(n_225)
);

BUFx12_ASAP7_75t_L g62 ( 
.A(n_4),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_5),
.A2(n_26),
.B1(n_33),
.B2(n_84),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_5),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_7),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_7),
.A2(n_42),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g168 ( 
.A1(n_7),
.A2(n_26),
.B1(n_33),
.B2(n_42),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_8),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g152 ( 
.A1(n_8),
.A2(n_56),
.B1(n_63),
.B2(n_64),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_8),
.A2(n_40),
.B1(n_41),
.B2(n_56),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_56),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_9),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_10),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_10),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_10),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_67),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_10),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_228)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_11),
.B(n_40),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_11),
.A2(n_26),
.B1(n_33),
.B2(n_46),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_11),
.B(n_26),
.Y(n_182)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_12),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_13),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_13),
.A2(n_26),
.B1(n_33),
.B2(n_50),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_13),
.A2(n_50),
.B1(n_63),
.B2(n_64),
.Y(n_129)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_15),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_15),
.A2(n_63),
.B1(n_64),
.B2(n_73),
.Y(n_77)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_133),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_132),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_111),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_21),
.B(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_87),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_22),
.B(n_81),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_23),
.B(n_54),
.C(n_68),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_38),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_24),
.B(n_38),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_25),
.A2(n_34),
.B1(n_36),
.B2(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_25),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g119 ( 
.A1(n_25),
.A2(n_34),
.B(n_83),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_25),
.A2(n_103),
.B1(n_168),
.B2(n_169),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_25),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_25),
.B(n_196),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_29),
.A2(n_201),
.B(n_209),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_31),
.A2(n_35),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g180 ( 
.A1(n_33),
.A2(n_41),
.A3(n_46),
.B1(n_181),
.B2(n_182),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_33),
.B(n_214),
.Y(n_213)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_34),
.Y(n_203)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx5_ASAP7_75t_SL g169 ( 
.A(n_35),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_35),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_35),
.A2(n_210),
.B(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_39),
.A2(n_51),
.B(n_144),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_45),
.B(n_47),
.C(n_48),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_40),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

AOI32xp33_ASAP7_75t_L g232 ( 
.A1(n_40),
.A2(n_63),
.A3(n_225),
.B1(n_233),
.B2(n_234),
.Y(n_232)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_41),
.B(n_74),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_43),
.A2(n_49),
.B1(n_51),
.B2(n_86),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g244 ( 
.A1(n_43),
.A2(n_245),
.B(n_246),
.Y(n_244)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_44),
.A2(n_48),
.B1(n_116),
.B2(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_44),
.B(n_145),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_44),
.A2(n_48),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_51),
.B(n_146),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_51),
.A2(n_144),
.B(n_191),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g207 ( 
.A(n_51),
.B(n_98),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_53),
.A2(n_54),
.B1(n_68),
.B2(n_69),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_55),
.A2(n_59),
.B1(n_60),
.B2(n_66),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_55),
.Y(n_91)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_57),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_58),
.B1(n_61),
.B2(n_62),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_59),
.B(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_59),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_59),
.A2(n_148),
.B(n_149),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_65),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_60),
.B(n_94),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g60 ( 
.A1(n_61),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_60)
);

OAI21xp33_ASAP7_75t_L g97 ( 
.A1(n_61),
.A2(n_64),
.B(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_63),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_66),
.Y(n_126)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_75),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_70),
.A2(n_71),
.B1(n_106),
.B2(n_129),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_71),
.B(n_79),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_71),
.A2(n_75),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_72),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_72),
.A2(n_76),
.B1(n_108),
.B2(n_151),
.Y(n_150)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx6_ASAP7_75t_L g233 ( 
.A(n_74),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_76),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_82),
.B(n_85),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_86),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_87),
.A2(n_88),
.B1(n_154),
.B2(n_155),
.Y(n_153)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_95),
.C(n_104),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_89),
.A2(n_90),
.B1(n_104),
.B2(n_105),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_93),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_95),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_99),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_96),
.A2(n_99),
.B1(n_100),
.B2(n_164),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_96),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_98),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_101),
.A2(n_200),
.B1(n_202),
.B2(n_203),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_109),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_131),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_118),
.B2(n_119),
.Y(n_113)
);

CKINVDCx14_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_123),
.B2(n_130),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_121),
.Y(n_130)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_SL g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B(n_127),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_127),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_173),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_156),
.B(n_172),
.Y(n_135)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_136),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_153),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_137),
.B(n_153),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_140),
.C(n_141),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_158),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_140),
.B(n_141),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_147),
.C(n_150),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_143),
.B1(n_150),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_147),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_150),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_154),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_157),
.B(n_159),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_163),
.C(n_165),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_160),
.B(n_251),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_163),
.B(n_165),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_167),
.C(n_170),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_166),
.B(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_167),
.A2(n_170),
.B1(n_171),
.B2(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_167),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_168),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

NOR3xp33_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_253),
.C(n_254),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_248),
.B(n_252),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_236),
.B(n_247),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_220),
.B(n_235),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_197),
.B(n_219),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_185),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_179),
.B(n_185),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_183),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_180),
.B(n_183),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_184),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_187),
.B(n_190),
.C(n_192),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_191),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_193),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_196),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_205),
.B(n_218),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_204),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_204),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_201),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_211),
.B(n_217),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_207),
.B(n_208),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_212),
.B(n_213),
.Y(n_211)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_221),
.B(n_222),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_229),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_224),
.B(n_226),
.C(n_229),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_232),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_230),
.B(n_232),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_237),
.B(n_238),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_242),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_239),
.B(n_243),
.C(n_244),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_250),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_249),
.B(n_250),
.Y(n_252)
);


endmodule