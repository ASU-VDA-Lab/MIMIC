module real_jpeg_31956_n_15 (n_123, n_8, n_116, n_0, n_2, n_114, n_10, n_9, n_12, n_6, n_121, n_11, n_14, n_120, n_7, n_117, n_3, n_119, n_5, n_4, n_115, n_122, n_1, n_118, n_13, n_113, n_15);

input n_123;
input n_8;
input n_116;
input n_0;
input n_2;
input n_114;
input n_10;
input n_9;
input n_12;
input n_6;
input n_121;
input n_11;
input n_14;
input n_120;
input n_7;
input n_117;
input n_3;
input n_119;
input n_5;
input n_4;
input n_115;
input n_122;
input n_1;
input n_118;
input n_13;
input n_113;

output n_15;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_68;
wire n_83;
wire n_78;
wire n_104;
wire n_64;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_0),
.B(n_79),
.Y(n_78)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_0),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_1),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_1),
.B(n_93),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_2),
.B(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_3),
.Y(n_85)
);

AOI322xp5_ASAP7_75t_L g105 ( 
.A1(n_3),
.A2(n_81),
.A3(n_83),
.B1(n_87),
.B2(n_106),
.C1(n_108),
.C2(n_123),
.Y(n_105)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_4),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_4),
.B(n_89),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_5),
.A2(n_17),
.B1(n_18),
.B2(n_26),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

AOI221xp5_ASAP7_75t_L g48 ( 
.A1(n_6),
.A2(n_14),
.B1(n_49),
.B2(n_56),
.C(n_58),
.Y(n_48)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_7),
.Y(n_67)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_8),
.Y(n_55)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_9),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_9),
.B(n_98),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_11),
.B(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_12),
.B(n_30),
.Y(n_111)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_14),
.B(n_49),
.C(n_56),
.Y(n_61)
);

XOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_27),
.Y(n_15)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NOR2xp67_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_20),
.Y(n_18)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_22),
.B(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_22),
.B(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

AOI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_36),
.B(n_111),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_35),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_99),
.Y(n_98)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_34),
.Y(n_66)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

AOI31xp33_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_75),
.A3(n_96),
.B(n_101),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_69),
.C(n_70),
.Y(n_38)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_62),
.B(n_68),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_41),
.A2(n_48),
.B1(n_60),
.B2(n_61),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_44),
.Y(n_42)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_46),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_50),
.B(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_52),
.B(n_53),
.Y(n_51)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_56),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_115),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_63),
.B(n_67),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_63),
.B(n_67),
.Y(n_68)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_73),
.Y(n_71)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NOR3xp33_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_86),
.C(n_92),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_102),
.B(n_105),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

NOR3xp33_ASAP7_75t_L g106 ( 
.A(n_78),
.B(n_92),
.C(n_107),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_79),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_119),
.Y(n_83)
);

OA21x2_ASAP7_75t_SL g102 ( 
.A1(n_86),
.A2(n_103),
.B(n_104),
.Y(n_102)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_97),
.B(n_100),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_113),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_114),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_116),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_117),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_118),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_120),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_121),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_122),
.Y(n_99)
);


endmodule