module fake_aes_12580_n_28 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_28);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_28;
wire n_20;
wire n_23;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
BUFx6f_ASAP7_75t_L g11 ( .A(n_1), .Y(n_11) );
CKINVDCx5p33_ASAP7_75t_R g12 ( .A(n_7), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
NOR2xp33_ASAP7_75t_L g14 ( .A(n_4), .B(n_2), .Y(n_14) );
HB1xp67_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
AND2x2_ASAP7_75t_L g16 ( .A(n_6), .B(n_10), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_15), .B(n_0), .Y(n_17) );
BUFx8_ASAP7_75t_L g18 ( .A(n_13), .Y(n_18) );
AOI22xp33_ASAP7_75t_L g19 ( .A1(n_17), .A2(n_16), .B1(n_12), .B2(n_11), .Y(n_19) );
AND2x4_ASAP7_75t_L g20 ( .A(n_18), .B(n_11), .Y(n_20) );
BUFx4f_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_21), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_19), .Y(n_24) );
AND3x2_ASAP7_75t_L g25 ( .A(n_23), .B(n_14), .C(n_0), .Y(n_25) );
CKINVDCx5p33_ASAP7_75t_R g26 ( .A(n_24), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_27), .A2(n_25), .B1(n_3), .B2(n_9), .Y(n_28) );
endmodule