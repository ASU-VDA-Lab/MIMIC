module fake_jpeg_2534_n_164 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_11;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_3),
.Y(n_11)
);

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_4),
.Y(n_12)
);

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

BUFx2_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_13),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_29),
.B(n_42),
.Y(n_67)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_20),
.B(n_1),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_31),
.B(n_33),
.Y(n_85)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_32),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_20),
.B(n_23),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_34),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_10),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_38),
.Y(n_74)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_11),
.B(n_19),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_12),
.B(n_9),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_12),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_46),
.Y(n_71)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_18),
.B(n_19),
.Y(n_46)
);

AO22x1_ASAP7_75t_L g47 ( 
.A1(n_17),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g86 ( 
.A(n_47),
.B(n_53),
.Y(n_86)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_52),
.Y(n_72)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_51),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_5),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_21),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

BUFx10_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_57),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_24),
.B(n_6),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_59),
.Y(n_80)
);

INVx4_ASAP7_75t_SL g59 ( 
.A(n_25),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_25),
.B(n_6),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_60),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_28),
.B(n_20),
.Y(n_61)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_62),
.B(n_63),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_65),
.Y(n_88)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_15),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_44),
.A2(n_52),
.B1(n_46),
.B2(n_60),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_76),
.A2(n_71),
.B1(n_80),
.B2(n_83),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_31),
.B(n_33),
.C(n_58),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_87),
.B(n_89),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_36),
.B(n_42),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_75),
.Y(n_94)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_47),
.B1(n_39),
.B2(n_54),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_95),
.Y(n_117)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_99),
.Y(n_122)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_77),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_110),
.B1(n_90),
.B2(n_79),
.Y(n_115)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_86),
.A2(n_85),
.B1(n_88),
.B2(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_103),
.B(n_105),
.Y(n_113)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_78),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_104),
.B(n_106),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_86),
.A2(n_85),
.B1(n_93),
.B2(n_68),
.Y(n_105)
);

INVx13_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_78),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_109),
.Y(n_124)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_90),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_68),
.A2(n_75),
.B1(n_72),
.B2(n_67),
.Y(n_110)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_111),
.B(n_112),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_81),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_115),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_91),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_81),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_91),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_126),
.B(n_101),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_95),
.B1(n_111),
.B2(n_110),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_113),
.B1(n_115),
.B2(n_119),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_116),
.Y(n_129)
);

NOR3xp33_ASAP7_75t_L g137 ( 
.A(n_129),
.B(n_133),
.C(n_118),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_117),
.A2(n_109),
.B1(n_69),
.B2(n_102),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_130),
.A2(n_126),
.B(n_124),
.Y(n_142)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_121),
.Y(n_131)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_104),
.C(n_69),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_134),
.B(n_120),
.C(n_123),
.Y(n_139)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_123),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_118),
.B(n_92),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_136),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_137),
.A2(n_142),
.B(n_132),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_138),
.B(n_143),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_139),
.B(n_124),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_134),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_145),
.B(n_148),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_129),
.B1(n_128),
.B2(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_146),
.Y(n_152)
);

XOR2x1_ASAP7_75t_SL g149 ( 
.A(n_143),
.B(n_128),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_149),
.A2(n_140),
.B(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_122),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_150),
.B(n_122),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_151),
.A2(n_147),
.B(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_155),
.A2(n_151),
.B(n_152),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_153),
.B(n_145),
.C(n_127),
.Y(n_156)
);

BUFx24_ASAP7_75t_SL g158 ( 
.A(n_156),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_114),
.B(n_120),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g160 ( 
.A1(n_158),
.A2(n_157),
.A3(n_141),
.B1(n_131),
.B2(n_116),
.C1(n_94),
.C2(n_121),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_160),
.A2(n_161),
.B(n_106),
.C(n_114),
.Y(n_162)
);

BUFx24_ASAP7_75t_SL g163 ( 
.A(n_162),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_92),
.Y(n_164)
);


endmodule