module fake_jpeg_11057_n_55 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_55);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_55;

wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_22;
wire n_51;
wire n_47;
wire n_40;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

BUFx5_ASAP7_75t_L g20 ( 
.A(n_17),
.Y(n_20)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_2),
.B(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_13),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_10),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_31),
.B1(n_25),
.B2(n_22),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_28),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_20),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g30 ( 
.A(n_23),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_3),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_22),
.A2(n_25),
.B1(n_24),
.B2(n_26),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_32),
.A2(n_34),
.B1(n_5),
.B2(n_6),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_33),
.A2(n_27),
.B(n_28),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_29),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_28),
.Y(n_35)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_35),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_4),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_42),
.C(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_6),
.Y(n_45)
);

A2O1A1O1Ixp25_ASAP7_75t_L g42 ( 
.A1(n_32),
.A2(n_12),
.B(n_7),
.C(n_8),
.D(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_38),
.C(n_16),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_49),
.C(n_19),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_38),
.C(n_15),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_51),
.B(n_47),
.C(n_42),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_53),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_54),
.B(n_50),
.Y(n_55)
);


endmodule