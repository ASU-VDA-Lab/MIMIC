module fake_jpeg_20886_n_287 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_287);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_287;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_91;
wire n_54;
wire n_33;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx10_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_21),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_SL g50 ( 
.A(n_36),
.Y(n_50)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_8),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g46 ( 
.A(n_37),
.B(n_20),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_39),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_43),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_22),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_54),
.Y(n_68)
);

AOI21xp33_ASAP7_75t_L g76 ( 
.A1(n_46),
.A2(n_30),
.B(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_22),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_57),
.Y(n_96)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_35),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_27),
.Y(n_53)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_37),
.B(n_27),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_55),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_39),
.B(n_20),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_59),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_30),
.Y(n_59)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_60),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_45),
.A2(n_32),
.B1(n_43),
.B2(n_28),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_61),
.A2(n_65),
.B1(n_75),
.B2(n_80),
.Y(n_124)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_62),
.Y(n_101)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_64),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_44),
.A2(n_45),
.B1(n_58),
.B2(n_48),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_36),
.C(n_22),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_91),
.C(n_96),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_32),
.B1(n_24),
.B2(n_28),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g113 ( 
.A(n_67),
.Y(n_113)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_32),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_70),
.B(n_79),
.Y(n_102)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_74),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_54),
.A2(n_43),
.B1(n_24),
.B2(n_28),
.Y(n_75)
);

BUFx24_ASAP7_75t_SL g107 ( 
.A(n_76),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_46),
.A2(n_17),
.B1(n_24),
.B2(n_30),
.Y(n_78)
);

AOI32xp33_ASAP7_75t_L g116 ( 
.A1(n_78),
.A2(n_87),
.A3(n_88),
.B1(n_33),
.B2(n_29),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_55),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_48),
.A2(n_19),
.B1(n_17),
.B2(n_23),
.Y(n_80)
);

AO22x2_ASAP7_75t_L g82 ( 
.A1(n_50),
.A2(n_42),
.B1(n_41),
.B2(n_22),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_82),
.B(n_84),
.Y(n_117)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_53),
.B(n_52),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_52),
.B(n_42),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_85),
.B(n_89),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_19),
.B1(n_23),
.B2(n_26),
.Y(n_86)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_95),
.B1(n_50),
.B2(n_56),
.Y(n_99)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_50),
.B(n_18),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_60),
.A2(n_26),
.B1(n_33),
.B2(n_22),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_57),
.B1(n_33),
.B2(n_22),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_51),
.B(n_57),
.C(n_56),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_56),
.Y(n_92)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_92),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_26),
.B1(n_18),
.B2(n_29),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_26),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_98),
.B(n_104),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_99),
.A2(n_93),
.B1(n_29),
.B2(n_18),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_0),
.B(n_1),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_100),
.A2(n_0),
.B(n_1),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_68),
.B(n_66),
.Y(n_104)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_105),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_57),
.C(n_29),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_97),
.Y(n_137)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_81),
.Y(n_112)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_112),
.Y(n_128)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_81),
.Y(n_115)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_115),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_116),
.A2(n_88),
.B1(n_82),
.B2(n_94),
.Y(n_126)
);

MAJx2_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_31),
.C(n_25),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_91),
.B(n_78),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_74),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_121),
.B(n_122),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_84),
.B(n_31),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_85),
.B(n_31),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_34),
.Y(n_141)
);

O2A1O1Ixp33_ASAP7_75t_L g125 ( 
.A1(n_117),
.A2(n_87),
.B(n_82),
.C(n_67),
.Y(n_125)
);

AO22x1_ASAP7_75t_L g177 ( 
.A1(n_125),
.A2(n_150),
.B1(n_2),
.B2(n_3),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_126),
.A2(n_132),
.B1(n_140),
.B2(n_152),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_127),
.B(n_141),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_113),
.A2(n_77),
.B1(n_63),
.B2(n_82),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_114),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_131),
.B(n_103),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_94),
.B1(n_69),
.B2(n_64),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_83),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_134),
.B(n_135),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_110),
.A2(n_73),
.B(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_137),
.B(n_147),
.Y(n_163)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_108),
.Y(n_138)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_108),
.Y(n_139)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_97),
.A2(n_71),
.B1(n_62),
.B2(n_90),
.Y(n_140)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_142),
.Y(n_165)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_115),
.Y(n_143)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_143),
.Y(n_167)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_111),
.Y(n_144)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_144),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_101),
.B1(n_109),
.B2(n_111),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_124),
.A2(n_93),
.B1(n_18),
.B2(n_10),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_146),
.A2(n_151),
.B1(n_153),
.B2(n_7),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_102),
.B(n_25),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g175 ( 
.A(n_148),
.B(n_1),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_104),
.B(n_34),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_122),
.A2(n_9),
.B1(n_16),
.B2(n_15),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_106),
.A2(n_34),
.B1(n_25),
.B2(n_3),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_123),
.A2(n_98),
.B1(n_118),
.B2(n_100),
.Y(n_153)
);

BUFx2_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_154),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_155),
.A2(n_174),
.B1(n_180),
.B2(n_181),
.Y(n_197)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_158),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_133),
.C(n_150),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_169),
.C(n_173),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_125),
.A2(n_101),
.B1(n_119),
.B2(n_114),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_166),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_205)
);

AND2x4_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_120),
.Y(n_168)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_143),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_133),
.B(n_120),
.C(n_119),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g171 ( 
.A(n_128),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_172),
.Y(n_198)
);

INVx13_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_153),
.B(n_8),
.C(n_14),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_177),
.Y(n_187)
);

AND2x6_ASAP7_75t_L g176 ( 
.A(n_140),
.B(n_127),
.Y(n_176)
);

A2O1A1O1Ixp25_ASAP7_75t_L g192 ( 
.A1(n_176),
.A2(n_136),
.B(n_9),
.C(n_5),
.D(n_6),
.Y(n_192)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_138),
.Y(n_178)
);

INVx1_ASAP7_75t_SL g202 ( 
.A(n_178),
.Y(n_202)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_139),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_179),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_146),
.A2(n_149),
.B1(n_145),
.B2(n_135),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_149),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_181)
);

INVx13_ASAP7_75t_L g182 ( 
.A(n_128),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_182),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_162),
.A2(n_148),
.B(n_129),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g213 ( 
.A1(n_183),
.A2(n_186),
.B(n_188),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_169),
.Y(n_184)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_162),
.A2(n_144),
.B(n_134),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_156),
.A2(n_151),
.B1(n_134),
.B2(n_142),
.Y(n_190)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_190),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_168),
.B(n_152),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_191),
.B(n_194),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_192),
.Y(n_217)
);

A2O1A1O1Ixp25_ASAP7_75t_L g193 ( 
.A1(n_176),
.A2(n_168),
.B(n_159),
.C(n_161),
.D(n_177),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_SL g220 ( 
.A(n_193),
.B(n_164),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_170),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_159),
.B(n_136),
.C(n_11),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_199),
.C(n_173),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_163),
.B(n_11),
.C(n_14),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_165),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_206),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_174),
.B(n_2),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_204),
.B(n_205),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_167),
.Y(n_206)
);

AOI22x1_ASAP7_75t_L g208 ( 
.A1(n_191),
.A2(n_168),
.B1(n_166),
.B2(n_156),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_200),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_203),
.B(n_172),
.Y(n_209)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_209),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_203),
.B(n_164),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_210),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_196),
.B1(n_183),
.B2(n_193),
.Y(n_228)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_192),
.Y(n_215)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_215),
.Y(n_230)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_160),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_219),
.A2(n_224),
.B(n_185),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_220),
.B(n_195),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_189),
.B(n_182),
.Y(n_221)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_221),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_195),
.B(n_157),
.C(n_180),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_187),
.C(n_188),
.Y(n_235)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_223),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g224 ( 
.A(n_186),
.B(n_175),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_197),
.A2(n_154),
.B1(n_181),
.B2(n_14),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_225),
.A2(n_205),
.B1(n_187),
.B2(n_197),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_226),
.B(n_228),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g229 ( 
.A(n_219),
.B(n_200),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_229),
.A2(n_185),
.B(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_231),
.A2(n_236),
.B1(n_213),
.B2(n_207),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_214),
.B(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_211),
.C(n_199),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_239),
.B(n_219),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_214),
.B(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_238),
.Y(n_244)
);

XNOR2x2_ASAP7_75t_SL g239 ( 
.A(n_216),
.B(n_202),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_212),
.A2(n_208),
.B1(n_222),
.B2(n_213),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_238),
.Y(n_245)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_245),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_246),
.A2(n_252),
.B1(n_229),
.B2(n_230),
.Y(n_264)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_247),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_248),
.A2(n_231),
.B1(n_243),
.B2(n_236),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_218),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_220),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_250),
.B(n_251),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_240),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_227),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_237),
.B(n_229),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_241),
.C(n_232),
.Y(n_262)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_247),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_258),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_253),
.B(n_217),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_262),
.B(n_242),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g263 ( 
.A(n_251),
.B(n_239),
.Y(n_263)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_263),
.A2(n_250),
.B(n_215),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_246),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_262),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_265),
.B(n_267),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_255),
.B(n_242),
.C(n_254),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_266),
.B(n_255),
.C(n_263),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_270),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_259),
.A2(n_256),
.B1(n_244),
.B2(n_257),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_269),
.B(n_272),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_276),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_271),
.B(n_233),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_274),
.B(n_266),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_279),
.B(n_281),
.Y(n_282)
);

NOR3xp33_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_269),
.C(n_225),
.Y(n_280)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_280),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_SL g281 ( 
.A1(n_273),
.A2(n_11),
.B(n_13),
.C(n_16),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_282),
.A2(n_278),
.B(n_277),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_284),
.B(n_283),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_285),
.A2(n_13),
.B(n_16),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_286),
.B(n_13),
.Y(n_287)
);


endmodule