module fake_jpeg_2402_n_196 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_196);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_196;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_11),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_44),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_12),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_4),
.B(n_8),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_10),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_15),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_9),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_1),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_10),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_67),
.B(n_0),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_73),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_71),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_59),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_58),
.B(n_0),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_1),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_74),
.B(n_76),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_2),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_77),
.Y(n_84)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_71),
.A2(n_69),
.B1(n_50),
.B2(n_59),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_82),
.B1(n_54),
.B2(n_65),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_81),
.B(n_68),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_77),
.A2(n_69),
.B1(n_50),
.B2(n_53),
.Y(n_82)
);

INVx13_ASAP7_75t_L g85 ( 
.A(n_75),
.Y(n_85)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_85),
.Y(n_101)
);

OA22x2_ASAP7_75t_L g87 ( 
.A1(n_75),
.A2(n_54),
.B1(n_64),
.B2(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_49),
.B1(n_60),
.B2(n_52),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g88 ( 
.A1(n_72),
.A2(n_64),
.B(n_60),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_88),
.B(n_65),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_74),
.Y(n_89)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_89),
.Y(n_105)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_76),
.Y(n_91)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_91),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_92),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_89),
.B(n_66),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_93),
.B(n_104),
.Y(n_119)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_84),
.Y(n_94)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_94),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_103),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_87),
.B1(n_49),
.B2(n_60),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_96),
.A2(n_98),
.B1(n_6),
.B2(n_7),
.Y(n_128)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g111 ( 
.A(n_100),
.B(n_88),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_86),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_102),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_85),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_66),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_57),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_108),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_82),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_63),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_109),
.B(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_111),
.B(n_7),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_27),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_87),
.C(n_79),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_114),
.B(n_117),
.C(n_19),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_100),
.A2(n_87),
.B1(n_86),
.B2(n_79),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_116),
.B1(n_120),
.B2(n_124),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_107),
.A2(n_55),
.B1(n_48),
.B2(n_78),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_105),
.B(n_106),
.Y(n_117)
);

AOI22x1_ASAP7_75t_SL g120 ( 
.A1(n_105),
.A2(n_94),
.B1(n_102),
.B2(n_101),
.Y(n_120)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_94),
.Y(n_122)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_97),
.B(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g137 ( 
.A(n_123),
.B(n_12),
.Y(n_137)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_99),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_129),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_99),
.A2(n_5),
.B(n_6),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_16),
.B(n_17),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_128),
.Y(n_130)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_94),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_134),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_133),
.A2(n_140),
.B(n_141),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_110),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_119),
.B(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_135),
.B(n_139),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_136),
.B(n_137),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_111),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_SL g140 ( 
.A1(n_126),
.A2(n_13),
.B(n_14),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_117),
.B(n_17),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_112),
.Y(n_144)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_18),
.Y(n_145)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_145),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_127),
.B(n_18),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_146),
.Y(n_158)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_120),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_115),
.B(n_118),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_148),
.Y(n_166)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_114),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_151),
.B(n_144),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_32),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_20),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_147),
.A2(n_149),
.B(n_132),
.Y(n_152)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_152),
.B(n_153),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_130),
.A2(n_21),
.B1(n_22),
.B2(n_23),
.Y(n_153)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_150),
.A2(n_24),
.B(n_25),
.C(n_28),
.D(n_31),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_162),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_161),
.B(n_168),
.Y(n_173)
);

A2O1A1O1Ixp25_ASAP7_75t_L g162 ( 
.A1(n_138),
.A2(n_33),
.B(n_34),
.C(n_36),
.D(n_37),
.Y(n_162)
);

AOI322xp5_ASAP7_75t_L g163 ( 
.A1(n_130),
.A2(n_39),
.A3(n_41),
.B1(n_43),
.B2(n_45),
.C1(n_46),
.C2(n_47),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

FAx1_ASAP7_75t_SL g164 ( 
.A(n_139),
.B(n_141),
.CI(n_143),
.CON(n_164),
.SN(n_164)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_168),
.A2(n_131),
.B1(n_134),
.B2(n_158),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_169),
.B(n_171),
.Y(n_180)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_160),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_167),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_172),
.B(n_173),
.Y(n_182)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

INVxp33_ASAP7_75t_SL g181 ( 
.A(n_174),
.Y(n_181)
);

AOI321xp33_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_154),
.A3(n_155),
.B1(n_166),
.B2(n_164),
.C(n_165),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_170),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_161),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_177),
.Y(n_187)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_180),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_184),
.B(n_185),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_182),
.B(n_183),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_186),
.B(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_159),
.Y(n_190)
);

OAI221xp5_ASAP7_75t_L g192 ( 
.A1(n_190),
.A2(n_175),
.B1(n_181),
.B2(n_164),
.C(n_162),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_177),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_191),
.B(n_192),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_193),
.A2(n_189),
.B(n_188),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_194),
.B(n_181),
.C(n_153),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_195),
.B(n_156),
.Y(n_196)
);


endmodule