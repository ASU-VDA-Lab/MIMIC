module fake_jpeg_3088_n_455 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_455);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx10_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx12_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_6),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_9),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx4f_ASAP7_75t_SL g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_5),
.Y(n_41)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_10),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_9),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_45),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_48),
.B(n_49),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_17),
.B(n_32),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g114 ( 
.A(n_50),
.Y(n_114)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

INVx2_ASAP7_75t_SL g139 ( 
.A(n_51),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_52),
.Y(n_127)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_53),
.Y(n_125)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_28),
.Y(n_54)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_54),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_55),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_57),
.Y(n_104)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_59),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_0),
.CON(n_62),
.SN(n_62)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_62),
.B(n_19),
.Y(n_123)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_33),
.B(n_15),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_63),
.B(n_69),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_17),
.B(n_32),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_64),
.B(n_65),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_33),
.B(n_14),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_66),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_22),
.B(n_15),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_67),
.B(n_11),
.Y(n_102)
);

BUFx12f_ASAP7_75t_L g68 ( 
.A(n_20),
.Y(n_68)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_68),
.Y(n_107)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_16),
.Y(n_71)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_71),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_20),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_38),
.Y(n_75)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_75),
.Y(n_136)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_41),
.Y(n_78)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_78),
.Y(n_112)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_79),
.B(n_80),
.Y(n_100)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_16),
.Y(n_81)
);

INVx6_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_82),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_26),
.B(n_14),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_47),
.Y(n_110)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_38),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_18),
.Y(n_85)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_35),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_86),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_87),
.Y(n_98)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_46),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_89),
.B(n_91),
.Y(n_131)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_90),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_35),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_20),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_19),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_93),
.A2(n_42),
.B1(n_31),
.B2(n_24),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_47),
.B1(n_37),
.B2(n_34),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_95),
.A2(n_119),
.B1(n_126),
.B2(n_56),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_102),
.B(n_105),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_63),
.B(n_26),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_110),
.B(n_137),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_55),
.A2(n_42),
.B1(n_26),
.B2(n_37),
.Y(n_113)
);

AO22x1_ASAP7_75t_SL g177 ( 
.A1(n_113),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_71),
.A2(n_44),
.B1(n_43),
.B2(n_18),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_115),
.A2(n_31),
.B1(n_24),
.B2(n_21),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_22),
.B1(n_34),
.B2(n_30),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_88),
.B(n_44),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_121),
.B(n_122),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_43),
.Y(n_122)
);

CKINVDCx14_ASAP7_75t_R g179 ( 
.A(n_123),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_30),
.B1(n_25),
.B2(n_23),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_50),
.B(n_36),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_132),
.B(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_58),
.B(n_29),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_73),
.B(n_23),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_1),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_62),
.A2(n_27),
.B1(n_29),
.B2(n_25),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_140),
.A2(n_19),
.B(n_31),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_50),
.B(n_27),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g152 ( 
.A(n_144),
.Y(n_152)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_70),
.B(n_78),
.C(n_21),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_SL g222 ( 
.A(n_147),
.B(n_157),
.Y(n_222)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_125),
.Y(n_149)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_150),
.Y(n_214)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g198 ( 
.A(n_153),
.Y(n_198)
);

O2A1O1Ixp33_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_59),
.B(n_91),
.C(n_93),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_154),
.A2(n_156),
.B(n_182),
.Y(n_209)
);

O2A1O1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_138),
.A2(n_54),
.B(n_24),
.C(n_19),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_82),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_113),
.A2(n_53),
.B1(n_74),
.B2(n_68),
.Y(n_158)
);

OAI21xp33_ASAP7_75t_SL g232 ( 
.A1(n_158),
.A2(n_164),
.B(n_167),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_130),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_159),
.Y(n_234)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_160),
.Y(n_197)
);

BUFx2_ASAP7_75t_SL g161 ( 
.A(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_109),
.Y(n_162)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_162),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_114),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_165),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_166),
.B(n_168),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_100),
.A2(n_74),
.B1(n_68),
.B2(n_52),
.Y(n_167)
);

AND2x2_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_52),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_122),
.A2(n_60),
.B1(n_61),
.B2(n_92),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_116),
.Y(n_205)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_135),
.Y(n_170)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_170),
.Y(n_230)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_103),
.A2(n_146),
.B1(n_98),
.B2(n_115),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_140),
.A2(n_118),
.B1(n_94),
.B2(n_90),
.Y(n_172)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_127),
.Y(n_173)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_139),
.B(n_1),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_174),
.B(n_175),
.Y(n_236)
);

OAI22xp33_ASAP7_75t_L g224 ( 
.A1(n_177),
.A2(n_107),
.B1(n_112),
.B2(n_19),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_117),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_180),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_131),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_120),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_181),
.B(n_184),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_99),
.A2(n_31),
.B(n_24),
.Y(n_182)
);

BUFx2_ASAP7_75t_SL g183 ( 
.A(n_134),
.Y(n_183)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_129),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_104),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_185),
.B(n_189),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g186 ( 
.A(n_104),
.B(n_136),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_186),
.A2(n_127),
.B(n_19),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_96),
.Y(n_187)
);

INVx8_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_139),
.B(n_11),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_13),
.Y(n_213)
);

INVx3_ASAP7_75t_L g189 ( 
.A(n_106),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_136),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_190),
.B(n_192),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_96),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_120),
.Y(n_192)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_97),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_193),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g194 ( 
.A(n_114),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_194),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_195),
.A2(n_21),
.B1(n_31),
.B2(n_24),
.Y(n_221)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_106),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_196),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_179),
.A2(n_101),
.B1(n_116),
.B2(n_145),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_200),
.B(n_202),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_128),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_205),
.B(n_224),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_101),
.B1(n_145),
.B2(n_97),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_210),
.A2(n_211),
.B1(n_237),
.B2(n_191),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_152),
.A2(n_142),
.B1(n_141),
.B2(n_129),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_159),
.B(n_124),
.C(n_111),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_212),
.B(n_217),
.C(n_238),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_213),
.B(n_148),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_142),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_216),
.B(n_220),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_147),
.B(n_111),
.C(n_133),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_151),
.B(n_12),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_219),
.B(n_149),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_174),
.B(n_141),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_221),
.A2(n_182),
.B1(n_108),
.B2(n_157),
.Y(n_255)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_223),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_152),
.A2(n_107),
.B1(n_111),
.B2(n_133),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g273 ( 
.A(n_225),
.B(n_2),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_L g237 ( 
.A1(n_171),
.A2(n_21),
.B1(n_133),
.B2(n_112),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_108),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g282 ( 
.A(n_240),
.B(n_244),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_236),
.B(n_156),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_241),
.B(n_251),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_166),
.B(n_154),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_242),
.A2(n_270),
.B(n_223),
.Y(n_280)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_197),
.Y(n_243)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_243),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_234),
.B(n_189),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_197),
.Y(n_245)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_245),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_181),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_250),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_168),
.C(n_157),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_249),
.B(n_262),
.C(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_236),
.B(n_168),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_236),
.B(n_190),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_207),
.Y(n_252)
);

INVx13_ASAP7_75t_L g281 ( 
.A(n_252),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_206),
.B(n_163),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_254),
.B(n_259),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_274),
.B1(n_228),
.B2(n_210),
.Y(n_289)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_231),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_256),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_257),
.A2(n_275),
.B1(n_235),
.B2(n_199),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_239),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_186),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_260),
.B(n_264),
.Y(n_293)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_261),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_186),
.C(n_196),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_222),
.B(n_186),
.C(n_170),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_219),
.B(n_153),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_265),
.Y(n_301)
);

BUFx12_ASAP7_75t_L g266 ( 
.A(n_229),
.Y(n_266)
);

CKINVDCx10_ASAP7_75t_R g287 ( 
.A(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_216),
.B(n_177),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_267),
.B(n_271),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_212),
.B(n_177),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_269),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_150),
.C(n_195),
.Y(n_269)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_209),
.A2(n_108),
.B(n_173),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_220),
.B(n_193),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_208),
.B(n_187),
.Y(n_272)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_272),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g295 ( 
.A1(n_273),
.A2(n_274),
.B1(n_255),
.B2(n_215),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_209),
.A2(n_21),
.B1(n_3),
.B2(n_4),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_228),
.B(n_10),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_217),
.B(n_2),
.Y(n_277)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_277),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_267),
.A2(n_221),
.B1(n_226),
.B2(n_232),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_278),
.A2(n_283),
.B1(n_289),
.B2(n_310),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_280),
.A2(n_295),
.B(n_270),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_276),
.A2(n_205),
.B1(n_200),
.B2(n_204),
.Y(n_283)
);

OA21x2_ASAP7_75t_L g286 ( 
.A1(n_241),
.A2(n_211),
.B(n_227),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_290),
.Y(n_317)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_242),
.A2(n_201),
.B(n_227),
.Y(n_290)
);

AND2x6_ASAP7_75t_L g292 ( 
.A(n_246),
.B(n_225),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_292),
.B(n_246),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_204),
.B1(n_203),
.B2(n_233),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_294),
.Y(n_320)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_243),
.Y(n_298)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_298),
.Y(n_332)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_245),
.Y(n_299)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_299),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_273),
.A2(n_203),
.B1(n_233),
.B2(n_215),
.Y(n_302)
);

NAND4xp25_ASAP7_75t_SL g341 ( 
.A(n_302),
.B(n_266),
.C(n_199),
.D(n_218),
.Y(n_341)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_261),
.Y(n_307)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_271),
.Y(n_308)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_308),
.Y(n_323)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_272),
.Y(n_309)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_309),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_253),
.A2(n_218),
.B1(n_198),
.B2(n_229),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_311),
.B(n_230),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_312),
.B(n_334),
.Y(n_349)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_287),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_313),
.B(n_329),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_213),
.Y(n_314)
);

NAND3xp33_ASAP7_75t_L g351 ( 
.A(n_314),
.B(n_301),
.C(n_285),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_279),
.B(n_249),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_315),
.B(n_324),
.C(n_327),
.Y(n_345)
);

AOI221xp5_ASAP7_75t_L g319 ( 
.A1(n_306),
.A2(n_251),
.B1(n_262),
.B2(n_263),
.C(n_260),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_319),
.A2(n_331),
.B1(n_335),
.B2(n_304),
.Y(n_366)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_321),
.A2(n_330),
.B(n_340),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_284),
.B(n_277),
.C(n_268),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_325),
.Y(n_346)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_299),
.Y(n_326)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_326),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_284),
.B(n_269),
.C(n_258),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_279),
.B(n_250),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_328),
.B(n_333),
.C(n_336),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_287),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g330 ( 
.A1(n_280),
.A2(n_273),
.B(n_247),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_278),
.A2(n_253),
.B1(n_247),
.B2(n_259),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_258),
.C(n_256),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_300),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g335 ( 
.A1(n_303),
.A2(n_253),
.B1(n_252),
.B2(n_275),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_198),
.C(n_230),
.Y(n_336)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_338),
.Y(n_352)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_291),
.Y(n_339)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_339),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_290),
.A2(n_266),
.B(n_235),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_341),
.Y(n_354)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_323),
.B(n_337),
.Y(n_342)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_342),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g343 ( 
.A(n_336),
.Y(n_343)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_343),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_322),
.A2(n_303),
.B1(n_290),
.B2(n_286),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_344),
.A2(n_348),
.B1(n_317),
.B2(n_335),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_333),
.B(n_309),
.Y(n_347)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_347),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_322),
.A2(n_289),
.B1(n_305),
.B2(n_288),
.Y(n_348)
);

FAx1_ASAP7_75t_SL g350 ( 
.A(n_327),
.B(n_293),
.CI(n_292),
.CON(n_350),
.SN(n_350)
);

FAx1_ASAP7_75t_SL g383 ( 
.A(n_350),
.B(n_310),
.CI(n_341),
.CON(n_383),
.SN(n_383)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_351),
.B(n_362),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_315),
.B(n_293),
.C(n_305),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_356),
.B(n_359),
.C(n_320),
.Y(n_372)
);

AND2x2_ASAP7_75t_SL g357 ( 
.A(n_317),
.B(n_308),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_357),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_324),
.B(n_297),
.C(n_307),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_339),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_360),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_328),
.B(n_294),
.Y(n_361)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_361),
.B(n_363),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_304),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_331),
.B(n_286),
.Y(n_363)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_318),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_365),
.B(n_316),
.Y(n_384)
);

XOR2x2_ASAP7_75t_L g379 ( 
.A(n_366),
.B(n_283),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_SL g368 ( 
.A(n_361),
.B(n_321),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_368),
.B(n_372),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_369),
.A2(n_371),
.B1(n_348),
.B2(n_367),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_344),
.A2(n_320),
.B1(n_330),
.B2(n_340),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g373 ( 
.A(n_345),
.B(n_326),
.C(n_325),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_373),
.B(n_376),
.C(n_378),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_349),
.B(n_296),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g389 ( 
.A(n_374),
.B(n_381),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_345),
.B(n_316),
.C(n_296),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_359),
.B(n_353),
.C(n_356),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g399 ( 
.A(n_379),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_347),
.B(n_291),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g400 ( 
.A1(n_383),
.A2(n_352),
.B1(n_354),
.B2(n_360),
.Y(n_400)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_384),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_SL g387 ( 
.A(n_353),
.B(n_332),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_387),
.B(n_364),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_350),
.B(n_332),
.C(n_281),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_388),
.B(n_346),
.C(n_358),
.Y(n_402)
);

A2O1A1Ixp33_ASAP7_75t_SL g391 ( 
.A1(n_371),
.A2(n_363),
.B(n_357),
.C(n_367),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_391),
.A2(n_370),
.B1(n_383),
.B2(n_386),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g419 ( 
.A1(n_392),
.A2(n_393),
.B1(n_404),
.B2(n_3),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_377),
.A2(n_352),
.B1(n_342),
.B2(n_362),
.Y(n_393)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_394),
.B(n_398),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_372),
.B(n_357),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_395),
.B(n_396),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_388),
.B(n_350),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_378),
.B(n_355),
.C(n_354),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_400),
.B(n_3),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g414 ( 
.A(n_402),
.B(n_2),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_376),
.B(n_218),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_403),
.B(n_405),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_380),
.A2(n_281),
.B1(n_266),
.B2(n_214),
.Y(n_404)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_382),
.Y(n_405)
);

AO32x1_ASAP7_75t_L g407 ( 
.A1(n_391),
.A2(n_370),
.A3(n_383),
.B1(n_379),
.B2(n_368),
.Y(n_407)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_407),
.B(n_408),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g408 ( 
.A(n_401),
.B(n_373),
.C(n_385),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_399),
.A2(n_380),
.B1(n_369),
.B2(n_375),
.Y(n_410)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_410),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_397),
.B(n_375),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g425 ( 
.A(n_411),
.B(n_395),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_412),
.B(n_414),
.Y(n_427)
);

FAx1_ASAP7_75t_SL g413 ( 
.A(n_391),
.B(n_386),
.CI(n_214),
.CON(n_413),
.SN(n_413)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_413),
.B(n_418),
.Y(n_421)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_415),
.Y(n_428)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_389),
.Y(n_416)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_416),
.Y(n_430)
);

INVxp33_ASAP7_75t_L g418 ( 
.A(n_402),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_4),
.Y(n_429)
);

BUFx24_ASAP7_75t_SL g422 ( 
.A(n_409),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_431),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_408),
.B(n_401),
.C(n_396),
.Y(n_423)
);

OR2x2_ASAP7_75t_L g439 ( 
.A(n_423),
.B(n_425),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g426 ( 
.A1(n_418),
.A2(n_390),
.B(n_391),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g432 ( 
.A(n_426),
.B(n_413),
.Y(n_432)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g431 ( 
.A(n_406),
.B(n_4),
.C(n_5),
.Y(n_431)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_432),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_420),
.B(n_406),
.C(n_414),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g445 ( 
.A(n_433),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_430),
.B(n_417),
.Y(n_434)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_434),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_427),
.B(n_412),
.Y(n_436)
);

INVxp33_ASAP7_75t_L g443 ( 
.A(n_436),
.Y(n_443)
);

AOI22xp5_ASAP7_75t_SL g437 ( 
.A1(n_424),
.A2(n_407),
.B1(n_415),
.B2(n_413),
.Y(n_437)
);

INVxp67_ASAP7_75t_L g442 ( 
.A(n_437),
.Y(n_442)
);

AOI21xp5_ASAP7_75t_L g438 ( 
.A1(n_427),
.A2(n_10),
.B(n_7),
.Y(n_438)
);

NOR2xp67_ASAP7_75t_L g441 ( 
.A(n_438),
.B(n_428),
.Y(n_441)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_441),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_445),
.B(n_439),
.C(n_434),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_448),
.B(n_449),
.C(n_443),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_446),
.A2(n_421),
.B1(n_432),
.B2(n_440),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_442),
.A2(n_421),
.B(n_435),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_450),
.A2(n_444),
.B(n_7),
.Y(n_452)
);

NAND3xp33_ASAP7_75t_L g453 ( 
.A(n_451),
.B(n_452),
.C(n_447),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_453),
.B(n_7),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_SL g455 ( 
.A(n_454),
.B(n_9),
.Y(n_455)
);


endmodule