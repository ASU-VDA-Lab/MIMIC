module fake_jpeg_18244_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx16f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx6_ASAP7_75t_SL g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx16_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_26),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g37 ( 
.A(n_20),
.B(n_0),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_26),
.B(n_0),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_39),
.B(n_40),
.Y(n_52)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_15),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_25),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_28),
.B1(n_20),
.B2(n_15),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_19),
.B1(n_44),
.B2(n_23),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_28),
.B1(n_33),
.B2(n_39),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_45),
.A2(n_49),
.B1(n_24),
.B2(n_16),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_46),
.B(n_32),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_36),
.A2(n_19),
.B1(n_22),
.B2(n_29),
.Y(n_49)
);

NOR2x1_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_40),
.Y(n_51)
);

O2A1O1Ixp33_ASAP7_75t_L g71 ( 
.A1(n_51),
.A2(n_24),
.B(n_27),
.C(n_23),
.Y(n_71)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_53),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_55),
.B(n_38),
.Y(n_58)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_66),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g77 ( 
.A1(n_59),
.A2(n_53),
.B(n_55),
.Y(n_77)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_56),
.Y(n_61)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_61),
.Y(n_79)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_62),
.Y(n_84)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_67),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g68 ( 
.A(n_49),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_52),
.B(n_31),
.C(n_35),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_76),
.C(n_50),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_52),
.A2(n_19),
.B1(n_29),
.B2(n_21),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_72),
.B1(n_73),
.B2(n_42),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_71),
.B(n_51),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_27),
.B1(n_31),
.B2(n_16),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_34),
.B1(n_16),
.B2(n_26),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_74),
.A2(n_75),
.B1(n_54),
.B2(n_50),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_47),
.A2(n_34),
.B1(n_35),
.B2(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_34),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_77),
.A2(n_76),
.B1(n_72),
.B2(n_63),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_35),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_78),
.A2(n_88),
.B(n_46),
.Y(n_113)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_58),
.B(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_94),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_91),
.B(n_46),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_92),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_93),
.A2(n_95),
.B1(n_74),
.B2(n_67),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_71),
.B(n_51),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_26),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_93),
.C(n_54),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_104),
.B1(n_100),
.B2(n_101),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_106),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_79),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_103),
.B(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_92),
.A2(n_42),
.B1(n_65),
.B2(n_54),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_105),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_83),
.B(n_84),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_80),
.B(n_16),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_108),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_81),
.Y(n_109)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_110),
.B(n_97),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_86),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_112),
.B(n_91),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g117 ( 
.A1(n_113),
.A2(n_82),
.B(n_88),
.C(n_78),
.D(n_86),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_114),
.B(n_118),
.Y(n_130)
);

OAI32xp33_ASAP7_75t_L g115 ( 
.A1(n_98),
.A2(n_77),
.A3(n_80),
.B1(n_89),
.B2(n_88),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_117),
.B(n_125),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_78),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_120),
.B(n_103),
.Y(n_138)
);

AOI322xp5_ASAP7_75t_SL g121 ( 
.A1(n_106),
.A2(n_82),
.A3(n_14),
.B1(n_13),
.B2(n_12),
.C1(n_11),
.C2(n_8),
.Y(n_121)
);

AOI322xp5_ASAP7_75t_SL g134 ( 
.A1(n_121),
.A2(n_10),
.A3(n_13),
.B1(n_9),
.B2(n_8),
.C1(n_6),
.C2(n_5),
.Y(n_134)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_122),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_99),
.C(n_107),
.Y(n_137)
);

INVx2_ASAP7_75t_SL g129 ( 
.A(n_120),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_127),
.B1(n_90),
.B2(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_126),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_133),
.B(n_134),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_123),
.A2(n_113),
.B1(n_100),
.B2(n_112),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_117),
.B(n_128),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_136),
.B(n_138),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_137),
.B(n_139),
.C(n_132),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_115),
.B(n_108),
.C(n_105),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_127),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_140),
.B(n_116),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_130),
.B(n_114),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_129),
.B1(n_131),
.B2(n_104),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_144),
.B(n_145),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_149),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_128),
.B(n_125),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_147),
.A2(n_135),
.B(n_137),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_119),
.C(n_110),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_151),
.A2(n_146),
.B1(n_149),
.B2(n_124),
.Y(n_157)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_148),
.B(n_131),
.C(n_129),
.Y(n_152)
);

AO21x1_ASAP7_75t_L g162 ( 
.A1(n_152),
.A2(n_18),
.B(n_2),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_153),
.B(n_156),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_124),
.B1(n_85),
.B2(n_65),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_157),
.B(n_161),
.C(n_1),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_154),
.B(n_17),
.C(n_46),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_160),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_150),
.B(n_10),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_152),
.A2(n_18),
.B1(n_17),
.B2(n_3),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_155),
.B(n_5),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_1),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_165),
.B(n_6),
.Y(n_169)
);

NOR2xp67_ASAP7_75t_SL g166 ( 
.A(n_158),
.B(n_1),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_166),
.A2(n_162),
.B(n_159),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_168),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_170),
.B(n_164),
.C(n_169),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_172),
.B(n_171),
.Y(n_173)
);


endmodule