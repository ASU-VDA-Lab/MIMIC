module fake_jpeg_26462_n_103 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_103);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_103;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_L g14 ( 
.A(n_4),
.B(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_3),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_24),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_0),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_12),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_25),
.B(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_14),
.B(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_16),
.Y(n_27)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_5),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_16),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_30),
.Y(n_31)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_24),
.B(n_21),
.Y(n_35)
);

AO21x1_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_36),
.B(n_38),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_30),
.Y(n_36)
);

NOR2x1_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_15),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_13),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_39),
.B(n_30),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_22),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_40),
.Y(n_48)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_39),
.Y(n_41)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_32),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_42),
.B(n_49),
.Y(n_55)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx2_ASAP7_75t_SL g44 ( 
.A(n_33),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_13),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_SL g58 ( 
.A(n_45),
.B(n_46),
.C(n_52),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_31),
.A2(n_12),
.B1(n_23),
.B2(n_16),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_43),
.B1(n_51),
.B2(n_48),
.Y(n_54)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_19),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_21),
.Y(n_62)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_52),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_12),
.B1(n_36),
.B2(n_35),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_53),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_54),
.A2(n_58),
.B(n_48),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_36),
.B1(n_35),
.B2(n_17),
.Y(n_59)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_59),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_21),
.B1(n_13),
.B2(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_65),
.B(n_66),
.Y(n_74)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_59),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_49),
.C(n_47),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_70),
.B(n_71),
.C(n_19),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_63),
.B(n_21),
.C(n_17),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_72),
.B(n_73),
.Y(n_81)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g88 ( 
.A(n_75),
.B(n_3),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_70),
.B(n_55),
.C(n_58),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_76),
.B(n_13),
.C(n_56),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_60),
.B1(n_11),
.B2(n_18),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_20),
.B1(n_22),
.B2(n_11),
.Y(n_85)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_71),
.Y(n_78)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_78),
.Y(n_83)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_64),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_69),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_80),
.A2(n_67),
.B1(n_60),
.B2(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_82),
.B(n_85),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_87),
.C(n_79),
.Y(n_90)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_86),
.B(n_88),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_87),
.C(n_9),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_83),
.A2(n_80),
.B(n_74),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_91),
.B(n_8),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_88),
.B(n_6),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_10),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_96),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_95),
.Y(n_100)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_89),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_97),
.A2(n_92),
.B(n_8),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_99),
.B(n_9),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_101),
.B(n_102),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_100),
.Y(n_102)
);


endmodule