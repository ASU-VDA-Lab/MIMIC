module fake_jpeg_12852_n_58 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_58);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_58;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx3_ASAP7_75t_L g8 ( 
.A(n_2),
.Y(n_8)
);

INVx6_ASAP7_75t_SL g9 ( 
.A(n_3),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

HB1xp67_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_5),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_0),
.Y(n_14)
);

INVx5_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx6_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_23),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_13),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_21),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx13_ASAP7_75t_L g32 ( 
.A(n_22),
.Y(n_32)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_1),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_24),
.B(n_20),
.Y(n_28)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_17),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_28),
.B(n_29),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_12),
.C(n_8),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g33 ( 
.A1(n_19),
.A2(n_17),
.B1(n_16),
.B2(n_15),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_21),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_27),
.Y(n_42)
);

CKINVDCx6p67_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_31),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_29),
.A2(n_25),
.B1(n_18),
.B2(n_23),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_26),
.B1(n_30),
.B2(n_25),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_R g46 ( 
.A(n_41),
.B(n_42),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_39),
.B(n_27),
.C(n_26),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_38),
.C(n_36),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_26),
.B1(n_30),
.B2(n_15),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_47)
);

OAI21x1_ASAP7_75t_L g50 ( 
.A1(n_47),
.A2(n_48),
.B(n_35),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_49),
.Y(n_51)
);

AO21x1_ASAP7_75t_L g54 ( 
.A1(n_50),
.A2(n_35),
.B(n_32),
.Y(n_54)
);

AOI322xp5_ASAP7_75t_L g53 ( 
.A1(n_51),
.A2(n_46),
.A3(n_48),
.B1(n_11),
.B2(n_16),
.C1(n_45),
.C2(n_9),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_53),
.A2(n_54),
.B(n_52),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_55),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_6),
.Y(n_56)
);

OAI321xp33_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_56),
.A3(n_6),
.B1(n_7),
.B2(n_11),
.C(n_1),
.Y(n_58)
);


endmodule