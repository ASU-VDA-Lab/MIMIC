module fake_jpeg_366_n_583 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_583);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_583;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_7),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_16),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_15),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_17),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx13_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_14),
.B(n_11),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_4),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_4),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_13),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_12),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_26),
.Y(n_57)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_57),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_19),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_58),
.B(n_61),
.Y(n_136)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_26),
.Y(n_59)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_59),
.Y(n_151)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_60),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_42),
.B(n_17),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_19),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_62),
.B(n_65),
.Y(n_165)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_63),
.Y(n_156)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_28),
.Y(n_64)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_64),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_20),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_66),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_28),
.B(n_56),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_67),
.B(n_68),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_11),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_24),
.B(n_11),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_69),
.B(n_70),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_20),
.Y(n_70)
);

BUFx12_ASAP7_75t_L g71 ( 
.A(n_36),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g180 ( 
.A(n_71),
.Y(n_180)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

INVx8_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_40),
.B(n_16),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_73),
.B(n_75),
.Y(n_176)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_27),
.Y(n_74)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_20),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_76),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g77 ( 
.A(n_35),
.Y(n_77)
);

BUFx2_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_79),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g146 ( 
.A(n_80),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_21),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_81),
.Y(n_158)
);

HB1xp67_ASAP7_75t_L g82 ( 
.A(n_23),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g154 ( 
.A(n_82),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_21),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g168 ( 
.A(n_83),
.Y(n_168)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_84),
.Y(n_134)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_85),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_86),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_27),
.Y(n_87)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_87),
.Y(n_127)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_88),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_33),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_89),
.Y(n_185)
);

INVx6_ASAP7_75t_L g90 ( 
.A(n_35),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_90),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_44),
.B(n_16),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_91),
.B(n_101),
.Y(n_199)
);

BUFx5_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

BUFx24_ASAP7_75t_L g126 ( 
.A(n_92),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_33),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_33),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_94),
.Y(n_133)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_27),
.Y(n_95)
);

INVx11_ASAP7_75t_L g179 ( 
.A(n_95),
.Y(n_179)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_56),
.Y(n_96)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_96),
.Y(n_164)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_27),
.Y(n_97)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_98),
.Y(n_167)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_25),
.Y(n_99)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_99),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_100),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_40),
.B(n_0),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_102),
.Y(n_141)
);

INVx4_ASAP7_75t_SL g103 ( 
.A(n_34),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g155 ( 
.A(n_103),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_54),
.B(n_0),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_104),
.B(n_106),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_55),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_105),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_55),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_30),
.Y(n_107)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_107),
.Y(n_143)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_34),
.Y(n_108)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_108),
.Y(n_153)
);

INVx4_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_109),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_55),
.Y(n_110)
);

INVx6_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_36),
.Y(n_111)
);

INVx6_ASAP7_75t_SL g147 ( 
.A(n_111),
.Y(n_147)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_34),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_34),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_113),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_51),
.B(n_1),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_114),
.B(n_119),
.Y(n_207)
);

BUFx12f_ASAP7_75t_L g115 ( 
.A(n_36),
.Y(n_115)
);

INVx8_ASAP7_75t_L g132 ( 
.A(n_115),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g116 ( 
.A(n_50),
.Y(n_116)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_116),
.Y(n_149)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx6_ASAP7_75t_L g145 ( 
.A(n_117),
.Y(n_145)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_54),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_25),
.Y(n_120)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_18),
.B(n_1),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_121),
.B(n_2),
.Y(n_208)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_122),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_18),
.B(n_9),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_123),
.B(n_22),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_51),
.Y(n_124)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_124),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_38),
.B1(n_52),
.B2(n_46),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_SL g240 ( 
.A1(n_142),
.A2(n_184),
.B1(n_29),
.B2(n_95),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_114),
.B(n_22),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g282 ( 
.A(n_148),
.B(n_192),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_157),
.B(n_190),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_90),
.Y(n_159)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_159),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g161 ( 
.A1(n_66),
.A2(n_39),
.B1(n_52),
.B2(n_46),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_161),
.A2(n_49),
.B1(n_47),
.B2(n_32),
.Y(n_220)
);

INVx6_ASAP7_75t_SL g162 ( 
.A(n_71),
.Y(n_162)
);

BUFx4f_ASAP7_75t_SL g272 ( 
.A(n_162),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_117),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_163),
.B(n_166),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_124),
.Y(n_166)
);

INVx3_ASAP7_75t_SL g169 ( 
.A(n_113),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g233 ( 
.A(n_169),
.Y(n_233)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_120),
.Y(n_177)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_177),
.Y(n_225)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_87),
.Y(n_178)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_178),
.Y(n_239)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_77),
.Y(n_181)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_181),
.Y(n_242)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_115),
.Y(n_182)
);

INVx4_ASAP7_75t_L g247 ( 
.A(n_182),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_SL g184 ( 
.A1(n_116),
.A2(n_38),
.B1(n_45),
.B2(n_43),
.Y(n_184)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_115),
.Y(n_187)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_187),
.Y(n_218)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_78),
.Y(n_189)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_189),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_102),
.B(n_53),
.Y(n_190)
);

BUFx12f_ASAP7_75t_L g191 ( 
.A(n_71),
.Y(n_191)
);

INVx11_ASAP7_75t_L g260 ( 
.A(n_191),
.Y(n_260)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_108),
.B(n_37),
.Y(n_192)
);

INVx3_ASAP7_75t_L g193 ( 
.A(n_84),
.Y(n_193)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_193),
.Y(n_219)
);

BUFx12f_ASAP7_75t_L g195 ( 
.A(n_97),
.Y(n_195)
);

INVx11_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_122),
.Y(n_196)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_196),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_80),
.B(n_37),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_208),
.Y(n_231)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_88),
.Y(n_201)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_201),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_60),
.B(n_39),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_202),
.B(n_72),
.Y(n_228)
);

BUFx5_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_205),
.Y(n_234)
);

BUFx12f_ASAP7_75t_L g209 ( 
.A(n_81),
.Y(n_209)
);

INVx11_ASAP7_75t_L g275 ( 
.A(n_209),
.Y(n_275)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_83),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_210),
.Y(n_223)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_92),
.Y(n_211)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_211),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_148),
.A2(n_107),
.B1(n_109),
.B2(n_43),
.Y(n_213)
);

OR2x2_ASAP7_75t_L g311 ( 
.A(n_213),
.B(n_215),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_190),
.A2(n_202),
.B1(n_207),
.B2(n_165),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_207),
.A2(n_41),
.B(n_53),
.Y(n_217)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_217),
.B(n_228),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_220),
.A2(n_245),
.B1(n_236),
.B2(n_267),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_154),
.A2(n_49),
.B1(n_47),
.B2(n_32),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g304 ( 
.A1(n_221),
.A2(n_267),
.B1(n_158),
.B2(n_168),
.Y(n_304)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_132),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g315 ( 
.A(n_224),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_165),
.B(n_45),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_226),
.B(n_229),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_154),
.B(n_72),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g331 ( 
.A(n_227),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_136),
.B(n_171),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_206),
.B(n_174),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_230),
.B(n_243),
.Y(n_328)
);

INVx6_ASAP7_75t_L g235 ( 
.A(n_144),
.Y(n_235)
);

INVx3_ASAP7_75t_SL g289 ( 
.A(n_235),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_169),
.B(n_41),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g336 ( 
.A(n_236),
.B(n_278),
.Y(n_336)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_155),
.Y(n_237)
);

INVxp67_ASAP7_75t_SL g306 ( 
.A(n_237),
.Y(n_306)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_129),
.Y(n_238)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_238),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_240),
.Y(n_327)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_135),
.Y(n_241)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_29),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_136),
.B(n_171),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_244),
.B(n_250),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_L g245 ( 
.A1(n_142),
.A2(n_86),
.B1(n_110),
.B2(n_105),
.Y(n_245)
);

INVx13_ASAP7_75t_L g246 ( 
.A(n_147),
.Y(n_246)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_246),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_144),
.Y(n_248)
);

INVx8_ASAP7_75t_L g303 ( 
.A(n_248),
.Y(n_303)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_161),
.A2(n_100),
.B1(n_94),
.B2(n_93),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_249),
.A2(n_284),
.B1(n_172),
.B2(n_185),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_203),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_175),
.A2(n_112),
.B1(n_74),
.B2(n_89),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g300 ( 
.A1(n_251),
.A2(n_254),
.B1(n_266),
.B2(n_280),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_174),
.B(n_2),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_252),
.B(n_258),
.Y(n_291)
);

AOI22xp33_ASAP7_75t_SL g254 ( 
.A1(n_134),
.A2(n_50),
.B1(n_3),
.B2(n_4),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_199),
.B(n_2),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_255),
.B(n_257),
.Y(n_297)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_150),
.Y(n_256)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_256),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_152),
.B(n_3),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_176),
.B(n_5),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_164),
.B(n_5),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_259),
.B(n_262),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_146),
.Y(n_261)
);

INVx3_ASAP7_75t_L g318 ( 
.A(n_261),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_176),
.B(n_5),
.Y(n_262)
);

INVx8_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_263),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_146),
.Y(n_265)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_265),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_143),
.A2(n_50),
.B1(n_7),
.B2(n_8),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_128),
.A2(n_151),
.B1(n_156),
.B2(n_167),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_188),
.Y(n_268)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_268),
.Y(n_295)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_127),
.Y(n_269)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_269),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_199),
.B(n_7),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_270),
.B(n_273),
.Y(n_330)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_203),
.Y(n_271)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_271),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_208),
.B(n_8),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_130),
.Y(n_274)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_274),
.Y(n_319)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_141),
.Y(n_276)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_194),
.B(n_8),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_138),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_279),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g280 ( 
.A1(n_160),
.A2(n_173),
.B1(n_153),
.B2(n_138),
.Y(n_280)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_149),
.A2(n_139),
.B1(n_200),
.B2(n_179),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g302 ( 
.A1(n_281),
.A2(n_180),
.B1(n_191),
.B2(n_125),
.Y(n_302)
);

OAI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_184),
.A2(n_204),
.B1(n_183),
.B2(n_140),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_145),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_285),
.B(n_233),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_288),
.B(n_304),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_215),
.A2(n_204),
.B1(n_137),
.B2(n_133),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_292),
.B(n_261),
.Y(n_348)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_282),
.A2(n_212),
.B1(n_185),
.B2(n_172),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_294),
.B(n_232),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_220),
.A2(n_212),
.B1(n_168),
.B2(n_158),
.Y(n_296)
);

INVxp67_ASAP7_75t_SL g344 ( 
.A(n_296),
.Y(n_344)
);

MAJx2_ASAP7_75t_L g301 ( 
.A(n_214),
.B(n_170),
.C(n_126),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_314),
.C(n_323),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_302),
.Y(n_342)
);

AOI32xp33_ASAP7_75t_L g305 ( 
.A1(n_230),
.A2(n_126),
.A3(n_198),
.B1(n_186),
.B2(n_180),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_305),
.B(n_272),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_231),
.A2(n_131),
.B1(n_195),
.B2(n_282),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_308),
.B(n_309),
.Y(n_379)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_235),
.Y(n_310)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_310),
.Y(n_346)
);

OA22x2_ASAP7_75t_L g312 ( 
.A1(n_213),
.A2(n_245),
.B1(n_232),
.B2(n_225),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_312),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_228),
.B(n_270),
.Y(n_314)
);

OAI22x1_ASAP7_75t_L g316 ( 
.A1(n_278),
.A2(n_252),
.B1(n_258),
.B2(n_273),
.Y(n_316)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_316),
.Y(n_341)
);

INVx2_ASAP7_75t_SL g317 ( 
.A(n_236),
.Y(n_317)
);

BUFx2_ASAP7_75t_L g350 ( 
.A(n_317),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_217),
.A2(n_278),
.B1(n_243),
.B2(n_227),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_320),
.A2(n_333),
.B1(n_253),
.B2(n_237),
.Y(n_351)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_223),
.Y(n_322)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_322),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_216),
.B(n_227),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_223),
.Y(n_324)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_324),
.Y(n_373)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_222),
.Y(n_326)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_326),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_225),
.B(n_239),
.C(n_277),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g377 ( 
.A(n_332),
.B(n_260),
.Y(n_377)
);

AOI22xp33_ASAP7_75t_L g333 ( 
.A1(n_253),
.A2(n_219),
.B1(n_239),
.B2(n_242),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_337),
.Y(n_376)
);

INVx2_ASAP7_75t_L g339 ( 
.A(n_219),
.Y(n_339)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_242),
.Y(n_340)
);

NAND2xp5_ASAP7_75t_SL g353 ( 
.A(n_340),
.B(n_283),
.Y(n_353)
);

INVxp67_ASAP7_75t_L g387 ( 
.A(n_343),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_345),
.A2(n_348),
.B1(n_381),
.B2(n_295),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_307),
.B(n_272),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_359),
.Y(n_385)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_322),
.Y(n_349)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_349),
.Y(n_400)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_351),
.Y(n_410)
);

INVx4_ASAP7_75t_L g352 ( 
.A(n_303),
.Y(n_352)
);

BUFx4f_ASAP7_75t_L g399 ( 
.A(n_352),
.Y(n_399)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_353),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_309),
.A2(n_265),
.B1(n_248),
.B2(n_283),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_355),
.A2(n_369),
.B1(n_327),
.B2(n_292),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_SL g356 ( 
.A(n_314),
.B(n_277),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g384 ( 
.A(n_356),
.B(n_368),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_291),
.B(n_272),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_357),
.B(n_358),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_328),
.B(n_247),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_307),
.B(n_247),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_334),
.B(n_218),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_362),
.Y(n_396)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_306),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_361),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g362 ( 
.A(n_334),
.B(n_218),
.Y(n_362)
);

AND2x6_ASAP7_75t_L g363 ( 
.A(n_311),
.B(n_246),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_363),
.B(n_364),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_321),
.B(n_224),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_334),
.B(n_234),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_365),
.B(n_378),
.Y(n_401)
);

INVx13_ASAP7_75t_L g367 ( 
.A(n_335),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g391 ( 
.A(n_367),
.Y(n_391)
);

AND2x2_ASAP7_75t_SL g368 ( 
.A(n_317),
.B(n_264),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_311),
.A2(n_263),
.B1(n_234),
.B2(n_275),
.Y(n_369)
);

BUFx5_ASAP7_75t_L g370 ( 
.A(n_339),
.Y(n_370)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_370),
.Y(n_390)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_264),
.Y(n_371)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_371),
.Y(n_415)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_329),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_372),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g406 ( 
.A(n_377),
.B(n_332),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_286),
.B(n_260),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_287),
.B(n_275),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_356),
.B(n_323),
.C(n_301),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_383),
.B(n_386),
.C(n_397),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_374),
.B(n_331),
.C(n_336),
.Y(n_386)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_392),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_375),
.A2(n_288),
.B1(n_327),
.B2(n_320),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_393),
.A2(n_398),
.B1(n_402),
.B2(n_404),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_375),
.A2(n_300),
.B(n_312),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g417 ( 
.A1(n_394),
.A2(n_342),
.B(n_366),
.Y(n_417)
);

OA22x2_ASAP7_75t_L g395 ( 
.A1(n_341),
.A2(n_312),
.B1(n_337),
.B2(n_318),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_395),
.B(n_411),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_374),
.B(n_336),
.C(n_290),
.Y(n_397)
);

OAI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_341),
.A2(n_312),
.B1(n_330),
.B2(n_291),
.Y(n_398)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_379),
.A2(n_316),
.B1(n_336),
.B2(n_330),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_379),
.A2(n_313),
.B1(n_297),
.B2(n_289),
.Y(n_404)
);

OA21x2_ASAP7_75t_L g405 ( 
.A1(n_379),
.A2(n_299),
.B(n_325),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_SL g435 ( 
.A1(n_405),
.A2(n_413),
.B(n_414),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g418 ( 
.A(n_406),
.B(n_362),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_408),
.A2(n_345),
.B1(n_348),
.B2(n_344),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_376),
.A2(n_289),
.B1(n_324),
.B2(n_310),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_377),
.B(n_319),
.C(n_298),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_412),
.B(n_368),
.C(n_369),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_376),
.A2(n_315),
.B(n_329),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_L g414 ( 
.A1(n_360),
.A2(n_315),
.B(n_293),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_366),
.A2(n_318),
.B1(n_293),
.B2(n_303),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_416),
.B(n_366),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_SL g463 ( 
.A1(n_417),
.A2(n_427),
.B(n_443),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_418),
.B(n_420),
.C(n_444),
.Y(n_453)
);

INVx13_ASAP7_75t_L g419 ( 
.A(n_407),
.Y(n_419)
);

AOI22xp33_ASAP7_75t_SL g472 ( 
.A1(n_419),
.A2(n_399),
.B1(n_352),
.B2(n_416),
.Y(n_472)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_357),
.Y(n_420)
);

INVxp67_ASAP7_75t_L g421 ( 
.A(n_385),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_421),
.B(n_433),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_391),
.B(n_380),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_422),
.B(n_428),
.Y(n_456)
);

NOR2x1_ASAP7_75t_L g423 ( 
.A(n_402),
.B(n_363),
.Y(n_423)
);

A2O1A1Ixp33_ASAP7_75t_L g455 ( 
.A1(n_423),
.A2(n_387),
.B(n_386),
.C(n_393),
.Y(n_455)
);

INVx6_ASAP7_75t_SL g426 ( 
.A(n_398),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_426),
.Y(n_459)
);

OAI21xp5_ASAP7_75t_L g427 ( 
.A1(n_396),
.A2(n_365),
.B(n_350),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g428 ( 
.A(n_415),
.B(n_358),
.Y(n_428)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_389),
.B(n_380),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_429),
.B(n_434),
.Y(n_449)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_411),
.Y(n_430)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_430),
.Y(n_450)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_400),
.Y(n_431)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_431),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_413),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g434 ( 
.A(n_401),
.B(n_382),
.Y(n_434)
);

BUFx12_ASAP7_75t_L g436 ( 
.A(n_399),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g476 ( 
.A(n_436),
.Y(n_476)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_400),
.Y(n_437)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_437),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_401),
.B(n_404),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g461 ( 
.A(n_438),
.B(n_388),
.Y(n_461)
);

AND2x6_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_367),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_439),
.B(n_441),
.Y(n_467)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_440),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_388),
.B(n_350),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g443 ( 
.A1(n_396),
.A2(n_350),
.B(n_342),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_405),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_410),
.Y(n_475)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_446),
.Y(n_465)
);

INVx3_ASAP7_75t_L g447 ( 
.A(n_390),
.Y(n_447)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_447),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_418),
.B(n_384),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g492 ( 
.A(n_448),
.B(n_435),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_420),
.B(n_397),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g478 ( 
.A(n_454),
.B(n_469),
.Y(n_478)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_455),
.A2(n_458),
.B(n_462),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_425),
.B(n_406),
.C(n_412),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_457),
.B(n_466),
.C(n_453),
.Y(n_483)
);

AO21x1_ASAP7_75t_L g458 ( 
.A1(n_432),
.A2(n_387),
.B(n_394),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_SL g499 ( 
.A1(n_458),
.A2(n_473),
.B(n_439),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g479 ( 
.A1(n_461),
.A2(n_472),
.B1(n_392),
.B2(n_442),
.Y(n_479)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_428),
.B(n_403),
.Y(n_464)
);

CKINVDCx14_ASAP7_75t_R g497 ( 
.A(n_464),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_425),
.B(n_384),
.C(n_405),
.Y(n_466)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_432),
.B(n_395),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g470 ( 
.A(n_421),
.B(n_382),
.Y(n_470)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_470),
.Y(n_477)
);

NAND2xp67_ASAP7_75t_L g471 ( 
.A(n_426),
.B(n_395),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_471),
.B(n_442),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_417),
.A2(n_414),
.B(n_395),
.Y(n_473)
);

AO22x2_ASAP7_75t_L g474 ( 
.A1(n_424),
.A2(n_410),
.B1(n_355),
.B2(n_351),
.Y(n_474)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_474),
.Y(n_480)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_475),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_L g507 ( 
.A1(n_479),
.A2(n_484),
.B1(n_465),
.B2(n_460),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_454),
.B(n_423),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_483),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_456),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_482),
.B(n_467),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_467),
.A2(n_424),
.B1(n_445),
.B2(n_430),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_456),
.Y(n_485)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_485),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_486),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_453),
.B(n_444),
.C(n_427),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g517 ( 
.A(n_487),
.B(n_489),
.C(n_495),
.Y(n_517)
);

XOR2x2_ASAP7_75t_L g488 ( 
.A(n_466),
.B(n_423),
.Y(n_488)
);

NOR2xp33_ASAP7_75t_L g519 ( 
.A(n_488),
.B(n_498),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_457),
.B(n_433),
.C(n_441),
.Y(n_489)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_455),
.B(n_443),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_490),
.B(n_492),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_435),
.Y(n_491)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_491),
.Y(n_514)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_451),
.Y(n_493)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_493),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_448),
.B(n_437),
.C(n_431),
.Y(n_495)
);

XOR2x2_ASAP7_75t_L g513 ( 
.A(n_496),
.B(n_500),
.Y(n_513)
);

XNOR2xp5_ASAP7_75t_SL g498 ( 
.A(n_469),
.B(n_440),
.Y(n_498)
);

AOI21xp5_ASAP7_75t_L g509 ( 
.A1(n_499),
.A2(n_501),
.B(n_463),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_460),
.B(n_368),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_SL g501 ( 
.A1(n_473),
.A2(n_447),
.B(n_419),
.Y(n_501)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_494),
.Y(n_505)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_505),
.Y(n_521)
);

AOI22xp5_ASAP7_75t_L g527 ( 
.A1(n_507),
.A2(n_489),
.B1(n_478),
.B2(n_500),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_L g508 ( 
.A1(n_491),
.A2(n_463),
.B(n_459),
.Y(n_508)
);

OAI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_508),
.A2(n_509),
.B(n_515),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_494),
.B(n_449),
.Y(n_510)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_510),
.Y(n_526)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_511),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_L g515 ( 
.A1(n_496),
.A2(n_459),
.B(n_465),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_486),
.Y(n_516)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_516),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_477),
.B(n_450),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_518),
.B(n_452),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_497),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_520),
.B(n_495),
.Y(n_528)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_508),
.A2(n_499),
.B(n_501),
.Y(n_522)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_522),
.Y(n_544)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_509),
.A2(n_490),
.B(n_480),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_524),
.B(n_514),
.Y(n_536)
);

AOI22xp33_ASAP7_75t_SL g525 ( 
.A1(n_505),
.A2(n_480),
.B1(n_450),
.B2(n_451),
.Y(n_525)
);

OAI22xp5_ASAP7_75t_SL g545 ( 
.A1(n_525),
.A2(n_527),
.B1(n_503),
.B2(n_504),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_528),
.B(n_531),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_506),
.B(n_478),
.Y(n_530)
);

XOR2xp5_ASAP7_75t_L g541 ( 
.A(n_530),
.B(n_534),
.Y(n_541)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_483),
.C(n_487),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_532),
.B(n_535),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g534 ( 
.A(n_506),
.B(n_481),
.Y(n_534)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_517),
.B(n_488),
.C(n_498),
.Y(n_535)
);

MAJx2_ASAP7_75t_L g553 ( 
.A(n_536),
.B(n_492),
.C(n_471),
.Y(n_553)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_532),
.B(n_510),
.C(n_502),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_538),
.B(n_539),
.Y(n_555)
);

NOR2xp33_ASAP7_75t_SL g539 ( 
.A(n_533),
.B(n_518),
.Y(n_539)
);

AOI22xp33_ASAP7_75t_SL g540 ( 
.A1(n_529),
.A2(n_516),
.B1(n_503),
.B2(n_515),
.Y(n_540)
);

OAI21xp5_ASAP7_75t_SL g551 ( 
.A1(n_540),
.A2(n_523),
.B(n_524),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g542 ( 
.A(n_530),
.B(n_513),
.C(n_512),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_542),
.B(n_546),
.Y(n_557)
);

XOR2xp5_ASAP7_75t_L g543 ( 
.A(n_534),
.B(n_513),
.Y(n_543)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_543),
.B(n_547),
.C(n_468),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_545),
.B(n_452),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_526),
.B(n_468),
.Y(n_546)
);

XOR2xp5_ASAP7_75t_L g547 ( 
.A(n_527),
.B(n_512),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_SL g549 ( 
.A1(n_544),
.A2(n_523),
.B(n_535),
.Y(n_549)
);

OAI22xp5_ASAP7_75t_L g561 ( 
.A1(n_549),
.A2(n_550),
.B1(n_552),
.B2(n_540),
.Y(n_561)
);

AOI31xp67_ASAP7_75t_L g550 ( 
.A1(n_542),
.A2(n_522),
.A3(n_529),
.B(n_521),
.Y(n_550)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_551),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g552 ( 
.A1(n_548),
.A2(n_519),
.B(n_531),
.Y(n_552)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_553),
.B(n_554),
.Y(n_563)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_537),
.B(n_476),
.C(n_504),
.Y(n_556)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_556),
.B(n_559),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_558),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_536),
.B(n_399),
.Y(n_559)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_561),
.Y(n_571)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_557),
.B(n_555),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g568 ( 
.A(n_562),
.B(n_565),
.Y(n_568)
);

XNOR2xp5_ASAP7_75t_L g564 ( 
.A(n_558),
.B(n_547),
.Y(n_564)
);

XOR2xp5_ASAP7_75t_L g572 ( 
.A(n_564),
.B(n_474),
.Y(n_572)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_553),
.B(n_541),
.Y(n_565)
);

AOI322xp5_ASAP7_75t_L g569 ( 
.A1(n_566),
.A2(n_436),
.A3(n_543),
.B1(n_419),
.B2(n_474),
.C1(n_541),
.C2(n_372),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_569),
.B(n_570),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_560),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_572),
.B(n_573),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_SL g573 ( 
.A1(n_564),
.A2(n_563),
.B(n_567),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_563),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_571),
.Y(n_577)
);

XOR2xp5_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_578),
.Y(n_579)
);

AOI322xp5_ASAP7_75t_L g578 ( 
.A1(n_574),
.A2(n_573),
.A3(n_436),
.B1(n_474),
.B2(n_354),
.C1(n_373),
.C2(n_361),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_L g580 ( 
.A1(n_579),
.A2(n_575),
.B(n_373),
.Y(n_580)
);

AOI221xp5_ASAP7_75t_L g581 ( 
.A1(n_580),
.A2(n_354),
.B1(n_436),
.B2(n_346),
.C(n_474),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_349),
.C(n_346),
.Y(n_582)
);

XOR2xp5_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_370),
.Y(n_583)
);


endmodule