module fake_ariane_3027_n_348 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_34, n_69, n_95, n_92, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_85, n_130, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_112, n_45, n_11, n_129, n_126, n_122, n_52, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_97, n_14, n_88, n_68, n_116, n_104, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_348);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_34;
input n_69;
input n_95;
input n_92;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_85;
input n_130;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_122;
input n_52;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_97;
input n_14;
input n_88;
input n_68;
input n_116;
input n_104;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_348;

wire n_295;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_307;
wire n_332;
wire n_294;
wire n_197;
wire n_176;
wire n_172;
wire n_347;
wire n_183;
wire n_299;
wire n_205;
wire n_341;
wire n_245;
wire n_319;
wire n_283;
wire n_187;
wire n_345;
wire n_318;
wire n_244;
wire n_226;
wire n_261;
wire n_220;
wire n_189;
wire n_286;
wire n_139;
wire n_346;
wire n_214;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_198;
wire n_232;
wire n_327;
wire n_279;
wire n_207;
wire n_140;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_336;
wire n_315;
wire n_311;
wire n_239;
wire n_272;
wire n_339;
wire n_167;
wire n_153;
wire n_269;
wire n_158;
wire n_259;
wire n_143;
wire n_152;
wire n_169;
wire n_173;
wire n_242;
wire n_309;
wire n_320;
wire n_331;
wire n_267;
wire n_335;
wire n_291;
wire n_344;
wire n_210;
wire n_200;
wire n_253;
wire n_166;
wire n_218;
wire n_271;
wire n_247;
wire n_240;
wire n_224;
wire n_222;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_330;
wire n_282;
wire n_328;
wire n_277;
wire n_248;
wire n_301;
wire n_293;
wire n_228;
wire n_325;
wire n_276;
wire n_303;
wire n_168;
wire n_206;
wire n_238;
wire n_136;
wire n_334;
wire n_192;
wire n_300;
wire n_163;
wire n_141;
wire n_314;
wire n_273;
wire n_305;
wire n_312;
wire n_233;
wire n_333;
wire n_221;
wire n_321;
wire n_149;
wire n_237;
wire n_175;
wire n_181;
wire n_260;
wire n_310;
wire n_236;
wire n_281;
wire n_209;
wire n_262;
wire n_225;
wire n_235;
wire n_297;
wire n_290;
wire n_199;
wire n_217;
wire n_178;
wire n_308;
wire n_201;
wire n_343;
wire n_287;
wire n_302;
wire n_284;
wire n_249;
wire n_212;
wire n_278;
wire n_255;
wire n_257;
wire n_148;
wire n_135;
wire n_171;
wire n_182;
wire n_316;
wire n_196;
wire n_254;
wire n_219;
wire n_231;
wire n_234;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_298;
wire n_216;
wire n_223;
wire n_288;
wire n_179;
wire n_195;
wire n_213;
wire n_304;
wire n_306;
wire n_313;
wire n_203;
wire n_150;
wire n_324;
wire n_337;
wire n_274;
wire n_296;
wire n_265;
wire n_208;
wire n_292;
wire n_156;
wire n_174;
wire n_275;
wire n_147;
wire n_204;
wire n_342;
wire n_246;
wire n_159;
wire n_263;
wire n_229;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_243;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_268;
wire n_266;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_258;
wire n_241;
wire n_191;
wire n_211;
wire n_322;
wire n_251;
wire n_155;

INVx1_ASAP7_75t_L g135 ( 
.A(n_25),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g136 ( 
.A(n_42),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_129),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_84),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_93),
.Y(n_139)
);

CKINVDCx5p33_ASAP7_75t_R g140 ( 
.A(n_96),
.Y(n_140)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_89),
.Y(n_141)
);

CKINVDCx5p33_ASAP7_75t_R g142 ( 
.A(n_115),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_14),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_85),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_63),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_R g146 ( 
.A(n_107),
.B(n_60),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_1),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_124),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_99),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_37),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_64),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_113),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_132),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_59),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_0),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_120),
.B(n_118),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_73),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_80),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_81),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

INVx1_ASAP7_75t_SL g161 ( 
.A(n_121),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_45),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_91),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_102),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_18),
.Y(n_166)
);

BUFx2_ASAP7_75t_SL g167 ( 
.A(n_128),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_39),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_69),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_53),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_127),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g173 ( 
.A(n_17),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_122),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_87),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_30),
.Y(n_176)
);

INVxp33_ASAP7_75t_SL g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_38),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_98),
.B(n_56),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_4),
.Y(n_180)
);

INVxp33_ASAP7_75t_SL g181 ( 
.A(n_119),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_82),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_44),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_105),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_5),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_32),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_66),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_108),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_92),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_49),
.B(n_19),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_40),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_61),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_55),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_3),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g196 ( 
.A(n_68),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_101),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_100),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_29),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_33),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_52),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_31),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_79),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_20),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_76),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_9),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_123),
.B(n_104),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_51),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_106),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_16),
.B(n_65),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_117),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_77),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_130),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_34),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_62),
.Y(n_217)
);

HB1xp67_ASAP7_75t_L g218 ( 
.A(n_125),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_116),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_75),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_54),
.Y(n_221)
);

INVxp67_ASAP7_75t_SL g222 ( 
.A(n_26),
.Y(n_222)
);

INVxp33_ASAP7_75t_L g223 ( 
.A(n_10),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_90),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_103),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_35),
.Y(n_226)
);

NOR2xp67_ASAP7_75t_L g227 ( 
.A(n_2),
.B(n_57),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_43),
.Y(n_228)
);

INVx1_ASAP7_75t_SL g229 ( 
.A(n_94),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_97),
.Y(n_230)
);

INVxp67_ASAP7_75t_SL g231 ( 
.A(n_95),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_8),
.Y(n_232)
);

OR2x6_ASAP7_75t_L g233 ( 
.A(n_196),
.B(n_6),
.Y(n_233)
);

NAND3xp33_ASAP7_75t_L g234 ( 
.A(n_218),
.B(n_11),
.C(n_12),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_147),
.Y(n_237)
);

INVx2_ASAP7_75t_SL g238 ( 
.A(n_213),
.Y(n_238)
);

AND2x6_ASAP7_75t_L g239 ( 
.A(n_157),
.B(n_13),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_137),
.B(n_15),
.Y(n_240)
);

AND2x6_ASAP7_75t_L g241 ( 
.A(n_208),
.B(n_21),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_144),
.B(n_22),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_138),
.B(n_139),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g244 ( 
.A(n_143),
.Y(n_244)
);

AND2x4_ASAP7_75t_L g245 ( 
.A(n_145),
.B(n_23),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_150),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_154),
.B(n_24),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_159),
.B(n_28),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_136),
.B(n_36),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_223),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_165),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_170),
.B(n_48),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_174),
.B(n_178),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_182),
.B(n_50),
.Y(n_254)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_140),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_149),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_177),
.A2(n_58),
.B1(n_70),
.B2(n_71),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_183),
.B(n_72),
.Y(n_258)
);

BUFx2_ASAP7_75t_L g259 ( 
.A(n_151),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_186),
.Y(n_260)
);

AND2x2_ASAP7_75t_SL g261 ( 
.A(n_215),
.B(n_74),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_187),
.B(n_190),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_192),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_195),
.Y(n_264)
);

INVx1_ASAP7_75t_SL g265 ( 
.A(n_155),
.Y(n_265)
);

AND2x2_ASAP7_75t_SL g266 ( 
.A(n_199),
.B(n_78),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_200),
.B(n_201),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_202),
.B(n_83),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_203),
.B(n_86),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_205),
.B(n_88),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_206),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_207),
.B(n_219),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_217),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_221),
.B(n_109),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_224),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g276 ( 
.A(n_225),
.B(n_111),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_249),
.B(n_181),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_261),
.B(n_229),
.Y(n_278)
);

NAND2xp33_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_162),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_266),
.B(n_245),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_276),
.B(n_244),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_173),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g283 ( 
.A(n_242),
.B(n_160),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_243),
.B(n_161),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_253),
.B(n_185),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_262),
.B(n_184),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_267),
.B(n_188),
.Y(n_287)
);

XNOR2x2_ASAP7_75t_L g288 ( 
.A(n_237),
.B(n_214),
.Y(n_288)
);

NAND2xp33_ASAP7_75t_SL g289 ( 
.A(n_247),
.B(n_168),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_238),
.B(n_167),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_189),
.Y(n_291)
);

NAND2xp33_ASAP7_75t_SL g292 ( 
.A(n_257),
.B(n_193),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_256),
.B(n_180),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_250),
.B(n_232),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_255),
.B(n_230),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_235),
.B(n_216),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_236),
.B(n_176),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_264),
.B(n_175),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_251),
.B(n_194),
.Y(n_299)
);

AND2x4_ASAP7_75t_L g300 ( 
.A(n_263),
.B(n_197),
.Y(n_300)
);

AND2x4_ASAP7_75t_L g301 ( 
.A(n_271),
.B(n_166),
.Y(n_301)
);

A2O1A1Ixp33_ASAP7_75t_L g302 ( 
.A1(n_280),
.A2(n_292),
.B(n_268),
.C(n_283),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_285),
.A2(n_252),
.B(n_274),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g304 ( 
.A1(n_286),
.A2(n_240),
.B(n_258),
.Y(n_304)
);

AO21x2_ASAP7_75t_L g305 ( 
.A1(n_278),
.A2(n_248),
.B(n_270),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_233),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_233),
.Y(n_307)
);

O2A1O1Ixp33_ASAP7_75t_L g308 ( 
.A1(n_277),
.A2(n_275),
.B(n_273),
.C(n_254),
.Y(n_308)
);

AOI22xp33_ASAP7_75t_SL g309 ( 
.A1(n_288),
.A2(n_259),
.B1(n_226),
.B2(n_158),
.Y(n_309)
);

AO21x2_ASAP7_75t_L g310 ( 
.A1(n_294),
.A2(n_234),
.B(n_227),
.Y(n_310)
);

OAI21x1_ASAP7_75t_SL g311 ( 
.A1(n_295),
.A2(n_156),
.B(n_209),
.Y(n_311)
);

AOI21x1_ASAP7_75t_L g312 ( 
.A1(n_287),
.A2(n_291),
.B(n_298),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_296),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_301),
.Y(n_314)
);

O2A1O1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_281),
.A2(n_260),
.B(n_246),
.C(n_284),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_282),
.B(n_164),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_315),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_300),
.Y(n_318)
);

NAND2xp33_ASAP7_75t_R g319 ( 
.A(n_316),
.B(n_299),
.Y(n_319)
);

AND2x2_ASAP7_75t_L g320 ( 
.A(n_314),
.B(n_293),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_307),
.B(n_289),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_312),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_L g323 ( 
.A(n_309),
.B(n_279),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_306),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_310),
.B(n_169),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_241),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_317),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_303),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_318),
.Y(n_329)
);

AO21x2_ASAP7_75t_L g330 ( 
.A1(n_326),
.A2(n_304),
.B(n_305),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_321),
.A2(n_308),
.B1(n_152),
.B2(n_231),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_322),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_324),
.Y(n_333)
);

INVx2_ASAP7_75t_L g334 ( 
.A(n_327),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_329),
.B(n_323),
.Y(n_335)
);

OAI22xp33_ASAP7_75t_L g336 ( 
.A1(n_333),
.A2(n_319),
.B1(n_222),
.B2(n_325),
.Y(n_336)
);

OAI22xp33_ASAP7_75t_L g337 ( 
.A1(n_328),
.A2(n_172),
.B1(n_211),
.B2(n_210),
.Y(n_337)
);

NOR4xp25_ASAP7_75t_SL g338 ( 
.A(n_332),
.B(n_163),
.C(n_204),
.D(n_198),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_334),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_335),
.A2(n_331),
.B1(n_330),
.B2(n_241),
.Y(n_340)
);

OAI221xp5_ASAP7_75t_L g341 ( 
.A1(n_336),
.A2(n_179),
.B1(n_212),
.B2(n_191),
.C(n_141),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_339),
.Y(n_342)
);

AOI22x1_ASAP7_75t_L g343 ( 
.A1(n_342),
.A2(n_311),
.B1(n_338),
.B2(n_228),
.Y(n_343)
);

NAND3xp33_ASAP7_75t_SL g344 ( 
.A(n_343),
.B(n_341),
.C(n_340),
.Y(n_344)
);

INVx1_ASAP7_75t_SL g345 ( 
.A(n_344),
.Y(n_345)
);

AOI31xp33_ASAP7_75t_L g346 ( 
.A1(n_345),
.A2(n_337),
.A3(n_171),
.B(n_220),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_346),
.A2(n_148),
.B1(n_142),
.B2(n_146),
.Y(n_347)
);

OAI221xp5_ASAP7_75t_R g348 ( 
.A1(n_347),
.A2(n_114),
.B1(n_126),
.B2(n_134),
.C(n_239),
.Y(n_348)
);


endmodule