module fake_jpeg_11552_n_139 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_139);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_139;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_22;
wire n_138;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_7),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g15 ( 
.A(n_5),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx12f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx4f_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

INVx1_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_11),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_30),
.B(n_32),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_18),
.B(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_33),
.Y(n_61)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_42),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_23),
.Y(n_43)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_27),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_46),
.Y(n_64)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_12),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_47),
.B(n_28),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_50),
.B(n_63),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_24),
.B1(n_22),
.B2(n_20),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_56),
.B1(n_66),
.B2(n_34),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_42),
.A2(n_26),
.B1(n_20),
.B2(n_24),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_36),
.B(n_22),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_68),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_65),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_43),
.A2(n_21),
.B1(n_26),
.B2(n_27),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_41),
.B(n_14),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_39),
.B(n_14),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_33),
.Y(n_83)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_64),
.Y(n_74)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_74),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_49),
.B(n_28),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_77),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_68),
.B(n_10),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_78),
.B(n_80),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_59),
.B(n_28),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_81),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_70),
.A2(n_38),
.B1(n_29),
.B2(n_19),
.Y(n_82)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_82),
.A2(n_90),
.B(n_91),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_86),
.Y(n_93)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_52),
.Y(n_84)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_51),
.A2(n_47),
.B1(n_37),
.B2(n_31),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_85),
.A2(n_87),
.B1(n_53),
.B2(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_19),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_54),
.Y(n_88)
);

INVx13_ASAP7_75t_L g105 ( 
.A(n_88),
.Y(n_105)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_89),
.B(n_62),
.C(n_69),
.Y(n_98)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_62),
.B(n_19),
.C(n_2),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_0),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_100),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_53),
.B1(n_48),
.B2(n_39),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_103),
.B1(n_104),
.B2(n_60),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_83),
.B(n_57),
.C(n_69),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_76),
.A2(n_71),
.B1(n_60),
.B2(n_61),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_100),
.A2(n_99),
.B1(n_94),
.B2(n_92),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_107),
.A2(n_111),
.B(n_116),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_101),
.A2(n_82),
.B1(n_76),
.B2(n_75),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_109),
.A2(n_112),
.B1(n_96),
.B2(n_97),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_110),
.B(n_114),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_101),
.A2(n_91),
.B(n_88),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_106),
.A2(n_90),
.B1(n_89),
.B2(n_84),
.Y(n_112)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_113),
.B(n_102),
.C(n_3),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_93),
.A2(n_81),
.B1(n_73),
.B2(n_71),
.Y(n_114)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_96),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_61),
.B(n_33),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_115),
.B(n_102),
.C(n_95),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_117),
.A2(n_107),
.B(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_114),
.B(n_95),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g126 ( 
.A(n_118),
.Y(n_126)
);

AOI322xp5_ASAP7_75t_SL g129 ( 
.A1(n_120),
.A2(n_1),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C1(n_124),
.C2(n_123),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_111),
.A2(n_106),
.B(n_97),
.Y(n_121)
);

AO221x1_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_124),
.B1(n_109),
.B2(n_105),
.C(n_108),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_122),
.A2(n_110),
.B1(n_96),
.B2(n_105),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_125),
.B(n_4),
.C(n_6),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_127),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_128),
.A2(n_129),
.B1(n_119),
.B2(n_5),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_130),
.B(n_131),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_132),
.A2(n_126),
.B1(n_127),
.B2(n_125),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_131),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_136),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_130),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_137),
.B(n_133),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_138),
.B(n_6),
.Y(n_139)
);


endmodule