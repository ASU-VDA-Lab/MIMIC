module real_aes_7409_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_319;
wire n_421;
wire n_555;
wire n_766;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_453;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_769;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_765;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g115 ( .A(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g490 ( .A(n_1), .Y(n_490) );
INVx1_ASAP7_75t_L g203 ( .A(n_2), .Y(n_203) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_3), .A2(n_37), .B1(n_164), .B2(n_520), .Y(n_535) );
AOI21xp33_ASAP7_75t_L g171 ( .A1(n_4), .A2(n_145), .B(n_172), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_5), .B(n_138), .Y(n_503) );
AND2x6_ASAP7_75t_L g150 ( .A(n_6), .B(n_151), .Y(n_150) );
AOI21xp5_ASAP7_75t_L g252 ( .A1(n_7), .A2(n_253), .B(n_254), .Y(n_252) );
NOR2xp33_ASAP7_75t_L g116 ( .A(n_8), .B(n_38), .Y(n_116) );
INVx1_ASAP7_75t_L g178 ( .A(n_9), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_10), .B(n_245), .Y(n_244) );
INVx1_ASAP7_75t_L g143 ( .A(n_11), .Y(n_143) );
INVx1_ASAP7_75t_L g484 ( .A(n_12), .Y(n_484) );
INVx1_ASAP7_75t_L g259 ( .A(n_13), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_14), .B(n_186), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_15), .B(n_139), .Y(n_561) );
AO32x2_ASAP7_75t_L g533 ( .A1(n_16), .A2(n_138), .A3(n_183), .B1(n_512), .B2(n_534), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_17), .A2(n_62), .B1(n_127), .B2(n_128), .Y(n_126) );
INVx1_ASAP7_75t_L g128 ( .A(n_17), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_18), .B(n_164), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_19), .B(n_159), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_20), .B(n_139), .Y(n_493) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_21), .A2(n_50), .B1(n_164), .B2(n_520), .Y(n_536) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_22), .B(n_145), .Y(n_215) );
AOI22xp33_ASAP7_75t_SL g521 ( .A1(n_23), .A2(n_78), .B1(n_164), .B2(n_186), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_24), .B(n_164), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_25), .B(n_167), .Y(n_166) );
A2O1A1Ixp33_ASAP7_75t_L g256 ( .A1(n_26), .A2(n_257), .B(n_258), .C(n_260), .Y(n_256) );
BUFx6f_ASAP7_75t_L g149 ( .A(n_27), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_28), .B(n_180), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_29), .B(n_176), .Y(n_205) );
INVx1_ASAP7_75t_L g192 ( .A(n_30), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g122 ( .A1(n_31), .A2(n_123), .B1(n_124), .B2(n_455), .Y(n_122) );
INVx1_ASAP7_75t_L g455 ( .A(n_31), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_32), .B(n_180), .Y(n_550) );
INVx2_ASAP7_75t_L g148 ( .A(n_33), .Y(n_148) );
NAND2xp5_ASAP7_75t_SL g507 ( .A(n_34), .B(n_164), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_35), .B(n_180), .Y(n_532) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_36), .A2(n_150), .B(n_154), .C(n_217), .Y(n_216) );
INVx1_ASAP7_75t_L g190 ( .A(n_39), .Y(n_190) );
OAI22xp5_ASAP7_75t_SL g764 ( .A1(n_40), .A2(n_765), .B1(n_768), .B2(n_769), .Y(n_764) );
CKINVDCx20_ASAP7_75t_R g769 ( .A(n_40), .Y(n_769) );
NAND2xp5_ASAP7_75t_SL g231 ( .A(n_41), .B(n_176), .Y(n_231) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_42), .B(n_164), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g519 ( .A1(n_43), .A2(n_89), .B1(n_222), .B2(n_520), .Y(n_519) );
NAND2xp5_ASAP7_75t_SL g501 ( .A(n_44), .B(n_164), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_45), .B(n_164), .Y(n_485) );
CKINVDCx16_ASAP7_75t_R g193 ( .A(n_46), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g765 ( .A1(n_47), .A2(n_71), .B1(n_766), .B2(n_767), .Y(n_765) );
CKINVDCx16_ASAP7_75t_R g767 ( .A(n_47), .Y(n_767) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_48), .B(n_489), .Y(n_502) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_49), .B(n_145), .Y(n_247) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_51), .A2(n_60), .B1(n_164), .B2(n_186), .Y(n_559) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_52), .A2(n_154), .B1(n_186), .B2(n_188), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g225 ( .A(n_53), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_54), .B(n_164), .Y(n_511) );
CKINVDCx16_ASAP7_75t_R g200 ( .A(n_55), .Y(n_200) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_56), .B(n_164), .Y(n_526) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_57), .A2(n_163), .B(n_175), .C(n_177), .Y(n_174) );
CKINVDCx20_ASAP7_75t_R g235 ( .A(n_58), .Y(n_235) );
INVx1_ASAP7_75t_L g173 ( .A(n_59), .Y(n_173) );
INVx1_ASAP7_75t_L g151 ( .A(n_61), .Y(n_151) );
INVx1_ASAP7_75t_L g127 ( .A(n_62), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g458 ( .A(n_63), .B(n_459), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_64), .B(n_164), .Y(n_491) );
INVx1_ASAP7_75t_L g142 ( .A(n_65), .Y(n_142) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_66), .Y(n_120) );
AO32x2_ASAP7_75t_L g517 ( .A1(n_67), .A2(n_138), .A3(n_239), .B1(n_512), .B2(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g510 ( .A(n_68), .Y(n_510) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_69), .A2(n_104), .B1(n_117), .B2(n_777), .Y(n_103) );
INVx1_ASAP7_75t_L g545 ( .A(n_70), .Y(n_545) );
INVx1_ASAP7_75t_L g766 ( .A(n_71), .Y(n_766) );
A2O1A1Ixp33_ASAP7_75t_SL g158 ( .A1(n_72), .A2(n_159), .B(n_160), .C(n_163), .Y(n_158) );
INVxp67_ASAP7_75t_L g161 ( .A(n_73), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g546 ( .A(n_74), .B(n_186), .Y(n_546) );
INVx1_ASAP7_75t_L g110 ( .A(n_75), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g196 ( .A(n_76), .Y(n_196) );
INVx1_ASAP7_75t_L g228 ( .A(n_77), .Y(n_228) );
AOI222xp33_ASAP7_75t_L g461 ( .A1(n_79), .A2(n_462), .B1(n_763), .B2(n_764), .C1(n_770), .C2(n_771), .Y(n_461) );
A2O1A1Ixp33_ASAP7_75t_L g229 ( .A1(n_80), .A2(n_150), .B(n_154), .C(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_81), .B(n_520), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_82), .B(n_186), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g218 ( .A(n_83), .B(n_204), .Y(n_218) );
INVx2_ASAP7_75t_L g140 ( .A(n_84), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_85), .B(n_159), .Y(n_219) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_86), .B(n_186), .Y(n_499) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_87), .A2(n_150), .B(n_154), .C(n_202), .Y(n_201) );
OR2x2_ASAP7_75t_L g112 ( .A(n_88), .B(n_113), .Y(n_112) );
OR2x2_ASAP7_75t_L g467 ( .A(n_88), .B(n_114), .Y(n_467) );
INVx2_ASAP7_75t_L g470 ( .A(n_88), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_90), .A2(n_102), .B1(n_186), .B2(n_187), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g179 ( .A(n_91), .B(n_180), .Y(n_179) );
CKINVDCx20_ASAP7_75t_R g208 ( .A(n_92), .Y(n_208) );
A2O1A1Ixp33_ASAP7_75t_L g241 ( .A1(n_93), .A2(n_150), .B(n_154), .C(n_242), .Y(n_241) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_94), .Y(n_249) );
INVx1_ASAP7_75t_L g157 ( .A(n_95), .Y(n_157) );
CKINVDCx16_ASAP7_75t_R g255 ( .A(n_96), .Y(n_255) );
NAND2xp5_ASAP7_75t_SL g243 ( .A(n_97), .B(n_204), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_98), .B(n_186), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_99), .B(n_138), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_100), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g144 ( .A1(n_101), .A2(n_145), .B(n_152), .Y(n_144) );
CKINVDCx20_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_106), .Y(n_105) );
CKINVDCx6p67_ASAP7_75t_R g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_L g778 ( .A(n_107), .Y(n_778) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_108), .B(n_111), .Y(n_107) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVx1_ASAP7_75t_SL g111 ( .A(n_112), .Y(n_111) );
HB1xp67_ASAP7_75t_L g457 ( .A(n_112), .Y(n_457) );
NOR2x2_ASAP7_75t_L g770 ( .A(n_113), .B(n_470), .Y(n_770) );
INVx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
OR2x2_ASAP7_75t_L g469 ( .A(n_114), .B(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
AO21x1_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_121), .B(n_460), .Y(n_117) );
INVx2_ASAP7_75t_SL g118 ( .A(n_119), .Y(n_118) );
BUFx2_ASAP7_75t_L g776 ( .A(n_119), .Y(n_776) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_456), .B(n_458), .Y(n_121) );
INVx1_ASAP7_75t_L g123 ( .A(n_124), .Y(n_123) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_126), .B1(n_129), .B2(n_454), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx2_ASAP7_75t_L g454 ( .A(n_129), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g463 ( .A1(n_129), .A2(n_464), .B1(n_468), .B2(n_471), .Y(n_463) );
INVx1_ASAP7_75t_SL g773 ( .A(n_129), .Y(n_773) );
INVx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
AND4x1_ASAP7_75t_L g130 ( .A(n_131), .B(n_372), .C(n_419), .D(n_439), .Y(n_130) );
NOR3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_302), .C(n_327), .Y(n_131) );
OAI211xp5_ASAP7_75t_SL g132 ( .A1(n_133), .A2(n_210), .B(n_262), .C(n_292), .Y(n_132) );
INVxp67_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g134 ( .A(n_135), .B(n_181), .Y(n_134) );
INVx3_ASAP7_75t_SL g344 ( .A(n_135), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_135), .B(n_275), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_135), .B(n_197), .Y(n_425) );
AND2x2_ASAP7_75t_L g448 ( .A(n_135), .B(n_314), .Y(n_448) );
AND2x4_ASAP7_75t_L g135 ( .A(n_136), .B(n_169), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_L g266 ( .A(n_137), .B(n_170), .Y(n_266) );
INVx3_ASAP7_75t_L g279 ( .A(n_137), .Y(n_279) );
AND2x2_ASAP7_75t_L g284 ( .A(n_137), .B(n_169), .Y(n_284) );
OR2x2_ASAP7_75t_L g335 ( .A(n_137), .B(n_276), .Y(n_335) );
BUFx2_ASAP7_75t_L g355 ( .A(n_137), .Y(n_355) );
AND2x2_ASAP7_75t_L g365 ( .A(n_137), .B(n_276), .Y(n_365) );
AND2x2_ASAP7_75t_L g371 ( .A(n_137), .B(n_182), .Y(n_371) );
OA21x2_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_144), .B(n_166), .Y(n_137) );
INVx4_ASAP7_75t_L g168 ( .A(n_138), .Y(n_168) );
OA21x2_ASAP7_75t_L g495 ( .A1(n_138), .A2(n_496), .B(n_503), .Y(n_495) );
BUFx6f_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx1_ASAP7_75t_L g183 ( .A(n_139), .Y(n_183) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_141), .Y(n_139) );
AND2x2_ASAP7_75t_SL g180 ( .A(n_140), .B(n_141), .Y(n_180) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_143), .Y(n_141) );
BUFx2_ASAP7_75t_L g253 ( .A(n_145), .Y(n_253) );
AND2x4_ASAP7_75t_L g145 ( .A(n_146), .B(n_150), .Y(n_145) );
NAND2x1p5_ASAP7_75t_L g194 ( .A(n_146), .B(n_150), .Y(n_194) );
AND2x2_ASAP7_75t_L g146 ( .A(n_147), .B(n_149), .Y(n_146) );
INVx1_ASAP7_75t_L g489 ( .A(n_147), .Y(n_489) );
INVx1_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g155 ( .A(n_148), .Y(n_155) );
INVx1_ASAP7_75t_L g187 ( .A(n_148), .Y(n_187) );
INVx1_ASAP7_75t_L g156 ( .A(n_149), .Y(n_156) );
INVx1_ASAP7_75t_L g159 ( .A(n_149), .Y(n_159) );
INVx3_ASAP7_75t_L g162 ( .A(n_149), .Y(n_162) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_149), .Y(n_176) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_149), .Y(n_189) );
INVx4_ASAP7_75t_SL g165 ( .A(n_150), .Y(n_165) );
OAI21xp5_ASAP7_75t_L g482 ( .A1(n_150), .A2(n_483), .B(n_487), .Y(n_482) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_150), .A2(n_497), .B(n_500), .Y(n_496) );
BUFx3_ASAP7_75t_L g512 ( .A(n_150), .Y(n_512) );
OAI21xp5_ASAP7_75t_L g524 ( .A1(n_150), .A2(n_525), .B(n_529), .Y(n_524) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_150), .A2(n_544), .B(n_547), .Y(n_543) );
O2A1O1Ixp33_ASAP7_75t_L g152 ( .A1(n_153), .A2(n_157), .B(n_158), .C(n_165), .Y(n_152) );
O2A1O1Ixp33_ASAP7_75t_L g172 ( .A1(n_153), .A2(n_165), .B(n_173), .C(n_174), .Y(n_172) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_153), .A2(n_165), .B(n_255), .C(n_256), .Y(n_254) );
INVx5_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
AND2x6_ASAP7_75t_L g154 ( .A(n_155), .B(n_156), .Y(n_154) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_155), .Y(n_164) );
BUFx3_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
INVx1_ASAP7_75t_L g520 ( .A(n_155), .Y(n_520) );
INVx1_ASAP7_75t_L g528 ( .A(n_159), .Y(n_528) );
NOR2xp33_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_L g177 ( .A(n_162), .B(n_178), .Y(n_177) );
INVx5_ASAP7_75t_L g204 ( .A(n_162), .Y(n_204) );
OAI22xp5_ASAP7_75t_SL g518 ( .A1(n_162), .A2(n_176), .B1(n_519), .B2(n_521), .Y(n_518) );
O2A1O1Ixp5_ASAP7_75t_SL g544 ( .A1(n_163), .A2(n_204), .B(n_545), .C(n_546), .Y(n_544) );
INVx3_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_164), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g184 ( .A1(n_165), .A2(n_185), .B1(n_193), .B2(n_194), .Y(n_184) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_167), .A2(n_171), .B(n_179), .Y(n_170) );
INVx3_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
NOR2xp33_ASAP7_75t_SL g224 ( .A(n_168), .B(n_225), .Y(n_224) );
AO21x1_ASAP7_75t_L g556 ( .A1(n_168), .A2(n_557), .B(n_560), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g575 ( .A(n_168), .B(n_512), .C(n_557), .Y(n_575) );
INVx1_ASAP7_75t_SL g169 ( .A(n_170), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_170), .B(n_276), .Y(n_290) );
INVx2_ASAP7_75t_L g300 ( .A(n_170), .Y(n_300) );
AND2x2_ASAP7_75t_L g313 ( .A(n_170), .B(n_279), .Y(n_313) );
OR2x2_ASAP7_75t_L g324 ( .A(n_170), .B(n_276), .Y(n_324) );
AND2x2_ASAP7_75t_SL g370 ( .A(n_170), .B(n_371), .Y(n_370) );
BUFx2_ASAP7_75t_L g382 ( .A(n_170), .Y(n_382) );
AND2x2_ASAP7_75t_L g428 ( .A(n_170), .B(n_182), .Y(n_428) );
O2A1O1Ixp5_ASAP7_75t_L g509 ( .A1(n_175), .A2(n_488), .B(n_510), .C(n_511), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_175), .A2(n_530), .B(n_531), .Y(n_529) );
INVx2_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx4_ASAP7_75t_L g245 ( .A(n_176), .Y(n_245) );
OAI22xp5_ASAP7_75t_L g534 ( .A1(n_176), .A2(n_492), .B1(n_535), .B2(n_536), .Y(n_534) );
OAI22xp5_ASAP7_75t_L g557 ( .A1(n_176), .A2(n_492), .B1(n_558), .B2(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g209 ( .A(n_180), .Y(n_209) );
INVx2_ASAP7_75t_L g239 ( .A(n_180), .Y(n_239) );
OA21x2_ASAP7_75t_L g251 ( .A1(n_180), .A2(n_252), .B(n_261), .Y(n_251) );
OA21x2_ASAP7_75t_L g523 ( .A1(n_180), .A2(n_524), .B(n_532), .Y(n_523) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_180), .A2(n_543), .B(n_550), .Y(n_542) );
INVx3_ASAP7_75t_SL g301 ( .A(n_181), .Y(n_301) );
OR2x2_ASAP7_75t_L g354 ( .A(n_181), .B(n_355), .Y(n_354) );
OR2x2_ASAP7_75t_L g181 ( .A(n_182), .B(n_197), .Y(n_181) );
INVx3_ASAP7_75t_L g276 ( .A(n_182), .Y(n_276) );
AND2x2_ASAP7_75t_L g343 ( .A(n_182), .B(n_198), .Y(n_343) );
HB1xp67_ASAP7_75t_L g411 ( .A(n_182), .Y(n_411) );
AOI33xp33_ASAP7_75t_L g415 ( .A1(n_182), .A2(n_344), .A3(n_351), .B1(n_360), .B2(n_416), .B3(n_417), .Y(n_415) );
AO21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_195), .Y(n_182) );
NOR2xp33_ASAP7_75t_L g195 ( .A(n_183), .B(n_196), .Y(n_195) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_183), .A2(n_199), .B(n_207), .Y(n_198) );
INVx2_ASAP7_75t_L g223 ( .A(n_183), .Y(n_223) );
INVx2_ASAP7_75t_L g206 ( .A(n_186), .Y(n_206) );
INVx3_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
OAI22xp5_ASAP7_75t_SL g188 ( .A1(n_189), .A2(n_190), .B1(n_191), .B2(n_192), .Y(n_188) );
INVx2_ASAP7_75t_L g191 ( .A(n_189), .Y(n_191) );
INVx4_ASAP7_75t_L g257 ( .A(n_189), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g199 ( .A1(n_194), .A2(n_200), .B(n_201), .Y(n_199) );
OAI21xp5_ASAP7_75t_L g227 ( .A1(n_194), .A2(n_228), .B(n_229), .Y(n_227) );
INVx1_ASAP7_75t_L g264 ( .A(n_197), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_197), .B(n_279), .Y(n_278) );
NOR3xp33_ASAP7_75t_L g338 ( .A(n_197), .B(n_339), .C(n_341), .Y(n_338) );
AND2x2_ASAP7_75t_L g364 ( .A(n_197), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_197), .B(n_371), .Y(n_374) );
AND2x2_ASAP7_75t_L g427 ( .A(n_197), .B(n_428), .Y(n_427) );
INVx3_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx3_ASAP7_75t_L g283 ( .A(n_198), .Y(n_283) );
OR2x2_ASAP7_75t_L g377 ( .A(n_198), .B(n_276), .Y(n_377) );
O2A1O1Ixp33_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .C(n_206), .Y(n_202) );
INVx2_ASAP7_75t_L g492 ( .A(n_204), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_204), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_204), .A2(n_507), .B(n_508), .Y(n_506) );
O2A1O1Ixp33_ASAP7_75t_L g483 ( .A1(n_206), .A2(n_484), .B(n_485), .C(n_486), .Y(n_483) );
NOR2xp33_ASAP7_75t_L g207 ( .A(n_208), .B(n_209), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g234 ( .A(n_209), .B(n_235), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_209), .B(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g210 ( .A(n_211), .B(n_236), .Y(n_210) );
AOI32xp33_ASAP7_75t_L g328 ( .A1(n_211), .A2(n_329), .A3(n_331), .B1(n_333), .B2(n_336), .Y(n_328) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_211), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g431 ( .A(n_211), .Y(n_431) );
INVx4_ASAP7_75t_L g211 ( .A(n_212), .Y(n_211) );
AND2x2_ASAP7_75t_L g363 ( .A(n_212), .B(n_347), .Y(n_363) );
AND2x2_ASAP7_75t_L g383 ( .A(n_212), .B(n_309), .Y(n_383) );
AND2x2_ASAP7_75t_L g451 ( .A(n_212), .B(n_369), .Y(n_451) );
AND2x2_ASAP7_75t_L g212 ( .A(n_213), .B(n_226), .Y(n_212) );
INVx3_ASAP7_75t_L g272 ( .A(n_213), .Y(n_272) );
AND2x2_ASAP7_75t_L g286 ( .A(n_213), .B(n_270), .Y(n_286) );
OR2x2_ASAP7_75t_L g291 ( .A(n_213), .B(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g298 ( .A(n_213), .Y(n_298) );
AND2x2_ASAP7_75t_L g306 ( .A(n_213), .B(n_280), .Y(n_306) );
AND2x2_ASAP7_75t_L g308 ( .A(n_213), .B(n_309), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_213), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g361 ( .A(n_213), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_213), .B(n_446), .Y(n_445) );
OR2x6_ASAP7_75t_L g213 ( .A(n_214), .B(n_224), .Y(n_213) );
AOI21xp5_ASAP7_75t_SL g214 ( .A1(n_215), .A2(n_216), .B(n_223), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_218), .A2(n_219), .B(n_220), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_220), .A2(n_231), .B(n_232), .Y(n_230) );
INVx2_ASAP7_75t_L g220 ( .A(n_221), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g260 ( .A(n_222), .Y(n_260) );
INVx1_ASAP7_75t_L g233 ( .A(n_223), .Y(n_233) );
OA21x2_ASAP7_75t_L g481 ( .A1(n_223), .A2(n_482), .B(n_493), .Y(n_481) );
OA21x2_ASAP7_75t_L g504 ( .A1(n_223), .A2(n_505), .B(n_513), .Y(n_504) );
INVx2_ASAP7_75t_L g270 ( .A(n_226), .Y(n_270) );
AND2x2_ASAP7_75t_L g316 ( .A(n_226), .B(n_237), .Y(n_316) );
AND2x2_ASAP7_75t_L g326 ( .A(n_226), .B(n_251), .Y(n_326) );
AO21x2_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_233), .B(n_234), .Y(n_226) );
INVx2_ASAP7_75t_L g446 ( .A(n_236), .Y(n_446) );
OR2x2_ASAP7_75t_L g236 ( .A(n_237), .B(n_250), .Y(n_236) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_237), .B(n_270), .Y(n_269) );
INVx1_ASAP7_75t_L g287 ( .A(n_237), .Y(n_287) );
AND2x2_ASAP7_75t_L g331 ( .A(n_237), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g347 ( .A(n_237), .B(n_310), .Y(n_347) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx1_ASAP7_75t_L g295 ( .A(n_238), .Y(n_295) );
AND2x2_ASAP7_75t_L g309 ( .A(n_238), .B(n_310), .Y(n_309) );
AND2x2_ASAP7_75t_L g360 ( .A(n_238), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g392 ( .A(n_238), .B(n_270), .Y(n_392) );
AO21x2_ASAP7_75t_L g238 ( .A1(n_239), .A2(n_240), .B(n_248), .Y(n_238) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_241), .B(n_247), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g242 ( .A1(n_243), .A2(n_244), .B(n_246), .Y(n_242) );
AND2x2_ASAP7_75t_L g271 ( .A(n_250), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g332 ( .A(n_250), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_250), .B(n_340), .Y(n_339) );
INVx1_ASAP7_75t_L g369 ( .A(n_250), .Y(n_369) );
INVx1_ASAP7_75t_L g402 ( .A(n_250), .Y(n_402) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
AND2x2_ASAP7_75t_L g280 ( .A(n_251), .B(n_270), .Y(n_280) );
INVx1_ASAP7_75t_L g310 ( .A(n_251), .Y(n_310) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_257), .B(n_259), .Y(n_258) );
INVx1_ASAP7_75t_L g486 ( .A(n_257), .Y(n_486) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_257), .A2(n_548), .B(n_549), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g262 ( .A1(n_263), .A2(n_267), .B1(n_273), .B2(n_280), .C(n_281), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_264), .B(n_265), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_264), .B(n_284), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_264), .B(n_347), .Y(n_424) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_266), .B(n_314), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_266), .B(n_275), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_266), .B(n_289), .Y(n_418) );
AND2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_271), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g340 ( .A(n_270), .Y(n_340) );
AND2x2_ASAP7_75t_L g315 ( .A(n_271), .B(n_316), .Y(n_315) );
INVx1_ASAP7_75t_L g393 ( .A(n_271), .Y(n_393) );
AND2x2_ASAP7_75t_L g325 ( .A(n_272), .B(n_326), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_272), .B(n_295), .Y(n_341) );
AND2x2_ASAP7_75t_L g405 ( .A(n_272), .B(n_331), .Y(n_405) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_275), .B(n_277), .Y(n_274) );
BUFx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g314 ( .A(n_276), .B(n_283), .Y(n_314) );
AND2x2_ASAP7_75t_L g410 ( .A(n_277), .B(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_279), .B(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_280), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_280), .B(n_287), .Y(n_375) );
AND2x2_ASAP7_75t_L g395 ( .A(n_280), .B(n_295), .Y(n_395) );
AND2x2_ASAP7_75t_L g416 ( .A(n_280), .B(n_360), .Y(n_416) );
OAI32xp33_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_285), .A3(n_287), .B1(n_288), .B2(n_291), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_284), .Y(n_282) );
INVx1_ASAP7_75t_SL g289 ( .A(n_283), .Y(n_289) );
NAND2x1_ASAP7_75t_L g330 ( .A(n_283), .B(n_313), .Y(n_330) );
OR2x2_ASAP7_75t_L g334 ( .A(n_283), .B(n_335), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_283), .B(n_382), .Y(n_435) );
INVx1_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
OAI221xp5_ASAP7_75t_SL g421 ( .A1(n_285), .A2(n_376), .B1(n_422), .B2(n_425), .C(n_426), .Y(n_421) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g293 ( .A(n_286), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g336 ( .A(n_286), .B(n_309), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_286), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g414 ( .A(n_286), .B(n_347), .Y(n_414) );
INVxp67_ASAP7_75t_L g350 ( .A(n_287), .Y(n_350) );
OR2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
AND2x2_ASAP7_75t_L g420 ( .A(n_289), .B(n_407), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_289), .B(n_370), .Y(n_443) );
INVx1_ASAP7_75t_L g318 ( .A(n_291), .Y(n_318) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_291), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g436 ( .A(n_291), .B(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_296), .B(n_299), .Y(n_292) );
AND2x2_ASAP7_75t_L g305 ( .A(n_294), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g389 ( .A(n_298), .B(n_309), .Y(n_389) );
AND2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_301), .Y(n_299) );
AND2x2_ASAP7_75t_L g407 ( .A(n_300), .B(n_365), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_300), .B(n_364), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_301), .B(n_313), .Y(n_387) );
OAI211xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_304), .B(n_307), .C(n_317), .Y(n_302) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_303), .A2(n_338), .B1(n_342), .B2(n_345), .C(n_348), .Y(n_337) );
AOI31xp33_ASAP7_75t_L g432 ( .A1(n_303), .A2(n_433), .A3(n_434), .B(n_436), .Y(n_432) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
AOI22xp5_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_311), .B1(n_313), .B2(n_315), .Y(n_307) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g433 ( .A(n_313), .Y(n_433) );
INVx1_ASAP7_75t_L g396 ( .A(n_314), .Y(n_396) );
O2A1O1Ixp33_ASAP7_75t_L g439 ( .A1(n_316), .A2(n_440), .B(n_442), .C(n_444), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_321), .B2(n_325), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_322), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
OAI221xp5_ASAP7_75t_SL g412 ( .A1(n_324), .A2(n_358), .B1(n_377), .B2(n_413), .C(n_415), .Y(n_412) );
INVx1_ASAP7_75t_L g408 ( .A(n_325), .Y(n_408) );
INVx1_ASAP7_75t_L g362 ( .A(n_326), .Y(n_362) );
NAND3xp33_ASAP7_75t_SL g327 ( .A(n_328), .B(n_337), .C(n_352), .Y(n_327) );
OAI21xp33_ASAP7_75t_L g378 ( .A1(n_329), .A2(n_379), .B(n_383), .Y(n_378) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_331), .B(n_431), .Y(n_430) );
INVxp67_ASAP7_75t_L g438 ( .A(n_332), .Y(n_438) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
OR2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_359), .Y(n_376) );
INVx1_ASAP7_75t_L g351 ( .A(n_340), .Y(n_351) );
AND2x2_ASAP7_75t_L g342 ( .A(n_343), .B(n_344), .Y(n_342) );
INVx1_ASAP7_75t_L g349 ( .A(n_343), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_343), .B(n_381), .Y(n_380) );
NOR4xp25_ASAP7_75t_L g348 ( .A(n_344), .B(n_349), .C(n_350), .D(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
AOI222xp33_ASAP7_75t_L g352 ( .A1(n_353), .A2(n_357), .B1(n_363), .B2(n_364), .C1(n_366), .C2(n_370), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_354), .B(n_356), .Y(n_353) );
INVx1_ASAP7_75t_L g450 ( .A(n_354), .Y(n_450) );
INVx1_ASAP7_75t_SL g357 ( .A(n_358), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_359), .B(n_362), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_366), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OAI21xp5_ASAP7_75t_SL g426 ( .A1(n_371), .A2(n_427), .B(n_429), .Y(n_426) );
NOR4xp25_ASAP7_75t_L g372 ( .A(n_373), .B(n_384), .C(n_397), .D(n_412), .Y(n_372) );
OAI221xp5_ASAP7_75t_SL g373 ( .A1(n_374), .A2(n_375), .B1(n_376), .B2(n_377), .C(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g453 ( .A(n_374), .Y(n_453) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_381), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_SL g381 ( .A(n_382), .Y(n_381) );
OAI222xp33_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_388), .B1(n_390), .B2(n_391), .C1(n_394), .C2(n_396), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI211xp5_ASAP7_75t_L g419 ( .A1(n_389), .A2(n_420), .B(n_421), .C(n_432), .Y(n_419) );
OR2x2_ASAP7_75t_L g391 ( .A(n_392), .B(n_393), .Y(n_391) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OAI222xp33_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_403), .B1(n_404), .B2(n_406), .C1(n_408), .C2(n_409), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx1_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g449 ( .A1(n_414), .A2(n_417), .B1(n_450), .B2(n_451), .Y(n_449) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
HB1xp67_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
OAI211xp5_ASAP7_75t_SL g444 ( .A1(n_445), .A2(n_447), .B(n_449), .C(n_452), .Y(n_444) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g459 ( .A(n_457), .Y(n_459) );
AOI21xp33_ASAP7_75t_L g460 ( .A1(n_458), .A2(n_461), .B(n_775), .Y(n_460) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
INVx1_ASAP7_75t_SL g464 ( .A(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g772 ( .A1(n_466), .A2(n_472), .B1(n_773), .B2(n_774), .Y(n_772) );
INVx1_ASAP7_75t_L g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx6_ASAP7_75t_L g774 ( .A(n_469), .Y(n_774) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
AND2x2_ASAP7_75t_SL g472 ( .A(n_473), .B(n_729), .Y(n_472) );
NOR3xp33_ASAP7_75t_L g473 ( .A(n_474), .B(n_633), .C(n_717), .Y(n_473) );
NAND4xp25_ASAP7_75t_L g474 ( .A(n_475), .B(n_576), .C(n_598), .D(n_614), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_514), .B1(n_537), .B2(n_555), .C(n_562), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_494), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_478), .B(n_555), .Y(n_588) );
NAND4xp25_ASAP7_75t_L g628 ( .A(n_478), .B(n_616), .C(n_629), .D(n_631), .Y(n_628) );
INVxp67_ASAP7_75t_L g745 ( .A(n_478), .Y(n_745) );
INVx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g627 ( .A(n_479), .B(n_565), .Y(n_627) );
AND2x2_ASAP7_75t_L g651 ( .A(n_479), .B(n_494), .Y(n_651) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g618 ( .A(n_480), .B(n_554), .Y(n_618) );
AND2x2_ASAP7_75t_L g658 ( .A(n_480), .B(n_639), .Y(n_658) );
AND2x2_ASAP7_75t_L g675 ( .A(n_480), .B(n_676), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_480), .B(n_495), .Y(n_699) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AND2x2_ASAP7_75t_L g553 ( .A(n_481), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g570 ( .A(n_481), .B(n_571), .Y(n_570) );
AND2x2_ASAP7_75t_L g582 ( .A(n_481), .B(n_495), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_481), .B(n_504), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_490), .B(n_491), .C(n_492), .Y(n_487) );
INVx2_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g500 ( .A1(n_492), .A2(n_501), .B(n_502), .Y(n_500) );
AND2x2_ASAP7_75t_L g585 ( .A(n_494), .B(n_586), .Y(n_585) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_494), .A2(n_635), .B1(n_638), .B2(n_640), .C(n_644), .Y(n_634) );
AND2x2_ASAP7_75t_L g693 ( .A(n_494), .B(n_658), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_494), .B(n_675), .Y(n_727) );
AND2x2_ASAP7_75t_L g494 ( .A(n_495), .B(n_504), .Y(n_494) );
INVx3_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
AND2x2_ASAP7_75t_L g602 ( .A(n_495), .B(n_603), .Y(n_602) );
AND2x2_ASAP7_75t_L g656 ( .A(n_495), .B(n_571), .Y(n_656) );
AND2x2_ASAP7_75t_L g714 ( .A(n_495), .B(n_715), .Y(n_714) );
AND2x2_ASAP7_75t_L g555 ( .A(n_504), .B(n_556), .Y(n_555) );
INVx2_ASAP7_75t_L g571 ( .A(n_504), .Y(n_571) );
INVx1_ASAP7_75t_L g626 ( .A(n_504), .Y(n_626) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_504), .Y(n_632) );
AND2x2_ASAP7_75t_L g677 ( .A(n_504), .B(n_554), .Y(n_677) );
OR2x2_ASAP7_75t_L g716 ( .A(n_504), .B(n_556), .Y(n_716) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_509), .B(n_512), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_514), .B(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_522), .Y(n_514) );
AND2x2_ASAP7_75t_L g712 ( .A(n_515), .B(n_709), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_515), .B(n_694), .Y(n_744) );
BUFx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
AND2x2_ASAP7_75t_L g643 ( .A(n_516), .B(n_567), .Y(n_643) );
AND2x2_ASAP7_75t_L g692 ( .A(n_516), .B(n_540), .Y(n_692) );
INVx1_ASAP7_75t_L g738 ( .A(n_516), .Y(n_738) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
BUFx6f_ASAP7_75t_L g552 ( .A(n_517), .Y(n_552) );
AND2x2_ASAP7_75t_L g593 ( .A(n_517), .B(n_567), .Y(n_593) );
INVx1_ASAP7_75t_L g610 ( .A(n_517), .Y(n_610) );
AND2x2_ASAP7_75t_L g616 ( .A(n_517), .B(n_533), .Y(n_616) );
AND2x2_ASAP7_75t_L g684 ( .A(n_522), .B(n_592), .Y(n_684) );
INVx2_ASAP7_75t_L g749 ( .A(n_522), .Y(n_749) );
AND2x2_ASAP7_75t_L g522 ( .A(n_523), .B(n_533), .Y(n_522) );
AND2x2_ASAP7_75t_L g566 ( .A(n_523), .B(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g579 ( .A(n_523), .B(n_541), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_523), .B(n_540), .Y(n_607) );
INVx1_ASAP7_75t_L g613 ( .A(n_523), .Y(n_613) );
INVx1_ASAP7_75t_L g630 ( .A(n_523), .Y(n_630) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_523), .Y(n_642) );
INVx2_ASAP7_75t_L g710 ( .A(n_523), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_526), .A2(n_527), .B(n_528), .Y(n_525) );
INVx2_ASAP7_75t_L g567 ( .A(n_533), .Y(n_567) );
BUFx2_ASAP7_75t_L g664 ( .A(n_533), .Y(n_664) );
AND2x2_ASAP7_75t_L g709 ( .A(n_533), .B(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_539), .B(n_551), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_539), .B(n_646), .Y(n_645) );
AOI21xp5_ASAP7_75t_L g732 ( .A1(n_539), .A2(n_708), .B(n_722), .Y(n_732) );
AND2x2_ASAP7_75t_L g757 ( .A(n_539), .B(n_643), .Y(n_757) );
BUFx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
INVx2_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
INVx1_ASAP7_75t_L g679 ( .A(n_541), .Y(n_679) );
AND2x2_ASAP7_75t_L g708 ( .A(n_541), .B(n_709), .Y(n_708) );
INVx2_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
HB1xp67_ASAP7_75t_L g592 ( .A(n_542), .Y(n_592) );
INVx2_ASAP7_75t_L g611 ( .A(n_542), .Y(n_611) );
OR2x2_ASAP7_75t_L g612 ( .A(n_542), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
INVx2_ASAP7_75t_L g565 ( .A(n_552), .Y(n_565) );
OR2x2_ASAP7_75t_L g578 ( .A(n_552), .B(n_579), .Y(n_578) );
AND2x2_ASAP7_75t_L g646 ( .A(n_552), .B(n_642), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_552), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g747 ( .A(n_552), .B(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_552), .B(n_684), .Y(n_759) );
AND2x2_ASAP7_75t_L g638 ( .A(n_553), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g661 ( .A(n_553), .B(n_555), .Y(n_661) );
INVx2_ASAP7_75t_L g573 ( .A(n_554), .Y(n_573) );
AND2x2_ASAP7_75t_L g601 ( .A(n_554), .B(n_574), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_554), .B(n_626), .Y(n_682) );
AND2x2_ASAP7_75t_L g596 ( .A(n_555), .B(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g743 ( .A(n_555), .Y(n_743) );
AND2x2_ASAP7_75t_L g755 ( .A(n_555), .B(n_618), .Y(n_755) );
AND2x2_ASAP7_75t_L g581 ( .A(n_556), .B(n_571), .Y(n_581) );
INVx1_ASAP7_75t_L g676 ( .A(n_556), .Y(n_676) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AND2x4_ASAP7_75t_L g574 ( .A(n_561), .B(n_575), .Y(n_574) );
INVxp67_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_564), .B(n_568), .Y(n_563) );
AND2x2_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .Y(n_564) );
NOR2xp33_ASAP7_75t_L g621 ( .A(n_565), .B(n_612), .Y(n_621) );
OR2x2_ASAP7_75t_L g753 ( .A(n_565), .B(n_754), .Y(n_753) );
AND2x2_ASAP7_75t_L g670 ( .A(n_566), .B(n_611), .Y(n_670) );
AND2x2_ASAP7_75t_L g678 ( .A(n_566), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g737 ( .A(n_566), .B(n_738), .Y(n_737) );
AND2x2_ASAP7_75t_L g761 ( .A(n_566), .B(n_608), .Y(n_761) );
NOR2xp67_ASAP7_75t_L g719 ( .A(n_567), .B(n_720), .Y(n_719) );
OR2x2_ASAP7_75t_L g748 ( .A(n_567), .B(n_611), .Y(n_748) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NAND2x1p5_ASAP7_75t_L g569 ( .A(n_570), .B(n_572), .Y(n_569) );
AND2x2_ASAP7_75t_L g600 ( .A(n_570), .B(n_601), .Y(n_600) );
INVxp67_ASAP7_75t_L g762 ( .A(n_570), .Y(n_762) );
NOR2x1_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
INVx1_ASAP7_75t_L g597 ( .A(n_573), .Y(n_597) );
AND2x2_ASAP7_75t_L g648 ( .A(n_573), .B(n_581), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g742 ( .A(n_573), .B(n_716), .Y(n_742) );
INVx2_ASAP7_75t_L g587 ( .A(n_574), .Y(n_587) );
INVx3_ASAP7_75t_L g639 ( .A(n_574), .Y(n_639) );
OR2x2_ASAP7_75t_L g667 ( .A(n_574), .B(n_668), .Y(n_667) );
AOI311xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .A3(n_582), .B(n_583), .C(n_594), .Y(n_576) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_577), .A2(n_615), .B(n_617), .C(n_619), .Y(n_614) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_SL g599 ( .A(n_579), .Y(n_599) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g617 ( .A(n_581), .B(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_581), .B(n_597), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g750 ( .A(n_581), .B(n_582), .Y(n_750) );
AND2x2_ASAP7_75t_L g672 ( .A(n_582), .B(n_586), .Y(n_672) );
AOI21xp33_ASAP7_75t_L g583 ( .A1(n_584), .A2(n_588), .B(n_589), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g730 ( .A(n_586), .B(n_618), .Y(n_730) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NOR2xp33_ASAP7_75t_L g603 ( .A(n_587), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g624 ( .A(n_587), .Y(n_624) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_593), .Y(n_590) );
AND2x2_ASAP7_75t_L g615 ( .A(n_591), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g660 ( .A(n_593), .Y(n_660) );
AND2x4_ASAP7_75t_L g722 ( .A(n_593), .B(n_691), .Y(n_722) );
INVx1_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
AOI222xp33_ASAP7_75t_L g673 ( .A1(n_596), .A2(n_662), .B1(n_674), .B2(n_678), .C1(n_680), .C2(n_684), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_602), .C(n_605), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_599), .B(n_643), .Y(n_666) );
INVx1_ASAP7_75t_L g688 ( .A(n_601), .Y(n_688) );
INVx1_ASAP7_75t_L g622 ( .A(n_603), .Y(n_622) );
OR2x2_ASAP7_75t_L g687 ( .A(n_604), .B(n_688), .Y(n_687) );
OAI21xp33_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_608), .B(n_612), .Y(n_605) );
NAND3xp33_ASAP7_75t_L g623 ( .A(n_606), .B(n_624), .C(n_625), .Y(n_623) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_606), .A2(n_643), .B(n_722), .Y(n_721) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
INVx1_ASAP7_75t_SL g608 ( .A(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_610), .Y(n_663) );
AND2x2_ASAP7_75t_SL g629 ( .A(n_611), .B(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g720 ( .A(n_611), .Y(n_720) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_611), .Y(n_736) );
INVx2_ASAP7_75t_L g694 ( .A(n_612), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_616), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g668 ( .A(n_618), .Y(n_668) );
OAI221xp5_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_622), .B1(n_623), .B2(n_627), .C(n_628), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_622), .B(n_702), .Y(n_701) );
INVx1_ASAP7_75t_SL g756 ( .A(n_622), .Y(n_756) );
INVx1_ASAP7_75t_L g625 ( .A(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g637 ( .A(n_629), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_629), .B(n_660), .Y(n_659) );
AND2x2_ASAP7_75t_L g695 ( .A(n_629), .B(n_643), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_629), .B(n_705), .Y(n_704) );
AND2x2_ASAP7_75t_L g728 ( .A(n_629), .B(n_663), .Y(n_728) );
BUFx3_ASAP7_75t_L g691 ( .A(n_630), .Y(n_691) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
NAND5xp2_ASAP7_75t_L g633 ( .A(n_634), .B(n_652), .C(n_673), .D(n_685), .E(n_700), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
AOI32xp33_ASAP7_75t_L g725 ( .A1(n_637), .A2(n_664), .A3(n_680), .B1(n_726), .B2(n_728), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_639), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_643), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
INVx1_ASAP7_75t_SL g649 ( .A(n_643), .Y(n_649) );
OAI22xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_647), .B1(n_649), .B2(n_650), .Y(n_644) );
INVx1_ASAP7_75t_L g647 ( .A(n_648), .Y(n_647) );
INVx1_ASAP7_75t_SL g650 ( .A(n_651), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_659), .B1(n_661), .B2(n_662), .C(n_665), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
OR2x2_ASAP7_75t_L g654 ( .A(n_655), .B(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g724 ( .A(n_656), .B(n_675), .Y(n_724) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g739 ( .A1(n_661), .A2(n_722), .B1(n_740), .B2(n_745), .C(n_746), .Y(n_739) );
AND2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
INVx2_ASAP7_75t_L g705 ( .A(n_664), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_667), .B1(n_669), .B2(n_671), .Y(n_665) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_677), .Y(n_674) );
INVx1_ASAP7_75t_L g683 ( .A(n_675), .Y(n_683) );
INVx1_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AOI222xp33_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_689), .B1(n_693), .B2(n_694), .C1(n_695), .C2(n_696), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_692), .Y(n_689) );
INVxp67_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
OAI22xp33_ASAP7_75t_L g740 ( .A1(n_694), .A2(n_741), .B1(n_743), .B2(n_744), .Y(n_740) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g698 ( .A(n_699), .Y(n_698) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_703), .B(n_706), .Y(n_700) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_711), .B(n_713), .Y(n_706) );
INVx2_ASAP7_75t_SL g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g754 ( .A(n_709), .Y(n_754) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_721), .B(n_723), .C(n_725), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_730), .A2(n_731), .B(n_733), .C(n_758), .Y(n_729) );
CKINVDCx16_ASAP7_75t_R g734 ( .A(n_730), .Y(n_734) );
INVxp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
OAI211xp5_ASAP7_75t_L g733 ( .A1(n_734), .A2(n_735), .B(n_739), .C(n_751), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_737), .Y(n_735) );
AOI21xp33_ASAP7_75t_L g746 ( .A1(n_747), .A2(n_749), .B(n_750), .Y(n_746) );
AOI22xp5_ASAP7_75t_L g751 ( .A1(n_752), .A2(n_755), .B1(n_756), .B2(n_757), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
AOI21xp33_ASAP7_75t_L g758 ( .A1(n_759), .A2(n_760), .B(n_762), .Y(n_758) );
INVx1_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g768 ( .A(n_765), .Y(n_768) );
INVx1_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx2_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
endmodule