module fake_jpeg_6086_n_293 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_293);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_293;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_259;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_155;
wire n_82;
wire n_258;
wire n_282;
wire n_96;

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx2_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_12),
.Y(n_24)
);

BUFx12_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx5_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_39),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_42),
.B(n_49),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.C(n_1),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_43),
.B(n_5),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_18),
.B(n_1),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_44),
.B(n_5),
.Y(n_97)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx5_ASAP7_75t_L g76 ( 
.A(n_45),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_20),
.B(n_2),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_48),
.B(n_52),
.Y(n_85)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_25),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_55),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_24),
.B(n_3),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_53),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_22),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_22),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_24),
.B(n_3),
.Y(n_58)
);

AOI21xp33_ASAP7_75t_L g62 ( 
.A1(n_58),
.A2(n_25),
.B(n_29),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_36),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_59),
.A2(n_60),
.B1(n_66),
.B2(n_75),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_36),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_50),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_64),
.Y(n_106)
);

A2O1A1Ixp33_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_103),
.B(n_89),
.C(n_100),
.Y(n_123)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVx3_ASAP7_75t_SL g65 ( 
.A(n_40),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g124 ( 
.A(n_65),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_51),
.A2(n_23),
.B1(n_35),
.B2(n_18),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_48),
.B(n_34),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g133 ( 
.A(n_69),
.B(n_72),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_83),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_34),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_78),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_23),
.B1(n_35),
.B2(n_32),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_58),
.B(n_26),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_77),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_80),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g80 ( 
.A(n_44),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_40),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_81),
.B(n_97),
.Y(n_116)
);

OR2x2_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_19),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_39),
.Y(n_84)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_84),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_43),
.B(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_41),
.B(n_32),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_47),
.A2(n_30),
.B1(n_21),
.B2(n_19),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_29),
.C(n_57),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_41),
.B(n_30),
.Y(n_90)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_21),
.Y(n_92)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_46),
.B(n_38),
.Y(n_93)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_54),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_98),
.B(n_102),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_38),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_99),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_42),
.B(n_6),
.Y(n_100)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

HAxp5_ASAP7_75t_SL g103 ( 
.A(n_53),
.B(n_31),
.CON(n_103),
.SN(n_103)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_63),
.A2(n_81),
.B1(n_101),
.B2(n_103),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_107),
.A2(n_125),
.B1(n_64),
.B2(n_73),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_109),
.B(n_118),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_111),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_101),
.Y(n_112)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_112),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_76),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_88),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_131),
.Y(n_151)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

INVxp33_ASAP7_75t_L g160 ( 
.A(n_120),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_83),
.A2(n_53),
.B1(n_39),
.B2(n_25),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_122),
.A2(n_29),
.B1(n_84),
.B2(n_96),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_123),
.B(n_129),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_63),
.A2(n_39),
.B1(n_7),
.B2(n_8),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_57),
.C(n_56),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_130),
.B(n_96),
.C(n_91),
.Y(n_145)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_85),
.B(n_6),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_134),
.B(n_80),
.Y(n_137)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_94),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_91),
.Y(n_157)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_136),
.B(n_138),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_137),
.B(n_126),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_79),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_139),
.B(n_140),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_132),
.B(n_78),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_98),
.B1(n_102),
.B2(n_70),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_141),
.A2(n_142),
.B1(n_167),
.B2(n_163),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_129),
.A2(n_70),
.B1(n_67),
.B2(n_68),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_146),
.Y(n_181)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_155),
.Y(n_187)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_114),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_123),
.B(n_115),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_150),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_115),
.B(n_7),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_152),
.B(n_154),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_84),
.C(n_74),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_161),
.C(n_108),
.Y(n_185)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_111),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_157),
.Y(n_196)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_124),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_158),
.B(n_159),
.Y(n_197)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_106),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_122),
.B(n_74),
.C(n_71),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_162),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_115),
.B(n_8),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_165),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_112),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_128),
.B(n_8),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_128),
.B(n_9),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_166),
.B(n_112),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_127),
.A2(n_71),
.B1(n_82),
.B2(n_29),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_133),
.B(n_82),
.Y(n_168)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_168),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_120),
.B(n_109),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_169),
.B(n_170),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_151),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_147),
.A2(n_127),
.B1(n_118),
.B2(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_139),
.B(n_134),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_178),
.B(n_180),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_140),
.A2(n_105),
.B(n_121),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_179),
.A2(n_199),
.B(n_154),
.Y(n_210)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_105),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_183),
.Y(n_211)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_185),
.B(n_186),
.C(n_104),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_108),
.C(n_131),
.Y(n_186)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_188),
.B(n_189),
.Y(n_218)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g200 ( 
.A1(n_190),
.A2(n_198),
.B1(n_158),
.B2(n_143),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_141),
.A2(n_147),
.B1(n_161),
.B2(n_142),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_192),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_150),
.B(n_16),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_193),
.B(n_9),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_137),
.B(n_9),
.Y(n_194)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_147),
.B(n_135),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_195),
.B(n_160),
.Y(n_201)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_165),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_166),
.B(n_112),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_L g239 ( 
.A1(n_200),
.A2(n_196),
.B1(n_188),
.B2(n_189),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_201),
.B(n_217),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_179),
.B(n_160),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_202),
.B(n_212),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_208),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_207),
.B(n_222),
.C(n_186),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_156),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_197),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_216),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_210),
.A2(n_169),
.B(n_177),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_172),
.Y(n_216)
);

INVxp67_ASAP7_75t_SL g217 ( 
.A(n_176),
.Y(n_217)
);

INVx6_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_219),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_175),
.B(n_104),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_220),
.B(n_221),
.Y(n_230)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_181),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_185),
.B(n_148),
.C(n_156),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_218),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_223),
.B(n_240),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_226),
.B(n_228),
.C(n_231),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_207),
.B(n_195),
.C(n_192),
.Y(n_228)
);

OAI21xp33_ASAP7_75t_L g229 ( 
.A1(n_213),
.A2(n_174),
.B(n_171),
.Y(n_229)
);

AOI321xp33_ASAP7_75t_L g248 ( 
.A1(n_229),
.A2(n_237),
.A3(n_205),
.B1(n_169),
.B2(n_199),
.C(n_203),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_213),
.B(n_174),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_211),
.A2(n_187),
.B1(n_184),
.B2(n_183),
.Y(n_232)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_232),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_187),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_233),
.B(n_235),
.C(n_236),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_187),
.C(n_182),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_216),
.B(n_211),
.C(n_219),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_177),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_198),
.C(n_173),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_239),
.A2(n_199),
.B1(n_215),
.B2(n_212),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_218),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_206),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_242),
.B(n_253),
.C(n_234),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_243),
.B(n_252),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_205),
.B(n_206),
.Y(n_245)
);

OAI21xp5_ASAP7_75t_SL g263 ( 
.A1(n_245),
.A2(n_248),
.B(n_255),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_230),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_250),
.B(n_251),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_236),
.Y(n_252)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_241),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_254),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_173),
.Y(n_255)
);

OA21x2_ASAP7_75t_SL g256 ( 
.A1(n_253),
.A2(n_229),
.B(n_238),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g269 ( 
.A(n_256),
.B(n_242),
.Y(n_269)
);

NAND4xp25_ASAP7_75t_SL g258 ( 
.A(n_244),
.B(n_224),
.C(n_148),
.D(n_221),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_258),
.B(n_259),
.Y(n_267)
);

NOR3xp33_ASAP7_75t_SL g259 ( 
.A(n_248),
.B(n_180),
.C(n_232),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_249),
.A2(n_224),
.B1(n_228),
.B2(n_235),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_260),
.B(n_264),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_249),
.A2(n_226),
.B1(n_214),
.B2(n_234),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_247),
.C(n_246),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_214),
.B1(n_193),
.B2(n_204),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_266),
.A2(n_247),
.B1(n_246),
.B2(n_255),
.Y(n_268)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_268),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_269),
.B(n_273),
.Y(n_282)
);

NAND2xp33_ASAP7_75t_SL g270 ( 
.A(n_263),
.B(n_251),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_270),
.A2(n_263),
.B1(n_259),
.B2(n_257),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_272),
.B(n_275),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_261),
.B(n_10),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_257),
.B(n_10),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g280 ( 
.A(n_274),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_10),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_13),
.C(n_282),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_258),
.B1(n_265),
.B2(n_260),
.Y(n_278)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_L g281 ( 
.A1(n_267),
.A2(n_264),
.B1(n_266),
.B2(n_11),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_281),
.B(n_13),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_280),
.B(n_271),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_283),
.A2(n_284),
.B(n_285),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_272),
.C(n_13),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g288 ( 
.A(n_286),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_287),
.B(n_277),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_290),
.B(n_276),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_291),
.B(n_292),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_289),
.B(n_280),
.C(n_288),
.Y(n_292)
);


endmodule