module fake_netlist_6_679_n_1778 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1778);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1778;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_851;
wire n_682;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_653;
wire n_236;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_73),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_15),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_144),
.Y(n_184)
);

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_101),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_166),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_180),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g188 ( 
.A(n_140),
.Y(n_188)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_64),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_176),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_118),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_108),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g193 ( 
.A(n_94),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_104),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_113),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_63),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_161),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_17),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_89),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_170),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_122),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_0),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_171),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_81),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_175),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_121),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_39),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_22),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_103),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_105),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_42),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_92),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_138),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_47),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_84),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_32),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_87),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_78),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_165),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_120),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_117),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_152),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_2),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_44),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_134),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_116),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_46),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_4),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_169),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_115),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_26),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_4),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_114),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_160),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_177),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_71),
.Y(n_237)
);

BUFx3_ASAP7_75t_L g238 ( 
.A(n_10),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_8),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_125),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_159),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_96),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_21),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_74),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_86),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_45),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_34),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_135),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_52),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_127),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_34),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_148),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_150),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_155),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_45),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_136),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_44),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_146),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_131),
.Y(n_261)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_124),
.Y(n_262)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g264 ( 
.A(n_130),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_1),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_99),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_76),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_47),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_8),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_145),
.Y(n_270)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_31),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_68),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_137),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_154),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_69),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_14),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_49),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_9),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_133),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_26),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_65),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_35),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_126),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_67),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_110),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_88),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_141),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_147),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_57),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_173),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_59),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_28),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_72),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_5),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_95),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_40),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_33),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_5),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_27),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_56),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_21),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_28),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_168),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_70),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_111),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_102),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_3),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_56),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_128),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_109),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_178),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_93),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_157),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_142),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_2),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_85),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_12),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_52),
.Y(n_318)
);

INVx1_ASAP7_75t_SL g319 ( 
.A(n_48),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_167),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_42),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_181),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_158),
.Y(n_323)
);

BUFx10_ASAP7_75t_L g324 ( 
.A(n_112),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_49),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_164),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_106),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_61),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_66),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_97),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_43),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_107),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_13),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_60),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_11),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_91),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_77),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_172),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_46),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_129),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_149),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_0),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_33),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_10),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_132),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_6),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_22),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_14),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_100),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_143),
.Y(n_350)
);

INVx1_ASAP7_75t_SL g351 ( 
.A(n_1),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_30),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_38),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_31),
.Y(n_354)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_139),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_39),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_51),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_90),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_98),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_6),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_83),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_80),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_27),
.Y(n_363)
);

BUFx2_ASAP7_75t_L g364 ( 
.A(n_119),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_50),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_23),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_43),
.Y(n_367)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_23),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_198),
.Y(n_369)
);

INVx2_ASAP7_75t_L g370 ( 
.A(n_263),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_198),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_214),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_187),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_263),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_225),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_263),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_183),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_238),
.Y(n_378)
);

INVxp67_ASAP7_75t_SL g379 ( 
.A(n_258),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_207),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_198),
.Y(n_382)
);

INVxp67_ASAP7_75t_SL g383 ( 
.A(n_188),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_229),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_297),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_206),
.Y(n_386)
);

INVxp67_ASAP7_75t_SL g387 ( 
.A(n_345),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_242),
.Y(n_388)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_198),
.Y(n_390)
);

INVxp33_ASAP7_75t_SL g391 ( 
.A(n_207),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_198),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_240),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_264),
.Y(n_394)
);

INVxp67_ASAP7_75t_SL g395 ( 
.A(n_364),
.Y(n_395)
);

BUFx3_ASAP7_75t_L g396 ( 
.A(n_324),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_355),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_240),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_240),
.Y(n_399)
);

INVxp33_ASAP7_75t_L g400 ( 
.A(n_202),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_312),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_238),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_196),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_271),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_200),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_271),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_240),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g408 ( 
.A(n_240),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_232),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_298),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_298),
.Y(n_411)
);

INVxp33_ASAP7_75t_SL g412 ( 
.A(n_208),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_298),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_298),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_233),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_298),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_368),
.Y(n_417)
);

CKINVDCx20_ASAP7_75t_R g418 ( 
.A(n_316),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_368),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_244),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_368),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_368),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_368),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_265),
.Y(n_424)
);

CKINVDCx16_ASAP7_75t_R g425 ( 
.A(n_204),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_211),
.Y(n_426)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_297),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_217),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_224),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_239),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_193),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_194),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_248),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_259),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_265),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_208),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_334),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_210),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_278),
.Y(n_439)
);

CKINVDCx20_ASAP7_75t_R g440 ( 
.A(n_212),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_278),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_315),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_315),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_213),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_268),
.Y(n_445)
);

INVxp33_ASAP7_75t_SL g446 ( 
.A(n_343),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_276),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_216),
.Y(n_448)
);

BUFx3_ASAP7_75t_L g449 ( 
.A(n_324),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_277),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_247),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_280),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_220),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_289),
.Y(n_454)
);

CKINVDCx16_ASAP7_75t_R g455 ( 
.A(n_324),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_302),
.Y(n_456)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_343),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_321),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_333),
.Y(n_459)
);

CKINVDCx20_ASAP7_75t_R g460 ( 
.A(n_221),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_296),
.Y(n_461)
);

CKINVDCx14_ASAP7_75t_R g462 ( 
.A(n_182),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_344),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_369),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_369),
.Y(n_465)
);

BUFx6f_ASAP7_75t_L g466 ( 
.A(n_403),
.Y(n_466)
);

INVx2_ASAP7_75t_L g467 ( 
.A(n_393),
.Y(n_467)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_403),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_371),
.Y(n_469)
);

INVx3_ASAP7_75t_L g470 ( 
.A(n_403),
.Y(n_470)
);

BUFx6f_ASAP7_75t_L g471 ( 
.A(n_403),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g472 ( 
.A(n_398),
.B(n_306),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_371),
.Y(n_473)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_373),
.Y(n_474)
);

INVxp67_ASAP7_75t_L g475 ( 
.A(n_380),
.Y(n_475)
);

BUFx6f_ASAP7_75t_L g476 ( 
.A(n_403),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_393),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_382),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g479 ( 
.A(n_386),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_382),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_438),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_390),
.Y(n_482)
);

BUFx6f_ASAP7_75t_L g483 ( 
.A(n_390),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_392),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_392),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_399),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_399),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_R g488 ( 
.A(n_462),
.B(n_222),
.Y(n_488)
);

INVx3_ASAP7_75t_L g489 ( 
.A(n_431),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_408),
.Y(n_490)
);

CKINVDCx20_ASAP7_75t_R g491 ( 
.A(n_388),
.Y(n_491)
);

BUFx12f_ASAP7_75t_L g492 ( 
.A(n_372),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_383),
.B(n_306),
.Y(n_493)
);

BUFx6f_ASAP7_75t_L g494 ( 
.A(n_370),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_410),
.Y(n_496)
);

AND2x4_ASAP7_75t_L g497 ( 
.A(n_370),
.B(n_189),
.Y(n_497)
);

INVx2_ASAP7_75t_L g498 ( 
.A(n_411),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_413),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_432),
.B(n_182),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_414),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_416),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_417),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_419),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_440),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_374),
.B(n_376),
.Y(n_506)
);

AND2x2_ASAP7_75t_L g507 ( 
.A(n_378),
.B(n_189),
.Y(n_507)
);

INVx2_ASAP7_75t_L g508 ( 
.A(n_421),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_422),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_402),
.B(n_262),
.Y(n_510)
);

NOR2xp67_ASAP7_75t_L g511 ( 
.A(n_431),
.B(n_201),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_423),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_445),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_444),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_445),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_447),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_447),
.Y(n_517)
);

AND2x4_ASAP7_75t_L g518 ( 
.A(n_404),
.B(n_262),
.Y(n_518)
);

CKINVDCx20_ASAP7_75t_R g519 ( 
.A(n_394),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_450),
.Y(n_521)
);

BUFx6f_ASAP7_75t_L g522 ( 
.A(n_424),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_406),
.B(n_267),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g524 ( 
.A(n_401),
.Y(n_524)
);

INVx3_ASAP7_75t_L g525 ( 
.A(n_424),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_452),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_452),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_435),
.Y(n_528)
);

NAND2xp5_ASAP7_75t_L g529 ( 
.A(n_397),
.B(n_184),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_463),
.B(n_184),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_454),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_454),
.Y(n_532)
);

BUFx8_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_372),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_435),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_456),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_439),
.B(n_267),
.Y(n_538)
);

NOR2x1_ASAP7_75t_L g539 ( 
.A(n_396),
.B(n_305),
.Y(n_539)
);

HB1xp67_ASAP7_75t_L g540 ( 
.A(n_461),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_458),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_439),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_498),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_489),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_488),
.B(n_405),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_490),
.B(n_425),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_529),
.B(n_455),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_489),
.Y(n_548)
);

AOI22xp33_ASAP7_75t_L g549 ( 
.A1(n_493),
.A2(n_379),
.B1(n_395),
.B2(n_387),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_SL g550 ( 
.A(n_529),
.B(n_427),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_464),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_489),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g553 ( 
.A(n_507),
.B(n_441),
.Y(n_553)
);

NOR3xp33_ASAP7_75t_L g554 ( 
.A(n_540),
.B(n_389),
.C(n_377),
.Y(n_554)
);

INVx2_ASAP7_75t_SL g555 ( 
.A(n_500),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_493),
.B(n_375),
.Y(n_556)
);

INVx2_ASAP7_75t_SL g557 ( 
.A(n_500),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_464),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_472),
.Y(n_559)
);

INVx2_ASAP7_75t_L g560 ( 
.A(n_498),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_466),
.Y(n_561)
);

BUFx3_ASAP7_75t_L g562 ( 
.A(n_490),
.Y(n_562)
);

OR2x6_ASAP7_75t_L g563 ( 
.A(n_492),
.B(n_305),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_466),
.Y(n_564)
);

OAI22xp33_ASAP7_75t_L g565 ( 
.A1(n_475),
.A2(n_351),
.B1(n_319),
.B2(n_253),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_465),
.Y(n_566)
);

INVx2_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_465),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_475),
.B(n_375),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_469),
.Y(n_570)
);

INVx3_ASAP7_75t_L g571 ( 
.A(n_466),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_469),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_SL g573 ( 
.A(n_534),
.B(n_381),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_499),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_473),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_481),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_499),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_499),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_473),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_502),
.Y(n_580)
);

NAND2xp33_ASAP7_75t_SL g581 ( 
.A(n_540),
.B(n_381),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_502),
.Y(n_582)
);

OAI22xp33_ASAP7_75t_L g583 ( 
.A1(n_530),
.A2(n_257),
.B1(n_269),
.B2(n_251),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_502),
.Y(n_584)
);

NOR2x1p5_ASAP7_75t_L g585 ( 
.A(n_492),
.B(n_396),
.Y(n_585)
);

INVx2_ASAP7_75t_SL g586 ( 
.A(n_472),
.Y(n_586)
);

CKINVDCx6p67_ASAP7_75t_R g587 ( 
.A(n_492),
.Y(n_587)
);

BUFx3_ASAP7_75t_L g588 ( 
.A(n_468),
.Y(n_588)
);

INVx6_ASAP7_75t_L g589 ( 
.A(n_483),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_489),
.Y(n_590)
);

OAI22xp33_ASAP7_75t_L g591 ( 
.A1(n_530),
.A2(n_282),
.B1(n_335),
.B2(n_331),
.Y(n_591)
);

INVx3_ASAP7_75t_L g592 ( 
.A(n_466),
.Y(n_592)
);

INVxp33_ASAP7_75t_L g593 ( 
.A(n_534),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_467),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_507),
.B(n_436),
.Y(n_595)
);

AOI22xp33_ASAP7_75t_L g596 ( 
.A1(n_518),
.A2(n_412),
.B1(n_391),
.B2(n_446),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_467),
.Y(n_597)
);

BUFx2_ASAP7_75t_L g598 ( 
.A(n_533),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_480),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_SL g600 ( 
.A(n_539),
.B(n_384),
.Y(n_600)
);

NAND2xp33_ASAP7_75t_L g601 ( 
.A(n_539),
.B(n_384),
.Y(n_601)
);

OR2x2_ASAP7_75t_L g602 ( 
.A(n_507),
.B(n_385),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_513),
.B(n_391),
.Y(n_603)
);

INVx3_ASAP7_75t_L g604 ( 
.A(n_466),
.Y(n_604)
);

INVx1_ASAP7_75t_SL g605 ( 
.A(n_474),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_518),
.A2(n_412),
.B1(n_446),
.B2(n_457),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_480),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_477),
.Y(n_608)
);

AND2x6_ASAP7_75t_L g609 ( 
.A(n_497),
.B(n_313),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_484),
.Y(n_610)
);

CKINVDCx5p33_ASAP7_75t_R g611 ( 
.A(n_505),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_508),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_484),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_508),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_508),
.Y(n_615)
);

INVx3_ASAP7_75t_L g616 ( 
.A(n_466),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_487),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_471),
.Y(n_618)
);

INVx5_ASAP7_75t_L g619 ( 
.A(n_471),
.Y(n_619)
);

BUFx6f_ASAP7_75t_SL g620 ( 
.A(n_518),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_487),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_495),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_468),
.B(n_409),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_509),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_509),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_SL g626 ( 
.A(n_533),
.B(n_409),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_506),
.B(n_313),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_533),
.B(n_415),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_495),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_510),
.Y(n_630)
);

BUFx3_ASAP7_75t_L g631 ( 
.A(n_468),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_509),
.Y(n_632)
);

INVx3_ASAP7_75t_L g633 ( 
.A(n_471),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_512),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_471),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_512),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_496),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_512),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_496),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_477),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_470),
.B(n_415),
.Y(n_641)
);

INVx2_ASAP7_75t_L g642 ( 
.A(n_477),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_471),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_470),
.B(n_420),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_514),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_501),
.Y(n_646)
);

AO21x2_ASAP7_75t_L g647 ( 
.A1(n_511),
.A2(n_218),
.B(n_215),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_470),
.B(n_420),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_478),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_470),
.B(n_451),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_510),
.B(n_441),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_501),
.B(n_451),
.Y(n_652)
);

NOR2xp33_ASAP7_75t_L g653 ( 
.A(n_513),
.B(n_457),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_503),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_503),
.B(n_449),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_533),
.B(n_448),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_471),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_478),
.Y(n_658)
);

INVx5_ASAP7_75t_L g659 ( 
.A(n_476),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_504),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_515),
.B(n_453),
.Y(n_661)
);

INVx4_ASAP7_75t_L g662 ( 
.A(n_483),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_504),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_SL g664 ( 
.A(n_518),
.B(n_460),
.Y(n_664)
);

BUFx10_ASAP7_75t_L g665 ( 
.A(n_506),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_482),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_506),
.B(n_449),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_506),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_497),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_482),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_497),
.Y(n_671)
);

NAND3xp33_ASAP7_75t_L g672 ( 
.A(n_510),
.B(n_428),
.C(n_426),
.Y(n_672)
);

NOR2xp33_ASAP7_75t_L g673 ( 
.A(n_516),
.B(n_400),
.Y(n_673)
);

HB1xp67_ASAP7_75t_L g674 ( 
.A(n_523),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_SL g675 ( 
.A(n_523),
.B(n_185),
.Y(n_675)
);

AOI22xp33_ASAP7_75t_L g676 ( 
.A1(n_523),
.A2(n_365),
.B1(n_352),
.B2(n_348),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_482),
.Y(n_677)
);

AND2x2_ASAP7_75t_SL g678 ( 
.A(n_538),
.B(n_329),
.Y(n_678)
);

INVx2_ASAP7_75t_SL g679 ( 
.A(n_538),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_485),
.Y(n_680)
);

NOR2xp33_ASAP7_75t_L g681 ( 
.A(n_516),
.B(n_418),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_486),
.Y(n_682)
);

AO21x2_ASAP7_75t_L g683 ( 
.A1(n_511),
.A2(n_231),
.B(n_219),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_517),
.B(n_437),
.Y(n_684)
);

OR2x6_ASAP7_75t_L g685 ( 
.A(n_517),
.B(n_329),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_486),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_555),
.B(n_494),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_555),
.B(n_185),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_L g689 ( 
.A(n_557),
.B(n_494),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_557),
.A2(n_349),
.B1(n_284),
.B2(n_273),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_595),
.Y(n_691)
);

INVx2_ASAP7_75t_SL g692 ( 
.A(n_595),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_669),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_602),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_559),
.B(n_186),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_559),
.A2(n_347),
.B1(n_366),
.B2(n_363),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_SL g697 ( 
.A(n_586),
.B(n_186),
.Y(n_697)
);

BUFx4f_ASAP7_75t_L g698 ( 
.A(n_587),
.Y(n_698)
);

AOI22xp5_ASAP7_75t_L g699 ( 
.A1(n_678),
.A2(n_341),
.B1(n_303),
.B2(n_291),
.Y(n_699)
);

AND2x2_ASAP7_75t_L g700 ( 
.A(n_673),
.B(n_520),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_L g701 ( 
.A(n_586),
.B(n_190),
.Y(n_701)
);

NAND3xp33_ASAP7_75t_L g702 ( 
.A(n_549),
.B(n_294),
.C(n_292),
.Y(n_702)
);

AOI22xp5_ASAP7_75t_L g703 ( 
.A1(n_678),
.A2(n_630),
.B1(n_679),
.B2(n_668),
.Y(n_703)
);

A2O1A1Ixp33_ASAP7_75t_L g704 ( 
.A1(n_679),
.A2(n_330),
.B(n_249),
.C(n_255),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_661),
.B(n_603),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_669),
.Y(n_706)
);

O2A1O1Ixp33_ASAP7_75t_L g707 ( 
.A1(n_674),
.A2(n_526),
.B(n_541),
.C(n_537),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_544),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_653),
.B(n_191),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_671),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_SL g711 ( 
.A(n_583),
.B(n_191),
.Y(n_711)
);

INVx5_ASAP7_75t_L g712 ( 
.A(n_609),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_576),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_562),
.B(n_494),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_562),
.B(n_525),
.Y(n_715)
);

INVx4_ASAP7_75t_L g716 ( 
.A(n_665),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_556),
.B(n_192),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_665),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_609),
.A2(n_330),
.B1(n_196),
.B2(n_283),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_611),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_652),
.B(n_192),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_593),
.B(n_520),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_665),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_562),
.B(n_525),
.Y(n_724)
);

BUFx4_ASAP7_75t_L g725 ( 
.A(n_587),
.Y(n_725)
);

NOR2xp33_ASAP7_75t_L g726 ( 
.A(n_602),
.B(n_195),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_SL g727 ( 
.A(n_591),
.B(n_195),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_547),
.B(n_197),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_SL g729 ( 
.A(n_596),
.B(n_197),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_L g730 ( 
.A1(n_609),
.A2(n_283),
.B1(n_196),
.B2(n_193),
.Y(n_730)
);

NOR2xp33_ASAP7_75t_L g731 ( 
.A(n_550),
.B(n_199),
.Y(n_731)
);

OAI221xp5_ASAP7_75t_L g732 ( 
.A1(n_676),
.A2(n_531),
.B1(n_541),
.B2(n_537),
.C(n_536),
.Y(n_732)
);

OR2x6_ASAP7_75t_L g733 ( 
.A(n_598),
.B(n_429),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_L g734 ( 
.A(n_546),
.B(n_199),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_681),
.B(n_521),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_553),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_553),
.Y(n_737)
);

AND2x2_ASAP7_75t_L g738 ( 
.A(n_684),
.B(n_521),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_569),
.B(n_203),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_651),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_SL g741 ( 
.A(n_606),
.B(n_203),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_551),
.A2(n_359),
.B(n_246),
.C(n_261),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_558),
.B(n_522),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_SL g744 ( 
.A(n_623),
.B(n_205),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_600),
.B(n_205),
.Y(n_745)
);

AOI22xp5_ASAP7_75t_L g746 ( 
.A1(n_601),
.A2(n_281),
.B1(n_274),
.B2(n_272),
.Y(n_746)
);

HB1xp67_ASAP7_75t_L g747 ( 
.A(n_685),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_566),
.B(n_522),
.Y(n_748)
);

O2A1O1Ixp33_ASAP7_75t_L g749 ( 
.A1(n_675),
.A2(n_527),
.B(n_536),
.C(n_526),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_548),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_568),
.B(n_522),
.Y(n_751)
);

AO22x2_ASAP7_75t_L g752 ( 
.A1(n_656),
.A2(n_234),
.B1(n_285),
.B2(n_293),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_651),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_622),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_641),
.B(n_209),
.Y(n_755)
);

A2O1A1Ixp33_ASAP7_75t_L g756 ( 
.A1(n_570),
.A2(n_295),
.B(n_309),
.C(n_337),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_570),
.B(n_522),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_572),
.B(n_575),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_629),
.Y(n_759)
);

BUFx2_ASAP7_75t_L g760 ( 
.A(n_581),
.Y(n_760)
);

INVxp67_ASAP7_75t_SL g761 ( 
.A(n_572),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_554),
.B(n_527),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_579),
.B(n_528),
.Y(n_763)
);

INVx4_ASAP7_75t_L g764 ( 
.A(n_665),
.Y(n_764)
);

BUFx5_ASAP7_75t_L g765 ( 
.A(n_609),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_645),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_548),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_609),
.B(n_193),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_644),
.B(n_209),
.Y(n_769)
);

NOR2xp33_ASAP7_75t_L g770 ( 
.A(n_648),
.B(n_350),
.Y(n_770)
);

AND2x2_ASAP7_75t_SL g771 ( 
.A(n_598),
.B(n_196),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_629),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_637),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_672),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_650),
.B(n_664),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_599),
.B(n_350),
.Y(n_776)
);

OAI22xp5_ASAP7_75t_L g777 ( 
.A1(n_685),
.A2(n_310),
.B1(n_311),
.B2(n_358),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_599),
.B(n_528),
.Y(n_778)
);

NOR2xp33_ASAP7_75t_L g779 ( 
.A(n_607),
.B(n_361),
.Y(n_779)
);

NAND2xp33_ASAP7_75t_L g780 ( 
.A(n_609),
.B(n_193),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_607),
.B(n_361),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_610),
.B(n_613),
.Y(n_782)
);

AOI22xp5_ASAP7_75t_L g783 ( 
.A1(n_620),
.A2(n_260),
.B1(n_235),
.B2(n_230),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_552),
.Y(n_784)
);

NOR2xp67_ASAP7_75t_L g785 ( 
.A(n_672),
.B(n_531),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_610),
.B(n_528),
.Y(n_786)
);

NOR2xp67_ASAP7_75t_L g787 ( 
.A(n_545),
.B(n_532),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_639),
.Y(n_788)
);

OAI22xp33_ASAP7_75t_L g789 ( 
.A1(n_685),
.A2(n_354),
.B1(n_346),
.B2(n_347),
.Y(n_789)
);

AOI22xp5_ASAP7_75t_L g790 ( 
.A1(n_620),
.A2(n_627),
.B1(n_667),
.B2(n_573),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_655),
.B(n_532),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_552),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_613),
.B(n_362),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_590),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_646),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_590),
.Y(n_796)
);

INVx2_ASAP7_75t_L g797 ( 
.A(n_594),
.Y(n_797)
);

OR2x6_ASAP7_75t_L g798 ( 
.A(n_563),
.B(n_430),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_617),
.B(n_528),
.Y(n_799)
);

CKINVDCx20_ASAP7_75t_R g800 ( 
.A(n_605),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_617),
.B(n_362),
.Y(n_801)
);

INVx2_ASAP7_75t_L g802 ( 
.A(n_594),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_563),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_597),
.Y(n_804)
);

INVx1_ASAP7_75t_L g805 ( 
.A(n_654),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_654),
.Y(n_806)
);

BUFx3_ASAP7_75t_L g807 ( 
.A(n_660),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_660),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_663),
.Y(n_809)
);

AND2x4_ASAP7_75t_L g810 ( 
.A(n_627),
.B(n_433),
.Y(n_810)
);

OAI22xp5_ASAP7_75t_L g811 ( 
.A1(n_685),
.A2(n_254),
.B1(n_250),
.B2(n_245),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_597),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_621),
.B(n_528),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_663),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_620),
.A2(n_256),
.B1(n_223),
.B2(n_226),
.Y(n_815)
);

INVxp33_ASAP7_75t_L g816 ( 
.A(n_626),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_588),
.B(n_483),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_565),
.B(n_227),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_563),
.B(n_434),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_588),
.Y(n_820)
);

INVxp67_ASAP7_75t_SL g821 ( 
.A(n_666),
.Y(n_821)
);

INVx1_ASAP7_75t_SL g822 ( 
.A(n_628),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_631),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_627),
.B(n_299),
.Y(n_824)
);

BUFx2_ASAP7_75t_R g825 ( 
.A(n_647),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_631),
.B(n_483),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_643),
.B(n_236),
.Y(n_827)
);

AND3x2_ASAP7_75t_SL g828 ( 
.A(n_825),
.B(n_353),
.C(n_346),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_693),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_706),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_807),
.B(n_563),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_738),
.B(n_585),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_710),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_761),
.B(n_627),
.Y(n_834)
);

OR2x2_ASAP7_75t_L g835 ( 
.A(n_691),
.B(n_627),
.Y(n_835)
);

OAI21xp33_ASAP7_75t_SL g836 ( 
.A1(n_703),
.A2(n_685),
.B(n_585),
.Y(n_836)
);

AOI22xp33_ASAP7_75t_L g837 ( 
.A1(n_736),
.A2(n_683),
.B1(n_647),
.B2(n_609),
.Y(n_837)
);

A2O1A1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_782),
.A2(n_458),
.B(n_459),
.C(n_356),
.Y(n_838)
);

NAND2x1p5_ASAP7_75t_L g839 ( 
.A(n_718),
.B(n_662),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_761),
.B(n_791),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_798),
.B(n_479),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_715),
.A2(n_724),
.B(n_821),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_713),
.Y(n_843)
);

INVx2_ASAP7_75t_L g844 ( 
.A(n_797),
.Y(n_844)
);

AND2x4_ASAP7_75t_SL g845 ( 
.A(n_800),
.B(n_491),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_722),
.B(n_519),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_737),
.A2(n_683),
.B1(n_647),
.B2(n_193),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_712),
.B(n_643),
.Y(n_848)
);

INVx5_ASAP7_75t_L g849 ( 
.A(n_718),
.Y(n_849)
);

AND2x2_ASAP7_75t_L g850 ( 
.A(n_692),
.B(n_524),
.Y(n_850)
);

INVxp67_ASAP7_75t_L g851 ( 
.A(n_694),
.Y(n_851)
);

NAND3xp33_ASAP7_75t_SL g852 ( 
.A(n_705),
.B(n_354),
.C(n_353),
.Y(n_852)
);

NOR2xp33_ASAP7_75t_R g853 ( 
.A(n_720),
.B(n_237),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_754),
.Y(n_854)
);

CKINVDCx20_ASAP7_75t_R g855 ( 
.A(n_766),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_740),
.B(n_459),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_700),
.B(n_561),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_782),
.B(n_695),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_SL g859 ( 
.A(n_712),
.B(n_643),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_759),
.Y(n_860)
);

OAI21xp33_ASAP7_75t_SL g861 ( 
.A1(n_772),
.A2(n_443),
.B(n_442),
.Y(n_861)
);

AND2x4_ASAP7_75t_L g862 ( 
.A(n_753),
.B(n_442),
.Y(n_862)
);

BUFx3_ASAP7_75t_L g863 ( 
.A(n_698),
.Y(n_863)
);

CKINVDCx14_ASAP7_75t_R g864 ( 
.A(n_698),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_712),
.B(n_643),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_773),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_712),
.B(n_765),
.Y(n_867)
);

INVx4_ASAP7_75t_L g868 ( 
.A(n_718),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_775),
.A2(n_683),
.B1(n_589),
.B2(n_564),
.Y(n_869)
);

NOR2xp33_ASAP7_75t_R g870 ( 
.A(n_803),
.B(n_241),
.Y(n_870)
);

OAI22xp33_ASAP7_75t_L g871 ( 
.A1(n_774),
.A2(n_363),
.B1(n_360),
.B2(n_367),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_739),
.B(n_443),
.Y(n_872)
);

AOI22xp33_ASAP7_75t_L g873 ( 
.A1(n_730),
.A2(n_193),
.B1(n_196),
.B2(n_283),
.Y(n_873)
);

OAI22xp5_ASAP7_75t_SL g874 ( 
.A1(n_822),
.A2(n_816),
.B1(n_760),
.B2(n_739),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_695),
.B(n_561),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_701),
.B(n_561),
.Y(n_876)
);

AOI22xp5_ASAP7_75t_L g877 ( 
.A1(n_721),
.A2(n_589),
.B1(n_564),
.B2(n_604),
.Y(n_877)
);

AOI22xp33_ASAP7_75t_L g878 ( 
.A1(n_730),
.A2(n_193),
.B1(n_283),
.B2(n_574),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_701),
.B(n_561),
.Y(n_879)
);

AOI22xp33_ASAP7_75t_L g880 ( 
.A1(n_719),
.A2(n_193),
.B1(n_283),
.B2(n_615),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_765),
.B(n_718),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_SL g882 ( 
.A(n_771),
.B(n_356),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_726),
.B(n_357),
.Y(n_883)
);

OR2x2_ASAP7_75t_SL g884 ( 
.A(n_702),
.B(n_357),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_770),
.B(n_564),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_770),
.B(n_571),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_802),
.Y(n_887)
);

INVx2_ASAP7_75t_L g888 ( 
.A(n_804),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_788),
.Y(n_889)
);

A2O1A1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_774),
.A2(n_360),
.B(n_366),
.C(n_367),
.Y(n_890)
);

BUFx10_ASAP7_75t_L g891 ( 
.A(n_728),
.Y(n_891)
);

INVx5_ASAP7_75t_L g892 ( 
.A(n_723),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_812),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_820),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_795),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_726),
.B(n_300),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_762),
.Y(n_897)
);

AND2x4_ASAP7_75t_L g898 ( 
.A(n_810),
.B(n_571),
.Y(n_898)
);

CKINVDCx20_ASAP7_75t_R g899 ( 
.A(n_733),
.Y(n_899)
);

BUFx3_ASAP7_75t_L g900 ( 
.A(n_819),
.Y(n_900)
);

INVx5_ASAP7_75t_L g901 ( 
.A(n_723),
.Y(n_901)
);

INVx3_ASAP7_75t_L g902 ( 
.A(n_823),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_734),
.B(n_571),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_765),
.B(n_643),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_805),
.Y(n_905)
);

AND2x4_ASAP7_75t_L g906 ( 
.A(n_810),
.B(n_571),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_806),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_723),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_808),
.Y(n_909)
);

INVx1_ASAP7_75t_L g910 ( 
.A(n_809),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_821),
.A2(n_662),
.B(n_543),
.Y(n_911)
);

INVx5_ASAP7_75t_L g912 ( 
.A(n_723),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_814),
.Y(n_913)
);

OAI22xp5_ASAP7_75t_SL g914 ( 
.A1(n_733),
.A2(n_317),
.B1(n_301),
.B2(n_307),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_747),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_709),
.B(n_308),
.Y(n_916)
);

INVx2_ASAP7_75t_SL g917 ( 
.A(n_688),
.Y(n_917)
);

NAND2xp33_ASAP7_75t_L g918 ( 
.A(n_765),
.B(n_719),
.Y(n_918)
);

INVxp67_ASAP7_75t_L g919 ( 
.A(n_776),
.Y(n_919)
);

NOR2xp33_ASAP7_75t_L g920 ( 
.A(n_717),
.B(n_318),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_733),
.Y(n_921)
);

INVx4_ASAP7_75t_L g922 ( 
.A(n_716),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_758),
.B(n_776),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_747),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_697),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_779),
.B(n_592),
.Y(n_926)
);

NAND3xp33_ASAP7_75t_SL g927 ( 
.A(n_717),
.B(n_339),
.C(n_325),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_798),
.Y(n_928)
);

INVx2_ASAP7_75t_SL g929 ( 
.A(n_752),
.Y(n_929)
);

INVx3_ASAP7_75t_L g930 ( 
.A(n_708),
.Y(n_930)
);

OAI22xp5_ASAP7_75t_L g931 ( 
.A1(n_790),
.A2(n_689),
.B1(n_687),
.B2(n_699),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_SL g932 ( 
.A(n_765),
.B(n_604),
.Y(n_932)
);

AOI22xp5_ASAP7_75t_L g933 ( 
.A1(n_745),
.A2(n_589),
.B1(n_604),
.B2(n_616),
.Y(n_933)
);

AND2x4_ASAP7_75t_L g934 ( 
.A(n_787),
.B(n_616),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_SL g935 ( 
.A(n_765),
.B(n_616),
.Y(n_935)
);

NOR2xp33_ASAP7_75t_L g936 ( 
.A(n_731),
.B(n_618),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_798),
.B(n_618),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_750),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_767),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_716),
.Y(n_940)
);

BUFx3_ASAP7_75t_L g941 ( 
.A(n_714),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_781),
.B(n_618),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_784),
.Y(n_943)
);

NAND3xp33_ASAP7_75t_L g944 ( 
.A(n_731),
.B(n_288),
.C(n_243),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_781),
.B(n_633),
.Y(n_945)
);

AND2x4_ASAP7_75t_L g946 ( 
.A(n_785),
.B(n_764),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_792),
.Y(n_947)
);

INVx2_ASAP7_75t_SL g948 ( 
.A(n_752),
.Y(n_948)
);

AOI22xp5_ASAP7_75t_L g949 ( 
.A1(n_745),
.A2(n_824),
.B1(n_769),
.B2(n_755),
.Y(n_949)
);

INVxp67_ASAP7_75t_L g950 ( 
.A(n_793),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_743),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_748),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_SL g953 ( 
.A(n_771),
.B(n_764),
.Y(n_953)
);

AND3x1_ASAP7_75t_L g954 ( 
.A(n_690),
.B(n_535),
.C(n_542),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_794),
.Y(n_955)
);

AND2x4_ASAP7_75t_L g956 ( 
.A(n_824),
.B(n_633),
.Y(n_956)
);

BUFx3_ASAP7_75t_L g957 ( 
.A(n_732),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_751),
.Y(n_958)
);

INVx2_ASAP7_75t_SL g959 ( 
.A(n_752),
.Y(n_959)
);

CKINVDCx11_ASAP7_75t_R g960 ( 
.A(n_725),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_757),
.Y(n_961)
);

CKINVDCx5p33_ASAP7_75t_R g962 ( 
.A(n_746),
.Y(n_962)
);

AND2x4_ASAP7_75t_L g963 ( 
.A(n_744),
.B(n_635),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_SL g964 ( 
.A(n_763),
.B(n_635),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_796),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_778),
.Y(n_966)
);

INVx2_ASAP7_75t_SL g967 ( 
.A(n_818),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_801),
.B(n_635),
.Y(n_968)
);

AOI22xp33_ASAP7_75t_SL g969 ( 
.A1(n_696),
.A2(n_287),
.B1(n_340),
.B2(n_338),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_786),
.Y(n_970)
);

AOI22xp33_ASAP7_75t_L g971 ( 
.A1(n_696),
.A2(n_634),
.B1(n_560),
.B2(n_567),
.Y(n_971)
);

INVx1_ASAP7_75t_SL g972 ( 
.A(n_711),
.Y(n_972)
);

BUFx4f_ASAP7_75t_L g973 ( 
.A(n_707),
.Y(n_973)
);

AOI211xp5_ASAP7_75t_L g974 ( 
.A1(n_729),
.A2(n_279),
.B(n_252),
.C(n_266),
.Y(n_974)
);

INVx5_ASAP7_75t_L g975 ( 
.A(n_768),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_799),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_749),
.B(n_635),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_813),
.B(n_657),
.Y(n_978)
);

INVx2_ASAP7_75t_L g979 ( 
.A(n_817),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_826),
.B(n_657),
.Y(n_980)
);

BUFx6f_ASAP7_75t_L g981 ( 
.A(n_827),
.Y(n_981)
);

OAI21xp33_ASAP7_75t_L g982 ( 
.A1(n_741),
.A2(n_275),
.B(n_270),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_919),
.B(n_727),
.Y(n_983)
);

OAI22xp5_ASAP7_75t_L g984 ( 
.A1(n_858),
.A2(n_789),
.B1(n_783),
.B2(n_815),
.Y(n_984)
);

NAND2x1p5_ASAP7_75t_L g985 ( 
.A(n_849),
.B(n_662),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_SL g986 ( 
.A1(n_855),
.A2(n_777),
.B1(n_789),
.B2(n_320),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_883),
.B(n_811),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_873),
.A2(n_840),
.B1(n_923),
.B2(n_878),
.Y(n_988)
);

AOI21x1_ASAP7_75t_L g989 ( 
.A1(n_875),
.A2(n_582),
.B(n_614),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_829),
.Y(n_990)
);

INVx3_ASAP7_75t_L g991 ( 
.A(n_908),
.Y(n_991)
);

OAI21x1_ASAP7_75t_L g992 ( 
.A1(n_842),
.A2(n_911),
.B(n_932),
.Y(n_992)
);

CKINVDCx14_ASAP7_75t_R g993 ( 
.A(n_855),
.Y(n_993)
);

AND2x6_ASAP7_75t_L g994 ( 
.A(n_908),
.B(n_666),
.Y(n_994)
);

A2O1A1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_920),
.A2(n_780),
.B(n_704),
.C(n_742),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_918),
.A2(n_975),
.B(n_892),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_833),
.Y(n_997)
);

AO32x2_ASAP7_75t_L g998 ( 
.A1(n_929),
.A2(n_662),
.A3(n_756),
.B1(n_9),
.B2(n_12),
.Y(n_998)
);

AND3x1_ASAP7_75t_SL g999 ( 
.A(n_828),
.B(n_3),
.C(n_7),
.Y(n_999)
);

BUFx6f_ASAP7_75t_L g1000 ( 
.A(n_908),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_919),
.B(n_649),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_850),
.Y(n_1002)
);

O2A1O1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_920),
.A2(n_636),
.B(n_577),
.C(n_578),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_950),
.B(n_649),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_950),
.B(n_658),
.Y(n_1005)
);

INVx2_ASAP7_75t_SL g1006 ( 
.A(n_845),
.Y(n_1006)
);

AOI21xp5_ASAP7_75t_L g1007 ( 
.A1(n_918),
.A2(n_619),
.B(n_659),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_896),
.B(n_542),
.Y(n_1008)
);

AOI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_927),
.A2(n_286),
.B1(n_304),
.B2(n_314),
.Y(n_1009)
);

AOI22xp33_ASAP7_75t_L g1010 ( 
.A1(n_927),
.A2(n_290),
.B1(n_322),
.B2(n_323),
.Y(n_1010)
);

HB1xp67_ASAP7_75t_L g1011 ( 
.A(n_915),
.Y(n_1011)
);

INVx4_ASAP7_75t_L g1012 ( 
.A(n_849),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_897),
.B(n_851),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_900),
.B(n_326),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_916),
.A2(n_657),
.B(n_580),
.C(n_636),
.Y(n_1015)
);

OAI22xp5_ASAP7_75t_L g1016 ( 
.A1(n_873),
.A2(n_878),
.B1(n_957),
.B2(n_880),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_844),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_975),
.A2(n_619),
.B(n_659),
.Y(n_1018)
);

NOR2xp67_ASAP7_75t_L g1019 ( 
.A(n_843),
.B(n_327),
.Y(n_1019)
);

O2A1O1Ixp33_ASAP7_75t_L g1020 ( 
.A1(n_852),
.A2(n_638),
.B(n_578),
.C(n_582),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_852),
.B(n_328),
.C(n_332),
.Y(n_1021)
);

CKINVDCx8_ASAP7_75t_R g1022 ( 
.A(n_872),
.Y(n_1022)
);

BUFx2_ASAP7_75t_L g1023 ( 
.A(n_841),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_851),
.B(n_657),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_830),
.Y(n_1025)
);

NOR3xp33_ASAP7_75t_SL g1026 ( 
.A(n_962),
.B(n_336),
.C(n_13),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_838),
.A2(n_638),
.B(n_612),
.C(n_614),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_832),
.B(n_584),
.Y(n_1028)
);

O2A1O1Ixp33_ASAP7_75t_L g1029 ( 
.A1(n_838),
.A2(n_624),
.B(n_625),
.C(n_632),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_887),
.Y(n_1030)
);

O2A1O1Ixp5_ASAP7_75t_L g1031 ( 
.A1(n_973),
.A2(n_624),
.B(n_625),
.C(n_632),
.Y(n_1031)
);

AND2x2_ASAP7_75t_L g1032 ( 
.A(n_856),
.B(n_612),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_854),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_853),
.Y(n_1034)
);

AO32x2_ASAP7_75t_L g1035 ( 
.A1(n_948),
.A2(n_7),
.A3(n_15),
.B1(n_16),
.B2(n_18),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_849),
.B(n_659),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_SL g1037 ( 
.A(n_891),
.B(n_686),
.Y(n_1037)
);

BUFx3_ASAP7_75t_L g1038 ( 
.A(n_863),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_928),
.Y(n_1039)
);

BUFx2_ASAP7_75t_SL g1040 ( 
.A(n_849),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_860),
.B(n_682),
.Y(n_1041)
);

OR2x6_ASAP7_75t_L g1042 ( 
.A(n_841),
.B(n_682),
.Y(n_1042)
);

NOR2xp33_ASAP7_75t_L g1043 ( 
.A(n_972),
.B(n_16),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_874),
.B(n_18),
.Y(n_1044)
);

INVx3_ASAP7_75t_SL g1045 ( 
.A(n_841),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_868),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_888),
.Y(n_1047)
);

AO22x1_ASAP7_75t_L g1048 ( 
.A1(n_831),
.A2(n_19),
.B1(n_20),
.B2(n_24),
.Y(n_1048)
);

OAI22xp5_ASAP7_75t_L g1049 ( 
.A1(n_880),
.A2(n_680),
.B1(n_677),
.B2(n_670),
.Y(n_1049)
);

NAND3xp33_ASAP7_75t_L g1050 ( 
.A(n_916),
.B(n_670),
.C(n_666),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_866),
.Y(n_1051)
);

OAI22xp5_ASAP7_75t_L g1052 ( 
.A1(n_969),
.A2(n_642),
.B1(n_640),
.B2(n_608),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_893),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_836),
.A2(n_967),
.B(n_936),
.C(n_925),
.Y(n_1054)
);

A2O1A1Ixp33_ASAP7_75t_L g1055 ( 
.A1(n_936),
.A2(n_642),
.B(n_640),
.C(n_608),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_889),
.B(n_483),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_895),
.B(n_19),
.Y(n_1057)
);

NAND3xp33_ASAP7_75t_SL g1058 ( 
.A(n_974),
.B(n_24),
.C(n_25),
.Y(n_1058)
);

AND2x4_ASAP7_75t_L g1059 ( 
.A(n_937),
.B(n_62),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_901),
.A2(n_476),
.B(n_58),
.Y(n_1060)
);

INVxp33_ASAP7_75t_L g1061 ( 
.A(n_853),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_905),
.B(n_25),
.Y(n_1062)
);

BUFx3_ASAP7_75t_L g1063 ( 
.A(n_960),
.Y(n_1063)
);

AND2x2_ASAP7_75t_L g1064 ( 
.A(n_856),
.B(n_29),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_L g1065 ( 
.A(n_907),
.B(n_29),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_959),
.A2(n_30),
.B1(n_32),
.B2(n_35),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_839),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_901),
.A2(n_79),
.B(n_174),
.Y(n_1068)
);

BUFx2_ASAP7_75t_L g1069 ( 
.A(n_915),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_917),
.B(n_36),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_912),
.A2(n_75),
.B(n_162),
.Y(n_1071)
);

AOI21xp33_ASAP7_75t_L g1072 ( 
.A1(n_882),
.A2(n_36),
.B(n_37),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_912),
.A2(n_82),
.B(n_153),
.Y(n_1073)
);

O2A1O1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_890),
.A2(n_953),
.B(n_871),
.C(n_931),
.Y(n_1074)
);

AND2x4_ASAP7_75t_L g1075 ( 
.A(n_937),
.B(n_179),
.Y(n_1075)
);

OR2x6_ASAP7_75t_L g1076 ( 
.A(n_921),
.B(n_151),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_909),
.B(n_37),
.Y(n_1077)
);

BUFx3_ASAP7_75t_L g1078 ( 
.A(n_960),
.Y(n_1078)
);

AO22x1_ASAP7_75t_L g1079 ( 
.A1(n_924),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_1079)
);

O2A1O1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_890),
.A2(n_41),
.B(n_48),
.C(n_50),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_834),
.A2(n_910),
.B(n_913),
.C(n_944),
.Y(n_1081)
);

O2A1O1Ixp33_ASAP7_75t_L g1082 ( 
.A1(n_871),
.A2(n_51),
.B(n_53),
.C(n_54),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_L g1083 ( 
.A1(n_884),
.A2(n_53),
.B1(n_55),
.B2(n_57),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_SL g1084 ( 
.A(n_835),
.B(n_123),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_L g1085 ( 
.A(n_924),
.B(n_55),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_951),
.A2(n_952),
.B(n_958),
.C(n_961),
.Y(n_1086)
);

INVxp67_ASAP7_75t_L g1087 ( 
.A(n_862),
.Y(n_1087)
);

NAND3xp33_ASAP7_75t_SL g1088 ( 
.A(n_870),
.B(n_982),
.C(n_899),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_864),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_867),
.A2(n_881),
.B(n_904),
.Y(n_1090)
);

NOR2xp33_ASAP7_75t_L g1091 ( 
.A(n_914),
.B(n_857),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_966),
.B(n_970),
.Y(n_1092)
);

AOI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_867),
.A2(n_881),
.B(n_904),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_976),
.B(n_979),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_903),
.B(n_941),
.Y(n_1095)
);

NOR3xp33_ASAP7_75t_L g1096 ( 
.A(n_861),
.B(n_898),
.C(n_906),
.Y(n_1096)
);

INVxp67_ASAP7_75t_L g1097 ( 
.A(n_954),
.Y(n_1097)
);

AOI21xp5_ASAP7_75t_L g1098 ( 
.A1(n_842),
.A2(n_839),
.B(n_885),
.Y(n_1098)
);

NAND2xp5_ASAP7_75t_L g1099 ( 
.A(n_876),
.B(n_879),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_886),
.A2(n_911),
.B(n_935),
.Y(n_1100)
);

BUFx2_ASAP7_75t_L g1101 ( 
.A(n_899),
.Y(n_1101)
);

AND2x2_ASAP7_75t_L g1102 ( 
.A(n_870),
.B(n_906),
.Y(n_1102)
);

NAND2xp5_ASAP7_75t_L g1103 ( 
.A(n_1092),
.B(n_956),
.Y(n_1103)
);

AO21x2_ASAP7_75t_L g1104 ( 
.A1(n_1100),
.A2(n_945),
.B(n_942),
.Y(n_1104)
);

O2A1O1Ixp33_ASAP7_75t_SL g1105 ( 
.A1(n_1054),
.A2(n_865),
.B(n_848),
.C(n_859),
.Y(n_1105)
);

AOI221x1_ASAP7_75t_L g1106 ( 
.A1(n_984),
.A2(n_1044),
.B1(n_1058),
.B2(n_1083),
.C(n_1072),
.Y(n_1106)
);

AOI221xp5_ASAP7_75t_SL g1107 ( 
.A1(n_984),
.A2(n_971),
.B1(n_847),
.B2(n_968),
.C(n_926),
.Y(n_1107)
);

AND2x4_ASAP7_75t_L g1108 ( 
.A(n_1102),
.B(n_898),
.Y(n_1108)
);

AOI211x1_ASAP7_75t_L g1109 ( 
.A1(n_1083),
.A2(n_977),
.B(n_828),
.C(n_964),
.Y(n_1109)
);

INVxp67_ASAP7_75t_SL g1110 ( 
.A(n_1011),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1091),
.A2(n_963),
.B1(n_946),
.B2(n_981),
.Y(n_1111)
);

INVxp67_ASAP7_75t_SL g1112 ( 
.A(n_1016),
.Y(n_1112)
);

NAND3xp33_ASAP7_75t_L g1113 ( 
.A(n_983),
.B(n_981),
.C(n_847),
.Y(n_1113)
);

INVx5_ASAP7_75t_L g1114 ( 
.A(n_994),
.Y(n_1114)
);

NAND2xp5_ASAP7_75t_SL g1115 ( 
.A(n_1002),
.B(n_981),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_990),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1025),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1015),
.A2(n_980),
.A3(n_978),
.B(n_938),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_1002),
.B(n_963),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_1092),
.B(n_894),
.Y(n_1120)
);

AOI221x1_ASAP7_75t_L g1121 ( 
.A1(n_1072),
.A2(n_1021),
.B1(n_988),
.B2(n_1066),
.C(n_995),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_1090),
.A2(n_1093),
.B(n_989),
.Y(n_1122)
);

BUFx10_ASAP7_75t_L g1123 ( 
.A(n_1013),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_1031),
.A2(n_902),
.B(n_837),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_1033),
.Y(n_1125)
);

OAI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1055),
.A2(n_869),
.B(n_837),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1016),
.A2(n_971),
.B1(n_922),
.B2(n_940),
.Y(n_1127)
);

AOI21x1_ASAP7_75t_L g1128 ( 
.A1(n_1095),
.A2(n_934),
.B(n_965),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1051),
.Y(n_1129)
);

INVx2_ASAP7_75t_SL g1130 ( 
.A(n_1038),
.Y(n_1130)
);

OA21x2_ASAP7_75t_L g1131 ( 
.A1(n_1095),
.A2(n_877),
.B(n_933),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_1007),
.A2(n_1029),
.B(n_1027),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_993),
.Y(n_1133)
);

OR2x2_ASAP7_75t_L g1134 ( 
.A(n_1069),
.B(n_947),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_997),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1018),
.A2(n_930),
.B(n_939),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_987),
.B(n_943),
.Y(n_1137)
);

OAI22xp5_ASAP7_75t_L g1138 ( 
.A1(n_988),
.A2(n_943),
.B1(n_955),
.B2(n_1094),
.Y(n_1138)
);

OA21x2_ASAP7_75t_L g1139 ( 
.A1(n_1081),
.A2(n_1086),
.B(n_1050),
.Y(n_1139)
);

INVx3_ASAP7_75t_SL g1140 ( 
.A(n_1089),
.Y(n_1140)
);

NAND3xp33_ASAP7_75t_L g1141 ( 
.A(n_1010),
.B(n_1009),
.C(n_1043),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1067),
.A2(n_985),
.B(n_1008),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_L g1143 ( 
.A(n_1028),
.B(n_1032),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1003),
.A2(n_1052),
.B(n_1020),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_1017),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_1000),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_L g1147 ( 
.A(n_1061),
.B(n_1097),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1087),
.B(n_1001),
.Y(n_1148)
);

NAND3xp33_ASAP7_75t_SL g1149 ( 
.A(n_1022),
.B(n_1026),
.C(n_1082),
.Y(n_1149)
);

INVxp67_ASAP7_75t_SL g1150 ( 
.A(n_1000),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1030),
.Y(n_1151)
);

HB1xp67_ASAP7_75t_L g1152 ( 
.A(n_1039),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_L g1153 ( 
.A(n_1004),
.B(n_1005),
.Y(n_1153)
);

OAI21xp5_ASAP7_75t_L g1154 ( 
.A1(n_1052),
.A2(n_1049),
.B(n_1041),
.Y(n_1154)
);

NAND2xp5_ASAP7_75t_SL g1155 ( 
.A(n_1034),
.B(n_1019),
.Y(n_1155)
);

AO22x2_ASAP7_75t_L g1156 ( 
.A1(n_1066),
.A2(n_1088),
.B1(n_1035),
.B2(n_1065),
.Y(n_1156)
);

A2O1A1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_1070),
.A2(n_1080),
.B(n_1096),
.C(n_1077),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_SL g1158 ( 
.A(n_986),
.B(n_1006),
.Y(n_1158)
);

AO31x2_ASAP7_75t_L g1159 ( 
.A1(n_1049),
.A2(n_1056),
.A3(n_1057),
.B(n_1062),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_1000),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_1063),
.Y(n_1161)
);

INVx1_ASAP7_75t_SL g1162 ( 
.A(n_1014),
.Y(n_1162)
);

OAI21xp5_ASAP7_75t_L g1163 ( 
.A1(n_1084),
.A2(n_1037),
.B(n_1060),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_1064),
.B(n_1085),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1059),
.B(n_1075),
.Y(n_1165)
);

NOR2xp67_ASAP7_75t_L g1166 ( 
.A(n_1047),
.B(n_1053),
.Y(n_1166)
);

AOI221x1_ASAP7_75t_L g1167 ( 
.A1(n_1068),
.A2(n_1071),
.B1(n_1073),
.B2(n_1024),
.C(n_998),
.Y(n_1167)
);

INVx6_ASAP7_75t_SL g1168 ( 
.A(n_1076),
.Y(n_1168)
);

BUFx12f_ASAP7_75t_L g1169 ( 
.A(n_1078),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1059),
.A2(n_1075),
.B(n_1046),
.C(n_991),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_1046),
.Y(n_1171)
);

NAND2xp33_ASAP7_75t_R g1172 ( 
.A(n_1023),
.B(n_1101),
.Y(n_1172)
);

INVx4_ASAP7_75t_L g1173 ( 
.A(n_991),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_1042),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_994),
.B(n_1042),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_1036),
.A2(n_1042),
.B(n_1040),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1036),
.A2(n_994),
.B(n_998),
.Y(n_1177)
);

AND2x2_ASAP7_75t_L g1178 ( 
.A(n_1076),
.B(n_1045),
.Y(n_1178)
);

INVx4_ASAP7_75t_L g1179 ( 
.A(n_994),
.Y(n_1179)
);

INVx3_ASAP7_75t_L g1180 ( 
.A(n_1076),
.Y(n_1180)
);

AOI21xp33_ASAP7_75t_L g1181 ( 
.A1(n_1035),
.A2(n_998),
.B(n_1079),
.Y(n_1181)
);

NAND2xp5_ASAP7_75t_L g1182 ( 
.A(n_1048),
.B(n_999),
.Y(n_1182)
);

NOR2xp67_ASAP7_75t_L g1183 ( 
.A(n_1035),
.B(n_843),
.Y(n_1183)
);

OAI21xp5_ASAP7_75t_SL g1184 ( 
.A1(n_1044),
.A2(n_920),
.B(n_705),
.Y(n_1184)
);

INVxp67_ASAP7_75t_L g1185 ( 
.A(n_1013),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_990),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1092),
.B(n_858),
.Y(n_1187)
);

NAND2xp5_ASAP7_75t_SL g1188 ( 
.A(n_1002),
.B(n_846),
.Y(n_1188)
);

NAND2xp5_ASAP7_75t_L g1189 ( 
.A(n_1092),
.B(n_858),
.Y(n_1189)
);

INVx4_ASAP7_75t_L g1190 ( 
.A(n_1000),
.Y(n_1190)
);

AOI211x1_ASAP7_75t_L g1191 ( 
.A1(n_1083),
.A2(n_1072),
.B(n_1079),
.C(n_984),
.Y(n_1191)
);

BUFx12f_ASAP7_75t_L g1192 ( 
.A(n_1089),
.Y(n_1192)
);

NAND2xp5_ASAP7_75t_L g1193 ( 
.A(n_1092),
.B(n_858),
.Y(n_1193)
);

OAI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1074),
.A2(n_1100),
.B(n_1099),
.Y(n_1194)
);

BUFx6f_ASAP7_75t_L g1195 ( 
.A(n_1000),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1092),
.B(n_858),
.Y(n_1196)
);

AOI21xp33_ASAP7_75t_L g1197 ( 
.A1(n_1074),
.A2(n_920),
.B(n_858),
.Y(n_1197)
);

NOR2xp33_ASAP7_75t_L g1198 ( 
.A(n_1002),
.B(n_373),
.Y(n_1198)
);

AO31x2_ASAP7_75t_L g1199 ( 
.A1(n_1098),
.A2(n_1054),
.A3(n_1015),
.B(n_1100),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_990),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_SL g1201 ( 
.A(n_1002),
.B(n_846),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1092),
.B(n_858),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1092),
.B(n_858),
.Y(n_1203)
);

INVx2_ASAP7_75t_SL g1204 ( 
.A(n_1038),
.Y(n_1204)
);

INVx5_ASAP7_75t_L g1205 ( 
.A(n_994),
.Y(n_1205)
);

INVx3_ASAP7_75t_L g1206 ( 
.A(n_1012),
.Y(n_1206)
);

AOI21x1_ASAP7_75t_L g1207 ( 
.A1(n_989),
.A2(n_1098),
.B(n_1100),
.Y(n_1207)
);

AOI21x1_ASAP7_75t_L g1208 ( 
.A1(n_989),
.A2(n_1098),
.B(n_1100),
.Y(n_1208)
);

INVx3_ASAP7_75t_L g1209 ( 
.A(n_1012),
.Y(n_1209)
);

NOR2xp67_ASAP7_75t_L g1210 ( 
.A(n_1034),
.B(n_843),
.Y(n_1210)
);

OR2x2_ASAP7_75t_L g1211 ( 
.A(n_1002),
.B(n_605),
.Y(n_1211)
);

NAND2x1p5_ASAP7_75t_L g1212 ( 
.A(n_1012),
.B(n_849),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1092),
.B(n_858),
.Y(n_1213)
);

AND2x2_ASAP7_75t_L g1214 ( 
.A(n_1002),
.B(n_735),
.Y(n_1214)
);

BUFx6f_ASAP7_75t_L g1215 ( 
.A(n_1000),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_SL g1216 ( 
.A1(n_996),
.A2(n_723),
.B(n_718),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_990),
.Y(n_1217)
);

OAI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1074),
.A2(n_1100),
.B(n_1099),
.Y(n_1218)
);

OA21x2_ASAP7_75t_L g1219 ( 
.A1(n_992),
.A2(n_1098),
.B(n_1100),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_1074),
.A2(n_920),
.B(n_949),
.C(n_983),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_990),
.Y(n_1221)
);

A2O1A1Ixp33_ASAP7_75t_L g1222 ( 
.A1(n_1074),
.A2(n_920),
.B(n_949),
.C(n_983),
.Y(n_1222)
);

OAI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_1074),
.A2(n_1100),
.B(n_1099),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1092),
.B(n_858),
.Y(n_1224)
);

A2O1A1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_1074),
.A2(n_920),
.B(n_949),
.C(n_983),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1038),
.Y(n_1226)
);

AO31x2_ASAP7_75t_L g1227 ( 
.A1(n_1098),
.A2(n_1054),
.A3(n_1015),
.B(n_1100),
.Y(n_1227)
);

BUFx8_ASAP7_75t_L g1228 ( 
.A(n_1063),
.Y(n_1228)
);

CKINVDCx20_ASAP7_75t_R g1229 ( 
.A(n_993),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_990),
.Y(n_1230)
);

A2O1A1Ixp33_ASAP7_75t_L g1231 ( 
.A1(n_1074),
.A2(n_920),
.B(n_949),
.C(n_983),
.Y(n_1231)
);

AND2x4_ASAP7_75t_L g1232 ( 
.A(n_1108),
.B(n_1180),
.Y(n_1232)
);

OAI22xp5_ASAP7_75t_L g1233 ( 
.A1(n_1184),
.A2(n_1203),
.B1(n_1224),
.B2(n_1196),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1234)
);

AOI21xp33_ASAP7_75t_SL g1235 ( 
.A1(n_1158),
.A2(n_1184),
.B(n_1141),
.Y(n_1235)
);

O2A1O1Ixp33_ASAP7_75t_L g1236 ( 
.A1(n_1220),
.A2(n_1231),
.B(n_1225),
.C(n_1222),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1164),
.B(n_1214),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_1187),
.B(n_1189),
.Y(n_1238)
);

INVx4_ASAP7_75t_L g1239 ( 
.A(n_1114),
.Y(n_1239)
);

NAND2xp5_ASAP7_75t_L g1240 ( 
.A(n_1202),
.B(n_1213),
.Y(n_1240)
);

OR2x2_ASAP7_75t_L g1241 ( 
.A(n_1211),
.B(n_1188),
.Y(n_1241)
);

AND2x4_ASAP7_75t_L g1242 ( 
.A(n_1108),
.B(n_1180),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_1193),
.B(n_1143),
.Y(n_1243)
);

OAI22xp5_ASAP7_75t_L g1244 ( 
.A1(n_1141),
.A2(n_1162),
.B1(n_1185),
.B2(n_1111),
.Y(n_1244)
);

BUFx6f_ASAP7_75t_L g1245 ( 
.A(n_1146),
.Y(n_1245)
);

INVx4_ASAP7_75t_L g1246 ( 
.A(n_1114),
.Y(n_1246)
);

AND2x4_ASAP7_75t_L g1247 ( 
.A(n_1165),
.B(n_1174),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1110),
.Y(n_1248)
);

AOI221xp5_ASAP7_75t_L g1249 ( 
.A1(n_1197),
.A2(n_1191),
.B1(n_1157),
.B2(n_1149),
.C(n_1156),
.Y(n_1249)
);

NOR2xp33_ASAP7_75t_R g1250 ( 
.A(n_1172),
.B(n_1133),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1197),
.A2(n_1112),
.B1(n_1156),
.B2(n_1181),
.Y(n_1251)
);

OR2x6_ASAP7_75t_L g1252 ( 
.A(n_1216),
.B(n_1142),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_1124),
.A2(n_1136),
.B(n_1128),
.Y(n_1253)
);

OAI22xp33_ASAP7_75t_L g1254 ( 
.A1(n_1106),
.A2(n_1183),
.B1(n_1121),
.B2(n_1182),
.Y(n_1254)
);

BUFx2_ASAP7_75t_R g1255 ( 
.A(n_1140),
.Y(n_1255)
);

INVx2_ASAP7_75t_L g1256 ( 
.A(n_1116),
.Y(n_1256)
);

INVx2_ASAP7_75t_L g1257 ( 
.A(n_1125),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1194),
.A2(n_1223),
.B(n_1218),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1194),
.A2(n_1223),
.B(n_1218),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1129),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_SL g1261 ( 
.A(n_1111),
.B(n_1113),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1181),
.A2(n_1113),
.B1(n_1201),
.B2(n_1126),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1186),
.Y(n_1263)
);

BUFx6f_ASAP7_75t_L g1264 ( 
.A(n_1146),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1200),
.Y(n_1265)
);

INVxp67_ASAP7_75t_L g1266 ( 
.A(n_1134),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1217),
.Y(n_1267)
);

NAND3xp33_ASAP7_75t_L g1268 ( 
.A(n_1109),
.B(n_1198),
.C(n_1147),
.Y(n_1268)
);

INVx3_ASAP7_75t_L g1269 ( 
.A(n_1179),
.Y(n_1269)
);

AO21x2_ASAP7_75t_L g1270 ( 
.A1(n_1126),
.A2(n_1154),
.B(n_1104),
.Y(n_1270)
);

AO21x2_ASAP7_75t_L g1271 ( 
.A1(n_1154),
.A2(n_1104),
.B(n_1163),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1221),
.Y(n_1272)
);

INVx2_ASAP7_75t_L g1273 ( 
.A(n_1230),
.Y(n_1273)
);

OAI21x1_ASAP7_75t_L g1274 ( 
.A1(n_1219),
.A2(n_1138),
.B(n_1177),
.Y(n_1274)
);

INVx3_ASAP7_75t_L g1275 ( 
.A(n_1179),
.Y(n_1275)
);

CKINVDCx20_ASAP7_75t_R g1276 ( 
.A(n_1229),
.Y(n_1276)
);

NAND2xp5_ASAP7_75t_L g1277 ( 
.A(n_1103),
.B(n_1148),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1168),
.A2(n_1137),
.B1(n_1119),
.B2(n_1135),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1120),
.B(n_1153),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1138),
.A2(n_1176),
.B(n_1127),
.Y(n_1280)
);

OAI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1127),
.A2(n_1107),
.B(n_1153),
.Y(n_1281)
);

BUFx6f_ASAP7_75t_L g1282 ( 
.A(n_1146),
.Y(n_1282)
);

NOR2xp33_ASAP7_75t_L g1283 ( 
.A(n_1115),
.B(n_1123),
.Y(n_1283)
);

INVxp67_ASAP7_75t_L g1284 ( 
.A(n_1152),
.Y(n_1284)
);

AND2x4_ASAP7_75t_L g1285 ( 
.A(n_1170),
.B(n_1178),
.Y(n_1285)
);

A2O1A1Ixp33_ASAP7_75t_L g1286 ( 
.A1(n_1107),
.A2(n_1114),
.B(n_1205),
.C(n_1151),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1167),
.A2(n_1175),
.B(n_1139),
.Y(n_1287)
);

INVxp67_ASAP7_75t_L g1288 ( 
.A(n_1145),
.Y(n_1288)
);

NOR2xp67_ASAP7_75t_L g1289 ( 
.A(n_1210),
.B(n_1204),
.Y(n_1289)
);

INVx1_ASAP7_75t_SL g1290 ( 
.A(n_1123),
.Y(n_1290)
);

NOR2xp67_ASAP7_75t_L g1291 ( 
.A(n_1130),
.B(n_1155),
.Y(n_1291)
);

AOI221xp5_ASAP7_75t_L g1292 ( 
.A1(n_1105),
.A2(n_1226),
.B1(n_1175),
.B2(n_1161),
.C(n_1171),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1139),
.A2(n_1131),
.B(n_1212),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1168),
.A2(n_1166),
.B1(n_1205),
.B2(n_1150),
.Y(n_1294)
);

NAND2xp5_ASAP7_75t_L g1295 ( 
.A(n_1159),
.B(n_1209),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1228),
.Y(n_1296)
);

NOR2xp33_ASAP7_75t_L g1297 ( 
.A(n_1192),
.B(n_1173),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1160),
.Y(n_1298)
);

NOR2x1_ASAP7_75t_R g1299 ( 
.A(n_1169),
.B(n_1190),
.Y(n_1299)
);

OAI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1205),
.A2(n_1131),
.B1(n_1173),
.B2(n_1206),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1160),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1212),
.A2(n_1227),
.B(n_1199),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1190),
.B(n_1195),
.Y(n_1303)
);

NAND2xp5_ASAP7_75t_L g1304 ( 
.A(n_1159),
.B(n_1160),
.Y(n_1304)
);

AOI22xp33_ASAP7_75t_L g1305 ( 
.A1(n_1228),
.A2(n_1195),
.B1(n_1215),
.B2(n_1199),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1118),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1215),
.B(n_1118),
.Y(n_1307)
);

NAND2xp5_ASAP7_75t_SL g1308 ( 
.A(n_1220),
.B(n_1225),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1220),
.A2(n_920),
.B(n_1222),
.Y(n_1309)
);

BUFx4f_ASAP7_75t_SL g1310 ( 
.A(n_1168),
.Y(n_1310)
);

CKINVDCx9p33_ASAP7_75t_R g1311 ( 
.A(n_1198),
.Y(n_1311)
);

AND2x2_ASAP7_75t_SL g1312 ( 
.A(n_1179),
.B(n_882),
.Y(n_1312)
);

OAI21x1_ASAP7_75t_L g1313 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1313)
);

HB1xp67_ASAP7_75t_L g1314 ( 
.A(n_1110),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1220),
.A2(n_920),
.B(n_1222),
.Y(n_1315)
);

O2A1O1Ixp33_ASAP7_75t_L g1316 ( 
.A1(n_1220),
.A2(n_1231),
.B(n_1225),
.C(n_1222),
.Y(n_1316)
);

OAI21x1_ASAP7_75t_L g1317 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1216),
.A2(n_996),
.B(n_918),
.Y(n_1318)
);

OR2x2_ASAP7_75t_L g1319 ( 
.A(n_1211),
.B(n_1214),
.Y(n_1319)
);

OAI21xp33_ASAP7_75t_SL g1320 ( 
.A1(n_1187),
.A2(n_873),
.B(n_1016),
.Y(n_1320)
);

NAND2x1p5_ASAP7_75t_L g1321 ( 
.A(n_1114),
.B(n_1205),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1211),
.Y(n_1322)
);

INVxp67_ASAP7_75t_L g1323 ( 
.A(n_1214),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1220),
.A2(n_920),
.B(n_1222),
.Y(n_1324)
);

OAI22xp33_ASAP7_75t_L g1325 ( 
.A1(n_1106),
.A2(n_882),
.B1(n_1184),
.B2(n_1083),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1152),
.Y(n_1326)
);

AO31x2_ASAP7_75t_L g1327 ( 
.A1(n_1121),
.A2(n_1167),
.A3(n_1222),
.B(n_1220),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1175),
.A2(n_948),
.B(n_929),
.Y(n_1328)
);

BUFx2_ASAP7_75t_L g1329 ( 
.A(n_1152),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1330)
);

OAI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1187),
.B(n_1189),
.Y(n_1332)
);

INVx3_ASAP7_75t_SL g1333 ( 
.A(n_1140),
.Y(n_1333)
);

OA21x2_ASAP7_75t_L g1334 ( 
.A1(n_1144),
.A2(n_1132),
.B(n_1194),
.Y(n_1334)
);

OA21x2_ASAP7_75t_L g1335 ( 
.A1(n_1144),
.A2(n_1132),
.B(n_1194),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1216),
.A2(n_996),
.B(n_918),
.Y(n_1336)
);

OAI21xp5_ASAP7_75t_L g1337 ( 
.A1(n_1220),
.A2(n_920),
.B(n_1222),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1164),
.B(n_1214),
.Y(n_1338)
);

OAI22xp33_ASAP7_75t_L g1339 ( 
.A1(n_1106),
.A2(n_882),
.B1(n_1184),
.B2(n_1083),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1117),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1117),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1220),
.A2(n_920),
.B(n_1222),
.Y(n_1342)
);

BUFx8_ASAP7_75t_L g1343 ( 
.A(n_1169),
.Y(n_1343)
);

BUFx2_ASAP7_75t_L g1344 ( 
.A(n_1152),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1117),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1164),
.B(n_1214),
.Y(n_1346)
);

NOR2xp33_ASAP7_75t_L g1347 ( 
.A(n_1184),
.B(n_920),
.Y(n_1347)
);

OAI22xp5_ASAP7_75t_L g1348 ( 
.A1(n_1184),
.A2(n_1189),
.B1(n_1196),
.B2(n_1187),
.Y(n_1348)
);

OAI21x1_ASAP7_75t_L g1349 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1349)
);

CKINVDCx8_ASAP7_75t_R g1350 ( 
.A(n_1146),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1122),
.A2(n_1208),
.B(n_1207),
.Y(n_1351)
);

INVx2_ASAP7_75t_SL g1352 ( 
.A(n_1226),
.Y(n_1352)
);

INVx1_ASAP7_75t_SL g1353 ( 
.A(n_1211),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1117),
.Y(n_1354)
);

NOR2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1210),
.B(n_713),
.Y(n_1355)
);

BUFx3_ASAP7_75t_L g1356 ( 
.A(n_1226),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1175),
.A2(n_948),
.B(n_929),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1277),
.B(n_1243),
.Y(n_1358)
);

O2A1O1Ixp33_ASAP7_75t_L g1359 ( 
.A1(n_1347),
.A2(n_1235),
.B(n_1337),
.C(n_1342),
.Y(n_1359)
);

O2A1O1Ixp33_ASAP7_75t_L g1360 ( 
.A1(n_1347),
.A2(n_1315),
.B(n_1309),
.C(n_1324),
.Y(n_1360)
);

AOI21xp5_ASAP7_75t_SL g1361 ( 
.A1(n_1321),
.A2(n_1240),
.B(n_1238),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1259),
.A2(n_1336),
.B(n_1318),
.Y(n_1362)
);

AOI21xp5_ASAP7_75t_SL g1363 ( 
.A1(n_1321),
.A2(n_1332),
.B(n_1316),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1232),
.B(n_1242),
.Y(n_1364)
);

OR2x6_ASAP7_75t_L g1365 ( 
.A(n_1252),
.B(n_1236),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1308),
.A2(n_1316),
.B(n_1236),
.Y(n_1366)
);

AOI21xp5_ASAP7_75t_SL g1367 ( 
.A1(n_1233),
.A2(n_1348),
.B(n_1252),
.Y(n_1367)
);

HB1xp67_ASAP7_75t_L g1368 ( 
.A(n_1248),
.Y(n_1368)
);

AND2x2_ASAP7_75t_L g1369 ( 
.A(n_1346),
.B(n_1323),
.Y(n_1369)
);

OA22x2_ASAP7_75t_L g1370 ( 
.A1(n_1244),
.A2(n_1357),
.B1(n_1328),
.B2(n_1247),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1322),
.B(n_1353),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_1314),
.Y(n_1372)
);

AOI21x1_ASAP7_75t_SL g1373 ( 
.A1(n_1304),
.A2(n_1295),
.B(n_1307),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_L g1374 ( 
.A(n_1266),
.B(n_1279),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1297),
.B(n_1241),
.Y(n_1375)
);

AOI21xp5_ASAP7_75t_L g1376 ( 
.A1(n_1252),
.A2(n_1258),
.B(n_1270),
.Y(n_1376)
);

O2A1O1Ixp5_ASAP7_75t_L g1377 ( 
.A1(n_1325),
.A2(n_1339),
.B(n_1261),
.C(n_1254),
.Y(n_1377)
);

O2A1O1Ixp5_ASAP7_75t_L g1378 ( 
.A1(n_1325),
.A2(n_1339),
.B(n_1261),
.C(n_1254),
.Y(n_1378)
);

CKINVDCx11_ASAP7_75t_R g1379 ( 
.A(n_1296),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1278),
.A2(n_1312),
.B1(n_1262),
.B2(n_1290),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1232),
.B(n_1242),
.Y(n_1381)
);

AOI31xp33_ASAP7_75t_L g1382 ( 
.A1(n_1249),
.A2(n_1292),
.A3(n_1299),
.B(n_1262),
.Y(n_1382)
);

AOI21xp5_ASAP7_75t_SL g1383 ( 
.A1(n_1239),
.A2(n_1246),
.B(n_1286),
.Y(n_1383)
);

NOR2xp67_ASAP7_75t_L g1384 ( 
.A(n_1297),
.B(n_1284),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_SL g1385 ( 
.A1(n_1239),
.A2(n_1246),
.B(n_1294),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1257),
.Y(n_1386)
);

OAI22xp5_ASAP7_75t_L g1387 ( 
.A1(n_1278),
.A2(n_1312),
.B1(n_1283),
.B2(n_1251),
.Y(n_1387)
);

O2A1O1Ixp33_ASAP7_75t_L g1388 ( 
.A1(n_1320),
.A2(n_1281),
.B(n_1288),
.C(n_1283),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1250),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1274),
.A2(n_1253),
.B(n_1351),
.Y(n_1390)
);

INVx3_ASAP7_75t_L g1391 ( 
.A(n_1350),
.Y(n_1391)
);

OA21x2_ASAP7_75t_L g1392 ( 
.A1(n_1234),
.A2(n_1313),
.B(n_1331),
.Y(n_1392)
);

NOR2xp67_ASAP7_75t_L g1393 ( 
.A(n_1289),
.B(n_1352),
.Y(n_1393)
);

HB1xp67_ASAP7_75t_L g1394 ( 
.A(n_1326),
.Y(n_1394)
);

INVx3_ASAP7_75t_SL g1395 ( 
.A(n_1333),
.Y(n_1395)
);

A2O1A1Ixp33_ASAP7_75t_L g1396 ( 
.A1(n_1280),
.A2(n_1251),
.B(n_1285),
.C(n_1291),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1305),
.A2(n_1310),
.B1(n_1344),
.B2(n_1329),
.Y(n_1397)
);

AND2x4_ASAP7_75t_L g1398 ( 
.A(n_1260),
.B(n_1267),
.Y(n_1398)
);

O2A1O1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1288),
.A2(n_1300),
.B(n_1272),
.C(n_1265),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1305),
.A2(n_1310),
.B1(n_1263),
.B2(n_1276),
.Y(n_1400)
);

OAI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1276),
.A2(n_1356),
.B1(n_1333),
.B2(n_1345),
.Y(n_1401)
);

INVxp33_ASAP7_75t_L g1402 ( 
.A(n_1250),
.Y(n_1402)
);

A2O1A1Ixp33_ASAP7_75t_L g1403 ( 
.A1(n_1287),
.A2(n_1302),
.B(n_1311),
.C(n_1340),
.Y(n_1403)
);

AND2x4_ASAP7_75t_L g1404 ( 
.A(n_1273),
.B(n_1269),
.Y(n_1404)
);

OA21x2_ASAP7_75t_L g1405 ( 
.A1(n_1317),
.A2(n_1349),
.B(n_1330),
.Y(n_1405)
);

AOI21xp5_ASAP7_75t_L g1406 ( 
.A1(n_1334),
.A2(n_1335),
.B(n_1271),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1341),
.B(n_1354),
.Y(n_1407)
);

AOI21xp5_ASAP7_75t_SL g1408 ( 
.A1(n_1334),
.A2(n_1335),
.B(n_1303),
.Y(n_1408)
);

AOI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1334),
.A2(n_1335),
.B(n_1271),
.Y(n_1409)
);

BUFx8_ASAP7_75t_SL g1410 ( 
.A(n_1296),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1298),
.B(n_1301),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1245),
.B(n_1264),
.Y(n_1412)
);

OR2x2_ASAP7_75t_L g1413 ( 
.A(n_1327),
.B(n_1306),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1293),
.A2(n_1303),
.B(n_1355),
.C(n_1327),
.Y(n_1414)
);

OR2x2_ASAP7_75t_L g1415 ( 
.A(n_1245),
.B(n_1264),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1264),
.A2(n_1282),
.B(n_1255),
.Y(n_1416)
);

AOI21xp5_ASAP7_75t_L g1417 ( 
.A1(n_1282),
.A2(n_1259),
.B(n_1309),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1282),
.A2(n_1347),
.B(n_1184),
.C(n_920),
.Y(n_1418)
);

AOI21xp5_ASAP7_75t_SL g1419 ( 
.A1(n_1343),
.A2(n_1222),
.B(n_1220),
.Y(n_1419)
);

NAND2xp5_ASAP7_75t_L g1420 ( 
.A(n_1343),
.B(n_1277),
.Y(n_1420)
);

HB1xp67_ASAP7_75t_L g1421 ( 
.A(n_1248),
.Y(n_1421)
);

O2A1O1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1347),
.A2(n_1184),
.B(n_1222),
.C(n_1220),
.Y(n_1422)
);

OAI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1347),
.A2(n_1184),
.B1(n_1141),
.B2(n_1268),
.Y(n_1423)
);

O2A1O1Ixp5_ASAP7_75t_L g1424 ( 
.A1(n_1309),
.A2(n_1315),
.B(n_1337),
.C(n_1324),
.Y(n_1424)
);

AND2x2_ASAP7_75t_L g1425 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1425)
);

BUFx3_ASAP7_75t_L g1426 ( 
.A(n_1356),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1347),
.A2(n_1184),
.B1(n_1141),
.B2(n_1268),
.Y(n_1427)
);

NOR2xp67_ASAP7_75t_L g1428 ( 
.A(n_1323),
.B(n_1185),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1429)
);

AOI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1259),
.A2(n_1315),
.B(n_1309),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1319),
.B(n_1241),
.Y(n_1431)
);

AND2x6_ASAP7_75t_L g1432 ( 
.A(n_1269),
.B(n_1275),
.Y(n_1432)
);

O2A1O1Ixp33_ASAP7_75t_L g1433 ( 
.A1(n_1347),
.A2(n_1184),
.B(n_1222),
.C(n_1220),
.Y(n_1433)
);

INVx1_ASAP7_75t_SL g1434 ( 
.A(n_1237),
.Y(n_1434)
);

AOI21xp5_ASAP7_75t_SL g1435 ( 
.A1(n_1309),
.A2(n_1222),
.B(n_1220),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1277),
.B(n_1243),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1347),
.A2(n_1184),
.B(n_920),
.C(n_1235),
.Y(n_1438)
);

AOI21xp5_ASAP7_75t_SL g1439 ( 
.A1(n_1309),
.A2(n_1222),
.B(n_1220),
.Y(n_1439)
);

AND2x2_ASAP7_75t_L g1440 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1440)
);

O2A1O1Ixp33_ASAP7_75t_L g1441 ( 
.A1(n_1347),
.A2(n_1184),
.B(n_1222),
.C(n_1220),
.Y(n_1441)
);

OA22x2_ASAP7_75t_L g1442 ( 
.A1(n_1309),
.A2(n_1184),
.B1(n_1106),
.B2(n_1315),
.Y(n_1442)
);

OA22x2_ASAP7_75t_L g1443 ( 
.A1(n_1309),
.A2(n_1184),
.B1(n_1106),
.B2(n_1315),
.Y(n_1443)
);

AND2x2_ASAP7_75t_L g1444 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1256),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1237),
.B(n_1338),
.Y(n_1449)
);

AOI21xp5_ASAP7_75t_SL g1450 ( 
.A1(n_1309),
.A2(n_1222),
.B(n_1220),
.Y(n_1450)
);

HB1xp67_ASAP7_75t_L g1451 ( 
.A(n_1248),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1326),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1413),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1448),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1442),
.A2(n_1443),
.B1(n_1423),
.B2(n_1427),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1430),
.B(n_1408),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1430),
.B(n_1376),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1406),
.B(n_1409),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1390),
.Y(n_1459)
);

BUFx2_ASAP7_75t_L g1460 ( 
.A(n_1368),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1406),
.B(n_1409),
.Y(n_1461)
);

OR2x2_ASAP7_75t_L g1462 ( 
.A(n_1372),
.B(n_1421),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1442),
.A2(n_1443),
.B1(n_1366),
.B2(n_1387),
.Y(n_1463)
);

AND2x2_ASAP7_75t_L g1464 ( 
.A(n_1362),
.B(n_1398),
.Y(n_1464)
);

INVxp67_ASAP7_75t_SL g1465 ( 
.A(n_1399),
.Y(n_1465)
);

INVx2_ASAP7_75t_L g1466 ( 
.A(n_1392),
.Y(n_1466)
);

INVx11_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1405),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1365),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_L g1470 ( 
.A(n_1438),
.B(n_1359),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1365),
.B(n_1403),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1424),
.A2(n_1378),
.B(n_1377),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1398),
.B(n_1417),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1386),
.B(n_1424),
.Y(n_1474)
);

INVx4_ASAP7_75t_SL g1475 ( 
.A(n_1432),
.Y(n_1475)
);

OA21x2_ASAP7_75t_L g1476 ( 
.A1(n_1414),
.A2(n_1396),
.B(n_1418),
.Y(n_1476)
);

AO21x2_ASAP7_75t_L g1477 ( 
.A1(n_1360),
.A2(n_1450),
.B(n_1439),
.Y(n_1477)
);

OR2x2_ASAP7_75t_L g1478 ( 
.A(n_1451),
.B(n_1431),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1360),
.A2(n_1435),
.B(n_1359),
.Y(n_1479)
);

OA21x2_ASAP7_75t_L g1480 ( 
.A1(n_1407),
.A2(n_1382),
.B(n_1404),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1367),
.A2(n_1422),
.B(n_1441),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1432),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1399),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1388),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1388),
.Y(n_1485)
);

INVx2_ASAP7_75t_L g1486 ( 
.A(n_1370),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1370),
.Y(n_1487)
);

AO21x2_ASAP7_75t_L g1488 ( 
.A1(n_1422),
.A2(n_1441),
.B(n_1433),
.Y(n_1488)
);

OAI21xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1363),
.A2(n_1419),
.B(n_1383),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1433),
.A2(n_1380),
.B(n_1400),
.Y(n_1490)
);

HB1xp67_ASAP7_75t_L g1491 ( 
.A(n_1394),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1358),
.B(n_1437),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1411),
.Y(n_1493)
);

INVx2_ASAP7_75t_L g1494 ( 
.A(n_1369),
.Y(n_1494)
);

NOR2x1_ASAP7_75t_L g1495 ( 
.A(n_1361),
.B(n_1385),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1374),
.Y(n_1496)
);

BUFx3_ASAP7_75t_L g1497 ( 
.A(n_1452),
.Y(n_1497)
);

OAI332xp33_ASAP7_75t_L g1498 ( 
.A1(n_1397),
.A2(n_1420),
.A3(n_1401),
.B1(n_1434),
.B2(n_1371),
.B3(n_1415),
.C1(n_1428),
.C2(n_1402),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1412),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1456),
.B(n_1449),
.Y(n_1500)
);

AND2x4_ASAP7_75t_L g1501 ( 
.A(n_1464),
.B(n_1375),
.Y(n_1501)
);

AND2x2_ASAP7_75t_L g1502 ( 
.A(n_1456),
.B(n_1447),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1496),
.B(n_1446),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1454),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1456),
.B(n_1445),
.Y(n_1505)
);

OAI222xp33_ASAP7_75t_L g1506 ( 
.A1(n_1455),
.A2(n_1416),
.B1(n_1389),
.B2(n_1440),
.C1(n_1436),
.C2(n_1429),
.Y(n_1506)
);

BUFx2_ASAP7_75t_L g1507 ( 
.A(n_1464),
.Y(n_1507)
);

OR2x2_ASAP7_75t_L g1508 ( 
.A(n_1462),
.B(n_1460),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1457),
.B(n_1444),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1457),
.B(n_1458),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1459),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1453),
.Y(n_1512)
);

CKINVDCx20_ASAP7_75t_R g1513 ( 
.A(n_1497),
.Y(n_1513)
);

AOI211xp5_ASAP7_75t_SL g1514 ( 
.A1(n_1470),
.A2(n_1498),
.B(n_1485),
.C(n_1484),
.Y(n_1514)
);

BUFx3_ASAP7_75t_L g1515 ( 
.A(n_1482),
.Y(n_1515)
);

OR2x2_ASAP7_75t_L g1516 ( 
.A(n_1462),
.B(n_1425),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1467),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1461),
.B(n_1473),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1496),
.B(n_1384),
.Y(n_1519)
);

AOI33xp33_ASAP7_75t_L g1520 ( 
.A1(n_1455),
.A2(n_1364),
.A3(n_1381),
.B1(n_1393),
.B2(n_1379),
.B3(n_1410),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1466),
.Y(n_1521)
);

INVx3_ASAP7_75t_SL g1522 ( 
.A(n_1475),
.Y(n_1522)
);

AND2x4_ASAP7_75t_L g1523 ( 
.A(n_1473),
.B(n_1416),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1496),
.B(n_1426),
.Y(n_1524)
);

AND2x2_ASAP7_75t_L g1525 ( 
.A(n_1461),
.B(n_1373),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1468),
.Y(n_1526)
);

AND2x4_ASAP7_75t_L g1527 ( 
.A(n_1473),
.B(n_1391),
.Y(n_1527)
);

AOI21xp33_ASAP7_75t_L g1528 ( 
.A1(n_1470),
.A2(n_1479),
.B(n_1477),
.Y(n_1528)
);

OR2x2_ASAP7_75t_L g1529 ( 
.A(n_1462),
.B(n_1395),
.Y(n_1529)
);

INVxp67_ASAP7_75t_SL g1530 ( 
.A(n_1474),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1474),
.B(n_1373),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1507),
.B(n_1494),
.Y(n_1532)
);

OAI33xp33_ASAP7_75t_L g1533 ( 
.A1(n_1519),
.A2(n_1492),
.A3(n_1485),
.B1(n_1484),
.B2(n_1483),
.B3(n_1478),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1511),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1512),
.Y(n_1535)
);

NAND3xp33_ASAP7_75t_L g1536 ( 
.A(n_1514),
.B(n_1463),
.C(n_1472),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1528),
.A2(n_1477),
.B1(n_1481),
.B2(n_1488),
.Y(n_1537)
);

HB1xp67_ASAP7_75t_L g1538 ( 
.A(n_1508),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1508),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1512),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1518),
.B(n_1494),
.Y(n_1542)
);

AND2x4_ASAP7_75t_L g1543 ( 
.A(n_1515),
.B(n_1471),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1522),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1504),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_R g1546 ( 
.A(n_1513),
.B(n_1391),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1547)
);

NOR3xp33_ASAP7_75t_SL g1548 ( 
.A(n_1506),
.B(n_1489),
.C(n_1465),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1509),
.B(n_1491),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1527),
.A2(n_1477),
.B1(n_1481),
.B2(n_1488),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1527),
.A2(n_1477),
.B1(n_1481),
.B2(n_1488),
.Y(n_1552)
);

INVx2_ASAP7_75t_SL g1553 ( 
.A(n_1529),
.Y(n_1553)
);

AOI221xp5_ASAP7_75t_L g1554 ( 
.A1(n_1506),
.A2(n_1463),
.B1(n_1498),
.B2(n_1465),
.C(n_1483),
.Y(n_1554)
);

OAI221xp5_ASAP7_75t_L g1555 ( 
.A1(n_1514),
.A2(n_1489),
.B1(n_1495),
.B2(n_1476),
.C(n_1472),
.Y(n_1555)
);

BUFx12f_ASAP7_75t_L g1556 ( 
.A(n_1529),
.Y(n_1556)
);

NAND3xp33_ASAP7_75t_L g1557 ( 
.A(n_1520),
.B(n_1472),
.C(n_1495),
.Y(n_1557)
);

AOI222xp33_ASAP7_75t_L g1558 ( 
.A1(n_1503),
.A2(n_1492),
.B1(n_1471),
.B2(n_1488),
.C1(n_1486),
.C2(n_1487),
.Y(n_1558)
);

OAI21xp5_ASAP7_75t_SL g1559 ( 
.A1(n_1520),
.A2(n_1471),
.B(n_1486),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1518),
.B(n_1499),
.Y(n_1560)
);

AOI33xp33_ASAP7_75t_L g1561 ( 
.A1(n_1525),
.A2(n_1487),
.A3(n_1486),
.B1(n_1474),
.B2(n_1461),
.B3(n_1493),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1508),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1527),
.A2(n_1477),
.B1(n_1481),
.B2(n_1488),
.Y(n_1563)
);

INVx2_ASAP7_75t_SL g1564 ( 
.A(n_1529),
.Y(n_1564)
);

BUFx4f_ASAP7_75t_SL g1565 ( 
.A(n_1513),
.Y(n_1565)
);

NOR2xp33_ASAP7_75t_R g1566 ( 
.A(n_1517),
.B(n_1497),
.Y(n_1566)
);

AOI31xp33_ASAP7_75t_L g1567 ( 
.A1(n_1519),
.A2(n_1471),
.A3(n_1487),
.B(n_1486),
.Y(n_1567)
);

BUFx3_ASAP7_75t_L g1568 ( 
.A(n_1522),
.Y(n_1568)
);

AOI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1527),
.A2(n_1481),
.B1(n_1479),
.B2(n_1490),
.Y(n_1569)
);

OAI31xp33_ASAP7_75t_L g1570 ( 
.A1(n_1525),
.A2(n_1487),
.A3(n_1471),
.B(n_1469),
.Y(n_1570)
);

AND2x6_ASAP7_75t_L g1571 ( 
.A(n_1544),
.B(n_1482),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1545),
.Y(n_1572)
);

AND2x4_ASAP7_75t_L g1573 ( 
.A(n_1544),
.B(n_1523),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1545),
.Y(n_1574)
);

NAND3xp33_ASAP7_75t_L g1575 ( 
.A(n_1536),
.B(n_1472),
.C(n_1476),
.Y(n_1575)
);

NOR3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1555),
.B(n_1531),
.C(n_1524),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1550),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1550),
.Y(n_1578)
);

OAI21xp5_ASAP7_75t_L g1579 ( 
.A1(n_1536),
.A2(n_1476),
.B(n_1472),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1534),
.A2(n_1526),
.B(n_1521),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1553),
.B(n_1564),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1538),
.B(n_1539),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1553),
.Y(n_1583)
);

INVx1_ASAP7_75t_SL g1584 ( 
.A(n_1546),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_SL g1585 ( 
.A(n_1557),
.B(n_1501),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1562),
.B(n_1530),
.Y(n_1586)
);

OR2x2_ASAP7_75t_L g1587 ( 
.A(n_1549),
.B(n_1530),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1564),
.B(n_1510),
.Y(n_1588)
);

INVx5_ASAP7_75t_L g1589 ( 
.A(n_1544),
.Y(n_1589)
);

INVx3_ASAP7_75t_L g1590 ( 
.A(n_1568),
.Y(n_1590)
);

BUFx2_ASAP7_75t_L g1591 ( 
.A(n_1566),
.Y(n_1591)
);

INVx4_ASAP7_75t_SL g1592 ( 
.A(n_1568),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1561),
.B(n_1509),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1542),
.B(n_1510),
.Y(n_1594)
);

INVx2_ASAP7_75t_L g1595 ( 
.A(n_1541),
.Y(n_1595)
);

NOR2x1p5_ASAP7_75t_L g1596 ( 
.A(n_1557),
.B(n_1517),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1542),
.B(n_1510),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1592),
.B(n_1568),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1576),
.B(n_1500),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1591),
.B(n_1543),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1571),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1591),
.B(n_1543),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1580),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1572),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1593),
.B(n_1535),
.Y(n_1605)
);

OAI21xp33_ASAP7_75t_L g1606 ( 
.A1(n_1579),
.A2(n_1537),
.B(n_1548),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1572),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1592),
.B(n_1543),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1585),
.B(n_1500),
.Y(n_1609)
);

INVx2_ASAP7_75t_L g1610 ( 
.A(n_1595),
.Y(n_1610)
);

AND2x4_ASAP7_75t_L g1611 ( 
.A(n_1592),
.B(n_1543),
.Y(n_1611)
);

NAND2xp33_ASAP7_75t_SL g1612 ( 
.A(n_1596),
.B(n_1522),
.Y(n_1612)
);

OAI31xp33_ASAP7_75t_SL g1613 ( 
.A1(n_1575),
.A2(n_1554),
.A3(n_1471),
.B(n_1500),
.Y(n_1613)
);

INVx1_ASAP7_75t_SL g1614 ( 
.A(n_1584),
.Y(n_1614)
);

OR2x2_ASAP7_75t_L g1615 ( 
.A(n_1582),
.B(n_1535),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1595),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1590),
.B(n_1502),
.Y(n_1617)
);

AND2x4_ASAP7_75t_SL g1618 ( 
.A(n_1590),
.B(n_1517),
.Y(n_1618)
);

INVx6_ASAP7_75t_L g1619 ( 
.A(n_1589),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1592),
.B(n_1547),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1590),
.B(n_1502),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1590),
.B(n_1502),
.Y(n_1623)
);

AND2x2_ASAP7_75t_L g1624 ( 
.A(n_1573),
.B(n_1581),
.Y(n_1624)
);

NAND4xp25_ASAP7_75t_L g1625 ( 
.A(n_1586),
.B(n_1558),
.C(n_1569),
.D(n_1559),
.Y(n_1625)
);

OR2x2_ASAP7_75t_L g1626 ( 
.A(n_1582),
.B(n_1540),
.Y(n_1626)
);

AND2x2_ASAP7_75t_L g1627 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1596),
.B(n_1505),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1573),
.B(n_1560),
.Y(n_1629)
);

INVx3_ASAP7_75t_L g1630 ( 
.A(n_1571),
.Y(n_1630)
);

AOI322xp5_ASAP7_75t_L g1631 ( 
.A1(n_1583),
.A2(n_1569),
.A3(n_1552),
.B1(n_1563),
.B2(n_1551),
.C1(n_1533),
.C2(n_1525),
.Y(n_1631)
);

NOR2xp33_ASAP7_75t_L g1632 ( 
.A(n_1573),
.B(n_1556),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1587),
.B(n_1505),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1581),
.B(n_1532),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1589),
.B(n_1532),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1574),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1574),
.Y(n_1637)
);

AOI22xp33_ASAP7_75t_L g1638 ( 
.A1(n_1571),
.A2(n_1479),
.B1(n_1490),
.B2(n_1476),
.Y(n_1638)
);

HB1xp67_ASAP7_75t_L g1639 ( 
.A(n_1577),
.Y(n_1639)
);

OR2x2_ASAP7_75t_L g1640 ( 
.A(n_1586),
.B(n_1540),
.Y(n_1640)
);

INVx3_ASAP7_75t_L g1641 ( 
.A(n_1571),
.Y(n_1641)
);

OR2x2_ASAP7_75t_L g1642 ( 
.A(n_1605),
.B(n_1588),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1608),
.B(n_1594),
.Y(n_1643)
);

AND2x4_ASAP7_75t_L g1644 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1639),
.Y(n_1645)
);

INVx1_ASAP7_75t_L g1646 ( 
.A(n_1604),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1647)
);

AND2x2_ASAP7_75t_SL g1648 ( 
.A(n_1613),
.B(n_1472),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1605),
.B(n_1577),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1604),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1633),
.B(n_1588),
.Y(n_1651)
);

NOR2xp67_ASAP7_75t_SL g1652 ( 
.A(n_1619),
.B(n_1589),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1598),
.B(n_1589),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1599),
.B(n_1578),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1607),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1608),
.B(n_1594),
.Y(n_1656)
);

AOI22xp5_ASAP7_75t_L g1657 ( 
.A1(n_1606),
.A2(n_1479),
.B1(n_1559),
.B2(n_1571),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1600),
.B(n_1602),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1631),
.B(n_1606),
.Y(n_1659)
);

NAND2x1p5_ASAP7_75t_L g1660 ( 
.A(n_1598),
.B(n_1480),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1619),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1601),
.B(n_1480),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1607),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1636),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1636),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1625),
.B(n_1516),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1637),
.Y(n_1667)
);

AND2x2_ASAP7_75t_L g1668 ( 
.A(n_1600),
.B(n_1597),
.Y(n_1668)
);

INVx2_ASAP7_75t_L g1669 ( 
.A(n_1619),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1602),
.B(n_1597),
.Y(n_1670)
);

AND2x4_ASAP7_75t_L g1671 ( 
.A(n_1611),
.B(n_1571),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1619),
.B(n_1517),
.Y(n_1672)
);

INVxp33_ASAP7_75t_L g1673 ( 
.A(n_1632),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1631),
.B(n_1578),
.Y(n_1674)
);

NAND3xp33_ASAP7_75t_SL g1675 ( 
.A(n_1614),
.B(n_1558),
.C(n_1570),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_SL g1676 ( 
.A(n_1625),
.B(n_1570),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1637),
.Y(n_1677)
);

NOR2x1_ASAP7_75t_L g1678 ( 
.A(n_1659),
.B(n_1601),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1646),
.Y(n_1679)
);

NAND3xp33_ASAP7_75t_L g1680 ( 
.A(n_1659),
.B(n_1638),
.C(n_1612),
.Y(n_1680)
);

AND2x2_ASAP7_75t_L g1681 ( 
.A(n_1658),
.B(n_1624),
.Y(n_1681)
);

NOR2x1_ASAP7_75t_L g1682 ( 
.A(n_1675),
.B(n_1601),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1644),
.B(n_1611),
.Y(n_1683)
);

INVx1_ASAP7_75t_SL g1684 ( 
.A(n_1644),
.Y(n_1684)
);

CKINVDCx16_ASAP7_75t_R g1685 ( 
.A(n_1676),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1647),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1645),
.B(n_1609),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1650),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1655),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1669),
.B(n_1634),
.Y(n_1690)
);

NOR2x1_ASAP7_75t_L g1691 ( 
.A(n_1675),
.B(n_1601),
.Y(n_1691)
);

INVx1_ASAP7_75t_SL g1692 ( 
.A(n_1647),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1663),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1664),
.Y(n_1694)
);

NOR2xp33_ASAP7_75t_L g1695 ( 
.A(n_1673),
.B(n_1628),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1643),
.Y(n_1696)
);

OAI22xp5_ASAP7_75t_L g1697 ( 
.A1(n_1657),
.A2(n_1630),
.B1(n_1641),
.B2(n_1611),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1676),
.B(n_1611),
.Y(n_1698)
);

INVx1_ASAP7_75t_SL g1699 ( 
.A(n_1653),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1665),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1667),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1668),
.B(n_1634),
.Y(n_1702)
);

AND3x1_ASAP7_75t_L g1703 ( 
.A(n_1674),
.B(n_1641),
.C(n_1630),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1679),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1678),
.Y(n_1705)
);

OAI211xp5_ASAP7_75t_L g1706 ( 
.A1(n_1682),
.A2(n_1674),
.B(n_1666),
.C(n_1661),
.Y(n_1706)
);

AND2x2_ASAP7_75t_L g1707 ( 
.A(n_1681),
.B(n_1656),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_SL g1708 ( 
.A(n_1685),
.B(n_1648),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1691),
.A2(n_1648),
.B1(n_1671),
.B2(n_1653),
.Y(n_1709)
);

NOR2x1_ASAP7_75t_L g1710 ( 
.A(n_1680),
.B(n_1661),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1688),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1683),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1703),
.A2(n_1671),
.B1(n_1652),
.B2(n_1672),
.Y(n_1713)
);

OAI22xp33_ASAP7_75t_L g1714 ( 
.A1(n_1698),
.A2(n_1660),
.B1(n_1567),
.B2(n_1662),
.Y(n_1714)
);

INVx1_ASAP7_75t_SL g1715 ( 
.A(n_1683),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_SL g1716 ( 
.A(n_1698),
.B(n_1630),
.Y(n_1716)
);

OAI21xp33_ASAP7_75t_L g1717 ( 
.A1(n_1695),
.A2(n_1654),
.B(n_1660),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1689),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1693),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1683),
.Y(n_1720)
);

AOI221x1_ASAP7_75t_L g1721 ( 
.A1(n_1697),
.A2(n_1677),
.B1(n_1654),
.B2(n_1641),
.C(n_1630),
.Y(n_1721)
);

INVxp67_ASAP7_75t_SL g1722 ( 
.A(n_1695),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1694),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1707),
.B(n_1684),
.Y(n_1724)
);

OAI221xp5_ASAP7_75t_L g1725 ( 
.A1(n_1706),
.A2(n_1686),
.B1(n_1699),
.B2(n_1692),
.C(n_1687),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1715),
.B(n_1696),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1705),
.Y(n_1727)
);

BUFx2_ASAP7_75t_L g1728 ( 
.A(n_1712),
.Y(n_1728)
);

INVxp67_ASAP7_75t_SL g1729 ( 
.A(n_1710),
.Y(n_1729)
);

INVx2_ASAP7_75t_L g1730 ( 
.A(n_1712),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1722),
.B(n_1696),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1720),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1720),
.B(n_1700),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_SL g1734 ( 
.A1(n_1704),
.A2(n_1701),
.B1(n_1662),
.B2(n_1479),
.Y(n_1734)
);

OAI22xp5_ASAP7_75t_L g1735 ( 
.A1(n_1729),
.A2(n_1709),
.B1(n_1708),
.B2(n_1713),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1729),
.B(n_1716),
.Y(n_1736)
);

NOR3xp33_ASAP7_75t_L g1737 ( 
.A(n_1731),
.B(n_1725),
.C(n_1726),
.Y(n_1737)
);

OAI21xp33_ASAP7_75t_L g1738 ( 
.A1(n_1724),
.A2(n_1708),
.B(n_1690),
.Y(n_1738)
);

AOI21xp5_ASAP7_75t_L g1739 ( 
.A1(n_1727),
.A2(n_1716),
.B(n_1717),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1728),
.Y(n_1740)
);

AOI211x1_ASAP7_75t_L g1741 ( 
.A1(n_1732),
.A2(n_1714),
.B(n_1711),
.C(n_1719),
.Y(n_1741)
);

AOI221xp5_ASAP7_75t_L g1742 ( 
.A1(n_1730),
.A2(n_1714),
.B1(n_1718),
.B2(n_1723),
.C(n_1702),
.Y(n_1742)
);

O2A1O1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1733),
.A2(n_1672),
.B(n_1649),
.C(n_1721),
.Y(n_1743)
);

AOI221xp5_ASAP7_75t_L g1744 ( 
.A1(n_1734),
.A2(n_1649),
.B1(n_1641),
.B2(n_1618),
.C(n_1670),
.Y(n_1744)
);

INVx3_ASAP7_75t_SL g1745 ( 
.A(n_1734),
.Y(n_1745)
);

OAI21xp33_ASAP7_75t_L g1746 ( 
.A1(n_1738),
.A2(n_1672),
.B(n_1618),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1740),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1736),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1741),
.Y(n_1749)
);

OAI21xp33_ASAP7_75t_SL g1750 ( 
.A1(n_1744),
.A2(n_1624),
.B(n_1642),
.Y(n_1750)
);

A2O1A1Ixp33_ASAP7_75t_L g1751 ( 
.A1(n_1743),
.A2(n_1618),
.B(n_1620),
.C(n_1621),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1749),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1748),
.B(n_1737),
.Y(n_1753)
);

XNOR2x1_ASAP7_75t_L g1754 ( 
.A(n_1747),
.B(n_1735),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1746),
.Y(n_1755)
);

NAND2x1p5_ASAP7_75t_L g1756 ( 
.A(n_1751),
.B(n_1739),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1750),
.Y(n_1757)
);

AOI22x1_ASAP7_75t_L g1758 ( 
.A1(n_1756),
.A2(n_1745),
.B1(n_1742),
.B2(n_1620),
.Y(n_1758)
);

NOR2xp33_ASAP7_75t_R g1759 ( 
.A(n_1753),
.B(n_1565),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1752),
.Y(n_1760)
);

AOI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1757),
.A2(n_1755),
.B1(n_1754),
.B2(n_1752),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1754),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1762),
.B(n_1635),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1761),
.B(n_1621),
.Y(n_1764)
);

AND3x2_ASAP7_75t_L g1765 ( 
.A(n_1760),
.B(n_1758),
.C(n_1759),
.Y(n_1765)
);

HB1xp67_ASAP7_75t_L g1766 ( 
.A(n_1764),
.Y(n_1766)
);

AOI322xp5_ASAP7_75t_L g1767 ( 
.A1(n_1766),
.A2(n_1763),
.A3(n_1765),
.B1(n_1603),
.B2(n_1635),
.C1(n_1622),
.C2(n_1623),
.Y(n_1767)
);

NOR3xp33_ASAP7_75t_SL g1768 ( 
.A(n_1767),
.B(n_1617),
.C(n_1524),
.Y(n_1768)
);

BUFx2_ASAP7_75t_L g1769 ( 
.A(n_1767),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1769),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1768),
.Y(n_1771)
);

OAI22x1_ASAP7_75t_L g1772 ( 
.A1(n_1770),
.A2(n_1610),
.B1(n_1616),
.B2(n_1603),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1772),
.Y(n_1773)
);

AOI21xp5_ASAP7_75t_L g1774 ( 
.A1(n_1773),
.A2(n_1771),
.B(n_1603),
.Y(n_1774)
);

NOR2xp67_ASAP7_75t_L g1775 ( 
.A(n_1774),
.B(n_1651),
.Y(n_1775)
);

AO21x2_ASAP7_75t_L g1776 ( 
.A1(n_1775),
.A2(n_1616),
.B(n_1610),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1776),
.A2(n_1629),
.B1(n_1627),
.B2(n_1626),
.Y(n_1777)
);

AOI211xp5_ASAP7_75t_L g1778 ( 
.A1(n_1777),
.A2(n_1615),
.B(n_1626),
.C(n_1640),
.Y(n_1778)
);


endmodule