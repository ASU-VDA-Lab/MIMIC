module fake_netlist_1_3802_n_514 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_75, n_19, n_61, n_21, n_6, n_4, n_74, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_514);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_75;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_74;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_514;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g76 ( .A(n_33), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_60), .Y(n_77) );
INVxp33_ASAP7_75t_SL g78 ( .A(n_41), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_12), .Y(n_79) );
INVxp67_ASAP7_75t_SL g80 ( .A(n_65), .Y(n_80) );
BUFx6f_ASAP7_75t_L g81 ( .A(n_48), .Y(n_81) );
BUFx2_ASAP7_75t_SL g82 ( .A(n_1), .Y(n_82) );
BUFx3_ASAP7_75t_L g83 ( .A(n_17), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_24), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_13), .Y(n_85) );
CKINVDCx5p33_ASAP7_75t_R g86 ( .A(n_22), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
CKINVDCx5p33_ASAP7_75t_R g88 ( .A(n_75), .Y(n_88) );
HB1xp67_ASAP7_75t_L g89 ( .A(n_14), .Y(n_89) );
INVx1_ASAP7_75t_L g90 ( .A(n_39), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_26), .Y(n_91) );
BUFx10_ASAP7_75t_L g92 ( .A(n_72), .Y(n_92) );
INVxp67_ASAP7_75t_SL g93 ( .A(n_13), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_35), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_54), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_36), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_67), .Y(n_97) );
INVxp67_ASAP7_75t_L g98 ( .A(n_34), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_12), .Y(n_99) );
BUFx2_ASAP7_75t_SL g100 ( .A(n_32), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_52), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_28), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_38), .Y(n_104) );
INVx2_ASAP7_75t_L g105 ( .A(n_49), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_27), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_11), .Y(n_107) );
BUFx2_ASAP7_75t_L g108 ( .A(n_10), .Y(n_108) );
INVxp33_ASAP7_75t_SL g109 ( .A(n_2), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_58), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_42), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_51), .Y(n_112) );
INVxp67_ASAP7_75t_L g113 ( .A(n_62), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_66), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_76), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_76), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_81), .Y(n_117) );
BUFx6f_ASAP7_75t_L g118 ( .A(n_81), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_77), .Y(n_119) );
INVx2_ASAP7_75t_L g120 ( .A(n_105), .Y(n_120) );
INVx2_ASAP7_75t_L g121 ( .A(n_105), .Y(n_121) );
INVx3_ASAP7_75t_L g122 ( .A(n_92), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_112), .Y(n_123) );
INVx2_ASAP7_75t_L g124 ( .A(n_81), .Y(n_124) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_81), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_92), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_81), .Y(n_127) );
HB1xp67_ASAP7_75t_L g128 ( .A(n_108), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_77), .Y(n_129) );
CKINVDCx20_ASAP7_75t_R g130 ( .A(n_108), .Y(n_130) );
NOR2xp67_ASAP7_75t_L g131 ( .A(n_98), .B(n_113), .Y(n_131) );
NOR2xp33_ASAP7_75t_L g132 ( .A(n_109), .B(n_0), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_89), .B(n_0), .Y(n_133) );
AND2x2_ASAP7_75t_L g134 ( .A(n_92), .B(n_1), .Y(n_134) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_92), .B(n_2), .Y(n_135) );
NAND2xp5_ASAP7_75t_SL g136 ( .A(n_115), .B(n_110), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_122), .B(n_83), .Y(n_137) );
NAND2x1p5_ASAP7_75t_L g138 ( .A(n_134), .B(n_79), .Y(n_138) );
AO22x2_ASAP7_75t_L g139 ( .A1(n_134), .A2(n_82), .B1(n_79), .B2(n_85), .Y(n_139) );
AOI22xp5_ASAP7_75t_L g140 ( .A1(n_128), .A2(n_85), .B1(n_103), .B2(n_99), .Y(n_140) );
CKINVDCx16_ASAP7_75t_R g141 ( .A(n_130), .Y(n_141) );
AND2x4_ASAP7_75t_L g142 ( .A(n_122), .B(n_83), .Y(n_142) );
INVx1_ASAP7_75t_L g143 ( .A(n_115), .Y(n_143) );
AND2x4_ASAP7_75t_L g144 ( .A(n_122), .B(n_99), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_116), .Y(n_145) );
INVxp67_ASAP7_75t_L g146 ( .A(n_133), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_116), .Y(n_147) );
BUFx3_ASAP7_75t_L g148 ( .A(n_122), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_131), .B(n_103), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_131), .B(n_86), .Y(n_150) );
AOI22xp5_ASAP7_75t_L g151 ( .A1(n_133), .A2(n_78), .B1(n_91), .B2(n_107), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_117), .Y(n_152) );
INVx1_ASAP7_75t_L g153 ( .A(n_119), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g154 ( .A1(n_126), .A2(n_93), .B1(n_82), .B2(n_84), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_119), .B(n_110), .Y(n_156) );
AND2x4_ASAP7_75t_L g157 ( .A(n_129), .B(n_97), .Y(n_157) );
NAND3x1_ASAP7_75t_L g158 ( .A(n_132), .B(n_84), .C(n_87), .Y(n_158) );
BUFx6f_ASAP7_75t_L g159 ( .A(n_118), .Y(n_159) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_143), .B(n_129), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_145), .Y(n_161) );
CKINVDCx5p33_ASAP7_75t_R g162 ( .A(n_141), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_157), .B(n_88), .Y(n_163) );
INVx2_ASAP7_75t_SL g164 ( .A(n_157), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_147), .Y(n_165) );
BUFx3_ASAP7_75t_L g166 ( .A(n_148), .Y(n_166) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_153), .B(n_144), .Y(n_167) );
OAI221xp5_ASAP7_75t_L g168 ( .A1(n_140), .A2(n_135), .B1(n_120), .B2(n_121), .C(n_80), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_152), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_148), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_144), .B(n_95), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_151), .Y(n_172) );
CKINVDCx5p33_ASAP7_75t_R g173 ( .A(n_154), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_159), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_155), .Y(n_176) );
INVx2_ASAP7_75t_SL g177 ( .A(n_138), .Y(n_177) );
AND2x4_ASAP7_75t_L g178 ( .A(n_144), .B(n_120), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_155), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_159), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_159), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
OR2x2_ASAP7_75t_L g183 ( .A(n_138), .B(n_146), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_146), .B(n_137), .Y(n_184) );
AND2x4_ASAP7_75t_L g185 ( .A(n_149), .B(n_121), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_159), .Y(n_186) );
NOR3xp33_ASAP7_75t_SL g187 ( .A(n_150), .B(n_123), .C(n_114), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_139), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_142), .Y(n_190) );
CKINVDCx11_ASAP7_75t_R g191 ( .A(n_162), .Y(n_191) );
BUFx2_ASAP7_75t_L g192 ( .A(n_177), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_177), .Y(n_193) );
INVx5_ASAP7_75t_L g194 ( .A(n_166), .Y(n_194) );
BUFx3_ASAP7_75t_L g195 ( .A(n_166), .Y(n_195) );
BUFx4_ASAP7_75t_SL g196 ( .A(n_183), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g197 ( .A(n_166), .B(n_136), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g198 ( .A(n_183), .B(n_149), .Y(n_198) );
AOI22xp5_ASAP7_75t_L g199 ( .A1(n_189), .A2(n_139), .B1(n_158), .B2(n_156), .Y(n_199) );
BUFx3_ASAP7_75t_L g200 ( .A(n_170), .Y(n_200) );
INVxp67_ASAP7_75t_L g201 ( .A(n_184), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_169), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_161), .Y(n_203) );
HB1xp67_ASAP7_75t_L g204 ( .A(n_164), .Y(n_204) );
BUFx10_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
CKINVDCx20_ASAP7_75t_R g206 ( .A(n_187), .Y(n_206) );
INVx1_ASAP7_75t_SL g207 ( .A(n_184), .Y(n_207) );
OAI22xp5_ASAP7_75t_L g208 ( .A1(n_167), .A2(n_139), .B1(n_156), .B2(n_136), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_160), .B(n_149), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g210 ( .A1(n_161), .A2(n_102), .B(n_87), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_174), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_174), .Y(n_212) );
BUFx2_ASAP7_75t_L g213 ( .A(n_178), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_165), .Y(n_214) );
BUFx3_ASAP7_75t_L g215 ( .A(n_170), .Y(n_215) );
BUFx3_ASAP7_75t_L g216 ( .A(n_188), .Y(n_216) );
BUFx6f_ASAP7_75t_L g217 ( .A(n_174), .Y(n_217) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_167), .B(n_101), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_169), .Y(n_219) );
AO21x2_ASAP7_75t_L g220 ( .A1(n_165), .A2(n_104), .B(n_90), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_188), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_194), .Y(n_222) );
INVx3_ASAP7_75t_L g223 ( .A(n_194), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_196), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_207), .B(n_185), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g226 ( .A(n_194), .B(n_178), .Y(n_226) );
AND2x2_ASAP7_75t_L g227 ( .A(n_207), .B(n_160), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_211), .Y(n_228) );
AO21x1_ASAP7_75t_L g229 ( .A1(n_208), .A2(n_203), .B(n_214), .Y(n_229) );
AND2x2_ASAP7_75t_L g230 ( .A(n_209), .B(n_178), .Y(n_230) );
OAI22xp5_ASAP7_75t_L g231 ( .A1(n_208), .A2(n_178), .B1(n_188), .B2(n_190), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_203), .Y(n_232) );
CKINVDCx5p33_ASAP7_75t_R g233 ( .A(n_191), .Y(n_233) );
INVx2_ASAP7_75t_L g234 ( .A(n_202), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_201), .B(n_185), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_214), .Y(n_236) );
BUFx2_ASAP7_75t_L g237 ( .A(n_192), .Y(n_237) );
INVx2_ASAP7_75t_SL g238 ( .A(n_205), .Y(n_238) );
AO22x2_ASAP7_75t_L g239 ( .A1(n_216), .A2(n_190), .B1(n_182), .B2(n_185), .Y(n_239) );
OR2x2_ASAP7_75t_L g240 ( .A(n_209), .B(n_172), .Y(n_240) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_192), .Y(n_241) );
AND2x4_ASAP7_75t_L g242 ( .A(n_193), .B(n_182), .Y(n_242) );
OAI22xp5_ASAP7_75t_L g243 ( .A1(n_199), .A2(n_185), .B1(n_168), .B2(n_90), .Y(n_243) );
AND2x2_ASAP7_75t_L g244 ( .A(n_202), .B(n_163), .Y(n_244) );
INVx4_ASAP7_75t_L g245 ( .A(n_194), .Y(n_245) );
AOI22xp33_ASAP7_75t_SL g246 ( .A1(n_193), .A2(n_173), .B1(n_171), .B2(n_100), .Y(n_246) );
OAI22xp5_ASAP7_75t_L g247 ( .A1(n_199), .A2(n_175), .B1(n_169), .B2(n_176), .Y(n_247) );
AND2x4_ASAP7_75t_L g248 ( .A(n_222), .B(n_213), .Y(n_248) );
AND2x2_ASAP7_75t_L g249 ( .A(n_240), .B(n_198), .Y(n_249) );
OAI221xp5_ASAP7_75t_L g250 ( .A1(n_240), .A2(n_204), .B1(n_218), .B2(n_213), .C(n_210), .Y(n_250) );
OAI22xp33_ASAP7_75t_L g251 ( .A1(n_224), .A2(n_206), .B1(n_202), .B2(n_219), .Y(n_251) );
AOI22xp33_ASAP7_75t_SL g252 ( .A1(n_237), .A2(n_220), .B1(n_100), .B2(n_205), .Y(n_252) );
OAI22xp5_ASAP7_75t_L g253 ( .A1(n_231), .A2(n_219), .B1(n_221), .B2(n_216), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g254 ( .A1(n_243), .A2(n_221), .B1(n_216), .B2(n_220), .Y(n_254) );
AND2x4_ASAP7_75t_L g255 ( .A(n_227), .B(n_194), .Y(n_255) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_229), .A2(n_220), .B(n_219), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_227), .B(n_221), .Y(n_257) );
OAI22xp5_ASAP7_75t_L g258 ( .A1(n_231), .A2(n_200), .B1(n_215), .B2(n_194), .Y(n_258) );
OAI211xp5_ASAP7_75t_SL g259 ( .A1(n_246), .A2(n_94), .B(n_96), .C(n_97), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_232), .Y(n_260) );
BUFx12f_ASAP7_75t_L g261 ( .A(n_233), .Y(n_261) );
INVx2_ASAP7_75t_L g262 ( .A(n_234), .Y(n_262) );
OAI22xp33_ASAP7_75t_L g263 ( .A1(n_237), .A2(n_215), .B1(n_200), .B2(n_194), .Y(n_263) );
AOI22xp5_ASAP7_75t_L g264 ( .A1(n_243), .A2(n_205), .B1(n_220), .B2(n_215), .Y(n_264) );
INVx2_ASAP7_75t_L g265 ( .A(n_234), .Y(n_265) );
AOI22xp5_ASAP7_75t_L g266 ( .A1(n_230), .A2(n_205), .B1(n_200), .B2(n_195), .Y(n_266) );
AOI22xp33_ASAP7_75t_L g267 ( .A1(n_229), .A2(n_195), .B1(n_197), .B2(n_96), .Y(n_267) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_230), .A2(n_195), .B1(n_197), .B2(n_179), .Y(n_268) );
NOR2xp33_ASAP7_75t_L g269 ( .A(n_235), .B(n_197), .Y(n_269) );
AND2x2_ASAP7_75t_L g270 ( .A(n_262), .B(n_234), .Y(n_270) );
AND2x4_ASAP7_75t_L g271 ( .A(n_262), .B(n_232), .Y(n_271) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_255), .Y(n_272) );
NAND4xp25_ASAP7_75t_SL g273 ( .A(n_250), .B(n_236), .C(n_102), .D(n_104), .Y(n_273) );
NAND4xp25_ASAP7_75t_SL g274 ( .A(n_249), .B(n_236), .C(n_106), .D(n_94), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_260), .Y(n_275) );
INVx2_ASAP7_75t_SL g276 ( .A(n_255), .Y(n_276) );
BUFx3_ASAP7_75t_L g277 ( .A(n_248), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g278 ( .A(n_251), .B(n_241), .Y(n_278) );
OAI221xp5_ASAP7_75t_L g279 ( .A1(n_259), .A2(n_225), .B1(n_226), .B2(n_244), .C(n_247), .Y(n_279) );
AND2x2_ASAP7_75t_L g280 ( .A(n_265), .B(n_239), .Y(n_280) );
OR2x2_ASAP7_75t_L g281 ( .A(n_257), .B(n_226), .Y(n_281) );
BUFx5_ASAP7_75t_L g282 ( .A(n_248), .Y(n_282) );
OAI21xp33_ASAP7_75t_SL g283 ( .A1(n_264), .A2(n_254), .B(n_267), .Y(n_283) );
OAI21x1_ASAP7_75t_L g284 ( .A1(n_267), .A2(n_223), .B(n_226), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_265), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_269), .B(n_244), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_248), .B(n_242), .Y(n_287) );
OR2x2_ASAP7_75t_L g288 ( .A(n_256), .B(n_242), .Y(n_288) );
AOI33xp33_ASAP7_75t_L g289 ( .A1(n_254), .A2(n_106), .A3(n_124), .B1(n_117), .B2(n_127), .B3(n_242), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_253), .A2(n_223), .B(n_124), .Y(n_290) );
OA21x2_ASAP7_75t_L g291 ( .A1(n_290), .A2(n_268), .B(n_269), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_275), .Y(n_292) );
OAI31xp33_ASAP7_75t_L g293 ( .A1(n_273), .A2(n_263), .A3(n_239), .B(n_258), .Y(n_293) );
OAI21xp33_ASAP7_75t_SL g294 ( .A1(n_284), .A2(n_222), .B(n_245), .Y(n_294) );
AND2x2_ASAP7_75t_L g295 ( .A(n_280), .B(n_256), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_275), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_280), .B(n_239), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_288), .Y(n_298) );
OAI31xp33_ASAP7_75t_L g299 ( .A1(n_274), .A2(n_239), .A3(n_242), .B(n_238), .Y(n_299) );
AOI21xp5_ASAP7_75t_L g300 ( .A1(n_285), .A2(n_228), .B(n_239), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_286), .B(n_252), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_285), .Y(n_302) );
AND2x2_ASAP7_75t_L g303 ( .A(n_270), .B(n_223), .Y(n_303) );
AOI211xp5_ASAP7_75t_L g304 ( .A1(n_278), .A2(n_81), .B(n_111), .C(n_266), .Y(n_304) );
AOI221xp5_ASAP7_75t_L g305 ( .A1(n_283), .A2(n_111), .B1(n_124), .B2(n_127), .C(n_125), .Y(n_305) );
AOI33xp33_ASAP7_75t_L g306 ( .A1(n_276), .A2(n_127), .A3(n_4), .B1(n_5), .B2(n_6), .B3(n_7), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_288), .Y(n_307) );
AND2x2_ASAP7_75t_L g308 ( .A(n_270), .B(n_223), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_271), .B(n_222), .Y(n_309) );
AND2x2_ASAP7_75t_L g310 ( .A(n_271), .B(n_222), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_271), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_271), .B(n_245), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_284), .Y(n_313) );
AND2x2_ASAP7_75t_L g314 ( .A(n_282), .B(n_245), .Y(n_314) );
OAI21xp5_ASAP7_75t_SL g315 ( .A1(n_279), .A2(n_238), .B(n_111), .Y(n_315) );
AND2x2_ASAP7_75t_L g316 ( .A(n_282), .B(n_245), .Y(n_316) );
INVx3_ASAP7_75t_L g317 ( .A(n_290), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_276), .B(n_261), .Y(n_318) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_289), .B(n_175), .C(n_176), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_295), .B(n_283), .Y(n_320) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_314), .Y(n_321) );
NOR2xp67_ASAP7_75t_L g322 ( .A(n_315), .B(n_261), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_292), .Y(n_323) );
NOR2xp33_ASAP7_75t_L g324 ( .A(n_318), .B(n_272), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_295), .B(n_282), .Y(n_325) );
AND2x2_ASAP7_75t_L g326 ( .A(n_298), .B(n_282), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_292), .B(n_286), .Y(n_327) );
NAND2xp33_ASAP7_75t_SL g328 ( .A(n_306), .B(n_281), .Y(n_328) );
OR2x2_ASAP7_75t_L g329 ( .A(n_298), .B(n_277), .Y(n_329) );
INVx5_ASAP7_75t_L g330 ( .A(n_317), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_307), .B(n_282), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_307), .B(n_282), .Y(n_332) );
OR2x2_ASAP7_75t_L g333 ( .A(n_311), .B(n_277), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_296), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_311), .B(n_282), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_302), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_302), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_297), .B(n_302), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_297), .B(n_277), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_301), .B(n_281), .Y(n_341) );
OR2x2_ASAP7_75t_L g342 ( .A(n_300), .B(n_287), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_313), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_303), .B(n_111), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_301), .B(n_3), .Y(n_345) );
NOR3xp33_ASAP7_75t_L g346 ( .A(n_315), .B(n_175), .C(n_176), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_317), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_317), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_317), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_303), .B(n_111), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_308), .B(n_111), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_309), .B(n_3), .Y(n_352) );
NOR2x1_ASAP7_75t_L g353 ( .A(n_300), .B(n_228), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_308), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_294), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_309), .B(n_125), .Y(n_356) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_314), .B(n_228), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_310), .Y(n_358) );
AOI21xp5_ASAP7_75t_L g359 ( .A1(n_304), .A2(n_228), .B(n_217), .Y(n_359) );
AOI22xp5_ASAP7_75t_L g360 ( .A1(n_304), .A2(n_228), .B1(n_179), .B2(n_118), .Y(n_360) );
AOI21xp33_ASAP7_75t_L g361 ( .A1(n_322), .A2(n_299), .B(n_293), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_336), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_320), .B(n_305), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_323), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_323), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_336), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_320), .B(n_305), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_334), .Y(n_368) );
AOI211xp5_ASAP7_75t_SL g369 ( .A1(n_346), .A2(n_316), .B(n_312), .C(n_310), .Y(n_369) );
OR2x2_ASAP7_75t_L g370 ( .A(n_358), .B(n_312), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g371 ( .A1(n_328), .A2(n_293), .B1(n_299), .B2(n_316), .Y(n_371) );
OR2x2_ASAP7_75t_L g372 ( .A(n_358), .B(n_291), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_344), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_334), .Y(n_374) );
OAI21xp5_ASAP7_75t_L g375 ( .A1(n_360), .A2(n_294), .B(n_319), .Y(n_375) );
OAI22xp5_ASAP7_75t_L g376 ( .A1(n_321), .A2(n_291), .B1(n_319), .B2(n_228), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_344), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_353), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_350), .Y(n_379) );
AOI32xp33_ASAP7_75t_L g380 ( .A1(n_350), .A2(n_4), .A3(n_5), .B1(n_6), .B2(n_8), .Y(n_380) );
NOR3xp33_ASAP7_75t_L g381 ( .A(n_345), .B(n_8), .C(n_9), .Y(n_381) );
AOI322xp5_ASAP7_75t_L g382 ( .A1(n_341), .A2(n_9), .A3(n_10), .B1(n_11), .B2(n_14), .C1(n_15), .C2(n_16), .Y(n_382) );
OR2x2_ASAP7_75t_L g383 ( .A(n_354), .B(n_291), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_351), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_327), .B(n_291), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g387 ( .A(n_338), .B(n_125), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_354), .Y(n_388) );
AOI21xp5_ASAP7_75t_L g389 ( .A1(n_359), .A2(n_217), .B(n_212), .Y(n_389) );
INVx2_ASAP7_75t_L g390 ( .A(n_337), .Y(n_390) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_338), .B(n_125), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_329), .Y(n_392) );
OAI22xp5_ASAP7_75t_L g393 ( .A1(n_321), .A2(n_15), .B1(n_16), .B2(n_17), .Y(n_393) );
OAI22xp5_ASAP7_75t_L g394 ( .A1(n_342), .A2(n_217), .B1(n_212), .B2(n_211), .Y(n_394) );
AOI221x1_ASAP7_75t_L g395 ( .A1(n_356), .A2(n_125), .B1(n_118), .B2(n_211), .C(n_217), .Y(n_395) );
AOI22xp5_ASAP7_75t_L g396 ( .A1(n_324), .A2(n_118), .B1(n_125), .B2(n_211), .Y(n_396) );
NAND3xp33_ASAP7_75t_L g397 ( .A(n_356), .B(n_118), .C(n_212), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_325), .B(n_118), .Y(n_398) );
NOR2xp33_ASAP7_75t_R g399 ( .A(n_352), .B(n_18), .Y(n_399) );
OAI21xp33_ASAP7_75t_L g400 ( .A1(n_355), .A2(n_179), .B(n_181), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_339), .B(n_19), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_339), .B(n_20), .Y(n_402) );
OA21x2_ASAP7_75t_L g403 ( .A1(n_355), .A2(n_181), .B(n_180), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_326), .Y(n_404) );
INVx3_ASAP7_75t_L g405 ( .A(n_330), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_326), .Y(n_406) );
OAI22xp33_ASAP7_75t_L g407 ( .A1(n_342), .A2(n_217), .B1(n_212), .B2(n_211), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_331), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_388), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_364), .Y(n_410) );
AOI21xp33_ASAP7_75t_SL g411 ( .A1(n_361), .A2(n_357), .B(n_333), .Y(n_411) );
OR2x2_ASAP7_75t_L g412 ( .A(n_370), .B(n_325), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_368), .Y(n_414) );
NOR4xp25_ASAP7_75t_SL g415 ( .A(n_361), .B(n_343), .C(n_353), .D(n_330), .Y(n_415) );
XOR2xp5_ASAP7_75t_L g416 ( .A(n_393), .B(n_340), .Y(n_416) );
XNOR2xp5_ASAP7_75t_L g417 ( .A(n_371), .B(n_340), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_374), .Y(n_418) );
XOR2x2_ASAP7_75t_L g419 ( .A(n_369), .B(n_357), .Y(n_419) );
INVxp67_ASAP7_75t_L g420 ( .A(n_398), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_399), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_392), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_387), .Y(n_423) );
XOR2xp5_ASAP7_75t_L g424 ( .A(n_404), .B(n_356), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_387), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_408), .B(n_331), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_391), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_391), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_377), .B(n_332), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_362), .Y(n_430) );
OAI211xp5_ASAP7_75t_L g431 ( .A1(n_380), .A2(n_330), .B(n_332), .C(n_335), .Y(n_431) );
NOR2xp33_ASAP7_75t_R g432 ( .A(n_405), .B(n_330), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_366), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_390), .Y(n_434) );
NAND2xp5_ASAP7_75t_SL g435 ( .A(n_405), .B(n_330), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_406), .B(n_335), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_373), .B(n_357), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_379), .B(n_343), .Y(n_438) );
NOR2xp33_ASAP7_75t_R g439 ( .A(n_363), .B(n_330), .Y(n_439) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_381), .A2(n_385), .B1(n_367), .B2(n_363), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_384), .Y(n_441) );
OAI311xp33_ASAP7_75t_L g442 ( .A1(n_382), .A2(n_356), .A3(n_349), .B1(n_348), .C1(n_347), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_383), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_372), .B(n_349), .Y(n_444) );
OAI21xp33_ASAP7_75t_L g445 ( .A1(n_386), .A2(n_348), .B(n_347), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_386), .B(n_21), .Y(n_446) );
NOR3xp33_ASAP7_75t_L g447 ( .A(n_381), .B(n_181), .C(n_180), .Y(n_447) );
INVx1_ASAP7_75t_SL g448 ( .A(n_397), .Y(n_448) );
AOI22xp33_ASAP7_75t_SL g449 ( .A1(n_375), .A2(n_217), .B1(n_212), .B2(n_211), .Y(n_449) );
AOI22xp5_ASAP7_75t_L g450 ( .A1(n_440), .A2(n_367), .B1(n_376), .B2(n_378), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g451 ( .A1(n_431), .A2(n_378), .B1(n_394), .B2(n_396), .Y(n_451) );
NOR2xp33_ASAP7_75t_L g452 ( .A(n_421), .B(n_402), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_443), .B(n_403), .Y(n_453) );
INVxp67_ASAP7_75t_SL g454 ( .A(n_420), .Y(n_454) );
NOR2xp33_ASAP7_75t_L g455 ( .A(n_417), .B(n_402), .Y(n_455) );
INVxp67_ASAP7_75t_SL g456 ( .A(n_420), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_431), .A2(n_400), .B1(n_407), .B2(n_401), .Y(n_457) );
AOI22xp33_ASAP7_75t_L g458 ( .A1(n_419), .A2(n_401), .B1(n_389), .B2(n_212), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_439), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_439), .Y(n_460) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_435), .B(n_389), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_409), .Y(n_462) );
NOR2x1p5_ASAP7_75t_L g463 ( .A(n_412), .B(n_395), .Y(n_463) );
AOI211xp5_ASAP7_75t_L g464 ( .A1(n_442), .A2(n_23), .B(n_25), .C(n_29), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_434), .Y(n_465) );
INVxp67_ASAP7_75t_L g466 ( .A(n_422), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g467 ( .A1(n_435), .A2(n_180), .B(n_31), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_410), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g469 ( .A(n_447), .B(n_30), .C(n_37), .D(n_40), .Y(n_469) );
NAND3xp33_ASAP7_75t_L g470 ( .A(n_411), .B(n_186), .C(n_174), .Y(n_470) );
AOI222xp33_ASAP7_75t_L g471 ( .A1(n_423), .A2(n_43), .B1(n_44), .B2(n_45), .C1(n_46), .C2(n_47), .Y(n_471) );
OR2x2_ASAP7_75t_L g472 ( .A(n_426), .B(n_50), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g473 ( .A1(n_415), .A2(n_55), .B(n_56), .Y(n_473) );
AOI22x1_ASAP7_75t_L g474 ( .A1(n_416), .A2(n_57), .B1(n_59), .B2(n_61), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_413), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_432), .B(n_186), .Y(n_476) );
NAND2xp5_ASAP7_75t_SL g477 ( .A(n_459), .B(n_432), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_460), .B(n_449), .Y(n_478) );
NOR2xp67_ASAP7_75t_L g479 ( .A(n_470), .B(n_445), .Y(n_479) );
INVxp67_ASAP7_75t_SL g480 ( .A(n_463), .Y(n_480) );
AOI221xp5_ASAP7_75t_L g481 ( .A1(n_454), .A2(n_447), .B1(n_441), .B2(n_414), .C(n_418), .Y(n_481) );
NAND2xp33_ASAP7_75t_SL g482 ( .A(n_458), .B(n_437), .Y(n_482) );
AOI22xp5_ASAP7_75t_L g483 ( .A1(n_455), .A2(n_424), .B1(n_429), .B2(n_428), .Y(n_483) );
BUFx2_ASAP7_75t_L g484 ( .A(n_465), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_456), .B(n_425), .Y(n_485) );
OAI22xp33_ASAP7_75t_L g486 ( .A1(n_450), .A2(n_448), .B1(n_427), .B2(n_438), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_462), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_466), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_476), .A2(n_449), .B(n_430), .Y(n_489) );
INVx1_ASAP7_75t_SL g490 ( .A(n_472), .Y(n_490) );
OAI211xp5_ASAP7_75t_SL g491 ( .A1(n_464), .A2(n_433), .B(n_446), .C(n_68), .Y(n_491) );
AOI22xp5_ASAP7_75t_L g492 ( .A1(n_452), .A2(n_444), .B1(n_436), .B2(n_186), .Y(n_492) );
NOR2x1_ASAP7_75t_L g493 ( .A(n_469), .B(n_63), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g494 ( .A(n_473), .B(n_64), .C(n_69), .Y(n_494) );
NAND4xp25_ASAP7_75t_SL g495 ( .A(n_461), .B(n_70), .C(n_71), .D(n_73), .Y(n_495) );
OAI322xp33_ASAP7_75t_L g496 ( .A1(n_453), .A2(n_74), .A3(n_174), .B1(n_186), .B2(n_475), .C1(n_468), .C2(n_451), .Y(n_496) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_473), .B(n_174), .C(n_186), .Y(n_497) );
OAI22xp5_ASAP7_75t_L g498 ( .A1(n_457), .A2(n_186), .B1(n_474), .B2(n_467), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_467), .A2(n_460), .B(n_459), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_471), .Y(n_500) );
OA22x2_ASAP7_75t_L g501 ( .A1(n_480), .A2(n_500), .B1(n_477), .B2(n_483), .Y(n_501) );
NAND4xp25_ASAP7_75t_L g502 ( .A(n_499), .B(n_493), .C(n_494), .D(n_491), .Y(n_502) );
HB1xp67_ASAP7_75t_L g503 ( .A(n_484), .Y(n_503) );
CKINVDCx5p33_ASAP7_75t_R g504 ( .A(n_488), .Y(n_504) );
NOR3xp33_ASAP7_75t_L g505 ( .A(n_498), .B(n_496), .C(n_478), .Y(n_505) );
AO22x2_ASAP7_75t_L g506 ( .A1(n_505), .A2(n_487), .B1(n_490), .B2(n_485), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g507 ( .A1(n_501), .A2(n_482), .B1(n_486), .B2(n_479), .Y(n_507) );
NOR3xp33_ASAP7_75t_L g508 ( .A(n_502), .B(n_495), .C(n_491), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_506), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_507), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_509), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g512 ( .A1(n_510), .A2(n_508), .B1(n_504), .B2(n_503), .Y(n_512) );
OAI211xp5_ASAP7_75t_L g513 ( .A1(n_512), .A2(n_481), .B(n_497), .C(n_492), .Y(n_513) );
AOI21xp5_ASAP7_75t_L g514 ( .A1(n_513), .A2(n_511), .B(n_489), .Y(n_514) );
endmodule