module fake_netlist_6_2880_n_915 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_915);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_915;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_853;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_909;
wire n_580;
wire n_762;
wire n_881;
wire n_875;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_760;
wire n_741;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_341;
wire n_362;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_671;
wire n_726;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_874;
wire n_724;
wire n_382;
wire n_673;
wire n_628;
wire n_883;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_898;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_865;
wire n_893;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_892;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_894;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_873;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_872;
wire n_198;
wire n_222;
wire n_300;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_852;
wire n_667;
wire n_229;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_901;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_510;
wire n_837;
wire n_836;
wire n_863;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_895;
wire n_866;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_761;
wire n_785;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_516;
wire n_720;
wire n_758;
wire n_525;
wire n_842;
wire n_611;
wire n_491;
wire n_878;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_899;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_844;
wire n_343;
wire n_448;
wire n_886;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_888;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_910;
wire n_486;
wire n_911;
wire n_381;
wire n_236;
wire n_653;
wire n_887;
wire n_752;
wire n_908;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_907;
wire n_854;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_870;
wire n_366;
wire n_904;
wire n_777;
wire n_407;
wire n_913;
wire n_450;
wire n_808;
wire n_867;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_552;
wire n_619;
wire n_885;
wire n_216;
wire n_455;
wire n_896;
wire n_521;
wire n_363;
wire n_572;
wire n_912;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_884;
wire n_599;
wire n_513;
wire n_855;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_868;
wire n_570;
wire n_731;
wire n_859;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_527;
wire n_474;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_394;
wire n_312;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_880;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_889;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_860;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_864;
wire n_879;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_905;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_386;
wire n_201;
wire n_249;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_849;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_882;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_861;
wire n_674;
wire n_857;
wire n_871;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_902;
wire n_333;
wire n_588;
wire n_215;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_914;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_497;
wire n_285;
wire n_780;
wire n_773;
wire n_675;
wire n_903;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_850;
wire n_401;
wire n_324;
wire n_766;
wire n_816;
wire n_743;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_877;
wire n_205;
wire n_604;
wire n_848;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_876;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_906;
wire n_722;
wire n_688;
wire n_862;
wire n_351;
wire n_869;
wire n_437;
wire n_259;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_697;
wire n_687;
wire n_364;
wire n_890;
wire n_637;
wire n_385;
wire n_295;
wire n_701;
wire n_817;
wire n_629;
wire n_388;
wire n_190;
wire n_858;
wire n_484;
wire n_262;
wire n_613;
wire n_736;
wire n_187;
wire n_897;
wire n_900;
wire n_846;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_332;
wire n_891;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx5p33_ASAP7_75t_R g185 ( 
.A(n_135),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_157),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_33),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_115),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_57),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_56),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_116),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_79),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_91),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_15),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_149),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_47),
.Y(n_196)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_177),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_97),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_62),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_131),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_167),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_166),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_76),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_172),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_28),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_19),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_109),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_77),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_68),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_159),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_160),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_125),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_22),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_27),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_70),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_3),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_95),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_144),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_119),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_72),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_105),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_64),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g225 ( 
.A(n_83),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_170),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_113),
.Y(n_227)
);

BUFx2_ASAP7_75t_L g228 ( 
.A(n_25),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_81),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_67),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_42),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_37),
.Y(n_232)
);

INVx1_ASAP7_75t_SL g233 ( 
.A(n_85),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_114),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_155),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_4),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_65),
.Y(n_237)
);

INVx1_ASAP7_75t_SL g238 ( 
.A(n_8),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_3),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_139),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_17),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_98),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_133),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_182),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g245 ( 
.A(n_43),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_143),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_18),
.Y(n_247)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_121),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_124),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_148),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_110),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_99),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_96),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_147),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_130),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_92),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_93),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_7),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_120),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_141),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_104),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_127),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_1),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_78),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_24),
.Y(n_267)
);

INVx1_ASAP7_75t_SL g268 ( 
.A(n_136),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_108),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_94),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_58),
.Y(n_271)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_180),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_163),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_129),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_71),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_32),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_0),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_50),
.Y(n_278)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_156),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_277),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_206),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_185),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_186),
.Y(n_283)
);

NOR2xp67_ASAP7_75t_L g284 ( 
.A(n_272),
.B(n_0),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_214),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_217),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_218),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_218),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_187),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_245),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_236),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_230),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_194),
.Y(n_293)
);

OR2x2_ASAP7_75t_L g294 ( 
.A(n_247),
.B(n_1),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_230),
.Y(n_295)
);

CKINVDCx16_ASAP7_75t_R g296 ( 
.A(n_198),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_194),
.Y(n_297)
);

CKINVDCx16_ASAP7_75t_R g298 ( 
.A(n_211),
.Y(n_298)
);

INVxp67_ASAP7_75t_SL g299 ( 
.A(n_190),
.Y(n_299)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_245),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g301 ( 
.A(n_248),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_279),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_279),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g304 ( 
.A(n_197),
.B(n_2),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_189),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g306 ( 
.A(n_248),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_197),
.B(n_5),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_272),
.B(n_5),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_195),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_191),
.Y(n_310)
);

INVxp33_ASAP7_75t_SL g311 ( 
.A(n_207),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_199),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_201),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_259),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_192),
.Y(n_316)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_272),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_196),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_200),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_209),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_202),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_238),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_210),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_R g324 ( 
.A(n_250),
.B(n_6),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_261),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_203),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_219),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_220),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_221),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_222),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_261),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_224),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_226),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_241),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_204),
.Y(n_335)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_278),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_229),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_278),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_205),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_235),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_242),
.Y(n_341)
);

HB1xp67_ASAP7_75t_L g342 ( 
.A(n_264),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_267),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_290),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_290),
.Y(n_345)
);

BUFx6f_ASAP7_75t_L g346 ( 
.A(n_290),
.Y(n_346)
);

CKINVDCx16_ASAP7_75t_R g347 ( 
.A(n_280),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_320),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_320),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_290),
.Y(n_350)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_330),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_284),
.B(n_307),
.Y(n_352)
);

BUFx2_ASAP7_75t_L g353 ( 
.A(n_322),
.Y(n_353)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_330),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_309),
.Y(n_355)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_315),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_313),
.Y(n_357)
);

NAND2xp33_ASAP7_75t_L g358 ( 
.A(n_294),
.B(n_193),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_225),
.Y(n_359)
);

NAND2xp33_ASAP7_75t_L g360 ( 
.A(n_300),
.B(n_193),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_314),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_317),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_317),
.Y(n_363)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_323),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g365 ( 
.A(n_334),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_327),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_283),
.B(n_228),
.Y(n_367)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_328),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_300),
.Y(n_369)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_329),
.Y(n_370)
);

AND2x2_ASAP7_75t_L g371 ( 
.A(n_302),
.B(n_188),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_332),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_303),
.B(n_188),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_333),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g375 ( 
.A(n_342),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_281),
.Y(n_376)
);

INVx2_ASAP7_75t_L g377 ( 
.A(n_337),
.Y(n_377)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_340),
.Y(n_378)
);

CKINVDCx14_ASAP7_75t_R g379 ( 
.A(n_343),
.Y(n_379)
);

AND2x2_ASAP7_75t_L g380 ( 
.A(n_299),
.B(n_188),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_293),
.B(n_239),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_341),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_311),
.B(n_233),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_285),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g385 ( 
.A(n_292),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_304),
.B(n_268),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_286),
.Y(n_387)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_291),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_308),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_308),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_304),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_296),
.A2(n_252),
.B1(n_212),
.B2(n_274),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_289),
.B(n_256),
.Y(n_393)
);

BUFx6f_ASAP7_75t_L g394 ( 
.A(n_305),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g395 ( 
.A(n_297),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_310),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_316),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_318),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

INVx3_ASAP7_75t_L g400 ( 
.A(n_346),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g401 ( 
.A(n_346),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_362),
.Y(n_402)
);

INVx5_ASAP7_75t_L g403 ( 
.A(n_348),
.Y(n_403)
);

HB1xp67_ASAP7_75t_L g404 ( 
.A(n_353),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_353),
.B(n_298),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_390),
.B(n_321),
.Y(n_406)
);

AND2x2_ASAP7_75t_L g407 ( 
.A(n_365),
.B(n_326),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_346),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_335),
.Y(n_409)
);

INVx4_ASAP7_75t_L g410 ( 
.A(n_346),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_386),
.B(n_339),
.Y(n_411)
);

NAND2x1p5_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_396),
.Y(n_412)
);

NOR3xp33_ASAP7_75t_L g413 ( 
.A(n_383),
.B(n_263),
.C(n_258),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_390),
.B(n_208),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_362),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_384),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_355),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_213),
.Y(n_418)
);

CKINVDCx11_ASAP7_75t_R g419 ( 
.A(n_347),
.Y(n_419)
);

BUFx6f_ASAP7_75t_L g420 ( 
.A(n_369),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_357),
.Y(n_421)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_359),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_363),
.Y(n_423)
);

AOI22xp33_ASAP7_75t_L g424 ( 
.A1(n_391),
.A2(n_265),
.B1(n_266),
.B2(n_269),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_369),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_361),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g427 ( 
.A(n_380),
.B(n_324),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_369),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_369),
.Y(n_429)
);

BUFx6f_ASAP7_75t_L g430 ( 
.A(n_348),
.Y(n_430)
);

NAND3xp33_ASAP7_75t_L g431 ( 
.A(n_358),
.B(n_216),
.C(n_215),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_363),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_394),
.B(n_393),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_348),
.Y(n_435)
);

INVx8_ASAP7_75t_L g436 ( 
.A(n_394),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_352),
.B(n_223),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_348),
.Y(n_439)
);

INVx2_ASAP7_75t_L g440 ( 
.A(n_349),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_349),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_356),
.B(n_227),
.Y(n_442)
);

AND2x2_ASAP7_75t_SL g443 ( 
.A(n_358),
.B(n_270),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_394),
.Y(n_444)
);

BUFx3_ASAP7_75t_L g445 ( 
.A(n_344),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_379),
.Y(n_446)
);

NAND3x1_ASAP7_75t_L g447 ( 
.A(n_392),
.B(n_275),
.C(n_324),
.Y(n_447)
);

BUFx4f_ASAP7_75t_L g448 ( 
.A(n_394),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_372),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_374),
.Y(n_450)
);

INVx3_ASAP7_75t_L g451 ( 
.A(n_376),
.Y(n_451)
);

INVx1_ASAP7_75t_SL g452 ( 
.A(n_367),
.Y(n_452)
);

INVx3_ASAP7_75t_L g453 ( 
.A(n_376),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_345),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_352),
.B(n_231),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_350),
.B(n_232),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_382),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_351),
.Y(n_458)
);

NAND2xp33_ASAP7_75t_L g459 ( 
.A(n_396),
.B(n_234),
.Y(n_459)
);

INVx3_ASAP7_75t_L g460 ( 
.A(n_376),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_379),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_375),
.B(n_237),
.Y(n_462)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_380),
.A2(n_271),
.B1(n_243),
.B2(n_244),
.Y(n_463)
);

INVx4_ASAP7_75t_L g464 ( 
.A(n_376),
.Y(n_464)
);

NAND2xp33_ASAP7_75t_R g465 ( 
.A(n_381),
.B(n_371),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_371),
.B(n_338),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_388),
.Y(n_467)
);

BUFx3_ASAP7_75t_L g468 ( 
.A(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_433),
.B(n_399),
.Y(n_470)
);

INVx2_ASAP7_75t_SL g471 ( 
.A(n_404),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_422),
.B(n_399),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_417),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_421),
.Y(n_474)
);

NAND2x1p5_ASAP7_75t_L g475 ( 
.A(n_448),
.B(n_397),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_426),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_433),
.B(n_398),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_434),
.Y(n_478)
);

AO22x2_ASAP7_75t_L g479 ( 
.A1(n_452),
.A2(n_381),
.B1(n_373),
.B2(n_287),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_449),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_450),
.Y(n_481)
);

AO22x2_ASAP7_75t_L g482 ( 
.A1(n_406),
.A2(n_373),
.B1(n_288),
.B2(n_287),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_402),
.Y(n_483)
);

INVxp67_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

OAI22xp33_ASAP7_75t_SL g485 ( 
.A1(n_409),
.A2(n_395),
.B1(n_385),
.B2(n_240),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_457),
.Y(n_486)
);

AO22x2_ASAP7_75t_L g487 ( 
.A1(n_406),
.A2(n_288),
.B1(n_331),
.B2(n_325),
.Y(n_487)
);

BUFx2_ASAP7_75t_L g488 ( 
.A(n_427),
.Y(n_488)
);

AO22x2_ASAP7_75t_L g489 ( 
.A1(n_413),
.A2(n_336),
.B1(n_312),
.B2(n_306),
.Y(n_489)
);

NAND2x1p5_ASAP7_75t_L g490 ( 
.A(n_448),
.B(n_370),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_445),
.B(n_387),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_407),
.B(n_295),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_440),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_440),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_441),
.Y(n_495)
);

OR2x6_ASAP7_75t_L g496 ( 
.A(n_446),
.B(n_387),
.Y(n_496)
);

NAND2xp33_ASAP7_75t_L g497 ( 
.A(n_436),
.B(n_246),
.Y(n_497)
);

OAI221xp5_ASAP7_75t_L g498 ( 
.A1(n_424),
.A2(n_360),
.B1(n_378),
.B2(n_377),
.C(n_368),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_441),
.Y(n_499)
);

AND2x4_ASAP7_75t_L g500 ( 
.A(n_445),
.B(n_364),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_458),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_458),
.Y(n_502)
);

BUFx6f_ASAP7_75t_SL g503 ( 
.A(n_443),
.Y(n_503)
);

INVxp33_ASAP7_75t_L g504 ( 
.A(n_405),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_402),
.Y(n_505)
);

BUFx8_ASAP7_75t_L g506 ( 
.A(n_466),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g507 ( 
.A(n_409),
.B(n_370),
.Y(n_507)
);

AND2x4_ASAP7_75t_L g508 ( 
.A(n_454),
.B(n_364),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

AND2x4_ASAP7_75t_L g510 ( 
.A(n_454),
.B(n_368),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_415),
.Y(n_511)
);

INVx2_ASAP7_75t_SL g512 ( 
.A(n_437),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g513 ( 
.A(n_411),
.B(n_370),
.Y(n_513)
);

AO22x2_ASAP7_75t_L g514 ( 
.A1(n_431),
.A2(n_301),
.B1(n_7),
.B2(n_8),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_423),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_423),
.Y(n_516)
);

AO22x2_ASAP7_75t_L g517 ( 
.A1(n_443),
.A2(n_6),
.B1(n_9),
.B2(n_10),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_432),
.Y(n_518)
);

INVx2_ASAP7_75t_SL g519 ( 
.A(n_455),
.Y(n_519)
);

AO22x2_ASAP7_75t_L g520 ( 
.A1(n_465),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_442),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_432),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_467),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_420),
.Y(n_524)
);

AO22x2_ASAP7_75t_L g525 ( 
.A1(n_465),
.A2(n_11),
.B1(n_12),
.B2(n_13),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_414),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_411),
.B(n_360),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_418),
.B(n_351),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_444),
.B(n_377),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_451),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_R g531 ( 
.A(n_461),
.B(n_249),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_436),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_451),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_412),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_453),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_453),
.Y(n_536)
);

INVxp67_ASAP7_75t_L g537 ( 
.A(n_442),
.Y(n_537)
);

NAND2xp5_ASAP7_75t_SL g538 ( 
.A(n_521),
.B(n_412),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_537),
.B(n_436),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_472),
.B(n_463),
.Y(n_540)
);

NAND2xp33_ASAP7_75t_SL g541 ( 
.A(n_503),
.B(n_463),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g542 ( 
.A(n_527),
.B(n_462),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_SL g543 ( 
.A(n_529),
.B(n_462),
.Y(n_543)
);

NAND2xp33_ASAP7_75t_SL g544 ( 
.A(n_531),
.B(n_424),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_512),
.B(n_519),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_477),
.B(n_488),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_488),
.B(n_456),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_526),
.B(n_459),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_507),
.B(n_464),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_SL g550 ( 
.A(n_504),
.B(n_251),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_SL g551 ( 
.A(n_513),
.B(n_464),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_471),
.B(n_468),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_470),
.B(n_528),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_532),
.B(n_468),
.Y(n_554)
);

NAND2xp33_ASAP7_75t_SL g555 ( 
.A(n_534),
.B(n_253),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_469),
.B(n_460),
.Y(n_556)
);

NAND2xp33_ASAP7_75t_SL g557 ( 
.A(n_492),
.B(n_254),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_491),
.B(n_460),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_491),
.B(n_420),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_500),
.B(n_420),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_500),
.B(n_420),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_SL g562 ( 
.A(n_508),
.B(n_425),
.Y(n_562)
);

NAND2xp33_ASAP7_75t_SL g563 ( 
.A(n_473),
.B(n_255),
.Y(n_563)
);

NAND2xp5_ASAP7_75t_SL g564 ( 
.A(n_508),
.B(n_425),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_510),
.B(n_425),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_510),
.B(n_425),
.Y(n_566)
);

AND2x4_ASAP7_75t_L g567 ( 
.A(n_474),
.B(n_378),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_SL g568 ( 
.A(n_475),
.B(n_428),
.Y(n_568)
);

NAND2xp33_ASAP7_75t_SL g569 ( 
.A(n_476),
.B(n_257),
.Y(n_569)
);

NOR2xp33_ASAP7_75t_SL g570 ( 
.A(n_506),
.B(n_484),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_478),
.B(n_428),
.Y(n_571)
);

NAND2xp33_ASAP7_75t_SL g572 ( 
.A(n_480),
.B(n_260),
.Y(n_572)
);

NAND2xp33_ASAP7_75t_SL g573 ( 
.A(n_481),
.B(n_262),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g574 ( 
.A(n_486),
.B(n_428),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g575 ( 
.A(n_485),
.B(n_429),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_490),
.B(n_429),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_523),
.B(n_429),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_496),
.B(n_524),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_530),
.B(n_273),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_SL g580 ( 
.A(n_533),
.B(n_429),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_496),
.B(n_419),
.Y(n_581)
);

NAND2xp5_ASAP7_75t_L g582 ( 
.A(n_493),
.B(n_435),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_SL g583 ( 
.A(n_536),
.B(n_430),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_535),
.B(n_430),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_494),
.B(n_435),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_495),
.B(n_430),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_499),
.B(n_430),
.Y(n_587)
);

NAND2xp5_ASAP7_75t_SL g588 ( 
.A(n_501),
.B(n_439),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_SL g589 ( 
.A(n_502),
.B(n_439),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_SL g590 ( 
.A(n_509),
.B(n_276),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_511),
.B(n_515),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_518),
.B(n_439),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_SL g593 ( 
.A(n_522),
.B(n_439),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_483),
.B(n_388),
.Y(n_594)
);

NAND2xp33_ASAP7_75t_SL g595 ( 
.A(n_517),
.B(n_447),
.Y(n_595)
);

OAI21xp5_ASAP7_75t_L g596 ( 
.A1(n_542),
.A2(n_505),
.B(n_516),
.Y(n_596)
);

OAI22x1_ASAP7_75t_L g597 ( 
.A1(n_540),
.A2(n_487),
.B1(n_517),
.B2(n_482),
.Y(n_597)
);

OAI21xp5_ASAP7_75t_L g598 ( 
.A1(n_553),
.A2(n_498),
.B(n_497),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_582),
.A2(n_438),
.B(n_408),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_548),
.B(n_479),
.Y(n_600)
);

OAI21xp5_ASAP7_75t_L g601 ( 
.A1(n_538),
.A2(n_546),
.B(n_549),
.Y(n_601)
);

BUFx8_ASAP7_75t_L g602 ( 
.A(n_581),
.Y(n_602)
);

CKINVDCx5p33_ASAP7_75t_R g603 ( 
.A(n_541),
.Y(n_603)
);

AOI21xp5_ASAP7_75t_L g604 ( 
.A1(n_551),
.A2(n_403),
.B(n_410),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_543),
.B(n_547),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_567),
.Y(n_606)
);

OAI21xp5_ASAP7_75t_L g607 ( 
.A1(n_591),
.A2(n_438),
.B(n_400),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_567),
.B(n_479),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_585),
.Y(n_609)
);

AND2x4_ASAP7_75t_L g610 ( 
.A(n_578),
.B(n_400),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_556),
.Y(n_611)
);

AOI21xp5_ASAP7_75t_L g612 ( 
.A1(n_559),
.A2(n_403),
.B(n_410),
.Y(n_612)
);

OA22x2_ASAP7_75t_L g613 ( 
.A1(n_545),
.A2(n_487),
.B1(n_482),
.B2(n_525),
.Y(n_613)
);

OAI21x1_ASAP7_75t_L g614 ( 
.A1(n_583),
.A2(n_584),
.B(n_580),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g615 ( 
.A1(n_539),
.A2(n_525),
.B1(n_520),
.B2(n_514),
.Y(n_615)
);

OAI21x1_ASAP7_75t_L g616 ( 
.A1(n_586),
.A2(n_408),
.B(n_354),
.Y(n_616)
);

OAI21x1_ASAP7_75t_L g617 ( 
.A1(n_587),
.A2(n_354),
.B(n_401),
.Y(n_617)
);

A2O1A1Ixp33_ASAP7_75t_L g618 ( 
.A1(n_544),
.A2(n_595),
.B(n_563),
.C(n_569),
.Y(n_618)
);

INVxp67_ASAP7_75t_L g619 ( 
.A(n_570),
.Y(n_619)
);

AO32x2_ASAP7_75t_L g620 ( 
.A1(n_575),
.A2(n_520),
.A3(n_514),
.B1(n_489),
.B2(n_15),
.Y(n_620)
);

O2A1O1Ixp33_ASAP7_75t_L g621 ( 
.A1(n_568),
.A2(n_489),
.B(n_13),
.C(n_14),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_560),
.A2(n_401),
.B1(n_403),
.B2(n_388),
.Y(n_622)
);

O2A1O1Ixp33_ASAP7_75t_SL g623 ( 
.A1(n_576),
.A2(n_100),
.B(n_184),
.C(n_183),
.Y(n_623)
);

A2O1A1Ixp33_ASAP7_75t_L g624 ( 
.A1(n_572),
.A2(n_401),
.B(n_403),
.C(n_419),
.Y(n_624)
);

NAND3x1_ASAP7_75t_L g625 ( 
.A(n_557),
.B(n_12),
.C(n_14),
.Y(n_625)
);

O2A1O1Ixp33_ASAP7_75t_SL g626 ( 
.A1(n_571),
.A2(n_90),
.B(n_181),
.C(n_179),
.Y(n_626)
);

NAND3xp33_ASAP7_75t_L g627 ( 
.A(n_573),
.B(n_401),
.C(n_17),
.Y(n_627)
);

BUFx12f_ASAP7_75t_L g628 ( 
.A(n_578),
.Y(n_628)
);

CKINVDCx16_ASAP7_75t_R g629 ( 
.A(n_550),
.Y(n_629)
);

OAI21x1_ASAP7_75t_L g630 ( 
.A1(n_588),
.A2(n_89),
.B(n_176),
.Y(n_630)
);

OAI22xp5_ASAP7_75t_L g631 ( 
.A1(n_561),
.A2(n_562),
.B1(n_564),
.B2(n_565),
.Y(n_631)
);

OR2x6_ASAP7_75t_L g632 ( 
.A(n_552),
.B(n_16),
.Y(n_632)
);

OAI21x1_ASAP7_75t_L g633 ( 
.A1(n_589),
.A2(n_88),
.B(n_175),
.Y(n_633)
);

AND2x4_ASAP7_75t_L g634 ( 
.A(n_558),
.B(n_26),
.Y(n_634)
);

BUFx3_ASAP7_75t_L g635 ( 
.A(n_555),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_L g636 ( 
.A(n_566),
.B(n_16),
.Y(n_636)
);

O2A1O1Ixp33_ASAP7_75t_L g637 ( 
.A1(n_574),
.A2(n_18),
.B(n_19),
.C(n_20),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g638 ( 
.A1(n_554),
.A2(n_101),
.B(n_174),
.Y(n_638)
);

AO21x1_ASAP7_75t_L g639 ( 
.A1(n_592),
.A2(n_20),
.B(n_21),
.Y(n_639)
);

AOI22xp5_ASAP7_75t_L g640 ( 
.A1(n_590),
.A2(n_87),
.B1(n_173),
.B2(n_171),
.Y(n_640)
);

OAI21xp5_ASAP7_75t_L g641 ( 
.A1(n_593),
.A2(n_86),
.B(n_169),
.Y(n_641)
);

OAI21x1_ASAP7_75t_L g642 ( 
.A1(n_599),
.A2(n_577),
.B(n_594),
.Y(n_642)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_617),
.A2(n_579),
.B(n_84),
.Y(n_643)
);

OAI21x1_ASAP7_75t_L g644 ( 
.A1(n_616),
.A2(n_82),
.B(n_168),
.Y(n_644)
);

AND2x4_ASAP7_75t_L g645 ( 
.A(n_606),
.B(n_29),
.Y(n_645)
);

AOI21x1_ASAP7_75t_L g646 ( 
.A1(n_604),
.A2(n_598),
.B(n_601),
.Y(n_646)
);

AND2x2_ASAP7_75t_L g647 ( 
.A(n_611),
.B(n_30),
.Y(n_647)
);

OA21x2_ASAP7_75t_L g648 ( 
.A1(n_596),
.A2(n_21),
.B(n_22),
.Y(n_648)
);

OAI21x1_ASAP7_75t_L g649 ( 
.A1(n_630),
.A2(n_103),
.B(n_31),
.Y(n_649)
);

OAI21x1_ASAP7_75t_SL g650 ( 
.A1(n_639),
.A2(n_106),
.B(n_34),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_605),
.B(n_23),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_636),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_609),
.Y(n_653)
);

AOI221xp5_ASAP7_75t_L g654 ( 
.A1(n_597),
.A2(n_23),
.B1(n_35),
.B2(n_36),
.C(n_38),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_611),
.Y(n_655)
);

OAI21x1_ASAP7_75t_L g656 ( 
.A1(n_633),
.A2(n_614),
.B(n_607),
.Y(n_656)
);

NOR2x1_ASAP7_75t_L g657 ( 
.A(n_627),
.B(n_39),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_600),
.Y(n_658)
);

BUFx12f_ASAP7_75t_L g659 ( 
.A(n_628),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_618),
.B(n_40),
.Y(n_660)
);

BUFx2_ASAP7_75t_L g661 ( 
.A(n_608),
.Y(n_661)
);

OAI21x1_ASAP7_75t_SL g662 ( 
.A1(n_621),
.A2(n_641),
.B(n_637),
.Y(n_662)
);

CKINVDCx6p67_ASAP7_75t_R g663 ( 
.A(n_635),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_610),
.Y(n_664)
);

INVx2_ASAP7_75t_L g665 ( 
.A(n_634),
.Y(n_665)
);

BUFx3_ASAP7_75t_L g666 ( 
.A(n_602),
.Y(n_666)
);

AND2x4_ASAP7_75t_L g667 ( 
.A(n_634),
.B(n_41),
.Y(n_667)
);

BUFx2_ASAP7_75t_L g668 ( 
.A(n_610),
.Y(n_668)
);

AOI22xp33_ASAP7_75t_L g669 ( 
.A1(n_613),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_631),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_620),
.Y(n_671)
);

OAI21x1_ASAP7_75t_L g672 ( 
.A1(n_612),
.A2(n_48),
.B(n_49),
.Y(n_672)
);

INVx3_ASAP7_75t_L g673 ( 
.A(n_629),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_622),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_620),
.Y(n_675)
);

AND2x2_ASAP7_75t_L g676 ( 
.A(n_620),
.B(n_51),
.Y(n_676)
);

A2O1A1Ixp33_ASAP7_75t_L g677 ( 
.A1(n_615),
.A2(n_640),
.B(n_638),
.C(n_624),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_632),
.B(n_603),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_SL g679 ( 
.A1(n_632),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_679)
);

BUFx2_ASAP7_75t_L g680 ( 
.A(n_619),
.Y(n_680)
);

NAND2x1_ASAP7_75t_L g681 ( 
.A(n_623),
.B(n_55),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_625),
.B(n_59),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_645),
.Y(n_683)
);

OA21x2_ASAP7_75t_L g684 ( 
.A1(n_671),
.A2(n_675),
.B(n_656),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_655),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g686 ( 
.A(n_652),
.B(n_602),
.Y(n_686)
);

AND2x4_ASAP7_75t_L g687 ( 
.A(n_665),
.B(n_60),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_653),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_670),
.Y(n_689)
);

A2O1A1Ixp33_ASAP7_75t_L g690 ( 
.A1(n_677),
.A2(n_626),
.B(n_63),
.C(n_66),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_680),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_676),
.B(n_61),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_648),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_668),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_658),
.B(n_178),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_648),
.Y(n_696)
);

CKINVDCx5p33_ASAP7_75t_R g697 ( 
.A(n_663),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_665),
.Y(n_698)
);

INVx3_ASAP7_75t_L g699 ( 
.A(n_645),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_661),
.B(n_69),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_661),
.B(n_164),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_648),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_647),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_663),
.Y(n_704)
);

NAND2x1p5_ASAP7_75t_L g705 ( 
.A(n_672),
.B(n_73),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_651),
.B(n_162),
.Y(n_706)
);

HB1xp67_ASAP7_75t_L g707 ( 
.A(n_680),
.Y(n_707)
);

AND2x2_ASAP7_75t_L g708 ( 
.A(n_676),
.B(n_647),
.Y(n_708)
);

HB1xp67_ASAP7_75t_L g709 ( 
.A(n_668),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_646),
.Y(n_710)
);

OAI21x1_ASAP7_75t_L g711 ( 
.A1(n_643),
.A2(n_74),
.B(n_75),
.Y(n_711)
);

INVx1_ASAP7_75t_L g712 ( 
.A(n_656),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_677),
.Y(n_713)
);

HB1xp67_ASAP7_75t_L g714 ( 
.A(n_664),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_672),
.Y(n_715)
);

AOI22xp33_ASAP7_75t_L g716 ( 
.A1(n_662),
.A2(n_80),
.B1(n_102),
.B2(n_107),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_642),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_644),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_642),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_667),
.B(n_161),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_644),
.Y(n_721)
);

HB1xp67_ASAP7_75t_L g722 ( 
.A(n_673),
.Y(n_722)
);

HB1xp67_ASAP7_75t_L g723 ( 
.A(n_673),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_667),
.B(n_111),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_649),
.Y(n_725)
);

AND2x2_ASAP7_75t_L g726 ( 
.A(n_667),
.B(n_158),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_643),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_649),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_645),
.B(n_112),
.Y(n_729)
);

CKINVDCx11_ASAP7_75t_R g730 ( 
.A(n_683),
.Y(n_730)
);

INVxp67_ASAP7_75t_L g731 ( 
.A(n_707),
.Y(n_731)
);

INVxp67_ASAP7_75t_L g732 ( 
.A(n_709),
.Y(n_732)
);

INVxp67_ASAP7_75t_L g733 ( 
.A(n_691),
.Y(n_733)
);

NOR2xp33_ASAP7_75t_R g734 ( 
.A(n_697),
.B(n_673),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_R g735 ( 
.A(n_697),
.B(n_678),
.Y(n_735)
);

INVxp67_ASAP7_75t_L g736 ( 
.A(n_722),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_723),
.Y(n_737)
);

CKINVDCx8_ASAP7_75t_R g738 ( 
.A(n_704),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_688),
.B(n_678),
.Y(n_739)
);

NOR2xp33_ASAP7_75t_R g740 ( 
.A(n_704),
.B(n_659),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_R g741 ( 
.A(n_699),
.B(n_659),
.Y(n_741)
);

INVxp67_ASAP7_75t_L g742 ( 
.A(n_686),
.Y(n_742)
);

CKINVDCx11_ASAP7_75t_R g743 ( 
.A(n_683),
.Y(n_743)
);

XOR2xp5_ASAP7_75t_L g744 ( 
.A(n_720),
.B(n_666),
.Y(n_744)
);

NAND2xp33_ASAP7_75t_R g745 ( 
.A(n_724),
.B(n_682),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_688),
.B(n_660),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_694),
.B(n_666),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_685),
.Y(n_748)
);

OR2x6_ASAP7_75t_L g749 ( 
.A(n_683),
.B(n_657),
.Y(n_749)
);

BUFx3_ASAP7_75t_L g750 ( 
.A(n_694),
.Y(n_750)
);

NAND2xp33_ASAP7_75t_SL g751 ( 
.A(n_724),
.B(n_669),
.Y(n_751)
);

AND2x2_ASAP7_75t_L g752 ( 
.A(n_708),
.B(n_654),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_708),
.B(n_674),
.Y(n_753)
);

INVxp67_ASAP7_75t_L g754 ( 
.A(n_714),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_713),
.B(n_679),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_726),
.B(n_118),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_R g757 ( 
.A(n_699),
.B(n_122),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_SL g758 ( 
.A(n_724),
.B(n_681),
.Y(n_758)
);

AND2x4_ASAP7_75t_L g759 ( 
.A(n_699),
.B(n_674),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_683),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_683),
.B(n_698),
.Y(n_761)
);

AND2x2_ASAP7_75t_L g762 ( 
.A(n_692),
.B(n_703),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_R g763 ( 
.A(n_726),
.B(n_123),
.Y(n_763)
);

INVxp67_ASAP7_75t_L g764 ( 
.A(n_700),
.Y(n_764)
);

NAND2xp33_ASAP7_75t_R g765 ( 
.A(n_729),
.B(n_126),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_R g766 ( 
.A(n_729),
.B(n_128),
.Y(n_766)
);

AND2x4_ASAP7_75t_L g767 ( 
.A(n_698),
.B(n_132),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_713),
.B(n_662),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_748),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_762),
.B(n_684),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_753),
.B(n_684),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_768),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_752),
.B(n_684),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_739),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_759),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_759),
.Y(n_776)
);

AOI22xp33_ASAP7_75t_L g777 ( 
.A1(n_751),
.A2(n_716),
.B1(n_706),
.B2(n_687),
.Y(n_777)
);

BUFx3_ASAP7_75t_L g778 ( 
.A(n_730),
.Y(n_778)
);

AND2x2_ASAP7_75t_L g779 ( 
.A(n_761),
.B(n_684),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_764),
.B(n_689),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_761),
.B(n_710),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_731),
.B(n_689),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_736),
.B(n_710),
.Y(n_783)
);

AND2x2_ASAP7_75t_L g784 ( 
.A(n_737),
.B(n_693),
.Y(n_784)
);

AND2x4_ASAP7_75t_L g785 ( 
.A(n_750),
.B(n_712),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_746),
.Y(n_786)
);

INVx3_ASAP7_75t_L g787 ( 
.A(n_767),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_742),
.A2(n_703),
.B1(n_700),
.B2(n_692),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_733),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_747),
.B(n_712),
.Y(n_790)
);

AND2x2_ASAP7_75t_L g791 ( 
.A(n_754),
.B(n_693),
.Y(n_791)
);

INVx2_ASAP7_75t_L g792 ( 
.A(n_732),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_755),
.B(n_696),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_747),
.B(n_696),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_740),
.Y(n_795)
);

BUFx3_ASAP7_75t_L g796 ( 
.A(n_760),
.Y(n_796)
);

AND2x4_ASAP7_75t_L g797 ( 
.A(n_767),
.B(n_717),
.Y(n_797)
);

INVxp67_ASAP7_75t_L g798 ( 
.A(n_792),
.Y(n_798)
);

BUFx2_ASAP7_75t_L g799 ( 
.A(n_790),
.Y(n_799)
);

INVx2_ASAP7_75t_L g800 ( 
.A(n_769),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_772),
.B(n_774),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_769),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_791),
.Y(n_803)
);

HB1xp67_ASAP7_75t_L g804 ( 
.A(n_772),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_773),
.B(n_702),
.Y(n_805)
);

INVxp67_ASAP7_75t_SL g806 ( 
.A(n_786),
.Y(n_806)
);

INVxp67_ASAP7_75t_L g807 ( 
.A(n_792),
.Y(n_807)
);

OR2x6_ASAP7_75t_L g808 ( 
.A(n_797),
.B(n_715),
.Y(n_808)
);

HB1xp67_ASAP7_75t_L g809 ( 
.A(n_779),
.Y(n_809)
);

OR2x2_ASAP7_75t_L g810 ( 
.A(n_770),
.B(n_702),
.Y(n_810)
);

OR2x2_ASAP7_75t_L g811 ( 
.A(n_770),
.B(n_717),
.Y(n_811)
);

NAND5xp2_ASAP7_75t_L g812 ( 
.A(n_777),
.B(n_756),
.C(n_745),
.D(n_705),
.E(n_690),
.Y(n_812)
);

NOR2x1_ASAP7_75t_L g813 ( 
.A(n_778),
.B(n_796),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_SL g814 ( 
.A(n_788),
.B(n_757),
.Y(n_814)
);

INVx2_ASAP7_75t_L g815 ( 
.A(n_779),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_778),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_815),
.Y(n_817)
);

AND2x2_ASAP7_75t_L g818 ( 
.A(n_809),
.B(n_793),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_801),
.B(n_793),
.Y(n_819)
);

AOI21xp33_ASAP7_75t_L g820 ( 
.A1(n_814),
.A2(n_765),
.B(n_766),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_798),
.B(n_786),
.Y(n_821)
);

OR2x2_ASAP7_75t_L g822 ( 
.A(n_815),
.B(n_773),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_806),
.B(n_791),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_799),
.B(n_794),
.Y(n_824)
);

AND3x2_ASAP7_75t_L g825 ( 
.A(n_804),
.B(n_789),
.C(n_735),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_807),
.B(n_794),
.Y(n_826)
);

INVxp67_ASAP7_75t_L g827 ( 
.A(n_813),
.Y(n_827)
);

INVx2_ASAP7_75t_L g828 ( 
.A(n_800),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_828),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_819),
.B(n_805),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_821),
.B(n_805),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_820),
.A2(n_814),
.B1(n_825),
.B2(n_827),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_820),
.A2(n_816),
.B1(n_758),
.B2(n_787),
.Y(n_833)
);

NAND2xp33_ASAP7_75t_SL g834 ( 
.A(n_818),
.B(n_734),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_829),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_832),
.B(n_823),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_831),
.B(n_824),
.Y(n_837)
);

INVx1_ASAP7_75t_SL g838 ( 
.A(n_834),
.Y(n_838)
);

AND2x2_ASAP7_75t_L g839 ( 
.A(n_830),
.B(n_816),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_833),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_835),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_836),
.A2(n_812),
.B(n_795),
.Y(n_842)
);

O2A1O1Ixp33_ASAP7_75t_L g843 ( 
.A1(n_840),
.A2(n_778),
.B(n_823),
.C(n_782),
.Y(n_843)
);

AND2x4_ASAP7_75t_L g844 ( 
.A(n_838),
.B(n_808),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_839),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_845),
.B(n_839),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_841),
.B(n_837),
.Y(n_847)
);

OR2x2_ASAP7_75t_L g848 ( 
.A(n_844),
.B(n_837),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_844),
.B(n_826),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_847),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_848),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_846),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_849),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_847),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_851),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_852),
.B(n_843),
.Y(n_856)
);

AOI221x1_ASAP7_75t_L g857 ( 
.A1(n_850),
.A2(n_842),
.B1(n_650),
.B2(n_695),
.C(n_701),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_852),
.B(n_817),
.Y(n_858)
);

AOI211x1_ASAP7_75t_L g859 ( 
.A1(n_853),
.A2(n_802),
.B(n_780),
.C(n_803),
.Y(n_859)
);

NOR3x1_ASAP7_75t_L g860 ( 
.A(n_854),
.B(n_738),
.C(n_744),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_851),
.B(n_796),
.C(n_687),
.Y(n_861)
);

NOR3x1_ASAP7_75t_SL g862 ( 
.A(n_851),
.B(n_763),
.C(n_741),
.Y(n_862)
);

INVxp67_ASAP7_75t_L g863 ( 
.A(n_856),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_855),
.Y(n_864)
);

AO22x1_ASAP7_75t_L g865 ( 
.A1(n_862),
.A2(n_687),
.B1(n_787),
.B2(n_685),
.Y(n_865)
);

NAND3xp33_ASAP7_75t_L g866 ( 
.A(n_857),
.B(n_783),
.C(n_784),
.Y(n_866)
);

A2O1A1Ixp33_ASAP7_75t_L g867 ( 
.A1(n_861),
.A2(n_858),
.B(n_860),
.C(n_859),
.Y(n_867)
);

AOI221xp5_ASAP7_75t_L g868 ( 
.A1(n_856),
.A2(n_650),
.B1(n_784),
.B2(n_785),
.C(n_790),
.Y(n_868)
);

NOR2x1_ASAP7_75t_L g869 ( 
.A(n_855),
.B(n_808),
.Y(n_869)
);

OAI31xp33_ASAP7_75t_L g870 ( 
.A1(n_862),
.A2(n_705),
.A3(n_787),
.B(n_822),
.Y(n_870)
);

AOI221xp5_ASAP7_75t_L g871 ( 
.A1(n_856),
.A2(n_785),
.B1(n_790),
.B2(n_800),
.C(n_783),
.Y(n_871)
);

O2A1O1Ixp33_ASAP7_75t_L g872 ( 
.A1(n_856),
.A2(n_705),
.B(n_749),
.C(n_808),
.Y(n_872)
);

INVxp67_ASAP7_75t_SL g873 ( 
.A(n_864),
.Y(n_873)
);

NAND4xp75_ASAP7_75t_L g874 ( 
.A(n_870),
.B(n_781),
.C(n_771),
.D(n_715),
.Y(n_874)
);

NOR2xp33_ASAP7_75t_L g875 ( 
.A(n_863),
.B(n_790),
.Y(n_875)
);

OAI22xp5_ASAP7_75t_L g876 ( 
.A1(n_867),
.A2(n_866),
.B1(n_869),
.B2(n_871),
.Y(n_876)
);

AO22x1_ASAP7_75t_L g877 ( 
.A1(n_865),
.A2(n_785),
.B1(n_797),
.B2(n_781),
.Y(n_877)
);

AOI22xp5_ASAP7_75t_L g878 ( 
.A1(n_868),
.A2(n_808),
.B1(n_785),
.B2(n_743),
.Y(n_878)
);

NOR2x1p5_ASAP7_75t_L g879 ( 
.A(n_872),
.B(n_810),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_863),
.B(n_810),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_864),
.Y(n_881)
);

XNOR2xp5_ASAP7_75t_L g882 ( 
.A(n_876),
.B(n_749),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_881),
.B(n_811),
.Y(n_883)
);

NAND2xp33_ASAP7_75t_SL g884 ( 
.A(n_879),
.B(n_811),
.Y(n_884)
);

NAND3xp33_ASAP7_75t_L g885 ( 
.A(n_873),
.B(n_727),
.C(n_776),
.Y(n_885)
);

NAND2xp33_ASAP7_75t_L g886 ( 
.A(n_874),
.B(n_776),
.Y(n_886)
);

NAND2xp33_ASAP7_75t_SL g887 ( 
.A(n_877),
.B(n_771),
.Y(n_887)
);

NOR2xp33_ASAP7_75t_R g888 ( 
.A(n_880),
.B(n_875),
.Y(n_888)
);

NOR2xp33_ASAP7_75t_R g889 ( 
.A(n_878),
.B(n_134),
.Y(n_889)
);

XOR2xp5_ASAP7_75t_L g890 ( 
.A(n_882),
.B(n_137),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_883),
.Y(n_891)
);

INVxp67_ASAP7_75t_SL g892 ( 
.A(n_886),
.Y(n_892)
);

INVx2_ASAP7_75t_L g893 ( 
.A(n_885),
.Y(n_893)
);

AO22x2_ASAP7_75t_L g894 ( 
.A1(n_888),
.A2(n_775),
.B1(n_797),
.B2(n_727),
.Y(n_894)
);

INVx2_ASAP7_75t_L g895 ( 
.A(n_887),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_884),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_889),
.B(n_775),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_896),
.A2(n_711),
.B(n_728),
.Y(n_898)
);

INVx2_ASAP7_75t_L g899 ( 
.A(n_895),
.Y(n_899)
);

OR4x1_ASAP7_75t_L g900 ( 
.A(n_890),
.B(n_721),
.C(n_719),
.D(n_142),
.Y(n_900)
);

INVx2_ASAP7_75t_L g901 ( 
.A(n_891),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_892),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_902),
.Y(n_903)
);

OAI21x1_ASAP7_75t_L g904 ( 
.A1(n_899),
.A2(n_893),
.B(n_897),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_901),
.B(n_894),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_903),
.A2(n_898),
.B1(n_900),
.B2(n_797),
.Y(n_906)
);

AOI31xp33_ASAP7_75t_L g907 ( 
.A1(n_905),
.A2(n_138),
.A3(n_140),
.B(n_145),
.Y(n_907)
);

AND3x1_ASAP7_75t_L g908 ( 
.A(n_906),
.B(n_904),
.C(n_150),
.Y(n_908)
);

AO21x1_ASAP7_75t_L g909 ( 
.A1(n_907),
.A2(n_146),
.B(n_151),
.Y(n_909)
);

XNOR2xp5_ASAP7_75t_L g910 ( 
.A(n_908),
.B(n_152),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_909),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_910),
.Y(n_912)
);

OAI222xp33_ASAP7_75t_L g913 ( 
.A1(n_911),
.A2(n_721),
.B1(n_728),
.B2(n_725),
.C1(n_719),
.C2(n_718),
.Y(n_913)
);

AOI22xp33_ASAP7_75t_L g914 ( 
.A1(n_912),
.A2(n_711),
.B1(n_725),
.B2(n_718),
.Y(n_914)
);

AOI211xp5_ASAP7_75t_L g915 ( 
.A1(n_914),
.A2(n_913),
.B(n_153),
.C(n_154),
.Y(n_915)
);


endmodule