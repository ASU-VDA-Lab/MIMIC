module fake_ariane_3160_n_96 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_38, n_2, n_18, n_32, n_28, n_37, n_9, n_11, n_34, n_26, n_3, n_14, n_0, n_36, n_33, n_19, n_30, n_39, n_40, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_35, n_10, n_25, n_96);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_38;
input n_2;
input n_18;
input n_32;
input n_28;
input n_37;
input n_9;
input n_11;
input n_34;
input n_26;
input n_3;
input n_14;
input n_0;
input n_36;
input n_33;
input n_19;
input n_30;
input n_39;
input n_40;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_35;
input n_10;
input n_25;

output n_96;

wire n_83;
wire n_56;
wire n_60;
wire n_64;
wire n_90;
wire n_47;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_69;
wire n_95;
wire n_92;
wire n_74;
wire n_53;
wire n_66;
wire n_71;
wire n_49;
wire n_50;
wire n_62;
wire n_51;
wire n_76;
wire n_79;
wire n_46;
wire n_84;
wire n_91;
wire n_72;
wire n_44;
wire n_82;
wire n_42;
wire n_57;
wire n_70;
wire n_85;
wire n_48;
wire n_94;
wire n_58;
wire n_65;
wire n_45;
wire n_52;
wire n_73;
wire n_77;
wire n_93;
wire n_61;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_55;
wire n_80;
wire n_88;
wire n_68;
wire n_78;
wire n_63;
wire n_59;
wire n_54;

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_11),
.B(n_0),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_40),
.Y(n_43)
);

OAI22x1_ASAP7_75t_R g44 ( 
.A1(n_2),
.A2(n_8),
.B1(n_29),
.B2(n_9),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_12),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_5),
.Y(n_48)
);

CKINVDCx5p33_ASAP7_75t_R g49 ( 
.A(n_21),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_35),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_15),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_6),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_1),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_19),
.B(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_0),
.B(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

NOR2xp67_ASAP7_75t_L g62 ( 
.A(n_58),
.B(n_13),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_54),
.A2(n_42),
.B1(n_51),
.B2(n_41),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_49),
.Y(n_64)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_60),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_16),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_43),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_57),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

BUFx4_ASAP7_75t_SL g72 ( 
.A(n_65),
.Y(n_72)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_59),
.B(n_52),
.C(n_55),
.Y(n_73)
);

AO31x2_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_44),
.A3(n_55),
.B(n_48),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_69),
.B(n_68),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_71),
.B(n_64),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_74),
.B(n_62),
.Y(n_79)
);

HB1xp67_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_77),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_72),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_73),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_82),
.B(n_79),
.Y(n_85)
);

NAND2x1p5_ASAP7_75t_L g86 ( 
.A(n_84),
.B(n_57),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_48),
.Y(n_87)
);

AOI211xp5_ASAP7_75t_SL g88 ( 
.A1(n_85),
.A2(n_81),
.B(n_83),
.C(n_23),
.Y(n_88)
);

AOI221xp5_ASAP7_75t_L g89 ( 
.A1(n_87),
.A2(n_56),
.B1(n_45),
.B2(n_25),
.C(n_27),
.Y(n_89)
);

NOR3xp33_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_86),
.C(n_20),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_88),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_18),
.Y(n_93)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_92),
.Y(n_94)
);

AOI222xp33_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_28),
.B1(n_31),
.B2(n_32),
.C1(n_33),
.C2(n_34),
.Y(n_95)
);

AOI221xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_94),
.B1(n_36),
.B2(n_37),
.C(n_39),
.Y(n_96)
);


endmodule