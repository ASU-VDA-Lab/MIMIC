module fake_netlist_6_384_n_2024 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_193, n_147, n_154, n_191, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_195, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_197, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_196, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_198, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_194, n_171, n_31, n_192, n_57, n_169, n_53, n_51, n_44, n_56, n_2024);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_193;
input n_147;
input n_154;
input n_191;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_195;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_197;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_196;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_194;
input n_171;
input n_31;
input n_192;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_2024;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1371;
wire n_1285;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1517;
wire n_1393;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_2019;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1912;
wire n_1563;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_2008;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_627;
wire n_595;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_851;
wire n_682;
wire n_644;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_1999;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_2002;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1993;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_2023;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_2016;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_575;
wire n_368;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_1997;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_2017;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_2021;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_2020;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_2005;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_2022;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_2015;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_2014;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_924;
wire n_475;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_2010;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_1996;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_2001;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1856;
wire n_1862;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx2_ASAP7_75t_SL g199 ( 
.A(n_27),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_156),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_76),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_188),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_136),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_149),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_178),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_145),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_59),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_9),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_117),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_140),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_194),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_74),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_80),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_161),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_135),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_124),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_7),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_64),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_86),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_109),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_61),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_24),
.Y(n_223)
);

BUFx10_ASAP7_75t_L g224 ( 
.A(n_163),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_0),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_57),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_92),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_123),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_41),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_63),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_114),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_73),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_111),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_72),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_198),
.Y(n_235)
);

BUFx5_ASAP7_75t_L g236 ( 
.A(n_98),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_81),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_187),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_142),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_32),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_174),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_8),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_147),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_78),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_12),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_83),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_89),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_191),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_110),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_61),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_40),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_12),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_67),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_134),
.Y(n_254)
);

BUFx10_ASAP7_75t_L g255 ( 
.A(n_26),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_18),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_175),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_52),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_35),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_159),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_96),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_84),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_7),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_59),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_168),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_154),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_26),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_43),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_126),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_91),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_57),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_50),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_100),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_36),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_94),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_53),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_193),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_190),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_166),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_5),
.Y(n_281)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_185),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_180),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_158),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_21),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_162),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_184),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_88),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_69),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_133),
.Y(n_290)
);

BUFx2_ASAP7_75t_L g291 ( 
.A(n_21),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_22),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_122),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_27),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_186),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_53),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_3),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_189),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_36),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_167),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_20),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_102),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_2),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_160),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g305 ( 
.A(n_129),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_66),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_22),
.Y(n_307)
);

INVx3_ASAP7_75t_L g308 ( 
.A(n_4),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_179),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_0),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_85),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_15),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_127),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_119),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_58),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_112),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g317 ( 
.A(n_196),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_60),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_70),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_82),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_152),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_153),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_79),
.Y(n_323)
);

INVx1_ASAP7_75t_SL g324 ( 
.A(n_115),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_28),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_146),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_71),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_177),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_68),
.Y(n_329)
);

BUFx6f_ASAP7_75t_L g330 ( 
.A(n_38),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_54),
.Y(n_331)
);

BUFx3_ASAP7_75t_L g332 ( 
.A(n_132),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_151),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_9),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_170),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_120),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_46),
.Y(n_337)
);

INVxp33_ASAP7_75t_SL g338 ( 
.A(n_40),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_143),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_14),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_4),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_35),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_2),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_75),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_19),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_43),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_107),
.Y(n_347)
);

BUFx5_ASAP7_75t_L g348 ( 
.A(n_65),
.Y(n_348)
);

INVxp33_ASAP7_75t_R g349 ( 
.A(n_17),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_20),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_41),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_49),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_169),
.Y(n_353)
);

INVxp33_ASAP7_75t_SL g354 ( 
.A(n_47),
.Y(n_354)
);

BUFx2_ASAP7_75t_L g355 ( 
.A(n_77),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_18),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_192),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_87),
.Y(n_358)
);

BUFx5_ASAP7_75t_L g359 ( 
.A(n_25),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_47),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_172),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_173),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_125),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_48),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_90),
.Y(n_365)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_44),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_37),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_56),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_183),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_121),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_104),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_39),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_137),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_15),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_105),
.Y(n_375)
);

INVx2_ASAP7_75t_SL g376 ( 
.A(n_11),
.Y(n_376)
);

BUFx3_ASAP7_75t_L g377 ( 
.A(n_118),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_138),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_139),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_11),
.Y(n_380)
);

BUFx8_ASAP7_75t_SL g381 ( 
.A(n_48),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_6),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_58),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_29),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_93),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_157),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_52),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_44),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_14),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_6),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_155),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_32),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_131),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_17),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_56),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_33),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_34),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_322),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_359),
.Y(n_399)
);

BUFx2_ASAP7_75t_SL g400 ( 
.A(n_217),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_217),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_359),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_359),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_232),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_359),
.Y(n_405)
);

INVxp67_ASAP7_75t_SL g406 ( 
.A(n_355),
.Y(n_406)
);

BUFx3_ASAP7_75t_L g407 ( 
.A(n_332),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

INVxp67_ASAP7_75t_SL g409 ( 
.A(n_308),
.Y(n_409)
);

HB1xp67_ASAP7_75t_L g410 ( 
.A(n_381),
.Y(n_410)
);

INVxp67_ASAP7_75t_SL g411 ( 
.A(n_308),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_308),
.Y(n_412)
);

CKINVDCx20_ASAP7_75t_R g413 ( 
.A(n_232),
.Y(n_413)
);

INVxp33_ASAP7_75t_SL g414 ( 
.A(n_218),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_359),
.Y(n_415)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_332),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_359),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_259),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_259),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_259),
.Y(n_420)
);

INVxp67_ASAP7_75t_SL g421 ( 
.A(n_377),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g422 ( 
.A(n_274),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_259),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_330),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_330),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_330),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_274),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_316),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_377),
.Y(n_429)
);

BUFx2_ASAP7_75t_L g430 ( 
.A(n_285),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_381),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_330),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_325),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_325),
.Y(n_434)
);

BUFx5_ASAP7_75t_L g435 ( 
.A(n_200),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_316),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_360),
.Y(n_437)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_236),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_360),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_218),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_211),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_245),
.Y(n_442)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_205),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_207),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_225),
.Y(n_445)
);

INVx1_ASAP7_75t_SL g446 ( 
.A(n_291),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_226),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_250),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g449 ( 
.A(n_206),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_252),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_294),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_296),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_236),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_297),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_301),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_307),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_337),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_340),
.Y(n_458)
);

BUFx2_ASAP7_75t_SL g459 ( 
.A(n_199),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_351),
.Y(n_460)
);

BUFx6f_ASAP7_75t_L g461 ( 
.A(n_201),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_352),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_256),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_364),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_236),
.Y(n_465)
);

INVxp67_ASAP7_75t_SL g466 ( 
.A(n_282),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_212),
.Y(n_467)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_366),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_382),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_397),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_389),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_202),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_203),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_236),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_199),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_236),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_376),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_376),
.Y(n_479)
);

HB1xp67_ASAP7_75t_L g480 ( 
.A(n_222),
.Y(n_480)
);

INVxp67_ASAP7_75t_SL g481 ( 
.A(n_282),
.Y(n_481)
);

BUFx3_ASAP7_75t_L g482 ( 
.A(n_224),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g483 ( 
.A(n_222),
.Y(n_483)
);

INVxp67_ASAP7_75t_SL g484 ( 
.A(n_282),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_213),
.Y(n_485)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_233),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_215),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_215),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_231),
.Y(n_489)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_231),
.Y(n_490)
);

BUFx6f_ASAP7_75t_L g491 ( 
.A(n_201),
.Y(n_491)
);

BUFx2_ASAP7_75t_L g492 ( 
.A(n_223),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_267),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_208),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_267),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_271),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_204),
.Y(n_497)
);

BUFx2_ASAP7_75t_L g498 ( 
.A(n_223),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g499 ( 
.A(n_461),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

OR2x2_ASAP7_75t_L g501 ( 
.A(n_446),
.B(n_277),
.Y(n_501)
);

AND2x4_ASAP7_75t_L g502 ( 
.A(n_466),
.B(n_271),
.Y(n_502)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_401),
.Y(n_503)
);

BUFx6f_ASAP7_75t_L g504 ( 
.A(n_461),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_409),
.B(n_280),
.Y(n_505)
);

AND2x4_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_280),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_484),
.B(n_338),
.Y(n_507)
);

AND2x2_ASAP7_75t_L g508 ( 
.A(n_411),
.B(n_335),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_399),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g510 ( 
.A(n_412),
.B(n_216),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_418),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_473),
.B(n_335),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_418),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_461),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_461),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_402),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_402),
.Y(n_517)
);

AND2x2_ASAP7_75t_SL g518 ( 
.A(n_461),
.B(n_393),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_403),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_419),
.Y(n_520)
);

HB1xp67_ASAP7_75t_L g521 ( 
.A(n_480),
.Y(n_521)
);

OA21x2_ASAP7_75t_L g522 ( 
.A1(n_487),
.A2(n_393),
.B(n_214),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_403),
.Y(n_523)
);

AND2x4_ASAP7_75t_L g524 ( 
.A(n_474),
.B(n_210),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_497),
.B(n_216),
.Y(n_525)
);

OAI21x1_ASAP7_75t_L g526 ( 
.A1(n_405),
.A2(n_243),
.B(n_228),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_405),
.Y(n_527)
);

CKINVDCx20_ASAP7_75t_R g528 ( 
.A(n_404),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_419),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_420),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

AND2x2_ASAP7_75t_L g532 ( 
.A(n_416),
.B(n_244),
.Y(n_532)
);

CKINVDCx8_ASAP7_75t_R g533 ( 
.A(n_400),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_420),
.Y(n_534)
);

INVx3_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

AND2x4_ASAP7_75t_L g536 ( 
.A(n_408),
.B(n_249),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_415),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_423),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_415),
.Y(n_539)
);

AND2x2_ASAP7_75t_L g540 ( 
.A(n_421),
.B(n_261),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_417),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_491),
.Y(n_542)
);

NAND2xp33_ASAP7_75t_L g543 ( 
.A(n_494),
.B(n_299),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_429),
.B(n_270),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_423),
.Y(n_545)
);

CKINVDCx20_ASAP7_75t_R g546 ( 
.A(n_413),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_424),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_407),
.B(n_288),
.Y(n_548)
);

CKINVDCx16_ASAP7_75t_R g549 ( 
.A(n_463),
.Y(n_549)
);

AND2x2_ASAP7_75t_L g550 ( 
.A(n_407),
.B(n_290),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_491),
.Y(n_551)
);

AOI22xp5_ASAP7_75t_L g552 ( 
.A1(n_468),
.A2(n_240),
.B1(n_251),
.B2(n_343),
.Y(n_552)
);

AND2x2_ASAP7_75t_SL g553 ( 
.A(n_491),
.B(n_201),
.Y(n_553)
);

BUFx6f_ASAP7_75t_L g554 ( 
.A(n_491),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_417),
.Y(n_555)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_459),
.B(n_209),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_438),
.Y(n_557)
);

HB1xp67_ASAP7_75t_L g558 ( 
.A(n_483),
.Y(n_558)
);

INVxp67_ASAP7_75t_L g559 ( 
.A(n_492),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g560 ( 
.A(n_459),
.B(n_300),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_422),
.A2(n_240),
.B1(n_251),
.B2(n_343),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_424),
.Y(n_562)
);

HB1xp67_ASAP7_75t_L g563 ( 
.A(n_492),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_425),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_425),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_438),
.Y(n_566)
);

HB1xp67_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_426),
.Y(n_568)
);

CKINVDCx20_ASAP7_75t_R g569 ( 
.A(n_427),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_426),
.Y(n_570)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_428),
.A2(n_387),
.B1(n_346),
.B2(n_392),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_453),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_432),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_453),
.Y(n_574)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_430),
.A2(n_346),
.B1(n_392),
.B2(n_390),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_443),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_432),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_449),
.Y(n_578)
);

AND2x6_ASAP7_75t_L g579 ( 
.A(n_465),
.B(n_201),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_487),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_505),
.B(n_435),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_516),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_569),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_SL g584 ( 
.A(n_556),
.B(n_494),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_SL g585 ( 
.A(n_556),
.B(n_442),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_556),
.B(n_442),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_516),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_500),
.Y(n_588)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_505),
.B(n_435),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_516),
.Y(n_590)
);

NOR2x1p5_ASAP7_75t_L g591 ( 
.A(n_501),
.B(n_431),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_517),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_500),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_517),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_500),
.Y(n_595)
);

INVx3_ASAP7_75t_L g596 ( 
.A(n_499),
.Y(n_596)
);

BUFx6f_ASAP7_75t_L g597 ( 
.A(n_499),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_509),
.Y(n_598)
);

AND2x6_ASAP7_75t_L g599 ( 
.A(n_502),
.B(n_260),
.Y(n_599)
);

INVx3_ASAP7_75t_L g600 ( 
.A(n_499),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_509),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_509),
.Y(n_602)
);

NAND3xp33_ASAP7_75t_L g603 ( 
.A(n_505),
.B(n_489),
.C(n_488),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_557),
.Y(n_604)
);

INVx3_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

NOR2x1p5_ASAP7_75t_L g606 ( 
.A(n_501),
.B(n_431),
.Y(n_606)
);

INVx3_ASAP7_75t_L g607 ( 
.A(n_499),
.Y(n_607)
);

INVx2_ASAP7_75t_L g608 ( 
.A(n_557),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_SL g609 ( 
.A(n_501),
.B(n_441),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_557),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_517),
.Y(n_611)
);

BUFx6f_ASAP7_75t_SL g612 ( 
.A(n_502),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_519),
.Y(n_613)
);

INVx8_ASAP7_75t_L g614 ( 
.A(n_502),
.Y(n_614)
);

INVx2_ASAP7_75t_SL g615 ( 
.A(n_560),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_519),
.Y(n_616)
);

BUFx6f_ASAP7_75t_SL g617 ( 
.A(n_502),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_502),
.A2(n_430),
.B1(n_406),
.B2(n_398),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_519),
.Y(n_619)
);

OAI22xp33_ASAP7_75t_L g620 ( 
.A1(n_559),
.A2(n_354),
.B1(n_338),
.B2(n_230),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_566),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_566),
.Y(n_622)
);

INVx2_ASAP7_75t_SL g623 ( 
.A(n_560),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_508),
.B(n_435),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_499),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_523),
.Y(n_626)
);

BUFx2_ASAP7_75t_L g627 ( 
.A(n_563),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_SL g628 ( 
.A(n_533),
.B(n_414),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_566),
.Y(n_629)
);

INVx3_ASAP7_75t_L g630 ( 
.A(n_499),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_523),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_574),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_523),
.Y(n_633)
);

CKINVDCx20_ASAP7_75t_R g634 ( 
.A(n_503),
.Y(n_634)
);

INVx3_ASAP7_75t_L g635 ( 
.A(n_504),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_504),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_527),
.Y(n_637)
);

AOI22xp33_ASAP7_75t_L g638 ( 
.A1(n_506),
.A2(n_498),
.B1(n_440),
.B2(n_354),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_536),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_527),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_574),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_504),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_536),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_574),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_527),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_533),
.B(n_440),
.Y(n_646)
);

BUFx3_ASAP7_75t_L g647 ( 
.A(n_536),
.Y(n_647)
);

NAND3xp33_ASAP7_75t_L g648 ( 
.A(n_508),
.B(n_489),
.C(n_488),
.Y(n_648)
);

NAND2xp5_ASAP7_75t_L g649 ( 
.A(n_506),
.B(n_435),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_531),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_531),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_531),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_537),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_SL g654 ( 
.A(n_510),
.B(n_467),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_504),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_537),
.Y(n_656)
);

INVx1_ASAP7_75t_L g657 ( 
.A(n_537),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_539),
.Y(n_658)
);

NAND3xp33_ASAP7_75t_L g659 ( 
.A(n_532),
.B(n_544),
.C(n_540),
.Y(n_659)
);

INVx3_ASAP7_75t_L g660 ( 
.A(n_504),
.Y(n_660)
);

INVx3_ASAP7_75t_L g661 ( 
.A(n_504),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_548),
.B(n_437),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_SL g663 ( 
.A(n_510),
.B(n_485),
.Y(n_663)
);

AOI21x1_ASAP7_75t_L g664 ( 
.A1(n_536),
.A2(n_493),
.B(n_490),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_576),
.Y(n_665)
);

NOR2xp33_ASAP7_75t_L g666 ( 
.A(n_507),
.B(n_486),
.Y(n_666)
);

AND2x2_ASAP7_75t_L g667 ( 
.A(n_548),
.B(n_439),
.Y(n_667)
);

NAND2xp33_ASAP7_75t_L g668 ( 
.A(n_560),
.B(n_260),
.Y(n_668)
);

NAND3xp33_ASAP7_75t_L g669 ( 
.A(n_532),
.B(n_493),
.C(n_490),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_539),
.Y(n_670)
);

INVx2_ASAP7_75t_SL g671 ( 
.A(n_506),
.Y(n_671)
);

INVxp33_ASAP7_75t_L g672 ( 
.A(n_563),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_539),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_541),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_541),
.Y(n_675)
);

INVx2_ASAP7_75t_SL g676 ( 
.A(n_506),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_SL g677 ( 
.A(n_507),
.B(n_482),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_SL g678 ( 
.A(n_553),
.B(n_482),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_L g679 ( 
.A1(n_559),
.A2(n_567),
.B1(n_525),
.B2(n_558),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_541),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_555),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_555),
.Y(n_682)
);

NOR2xp33_ASAP7_75t_L g683 ( 
.A(n_543),
.B(n_410),
.Y(n_683)
);

INVx4_ASAP7_75t_L g684 ( 
.A(n_579),
.Y(n_684)
);

AND2x2_ASAP7_75t_SL g685 ( 
.A(n_518),
.B(n_260),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_555),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_506),
.B(n_435),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_572),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_578),
.Y(n_689)
);

AND3x2_ASAP7_75t_L g690 ( 
.A(n_567),
.B(n_221),
.C(n_302),
.Y(n_690)
);

NOR2xp33_ASAP7_75t_L g691 ( 
.A(n_532),
.B(n_400),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_548),
.B(n_495),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_572),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_572),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_572),
.Y(n_695)
);

INVx2_ASAP7_75t_L g696 ( 
.A(n_572),
.Y(n_696)
);

INVx6_ASAP7_75t_L g697 ( 
.A(n_536),
.Y(n_697)
);

OR2x2_ASAP7_75t_L g698 ( 
.A(n_521),
.B(n_444),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_511),
.Y(n_699)
);

AOI21x1_ASAP7_75t_L g700 ( 
.A1(n_522),
.A2(n_496),
.B(n_495),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_511),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_540),
.B(n_544),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_513),
.Y(n_703)
);

NOR2xp33_ASAP7_75t_L g704 ( 
.A(n_540),
.B(n_436),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_513),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_550),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_504),
.Y(n_707)
);

INVx2_ASAP7_75t_L g708 ( 
.A(n_520),
.Y(n_708)
);

INVx2_ASAP7_75t_L g709 ( 
.A(n_520),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_553),
.B(n_224),
.Y(n_710)
);

OAI22xp33_ASAP7_75t_L g711 ( 
.A1(n_552),
.A2(n_242),
.B1(n_258),
.B2(n_229),
.Y(n_711)
);

AO22x2_ASAP7_75t_L g712 ( 
.A1(n_544),
.A2(n_309),
.B1(n_311),
.B2(n_304),
.Y(n_712)
);

NOR2xp33_ASAP7_75t_L g713 ( 
.A(n_525),
.B(n_521),
.Y(n_713)
);

BUFx4f_ASAP7_75t_L g714 ( 
.A(n_518),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_529),
.Y(n_715)
);

INVx3_ASAP7_75t_L g716 ( 
.A(n_514),
.Y(n_716)
);

AOI22xp33_ASAP7_75t_L g717 ( 
.A1(n_518),
.A2(n_496),
.B1(n_435),
.B2(n_447),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_518),
.B(n_435),
.Y(n_718)
);

AOI22xp33_ASAP7_75t_L g719 ( 
.A1(n_524),
.A2(n_454),
.B1(n_445),
.B2(n_448),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_553),
.B(n_220),
.Y(n_720)
);

HB1xp67_ASAP7_75t_L g721 ( 
.A(n_558),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_553),
.B(n_262),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_529),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_550),
.B(n_320),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_530),
.Y(n_725)
);

AO21x2_ASAP7_75t_L g726 ( 
.A1(n_526),
.A2(n_327),
.B(n_323),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_530),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_549),
.B(n_550),
.Y(n_728)
);

BUFx6f_ASAP7_75t_SL g729 ( 
.A(n_524),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_534),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_534),
.Y(n_731)
);

NAND2xp33_ASAP7_75t_SL g732 ( 
.A(n_591),
.B(n_387),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_714),
.B(n_549),
.Y(n_733)
);

O2A1O1Ixp33_ASAP7_75t_L g734 ( 
.A1(n_702),
.A2(n_524),
.B(n_512),
.C(n_580),
.Y(n_734)
);

NAND2xp33_ASAP7_75t_L g735 ( 
.A(n_614),
.B(n_236),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_671),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_676),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_676),
.B(n_524),
.Y(n_738)
);

BUFx3_ASAP7_75t_L g739 ( 
.A(n_639),
.Y(n_739)
);

NAND2xp33_ASAP7_75t_L g740 ( 
.A(n_614),
.B(n_236),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_615),
.B(n_623),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_639),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_627),
.B(n_575),
.Y(n_743)
);

INVxp67_ASAP7_75t_L g744 ( 
.A(n_713),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_639),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_643),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_SL g747 ( 
.A(n_714),
.B(n_260),
.Y(n_747)
);

AOI22xp33_ASAP7_75t_L g748 ( 
.A1(n_685),
.A2(n_522),
.B1(n_526),
.B2(n_512),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_714),
.B(n_286),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_615),
.B(n_512),
.Y(n_750)
);

AOI22xp33_ASAP7_75t_L g751 ( 
.A1(n_685),
.A2(n_522),
.B1(n_526),
.B2(n_512),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_588),
.Y(n_752)
);

INVx2_ASAP7_75t_SL g753 ( 
.A(n_698),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_685),
.B(n_286),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_623),
.B(n_286),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_643),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_706),
.B(n_512),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_593),
.Y(n_758)
);

AOI22xp5_ASAP7_75t_L g759 ( 
.A1(n_691),
.A2(n_324),
.B1(n_235),
.B2(n_237),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_SL g760 ( 
.A(n_659),
.B(n_286),
.Y(n_760)
);

AOI22xp33_ASAP7_75t_L g761 ( 
.A1(n_712),
.A2(n_522),
.B1(n_390),
.B2(n_339),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_701),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_720),
.B(n_538),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_643),
.Y(n_764)
);

INVxp33_ASAP7_75t_L g765 ( 
.A(n_721),
.Y(n_765)
);

NOR2xp33_ASAP7_75t_L g766 ( 
.A(n_659),
.B(n_219),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_647),
.Y(n_767)
);

NAND2xp33_ASAP7_75t_L g768 ( 
.A(n_614),
.B(n_348),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_722),
.B(n_545),
.Y(n_769)
);

INVx3_ASAP7_75t_L g770 ( 
.A(n_647),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_581),
.B(n_545),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_647),
.Y(n_772)
);

NOR2xp67_ASAP7_75t_L g773 ( 
.A(n_666),
.B(n_580),
.Y(n_773)
);

NAND3xp33_ASAP7_75t_L g774 ( 
.A(n_638),
.B(n_552),
.C(n_575),
.Y(n_774)
);

OR2x2_ASAP7_75t_SL g775 ( 
.A(n_698),
.B(n_349),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_SL g776 ( 
.A(n_589),
.B(n_287),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_SL g777 ( 
.A(n_624),
.B(n_287),
.Y(n_777)
);

NOR2xp33_ASAP7_75t_L g778 ( 
.A(n_677),
.B(n_219),
.Y(n_778)
);

AOI22xp33_ASAP7_75t_L g779 ( 
.A1(n_712),
.A2(n_522),
.B1(n_353),
.B2(n_386),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_614),
.B(n_547),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_614),
.B(n_547),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_593),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_718),
.B(n_287),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_595),
.Y(n_784)
);

NOR2xp33_ASAP7_75t_L g785 ( 
.A(n_679),
.B(n_227),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_627),
.B(n_561),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_584),
.B(n_227),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_649),
.B(n_305),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_704),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_SL g790 ( 
.A(n_665),
.B(n_561),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_SL g791 ( 
.A(n_665),
.B(n_689),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_692),
.B(n_699),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_672),
.B(n_476),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_697),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_SL g795 ( 
.A(n_687),
.B(n_305),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_684),
.B(n_717),
.Y(n_796)
);

BUFx6f_ASAP7_75t_L g797 ( 
.A(n_697),
.Y(n_797)
);

AND2x2_ASAP7_75t_L g798 ( 
.A(n_662),
.B(n_476),
.Y(n_798)
);

INVx2_ASAP7_75t_L g799 ( 
.A(n_703),
.Y(n_799)
);

INVx8_ASAP7_75t_L g800 ( 
.A(n_729),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_654),
.B(n_663),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_699),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_697),
.Y(n_803)
);

NOR3xp33_ASAP7_75t_L g804 ( 
.A(n_609),
.B(n_571),
.C(n_451),
.Y(n_804)
);

INVx4_ASAP7_75t_L g805 ( 
.A(n_697),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_SL g806 ( 
.A(n_684),
.B(n_305),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_L g807 ( 
.A(n_692),
.B(n_562),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_712),
.A2(n_333),
.B1(n_348),
.B2(n_305),
.Y(n_808)
);

INVx2_ASAP7_75t_L g809 ( 
.A(n_703),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_585),
.B(n_328),
.Y(n_810)
);

AND2x4_ASAP7_75t_L g811 ( 
.A(n_662),
.B(n_450),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_715),
.B(n_562),
.Y(n_812)
);

OR2x2_ASAP7_75t_L g813 ( 
.A(n_618),
.B(n_571),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_715),
.Y(n_814)
);

HB1xp67_ASAP7_75t_L g815 ( 
.A(n_728),
.Y(n_815)
);

INVxp67_ASAP7_75t_SL g816 ( 
.A(n_597),
.Y(n_816)
);

NOR2xp67_ASAP7_75t_L g817 ( 
.A(n_669),
.B(n_564),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_684),
.B(n_317),
.Y(n_818)
);

AOI22xp5_ASAP7_75t_L g819 ( 
.A1(n_612),
.A2(n_347),
.B1(n_336),
.B2(n_329),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_723),
.B(n_727),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_727),
.B(n_564),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_667),
.B(n_478),
.Y(n_822)
);

INVx8_ASAP7_75t_L g823 ( 
.A(n_729),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_667),
.B(n_452),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_684),
.B(n_678),
.Y(n_825)
);

NOR3xp33_ASAP7_75t_L g826 ( 
.A(n_586),
.B(n_456),
.C(n_455),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_L g827 ( 
.A(n_730),
.B(n_724),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_SL g829 ( 
.A(n_710),
.B(n_317),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_705),
.Y(n_830)
);

NAND3xp33_ASAP7_75t_L g831 ( 
.A(n_669),
.B(n_264),
.C(n_263),
.Y(n_831)
);

HB1xp67_ASAP7_75t_L g832 ( 
.A(n_634),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_628),
.B(n_478),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_598),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_646),
.B(n_479),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_708),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_L g837 ( 
.A(n_708),
.B(n_565),
.Y(n_837)
);

AOI22xp5_ASAP7_75t_L g838 ( 
.A1(n_612),
.A2(n_357),
.B1(n_248),
.B2(n_247),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_683),
.B(n_328),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_612),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_591),
.B(n_479),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_709),
.B(n_317),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_709),
.B(n_568),
.Y(n_843)
);

NAND2xp33_ASAP7_75t_L g844 ( 
.A(n_599),
.B(n_348),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_725),
.B(n_568),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_725),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_731),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_598),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_617),
.Y(n_849)
);

AND2x4_ASAP7_75t_L g850 ( 
.A(n_603),
.B(n_457),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_731),
.Y(n_851)
);

NOR2xp67_ASAP7_75t_L g852 ( 
.A(n_603),
.B(n_570),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_SL g853 ( 
.A(n_645),
.B(n_317),
.Y(n_853)
);

INVx2_ASAP7_75t_SL g854 ( 
.A(n_690),
.Y(n_854)
);

INVx2_ASAP7_75t_SL g855 ( 
.A(n_606),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_L g856 ( 
.A(n_668),
.B(n_570),
.Y(n_856)
);

OR2x6_ASAP7_75t_L g857 ( 
.A(n_606),
.B(n_458),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_620),
.B(n_391),
.Y(n_858)
);

NAND2xp5_ASAP7_75t_L g859 ( 
.A(n_693),
.B(n_573),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_693),
.B(n_573),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_694),
.B(n_577),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_648),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_694),
.B(n_577),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_601),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_SL g865 ( 
.A(n_645),
.B(n_326),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_601),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_653),
.B(n_326),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_582),
.B(n_515),
.Y(n_868)
);

NOR2xp33_ASAP7_75t_R g869 ( 
.A(n_689),
.B(n_503),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_602),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_582),
.B(n_515),
.Y(n_871)
);

BUFx3_ASAP7_75t_L g872 ( 
.A(n_583),
.Y(n_872)
);

INVx3_ASAP7_75t_L g873 ( 
.A(n_617),
.Y(n_873)
);

BUFx8_ASAP7_75t_L g874 ( 
.A(n_729),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_587),
.B(n_515),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_602),
.Y(n_876)
);

NOR2xp33_ASAP7_75t_L g877 ( 
.A(n_711),
.B(n_617),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_587),
.B(n_515),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_590),
.B(n_515),
.Y(n_879)
);

INVx2_ASAP7_75t_L g880 ( 
.A(n_604),
.Y(n_880)
);

INVx2_ASAP7_75t_L g881 ( 
.A(n_604),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_590),
.B(n_535),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_592),
.B(n_535),
.Y(n_883)
);

INVx2_ASAP7_75t_L g884 ( 
.A(n_608),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_648),
.B(n_391),
.Y(n_885)
);

OAI22xp5_ASAP7_75t_L g886 ( 
.A1(n_712),
.A2(n_719),
.B1(n_594),
.B2(n_611),
.Y(n_886)
);

OR2x2_ASAP7_75t_L g887 ( 
.A(n_726),
.B(n_460),
.Y(n_887)
);

OAI22xp33_ASAP7_75t_L g888 ( 
.A1(n_700),
.A2(n_299),
.B1(n_388),
.B2(n_394),
.Y(n_888)
);

AO22x2_ASAP7_75t_L g889 ( 
.A1(n_592),
.A2(n_471),
.B1(n_470),
.B2(n_464),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_594),
.B(n_535),
.Y(n_890)
);

NOR3xp33_ASAP7_75t_L g891 ( 
.A(n_664),
.B(n_469),
.C(n_462),
.Y(n_891)
);

NAND2xp5_ASAP7_75t_L g892 ( 
.A(n_611),
.B(n_535),
.Y(n_892)
);

AND2x4_ASAP7_75t_L g893 ( 
.A(n_664),
.B(n_472),
.Y(n_893)
);

NAND2xp33_ASAP7_75t_L g894 ( 
.A(n_599),
.B(n_348),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_613),
.B(n_535),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_762),
.Y(n_896)
);

INVx2_ASAP7_75t_SL g897 ( 
.A(n_793),
.Y(n_897)
);

AND2x6_ASAP7_75t_L g898 ( 
.A(n_862),
.B(n_840),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_798),
.Y(n_899)
);

BUFx6f_ASAP7_75t_L g900 ( 
.A(n_797),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_827),
.B(n_613),
.Y(n_901)
);

BUFx6f_ASAP7_75t_L g902 ( 
.A(n_797),
.Y(n_902)
);

HB1xp67_ASAP7_75t_L g903 ( 
.A(n_815),
.Y(n_903)
);

AND2x4_ASAP7_75t_L g904 ( 
.A(n_739),
.B(n_464),
.Y(n_904)
);

INVx2_ASAP7_75t_SL g905 ( 
.A(n_822),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_744),
.B(n_528),
.Y(n_906)
);

INVx2_ASAP7_75t_SL g907 ( 
.A(n_811),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_799),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_741),
.B(n_616),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_773),
.B(n_234),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_801),
.A2(n_599),
.B1(n_726),
.B2(n_619),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_763),
.B(n_616),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_809),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_769),
.B(n_619),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_820),
.B(n_792),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_870),
.Y(n_916)
);

INVx1_ASAP7_75t_SL g917 ( 
.A(n_869),
.Y(n_917)
);

NOR2xp33_ASAP7_75t_L g918 ( 
.A(n_839),
.B(n_528),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_802),
.B(n_626),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_796),
.A2(n_631),
.B(n_626),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_736),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_801),
.A2(n_839),
.B1(n_733),
.B2(n_745),
.Y(n_922)
);

AND2x4_ASAP7_75t_L g923 ( 
.A(n_739),
.B(n_470),
.Y(n_923)
);

INVx2_ASAP7_75t_L g924 ( 
.A(n_870),
.Y(n_924)
);

CKINVDCx20_ASAP7_75t_R g925 ( 
.A(n_869),
.Y(n_925)
);

NOR2x1p5_ASAP7_75t_L g926 ( 
.A(n_774),
.B(n_388),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_880),
.Y(n_927)
);

INVx2_ASAP7_75t_L g928 ( 
.A(n_880),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_737),
.Y(n_929)
);

BUFx3_ASAP7_75t_L g930 ( 
.A(n_872),
.Y(n_930)
);

BUFx6f_ASAP7_75t_L g931 ( 
.A(n_797),
.Y(n_931)
);

AOI22xp5_ASAP7_75t_L g932 ( 
.A1(n_733),
.A2(n_599),
.B1(n_726),
.B2(n_658),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_830),
.Y(n_933)
);

NOR2xp33_ASAP7_75t_L g934 ( 
.A(n_765),
.B(n_546),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_881),
.Y(n_935)
);

BUFx6f_ASAP7_75t_L g936 ( 
.A(n_803),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_770),
.Y(n_937)
);

INVx2_ASAP7_75t_SL g938 ( 
.A(n_811),
.Y(n_938)
);

INVx3_ASAP7_75t_L g939 ( 
.A(n_770),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_836),
.Y(n_940)
);

NAND2x1p5_ASAP7_75t_L g941 ( 
.A(n_805),
.B(n_600),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_846),
.Y(n_942)
);

CKINVDCx5p33_ASAP7_75t_R g943 ( 
.A(n_872),
.Y(n_943)
);

NAND2xp5_ASAP7_75t_L g944 ( 
.A(n_814),
.B(n_631),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_800),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_881),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_884),
.Y(n_947)
);

AND2x4_ASAP7_75t_L g948 ( 
.A(n_824),
.B(n_849),
.Y(n_948)
);

INVx4_ASAP7_75t_L g949 ( 
.A(n_803),
.Y(n_949)
);

INVx2_ASAP7_75t_L g950 ( 
.A(n_884),
.Y(n_950)
);

INVx4_ASAP7_75t_L g951 ( 
.A(n_803),
.Y(n_951)
);

INVxp67_ASAP7_75t_SL g952 ( 
.A(n_803),
.Y(n_952)
);

AND2x2_ASAP7_75t_L g953 ( 
.A(n_753),
.B(n_546),
.Y(n_953)
);

INVx2_ASAP7_75t_SL g954 ( 
.A(n_824),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_847),
.Y(n_955)
);

OR2x2_ASAP7_75t_L g956 ( 
.A(n_743),
.B(n_471),
.Y(n_956)
);

OR2x6_ASAP7_75t_L g957 ( 
.A(n_800),
.B(n_433),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_766),
.A2(n_599),
.B1(n_658),
.B2(n_657),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_800),
.B(n_433),
.Y(n_959)
);

BUFx12f_ASAP7_75t_SL g960 ( 
.A(n_857),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_828),
.B(n_633),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_851),
.Y(n_962)
);

NAND2xp33_ASAP7_75t_L g963 ( 
.A(n_887),
.B(n_599),
.Y(n_963)
);

AND2x4_ASAP7_75t_L g964 ( 
.A(n_849),
.B(n_434),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_742),
.Y(n_965)
);

AOI22xp33_ASAP7_75t_L g966 ( 
.A1(n_766),
.A2(n_675),
.B1(n_637),
.B2(n_651),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_746),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_756),
.Y(n_968)
);

BUFx2_ASAP7_75t_SL g969 ( 
.A(n_840),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_794),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_771),
.B(n_637),
.Y(n_971)
);

AND2x6_ASAP7_75t_L g972 ( 
.A(n_873),
.B(n_640),
.Y(n_972)
);

AND2x6_ASAP7_75t_L g973 ( 
.A(n_873),
.B(n_640),
.Y(n_973)
);

AO22x1_ASAP7_75t_L g974 ( 
.A1(n_858),
.A2(n_394),
.B1(n_395),
.B2(n_396),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_841),
.Y(n_975)
);

INVx3_ASAP7_75t_L g976 ( 
.A(n_794),
.Y(n_976)
);

OR2x2_ASAP7_75t_L g977 ( 
.A(n_786),
.B(n_395),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_823),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_764),
.Y(n_979)
);

BUFx3_ASAP7_75t_L g980 ( 
.A(n_832),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_750),
.B(n_650),
.Y(n_981)
);

INVx1_ASAP7_75t_L g982 ( 
.A(n_767),
.Y(n_982)
);

INVx1_ASAP7_75t_L g983 ( 
.A(n_772),
.Y(n_983)
);

OAI22xp33_ASAP7_75t_SL g984 ( 
.A1(n_813),
.A2(n_396),
.B1(n_275),
.B2(n_273),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_837),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_L g986 ( 
.A(n_760),
.B(n_651),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_757),
.B(n_652),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_738),
.A2(n_656),
.B(n_653),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_843),
.Y(n_989)
);

INVx5_ASAP7_75t_L g990 ( 
.A(n_805),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_L g991 ( 
.A(n_850),
.B(n_807),
.Y(n_991)
);

NOR2xp33_ASAP7_75t_L g992 ( 
.A(n_787),
.B(n_265),
.Y(n_992)
);

INVx2_ASAP7_75t_L g993 ( 
.A(n_752),
.Y(n_993)
);

NOR2xp33_ASAP7_75t_SL g994 ( 
.A(n_823),
.B(n_224),
.Y(n_994)
);

INVx3_ASAP7_75t_L g995 ( 
.A(n_758),
.Y(n_995)
);

AOI22xp5_ASAP7_75t_L g996 ( 
.A1(n_877),
.A2(n_829),
.B1(n_787),
.B2(n_810),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_874),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_782),
.Y(n_998)
);

BUFx3_ASAP7_75t_L g999 ( 
.A(n_874),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_850),
.B(n_652),
.Y(n_1000)
);

INVx5_ASAP7_75t_L g1001 ( 
.A(n_823),
.Y(n_1001)
);

AOI22xp33_ASAP7_75t_L g1002 ( 
.A1(n_761),
.A2(n_657),
.B1(n_673),
.B2(n_675),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_732),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_893),
.B(n_673),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_893),
.B(n_680),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_845),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_748),
.B(n_680),
.Y(n_1007)
);

INVx2_ASAP7_75t_L g1008 ( 
.A(n_784),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_812),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_748),
.B(n_681),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_751),
.B(n_681),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_785),
.B(n_269),
.C(n_268),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_825),
.A2(n_670),
.B(n_656),
.Y(n_1013)
);

AND2x2_ASAP7_75t_L g1014 ( 
.A(n_833),
.B(n_255),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_821),
.Y(n_1015)
);

BUFx4f_ASAP7_75t_L g1016 ( 
.A(n_857),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_835),
.B(n_255),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_791),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_SL g1019 ( 
.A(n_810),
.B(n_238),
.Y(n_1019)
);

AO22x1_ASAP7_75t_L g1020 ( 
.A1(n_858),
.A2(n_785),
.B1(n_877),
.B2(n_804),
.Y(n_1020)
);

AND2x4_ASAP7_75t_L g1021 ( 
.A(n_855),
.B(n_434),
.Y(n_1021)
);

OAI22xp33_ASAP7_75t_L g1022 ( 
.A1(n_759),
.A2(n_326),
.B1(n_310),
.B2(n_303),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_857),
.Y(n_1023)
);

INVx2_ASAP7_75t_SL g1024 ( 
.A(n_854),
.Y(n_1024)
);

NAND3xp33_ASAP7_75t_L g1025 ( 
.A(n_891),
.B(n_682),
.C(n_674),
.Y(n_1025)
);

AND2x4_ASAP7_75t_L g1026 ( 
.A(n_826),
.B(n_600),
.Y(n_1026)
);

AOI22xp33_ASAP7_75t_L g1027 ( 
.A1(n_761),
.A2(n_682),
.B1(n_674),
.B2(n_686),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_SL g1028 ( 
.A(n_790),
.B(n_255),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_SL g1029 ( 
.A(n_778),
.B(n_239),
.Y(n_1029)
);

INVx4_ASAP7_75t_L g1030 ( 
.A(n_889),
.Y(n_1030)
);

AND2x4_ASAP7_75t_L g1031 ( 
.A(n_831),
.B(n_600),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_834),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_859),
.Y(n_1033)
);

OAI22xp5_ASAP7_75t_SL g1034 ( 
.A1(n_775),
.A2(n_331),
.B1(n_272),
.B2(n_384),
.Y(n_1034)
);

AOI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_829),
.A2(n_686),
.B1(n_670),
.B2(n_695),
.Y(n_1035)
);

NAND2xp33_ASAP7_75t_L g1036 ( 
.A(n_808),
.B(n_779),
.Y(n_1036)
);

AND2x4_ASAP7_75t_L g1037 ( 
.A(n_817),
.B(n_600),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_SL g1038 ( 
.A(n_778),
.B(n_241),
.Y(n_1038)
);

INVx2_ASAP7_75t_L g1039 ( 
.A(n_848),
.Y(n_1039)
);

AND2x6_ASAP7_75t_SL g1040 ( 
.A(n_885),
.B(n_281),
.Y(n_1040)
);

NOR3xp33_ASAP7_75t_SL g1041 ( 
.A(n_888),
.B(n_312),
.C(n_292),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_751),
.B(n_608),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_864),
.Y(n_1043)
);

NOR2xp33_ASAP7_75t_L g1044 ( 
.A(n_885),
.B(n_315),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_860),
.Y(n_1045)
);

INVx3_ASAP7_75t_L g1046 ( 
.A(n_866),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_861),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_SL g1048 ( 
.A(n_808),
.B(n_246),
.Y(n_1048)
);

O2A1O1Ixp33_ASAP7_75t_L g1049 ( 
.A1(n_888),
.A2(n_629),
.B(n_610),
.C(n_641),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_852),
.B(n_318),
.Y(n_1050)
);

BUFx8_ASAP7_75t_L g1051 ( 
.A(n_876),
.Y(n_1051)
);

INVx2_ASAP7_75t_L g1052 ( 
.A(n_868),
.Y(n_1052)
);

OAI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_779),
.A2(n_367),
.B1(n_374),
.B2(n_334),
.Y(n_1053)
);

OR2x4_ASAP7_75t_L g1054 ( 
.A(n_856),
.B(n_326),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_863),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_889),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_889),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_780),
.Y(n_1058)
);

BUFx2_ASAP7_75t_L g1059 ( 
.A(n_819),
.Y(n_1059)
);

INVx1_ASAP7_75t_L g1060 ( 
.A(n_871),
.Y(n_1060)
);

INVx2_ASAP7_75t_L g1061 ( 
.A(n_875),
.Y(n_1061)
);

OAI22xp5_ASAP7_75t_L g1062 ( 
.A1(n_754),
.A2(n_341),
.B1(n_372),
.B2(n_342),
.Y(n_1062)
);

NOR3xp33_ASAP7_75t_SL g1063 ( 
.A(n_886),
.B(n_345),
.C(n_350),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_825),
.B(n_747),
.Y(n_1064)
);

INVx1_ASAP7_75t_L g1065 ( 
.A(n_878),
.Y(n_1065)
);

NOR2xp33_ASAP7_75t_L g1066 ( 
.A(n_747),
.B(n_356),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_879),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_838),
.Y(n_1068)
);

NAND2xp5_ASAP7_75t_L g1069 ( 
.A(n_749),
.B(n_621),
.Y(n_1069)
);

INVx2_ASAP7_75t_SL g1070 ( 
.A(n_755),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_SL g1071 ( 
.A(n_755),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_882),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_996),
.B(n_781),
.Y(n_1073)
);

INVx1_ASAP7_75t_SL g1074 ( 
.A(n_953),
.Y(n_1074)
);

O2A1O1Ixp33_ASAP7_75t_L g1075 ( 
.A1(n_1044),
.A2(n_749),
.B(n_783),
.C(n_734),
.Y(n_1075)
);

OAI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1064),
.A2(n_783),
.B(n_777),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_990),
.A2(n_740),
.B(n_735),
.Y(n_1077)
);

AND2x2_ASAP7_75t_L g1078 ( 
.A(n_1014),
.B(n_776),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_SL g1079 ( 
.A(n_899),
.B(n_905),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_943),
.Y(n_1080)
);

OAI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_1064),
.A2(n_1042),
.B(n_920),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_915),
.B(n_816),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_R g1083 ( 
.A(n_925),
.B(n_768),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_930),
.Y(n_1084)
);

AND2x2_ASAP7_75t_L g1085 ( 
.A(n_1017),
.B(n_368),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_1009),
.B(n_883),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_916),
.Y(n_1087)
);

BUFx12f_ASAP7_75t_L g1088 ( 
.A(n_978),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_R g1089 ( 
.A(n_1003),
.B(n_844),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_990),
.A2(n_818),
.B(n_806),
.Y(n_1090)
);

AOI21xp5_ASAP7_75t_L g1091 ( 
.A1(n_990),
.A2(n_818),
.B(n_806),
.Y(n_1091)
);

NOR3xp33_ASAP7_75t_L g1092 ( 
.A(n_918),
.B(n_383),
.C(n_894),
.Y(n_1092)
);

O2A1O1Ixp33_ASAP7_75t_L g1093 ( 
.A1(n_1022),
.A2(n_842),
.B(n_788),
.C(n_795),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_924),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_906),
.B(n_890),
.Y(n_1095)
);

INVx2_ASAP7_75t_L g1096 ( 
.A(n_927),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_963),
.A2(n_915),
.B(n_971),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_SL g1098 ( 
.A(n_897),
.B(n_253),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_1066),
.A2(n_895),
.B(n_892),
.C(n_842),
.Y(n_1099)
);

NOR2xp33_ASAP7_75t_L g1100 ( 
.A(n_1020),
.B(n_596),
.Y(n_1100)
);

NAND2xp5_ASAP7_75t_L g1101 ( 
.A(n_1015),
.B(n_621),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_975),
.B(n_596),
.Y(n_1102)
);

BUFx6f_ASAP7_75t_L g1103 ( 
.A(n_978),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_928),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_991),
.B(n_622),
.Y(n_1105)
);

OR2x6_ASAP7_75t_L g1106 ( 
.A(n_978),
.B(n_867),
.Y(n_1106)
);

A2O1A1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_922),
.A2(n_867),
.B(n_865),
.C(n_853),
.Y(n_1107)
);

BUFx8_ASAP7_75t_L g1108 ( 
.A(n_997),
.Y(n_1108)
);

O2A1O1Ixp33_ASAP7_75t_L g1109 ( 
.A1(n_984),
.A2(n_865),
.B(n_853),
.C(n_632),
.Y(n_1109)
);

OAI21xp33_ASAP7_75t_L g1110 ( 
.A1(n_1028),
.A2(n_278),
.B(n_254),
.Y(n_1110)
);

INVx4_ASAP7_75t_L g1111 ( 
.A(n_1001),
.Y(n_1111)
);

OAI22xp5_ASAP7_75t_L g1112 ( 
.A1(n_991),
.A2(n_700),
.B1(n_632),
.B2(n_622),
.Y(n_1112)
);

OAI22xp5_ASAP7_75t_L g1113 ( 
.A1(n_901),
.A2(n_629),
.B1(n_641),
.B2(n_644),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_907),
.B(n_257),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_934),
.B(n_596),
.Y(n_1115)
);

NOR2xp33_ASAP7_75t_L g1116 ( 
.A(n_903),
.B(n_917),
.Y(n_1116)
);

AOI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_1042),
.A2(n_1036),
.B(n_1010),
.Y(n_1117)
);

HB1xp67_ASAP7_75t_L g1118 ( 
.A(n_980),
.Y(n_1118)
);

AO32x2_ASAP7_75t_L g1119 ( 
.A1(n_1030),
.A2(n_1),
.A3(n_5),
.B1(n_8),
.B2(n_10),
.Y(n_1119)
);

OAI22x1_ASAP7_75t_L g1120 ( 
.A1(n_1018),
.A2(n_276),
.B1(n_385),
.B2(n_379),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_917),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1033),
.B(n_644),
.Y(n_1122)
);

INVx2_ASAP7_75t_SL g1123 ( 
.A(n_1024),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_960),
.Y(n_1124)
);

NOR2x1_ASAP7_75t_L g1125 ( 
.A(n_949),
.B(n_605),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1045),
.B(n_605),
.Y(n_1126)
);

BUFx4f_ASAP7_75t_L g1127 ( 
.A(n_957),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_1007),
.A2(n_707),
.B(n_597),
.Y(n_1128)
);

AND2x2_ASAP7_75t_SL g1129 ( 
.A(n_994),
.B(n_688),
.Y(n_1129)
);

O2A1O1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_1012),
.A2(n_696),
.B(n_695),
.C(n_688),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1047),
.B(n_605),
.Y(n_1131)
);

AOI21xp5_ASAP7_75t_L g1132 ( 
.A1(n_1007),
.A2(n_1011),
.B(n_1010),
.Y(n_1132)
);

BUFx6f_ASAP7_75t_L g1133 ( 
.A(n_900),
.Y(n_1133)
);

INVx4_ASAP7_75t_L g1134 ( 
.A(n_1001),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_913),
.Y(n_1135)
);

AND2x2_ASAP7_75t_L g1136 ( 
.A(n_956),
.B(n_266),
.Y(n_1136)
);

NOR2xp33_ASAP7_75t_L g1137 ( 
.A(n_1018),
.B(n_655),
.Y(n_1137)
);

AOI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_1011),
.A2(n_707),
.B(n_597),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_900),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_896),
.Y(n_1140)
);

INVx3_ASAP7_75t_SL g1141 ( 
.A(n_1023),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_981),
.A2(n_707),
.B(n_636),
.Y(n_1142)
);

NOR2x1p5_ASAP7_75t_SL g1143 ( 
.A(n_1052),
.B(n_696),
.Y(n_1143)
);

A2O1A1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_1049),
.A2(n_635),
.B(n_605),
.C(n_661),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_900),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_1055),
.B(n_607),
.Y(n_1146)
);

O2A1O1Ixp33_ASAP7_75t_L g1147 ( 
.A1(n_1019),
.A2(n_465),
.B(n_475),
.C(n_477),
.Y(n_1147)
);

O2A1O1Ixp5_ASAP7_75t_L g1148 ( 
.A1(n_1029),
.A2(n_716),
.B(n_655),
.C(n_660),
.Y(n_1148)
);

AND2x2_ASAP7_75t_L g1149 ( 
.A(n_904),
.B(n_279),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_1040),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_SL g1151 ( 
.A(n_938),
.B(n_283),
.Y(n_1151)
);

NAND2x1p5_ASAP7_75t_L g1152 ( 
.A(n_1001),
.B(n_607),
.Y(n_1152)
);

AND2x2_ASAP7_75t_L g1153 ( 
.A(n_904),
.B(n_284),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1013),
.A2(n_630),
.B(n_607),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_977),
.B(n_655),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_1028),
.B(n_289),
.C(n_293),
.Y(n_1156)
);

INVx2_ASAP7_75t_L g1157 ( 
.A(n_935),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_954),
.B(n_295),
.Y(n_1158)
);

OAI22xp5_ASAP7_75t_L g1159 ( 
.A1(n_901),
.A2(n_1057),
.B1(n_1056),
.B2(n_912),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_908),
.Y(n_1160)
);

AND2x2_ASAP7_75t_L g1161 ( 
.A(n_923),
.B(n_298),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_SL g1162 ( 
.A(n_948),
.B(n_306),
.Y(n_1162)
);

AND2x4_ASAP7_75t_L g1163 ( 
.A(n_948),
.B(n_716),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_985),
.B(n_625),
.Y(n_1164)
);

NOR2xp33_ASAP7_75t_L g1165 ( 
.A(n_1059),
.B(n_716),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1063),
.A2(n_625),
.B(n_661),
.C(n_660),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_946),
.Y(n_1167)
);

INVx2_ASAP7_75t_L g1168 ( 
.A(n_947),
.Y(n_1168)
);

BUFx8_ASAP7_75t_SL g1169 ( 
.A(n_999),
.Y(n_1169)
);

INVx3_ASAP7_75t_L g1170 ( 
.A(n_902),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_950),
.Y(n_1171)
);

NOR2xp67_ASAP7_75t_SL g1172 ( 
.A(n_1001),
.B(n_313),
.Y(n_1172)
);

AOI22xp5_ASAP7_75t_L g1173 ( 
.A1(n_1068),
.A2(n_375),
.B1(n_319),
.B2(n_321),
.Y(n_1173)
);

CKINVDCx5p33_ASAP7_75t_R g1174 ( 
.A(n_945),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_987),
.A2(n_914),
.B(n_912),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_923),
.Y(n_1176)
);

OR2x6_ASAP7_75t_L g1177 ( 
.A(n_957),
.B(n_959),
.Y(n_1177)
);

NAND3xp33_ASAP7_75t_SL g1178 ( 
.A(n_994),
.B(n_314),
.C(n_344),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_1021),
.Y(n_1179)
);

NOR2x1_ASAP7_75t_L g1180 ( 
.A(n_949),
.B(n_625),
.Y(n_1180)
);

NAND2xp5_ASAP7_75t_L g1181 ( 
.A(n_989),
.B(n_625),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_945),
.Y(n_1182)
);

A2O1A1Ixp33_ASAP7_75t_SL g1183 ( 
.A1(n_1006),
.A2(n_635),
.B(n_661),
.C(n_660),
.Y(n_1183)
);

NOR2xp33_ASAP7_75t_L g1184 ( 
.A(n_921),
.B(n_630),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1058),
.B(n_358),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_933),
.Y(n_1186)
);

NAND2xp5_ASAP7_75t_L g1187 ( 
.A(n_1050),
.B(n_909),
.Y(n_1187)
);

INVx3_ASAP7_75t_L g1188 ( 
.A(n_902),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1051),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_929),
.B(n_630),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_995),
.Y(n_1191)
);

AOI22x1_ASAP7_75t_L g1192 ( 
.A1(n_1061),
.A2(n_660),
.B1(n_635),
.B2(n_630),
.Y(n_1192)
);

O2A1O1Ixp33_ASAP7_75t_L g1193 ( 
.A1(n_1038),
.A2(n_475),
.B(n_477),
.C(n_542),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_902),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_SL g1195 ( 
.A(n_1058),
.B(n_361),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_L g1196 ( 
.A1(n_1062),
.A2(n_542),
.B(n_551),
.C(n_16),
.Y(n_1196)
);

INVx3_ASAP7_75t_L g1197 ( 
.A(n_931),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1030),
.A2(n_362),
.B1(n_363),
.B2(n_365),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_940),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_942),
.Y(n_1200)
);

NOR2xp33_ASAP7_75t_R g1201 ( 
.A(n_1016),
.B(n_369),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_926),
.A2(n_370),
.B1(n_371),
.B2(n_373),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_995),
.Y(n_1203)
);

NOR2xp33_ASAP7_75t_L g1204 ( 
.A(n_1071),
.B(n_378),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_L g1205 ( 
.A1(n_1062),
.A2(n_542),
.B(n_551),
.C(n_16),
.Y(n_1205)
);

BUFx2_ASAP7_75t_L g1206 ( 
.A(n_1051),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_955),
.Y(n_1207)
);

OAI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1000),
.A2(n_707),
.B1(n_642),
.B2(n_551),
.Y(n_1208)
);

OAI21xp33_ASAP7_75t_L g1209 ( 
.A1(n_1053),
.A2(n_551),
.B(n_542),
.Y(n_1209)
);

NOR2xp33_ASAP7_75t_L g1210 ( 
.A(n_1071),
.B(n_642),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_909),
.B(n_642),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_L g1212 ( 
.A(n_931),
.Y(n_1212)
);

NAND2xp5_ASAP7_75t_L g1213 ( 
.A(n_1000),
.B(n_348),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_962),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1002),
.A2(n_542),
.B1(n_551),
.B2(n_19),
.Y(n_1215)
);

BUFx2_ASAP7_75t_L g1216 ( 
.A(n_957),
.Y(n_1216)
);

NOR2xp33_ASAP7_75t_L g1217 ( 
.A(n_1021),
.B(n_1),
.Y(n_1217)
);

INVx5_ASAP7_75t_L g1218 ( 
.A(n_898),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_919),
.Y(n_1219)
);

OAI22xp5_ASAP7_75t_L g1220 ( 
.A1(n_958),
.A2(n_13),
.B1(n_23),
.B2(n_24),
.Y(n_1220)
);

A2O1A1Ixp33_ASAP7_75t_L g1221 ( 
.A1(n_1070),
.A2(n_348),
.B(n_514),
.C(n_554),
.Y(n_1221)
);

OR2x2_ASAP7_75t_L g1222 ( 
.A(n_1074),
.B(n_1053),
.Y(n_1222)
);

OAI21x1_ASAP7_75t_L g1223 ( 
.A1(n_1154),
.A2(n_1013),
.B(n_988),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1219),
.B(n_1072),
.Y(n_1224)
);

NAND2xp5_ASAP7_75t_SL g1225 ( 
.A(n_1121),
.B(n_1016),
.Y(n_1225)
);

OR2x2_ASAP7_75t_L g1226 ( 
.A(n_1074),
.B(n_965),
.Y(n_1226)
);

AOI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1073),
.A2(n_988),
.B(n_1069),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1186),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1128),
.A2(n_1069),
.B(n_986),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1199),
.Y(n_1230)
);

BUFx2_ASAP7_75t_L g1231 ( 
.A(n_1118),
.Y(n_1231)
);

O2A1O1Ixp5_ASAP7_75t_L g1232 ( 
.A1(n_1166),
.A2(n_910),
.B(n_1048),
.C(n_1031),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_L g1233 ( 
.A(n_1174),
.B(n_898),
.Y(n_1233)
);

INVx1_ASAP7_75t_SL g1234 ( 
.A(n_1176),
.Y(n_1234)
);

CKINVDCx11_ASAP7_75t_R g1235 ( 
.A(n_1080),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1200),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1085),
.B(n_964),
.Y(n_1237)
);

INVx1_ASAP7_75t_L g1238 ( 
.A(n_1207),
.Y(n_1238)
);

AND2x2_ASAP7_75t_L g1239 ( 
.A(n_1136),
.B(n_964),
.Y(n_1239)
);

AO31x2_ASAP7_75t_L g1240 ( 
.A1(n_1159),
.A2(n_1221),
.A3(n_1112),
.B(n_1107),
.Y(n_1240)
);

NAND2x1p5_ASAP7_75t_L g1241 ( 
.A(n_1111),
.B(n_951),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1177),
.B(n_969),
.Y(n_1242)
);

NAND2x1_ASAP7_75t_L g1243 ( 
.A(n_1111),
.B(n_937),
.Y(n_1243)
);

NAND2xp33_ASAP7_75t_L g1244 ( 
.A(n_1182),
.B(n_898),
.Y(n_1244)
);

OAI21xp5_ASAP7_75t_L g1245 ( 
.A1(n_1117),
.A2(n_911),
.B(n_1025),
.Y(n_1245)
);

AOI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1077),
.A2(n_1005),
.B(n_1004),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_1214),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_L g1248 ( 
.A(n_1187),
.B(n_1060),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1169),
.Y(n_1249)
);

AOI21xp5_ASAP7_75t_L g1250 ( 
.A1(n_1082),
.A2(n_944),
.B(n_961),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1095),
.B(n_1041),
.C(n_974),
.Y(n_1251)
);

A2O1A1Ixp33_ASAP7_75t_L g1252 ( 
.A1(n_1075),
.A2(n_1026),
.B(n_932),
.C(n_982),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_1220),
.A2(n_1065),
.B(n_961),
.C(n_944),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1082),
.A2(n_919),
.B(n_952),
.Y(n_1254)
);

OR2x2_ASAP7_75t_L g1255 ( 
.A(n_1176),
.B(n_967),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1192),
.A2(n_941),
.B(n_966),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_L g1257 ( 
.A(n_1086),
.B(n_1067),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1142),
.A2(n_941),
.B(n_1035),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_SL g1259 ( 
.A(n_1116),
.B(n_1034),
.Y(n_1259)
);

AOI221x1_ASAP7_75t_L g1260 ( 
.A1(n_1159),
.A2(n_1025),
.B1(n_968),
.B2(n_983),
.C(n_979),
.Y(n_1260)
);

CKINVDCx8_ASAP7_75t_R g1261 ( 
.A(n_1103),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1087),
.Y(n_1262)
);

O2A1O1Ixp5_ASAP7_75t_SL g1263 ( 
.A1(n_1220),
.A2(n_1046),
.B(n_1032),
.C(n_939),
.Y(n_1263)
);

INVx1_ASAP7_75t_SL g1264 ( 
.A(n_1084),
.Y(n_1264)
);

BUFx3_ASAP7_75t_L g1265 ( 
.A(n_1088),
.Y(n_1265)
);

HB1xp67_ASAP7_75t_L g1266 ( 
.A(n_1179),
.Y(n_1266)
);

NOR2xp67_ASAP7_75t_L g1267 ( 
.A(n_1123),
.B(n_970),
.Y(n_1267)
);

BUFx3_ASAP7_75t_L g1268 ( 
.A(n_1103),
.Y(n_1268)
);

OAI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1132),
.A2(n_1027),
.B(n_1037),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1078),
.B(n_1032),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1090),
.A2(n_1091),
.B(n_1211),
.Y(n_1271)
);

AOI211x1_ASAP7_75t_L g1272 ( 
.A1(n_1215),
.A2(n_1054),
.B(n_23),
.C(n_25),
.Y(n_1272)
);

OA22x2_ASAP7_75t_L g1273 ( 
.A1(n_1177),
.A2(n_959),
.B1(n_1037),
.B2(n_1043),
.Y(n_1273)
);

INVx8_ASAP7_75t_L g1274 ( 
.A(n_1103),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_L g1275 ( 
.A1(n_1076),
.A2(n_970),
.B(n_976),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1134),
.Y(n_1276)
);

OA21x2_ASAP7_75t_L g1277 ( 
.A1(n_1076),
.A2(n_1081),
.B(n_1148),
.Y(n_1277)
);

AND2x2_ASAP7_75t_L g1278 ( 
.A(n_1149),
.B(n_959),
.Y(n_1278)
);

INVx1_ASAP7_75t_SL g1279 ( 
.A(n_1089),
.Y(n_1279)
);

NOR2xp67_ASAP7_75t_L g1280 ( 
.A(n_1178),
.B(n_976),
.Y(n_1280)
);

NOR2xp67_ASAP7_75t_L g1281 ( 
.A(n_1156),
.B(n_951),
.Y(n_1281)
);

NOR4xp25_ASAP7_75t_L g1282 ( 
.A(n_1196),
.B(n_1008),
.C(n_993),
.D(n_1039),
.Y(n_1282)
);

BUFx6f_ASAP7_75t_L g1283 ( 
.A(n_1133),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1081),
.B(n_1046),
.Y(n_1284)
);

A2O1A1Ixp33_ASAP7_75t_L g1285 ( 
.A1(n_1093),
.A2(n_998),
.B(n_931),
.C(n_936),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1124),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1153),
.B(n_1161),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_1105),
.B(n_1101),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1135),
.Y(n_1289)
);

OAI21x1_ASAP7_75t_L g1290 ( 
.A1(n_1112),
.A2(n_898),
.B(n_973),
.Y(n_1290)
);

INVxp67_ASAP7_75t_L g1291 ( 
.A(n_1079),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1099),
.A2(n_936),
.B(n_1054),
.Y(n_1292)
);

AO32x2_ASAP7_75t_L g1293 ( 
.A1(n_1215),
.A2(n_973),
.A3(n_972),
.B1(n_936),
.B2(n_30),
.Y(n_1293)
);

AOI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1204),
.A2(n_973),
.B1(n_972),
.B2(n_348),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1217),
.Y(n_1295)
);

O2A1O1Ixp5_ASAP7_75t_L g1296 ( 
.A1(n_1115),
.A2(n_973),
.B(n_972),
.C(n_29),
.Y(n_1296)
);

OAI21x1_ASAP7_75t_L g1297 ( 
.A1(n_1113),
.A2(n_108),
.B(n_197),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_1108),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1113),
.A2(n_106),
.B(n_195),
.Y(n_1299)
);

O2A1O1Ixp33_ASAP7_75t_L g1300 ( 
.A1(n_1205),
.A2(n_13),
.B(n_28),
.C(n_30),
.Y(n_1300)
);

AOI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1134),
.A2(n_514),
.B(n_554),
.Y(n_1301)
);

BUFx12f_ASAP7_75t_L g1302 ( 
.A(n_1108),
.Y(n_1302)
);

AOI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1213),
.A2(n_579),
.B(n_554),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1140),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1155),
.B(n_31),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1105),
.B(n_31),
.Y(n_1306)
);

NAND2xp5_ASAP7_75t_L g1307 ( 
.A(n_1122),
.B(n_579),
.Y(n_1307)
);

OR2x2_ASAP7_75t_L g1308 ( 
.A(n_1158),
.B(n_33),
.Y(n_1308)
);

BUFx4_ASAP7_75t_SL g1309 ( 
.A(n_1189),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_1141),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1165),
.B(n_34),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_SL g1312 ( 
.A1(n_1109),
.A2(n_1164),
.B(n_1130),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1100),
.A2(n_579),
.A3(n_39),
.B(n_42),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1137),
.B(n_38),
.Y(n_1314)
);

OAI21xp5_ASAP7_75t_L g1315 ( 
.A1(n_1209),
.A2(n_579),
.B(n_130),
.Y(n_1315)
);

AND2x2_ASAP7_75t_L g1316 ( 
.A(n_1083),
.B(n_42),
.Y(n_1316)
);

NOR3xp33_ASAP7_75t_SL g1317 ( 
.A(n_1150),
.B(n_45),
.C(n_46),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_1160),
.Y(n_1318)
);

AO31x2_ASAP7_75t_L g1319 ( 
.A1(n_1208),
.A2(n_579),
.A3(n_49),
.B(n_51),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1167),
.Y(n_1320)
);

NAND2xp5_ASAP7_75t_L g1321 ( 
.A(n_1164),
.B(n_579),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1092),
.A2(n_514),
.B(n_554),
.C(n_55),
.Y(n_1322)
);

A2O1A1Ixp33_ASAP7_75t_L g1323 ( 
.A1(n_1110),
.A2(n_1129),
.B(n_1143),
.C(n_1173),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1144),
.A2(n_579),
.B(n_128),
.Y(n_1324)
);

NAND3xp33_ASAP7_75t_L g1325 ( 
.A(n_1202),
.B(n_514),
.C(n_54),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1094),
.B(n_579),
.Y(n_1326)
);

AOI31xp67_ASAP7_75t_L g1327 ( 
.A1(n_1183),
.A2(n_116),
.A3(n_182),
.B(n_181),
.Y(n_1327)
);

OAI21xp5_ASAP7_75t_L g1328 ( 
.A1(n_1181),
.A2(n_113),
.B(n_176),
.Y(n_1328)
);

OAI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1126),
.A2(n_103),
.B(n_171),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1125),
.A2(n_101),
.B(n_165),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1171),
.Y(n_1331)
);

AND2x4_ASAP7_75t_L g1332 ( 
.A(n_1163),
.B(n_1177),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_1133),
.Y(n_1333)
);

NAND2xp5_ASAP7_75t_L g1334 ( 
.A(n_1096),
.B(n_45),
.Y(n_1334)
);

OAI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1218),
.A2(n_55),
.B1(n_60),
.B2(n_62),
.Y(n_1335)
);

A2O1A1Ixp33_ASAP7_75t_L g1336 ( 
.A1(n_1184),
.A2(n_514),
.B(n_63),
.C(n_62),
.Y(n_1336)
);

NOR2x1_ASAP7_75t_SL g1337 ( 
.A(n_1218),
.B(n_95),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1104),
.B(n_97),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1157),
.Y(n_1339)
);

A2O1A1Ixp33_ASAP7_75t_L g1340 ( 
.A1(n_1190),
.A2(n_99),
.B(n_141),
.C(n_144),
.Y(n_1340)
);

AOI21x1_ASAP7_75t_L g1341 ( 
.A1(n_1185),
.A2(n_148),
.B(n_150),
.Y(n_1341)
);

OA21x2_ASAP7_75t_L g1342 ( 
.A1(n_1131),
.A2(n_164),
.B(n_1146),
.Y(n_1342)
);

AOI21xp33_ASAP7_75t_L g1343 ( 
.A1(n_1198),
.A2(n_1120),
.B(n_1195),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1218),
.A2(n_1162),
.B(n_1098),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1180),
.A2(n_1152),
.B(n_1193),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1218),
.A2(n_1151),
.B(n_1114),
.Y(n_1346)
);

O2A1O1Ixp5_ASAP7_75t_SL g1347 ( 
.A1(n_1139),
.A2(n_1197),
.B(n_1188),
.C(n_1145),
.Y(n_1347)
);

NOR2xp67_ASAP7_75t_L g1348 ( 
.A(n_1191),
.B(n_1203),
.Y(n_1348)
);

AOI221x1_ASAP7_75t_L g1349 ( 
.A1(n_1210),
.A2(n_1102),
.B1(n_1119),
.B2(n_1168),
.C(n_1170),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1133),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_1206),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1216),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1163),
.A2(n_1147),
.B(n_1106),
.Y(n_1353)
);

AOI21xp33_ASAP7_75t_L g1354 ( 
.A1(n_1127),
.A2(n_1172),
.B(n_1106),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1201),
.A2(n_1119),
.B(n_1106),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1139),
.Y(n_1356)
);

OAI22xp5_ASAP7_75t_L g1357 ( 
.A1(n_1127),
.A2(n_1119),
.B1(n_1152),
.B2(n_1145),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1170),
.B(n_1188),
.Y(n_1358)
);

AOI21xp5_ASAP7_75t_SL g1359 ( 
.A1(n_1194),
.A2(n_1212),
.B(n_1197),
.Y(n_1359)
);

AND2x2_ASAP7_75t_L g1360 ( 
.A(n_1194),
.B(n_1212),
.Y(n_1360)
);

INVx2_ASAP7_75t_SL g1361 ( 
.A(n_1212),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1175),
.A2(n_990),
.B(n_714),
.Y(n_1362)
);

INVx2_ASAP7_75t_SL g1363 ( 
.A(n_1084),
.Y(n_1363)
);

AND2x4_ASAP7_75t_L g1364 ( 
.A(n_1176),
.B(n_948),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1219),
.B(n_744),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1175),
.A2(n_990),
.B(n_714),
.Y(n_1366)
);

OAI21x1_ASAP7_75t_L g1367 ( 
.A1(n_1154),
.A2(n_1138),
.B(n_1128),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1186),
.Y(n_1368)
);

OAI21xp33_ASAP7_75t_L g1369 ( 
.A1(n_1085),
.A2(n_992),
.B(n_1044),
.Y(n_1369)
);

OAI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1097),
.A2(n_1117),
.B(n_1175),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1219),
.B(n_915),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1118),
.Y(n_1372)
);

AO22x1_ASAP7_75t_L g1373 ( 
.A1(n_1121),
.A2(n_992),
.B1(n_918),
.B2(n_1044),
.Y(n_1373)
);

AOI21xp5_ASAP7_75t_L g1374 ( 
.A1(n_1175),
.A2(n_990),
.B(n_714),
.Y(n_1374)
);

AND2x4_ASAP7_75t_L g1375 ( 
.A(n_1176),
.B(n_948),
.Y(n_1375)
);

INVxp67_ASAP7_75t_L g1376 ( 
.A(n_1118),
.Y(n_1376)
);

INVx3_ASAP7_75t_L g1377 ( 
.A(n_1276),
.Y(n_1377)
);

BUFx2_ASAP7_75t_L g1378 ( 
.A(n_1231),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1230),
.Y(n_1380)
);

NOR2x2_ASAP7_75t_L g1381 ( 
.A(n_1242),
.B(n_1236),
.Y(n_1381)
);

INVx3_ASAP7_75t_L g1382 ( 
.A(n_1276),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1371),
.A2(n_1295),
.B1(n_1369),
.B2(n_1365),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1248),
.B(n_1373),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1247),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1274),
.Y(n_1386)
);

AND2x4_ASAP7_75t_L g1387 ( 
.A(n_1332),
.B(n_1242),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1309),
.Y(n_1388)
);

BUFx2_ASAP7_75t_L g1389 ( 
.A(n_1372),
.Y(n_1389)
);

INVx2_ASAP7_75t_L g1390 ( 
.A(n_1368),
.Y(n_1390)
);

INVx6_ASAP7_75t_L g1391 ( 
.A(n_1274),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1371),
.B(n_1257),
.Y(n_1392)
);

NAND2xp5_ASAP7_75t_L g1393 ( 
.A(n_1224),
.B(n_1222),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1228),
.Y(n_1394)
);

BUFx2_ASAP7_75t_L g1395 ( 
.A(n_1352),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1246),
.A2(n_1227),
.B(n_1362),
.Y(n_1396)
);

NAND2xp5_ASAP7_75t_L g1397 ( 
.A(n_1224),
.B(n_1279),
.Y(n_1397)
);

CKINVDCx20_ASAP7_75t_R g1398 ( 
.A(n_1235),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1238),
.Y(n_1399)
);

OAI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1251),
.A2(n_1259),
.B1(n_1234),
.B2(n_1291),
.Y(n_1400)
);

AOI221xp5_ASAP7_75t_L g1401 ( 
.A1(n_1300),
.A2(n_1253),
.B1(n_1272),
.B2(n_1343),
.C(n_1325),
.Y(n_1401)
);

A2O1A1Ixp33_ASAP7_75t_L g1402 ( 
.A1(n_1315),
.A2(n_1250),
.B(n_1328),
.C(n_1329),
.Y(n_1402)
);

AO21x2_ASAP7_75t_L g1403 ( 
.A1(n_1370),
.A2(n_1245),
.B(n_1312),
.Y(n_1403)
);

AO31x2_ASAP7_75t_L g1404 ( 
.A1(n_1349),
.A2(n_1260),
.A3(n_1252),
.B(n_1285),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1229),
.A2(n_1256),
.B(n_1370),
.Y(n_1405)
);

BUFx4f_ASAP7_75t_SL g1406 ( 
.A(n_1298),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1274),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1303),
.A2(n_1275),
.B(n_1290),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1226),
.A2(n_1273),
.B1(n_1255),
.B2(n_1242),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1232),
.A2(n_1269),
.B(n_1292),
.Y(n_1410)
);

AO31x2_ASAP7_75t_L g1411 ( 
.A1(n_1357),
.A2(n_1284),
.A3(n_1323),
.B(n_1254),
.Y(n_1411)
);

AOI22xp5_ASAP7_75t_L g1412 ( 
.A1(n_1287),
.A2(n_1239),
.B1(n_1237),
.B2(n_1278),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1289),
.Y(n_1413)
);

AO21x2_ASAP7_75t_L g1414 ( 
.A1(n_1324),
.A2(n_1282),
.B(n_1315),
.Y(n_1414)
);

NAND3xp33_ASAP7_75t_L g1415 ( 
.A(n_1322),
.B(n_1343),
.C(n_1317),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1304),
.Y(n_1416)
);

OAI21x1_ASAP7_75t_L g1417 ( 
.A1(n_1297),
.A2(n_1299),
.B(n_1345),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1318),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1320),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1270),
.B(n_1266),
.Y(n_1420)
);

OAI21xp5_ASAP7_75t_L g1421 ( 
.A1(n_1269),
.A2(n_1296),
.B(n_1263),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1273),
.A2(n_1376),
.B1(n_1225),
.B2(n_1279),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_SL g1423 ( 
.A1(n_1335),
.A2(n_1355),
.B1(n_1311),
.B2(n_1314),
.Y(n_1423)
);

OAI21x1_ASAP7_75t_L g1424 ( 
.A1(n_1353),
.A2(n_1330),
.B(n_1347),
.Y(n_1424)
);

OAI21x1_ASAP7_75t_L g1425 ( 
.A1(n_1284),
.A2(n_1341),
.B(n_1342),
.Y(n_1425)
);

BUFx6f_ASAP7_75t_L g1426 ( 
.A(n_1283),
.Y(n_1426)
);

O2A1O1Ixp33_ASAP7_75t_SL g1427 ( 
.A1(n_1336),
.A2(n_1340),
.B(n_1335),
.C(n_1328),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1316),
.B(n_1332),
.Y(n_1428)
);

AOI21xp5_ASAP7_75t_L g1429 ( 
.A1(n_1288),
.A2(n_1344),
.B(n_1233),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1331),
.Y(n_1430)
);

OAI21x1_ASAP7_75t_L g1431 ( 
.A1(n_1342),
.A2(n_1277),
.B(n_1329),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1277),
.A2(n_1346),
.B(n_1288),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1305),
.B(n_1364),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1249),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1339),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1262),
.Y(n_1436)
);

NOR2x1_ASAP7_75t_SL g1437 ( 
.A(n_1355),
.B(n_1357),
.Y(n_1437)
);

AOI21x1_ASAP7_75t_L g1438 ( 
.A1(n_1306),
.A2(n_1281),
.B(n_1280),
.Y(n_1438)
);

INVx2_ASAP7_75t_SL g1439 ( 
.A(n_1363),
.Y(n_1439)
);

AO21x1_ASAP7_75t_L g1440 ( 
.A1(n_1334),
.A2(n_1338),
.B(n_1270),
.Y(n_1440)
);

CKINVDCx20_ASAP7_75t_R g1441 ( 
.A(n_1310),
.Y(n_1441)
);

AOI21xp5_ASAP7_75t_L g1442 ( 
.A1(n_1244),
.A2(n_1301),
.B(n_1282),
.Y(n_1442)
);

OAI21xp5_ASAP7_75t_L g1443 ( 
.A1(n_1294),
.A2(n_1338),
.B(n_1307),
.Y(n_1443)
);

NAND2xp5_ASAP7_75t_L g1444 ( 
.A(n_1375),
.B(n_1264),
.Y(n_1444)
);

OAI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1308),
.A2(n_1334),
.B1(n_1293),
.B2(n_1264),
.Y(n_1445)
);

AOI21xp5_ASAP7_75t_L g1446 ( 
.A1(n_1321),
.A2(n_1337),
.B(n_1354),
.Y(n_1446)
);

OAI21xp5_ASAP7_75t_L g1447 ( 
.A1(n_1307),
.A2(n_1321),
.B(n_1354),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1375),
.B(n_1348),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1326),
.A2(n_1240),
.B(n_1327),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1243),
.A2(n_1326),
.B(n_1241),
.Y(n_1450)
);

AOI21xp33_ASAP7_75t_SL g1451 ( 
.A1(n_1286),
.A2(n_1361),
.B(n_1356),
.Y(n_1451)
);

OAI21x1_ASAP7_75t_L g1452 ( 
.A1(n_1241),
.A2(n_1358),
.B(n_1359),
.Y(n_1452)
);

AND2x4_ASAP7_75t_L g1453 ( 
.A(n_1360),
.B(n_1358),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1267),
.A2(n_1240),
.B(n_1293),
.Y(n_1454)
);

OA21x2_ASAP7_75t_L g1455 ( 
.A1(n_1240),
.A2(n_1293),
.B(n_1319),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1268),
.B(n_1261),
.Y(n_1456)
);

INVx2_ASAP7_75t_SL g1457 ( 
.A(n_1265),
.Y(n_1457)
);

INVx2_ASAP7_75t_SL g1458 ( 
.A(n_1351),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1302),
.B(n_1350),
.Y(n_1459)
);

OAI21x1_ASAP7_75t_L g1460 ( 
.A1(n_1319),
.A2(n_1313),
.B(n_1350),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_SL g1461 ( 
.A(n_1283),
.B(n_1333),
.Y(n_1461)
);

INVx3_ASAP7_75t_L g1462 ( 
.A(n_1283),
.Y(n_1462)
);

OAI21x1_ASAP7_75t_L g1463 ( 
.A1(n_1319),
.A2(n_1313),
.B(n_1333),
.Y(n_1463)
);

NAND2xp5_ASAP7_75t_L g1464 ( 
.A(n_1333),
.B(n_1248),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1230),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1369),
.A2(n_992),
.B(n_1044),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_L g1467 ( 
.A(n_1248),
.B(n_744),
.Y(n_1467)
);

OAI21x1_ASAP7_75t_L g1468 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_SL g1469 ( 
.A1(n_1315),
.A2(n_1336),
.B(n_1340),
.C(n_1322),
.Y(n_1469)
);

AO31x2_ASAP7_75t_L g1470 ( 
.A1(n_1349),
.A2(n_1260),
.A3(n_1252),
.B(n_1271),
.Y(n_1470)
);

AOI21xp5_ASAP7_75t_L g1471 ( 
.A1(n_1370),
.A2(n_1175),
.B(n_1250),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1230),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1248),
.B(n_744),
.Y(n_1474)
);

INVx2_ASAP7_75t_L g1475 ( 
.A(n_1230),
.Y(n_1475)
);

OAI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1476)
);

OAI21x1_ASAP7_75t_L g1477 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1477)
);

AND2x4_ASAP7_75t_L g1478 ( 
.A(n_1332),
.B(n_1242),
.Y(n_1478)
);

AOI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1369),
.A2(n_918),
.B1(n_992),
.B2(n_1044),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1369),
.A2(n_992),
.B(n_1044),
.Y(n_1480)
);

AOI221xp5_ASAP7_75t_L g1481 ( 
.A1(n_1369),
.A2(n_1020),
.B1(n_992),
.B2(n_785),
.C(n_1044),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1230),
.Y(n_1482)
);

OR2x2_ASAP7_75t_L g1483 ( 
.A(n_1222),
.B(n_1226),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1370),
.A2(n_1245),
.B(n_1271),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1230),
.Y(n_1485)
);

BUFx2_ASAP7_75t_SL g1486 ( 
.A(n_1310),
.Y(n_1486)
);

AO21x2_ASAP7_75t_L g1487 ( 
.A1(n_1370),
.A2(n_1245),
.B(n_1271),
.Y(n_1487)
);

CKINVDCx5p33_ASAP7_75t_R g1488 ( 
.A(n_1309),
.Y(n_1488)
);

AO21x2_ASAP7_75t_L g1489 ( 
.A1(n_1370),
.A2(n_1245),
.B(n_1271),
.Y(n_1489)
);

AOI21xp5_ASAP7_75t_L g1490 ( 
.A1(n_1370),
.A2(n_1175),
.B(n_1250),
.Y(n_1490)
);

CKINVDCx11_ASAP7_75t_R g1491 ( 
.A(n_1298),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1230),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1335),
.A2(n_401),
.B1(n_413),
.B2(n_404),
.Y(n_1493)
);

AOI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1362),
.A2(n_1374),
.B(n_1366),
.Y(n_1494)
);

INVx1_ASAP7_75t_L g1495 ( 
.A(n_1230),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1369),
.B(n_789),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1497)
);

NAND2x1p5_ASAP7_75t_L g1498 ( 
.A(n_1276),
.B(n_1218),
.Y(n_1498)
);

A2O1A1Ixp33_ASAP7_75t_L g1499 ( 
.A1(n_1369),
.A2(n_1036),
.B(n_1315),
.C(n_996),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1287),
.B(n_1237),
.Y(n_1500)
);

INVx1_ASAP7_75t_L g1501 ( 
.A(n_1230),
.Y(n_1501)
);

NOR2xp33_ASAP7_75t_SL g1502 ( 
.A(n_1249),
.B(n_791),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1230),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1287),
.B(n_1237),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1287),
.B(n_1237),
.Y(n_1505)
);

AOI21x1_ASAP7_75t_L g1506 ( 
.A1(n_1362),
.A2(n_1374),
.B(n_1366),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1248),
.B(n_744),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1230),
.Y(n_1508)
);

CKINVDCx14_ASAP7_75t_R g1509 ( 
.A(n_1235),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1276),
.B(n_1218),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1309),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_SL g1512 ( 
.A(n_1369),
.B(n_996),
.Y(n_1512)
);

OA21x2_ASAP7_75t_L g1513 ( 
.A1(n_1370),
.A2(n_1367),
.B(n_1260),
.Y(n_1513)
);

OAI21x1_ASAP7_75t_L g1514 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1514)
);

OAI21x1_ASAP7_75t_L g1515 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1248),
.B(n_744),
.Y(n_1516)
);

INVx1_ASAP7_75t_SL g1517 ( 
.A(n_1231),
.Y(n_1517)
);

AOI21xp5_ASAP7_75t_L g1518 ( 
.A1(n_1370),
.A2(n_1175),
.B(n_1250),
.Y(n_1518)
);

OAI21xp5_ASAP7_75t_L g1519 ( 
.A1(n_1369),
.A2(n_992),
.B(n_1044),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1230),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1230),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1370),
.A2(n_1367),
.B(n_1260),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1230),
.Y(n_1523)
);

INVx6_ASAP7_75t_L g1524 ( 
.A(n_1274),
.Y(n_1524)
);

OA21x2_ASAP7_75t_L g1525 ( 
.A1(n_1370),
.A2(n_1367),
.B(n_1260),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1230),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1230),
.Y(n_1527)
);

A2O1A1Ixp33_ASAP7_75t_L g1528 ( 
.A1(n_1369),
.A2(n_1036),
.B(n_1315),
.C(n_996),
.Y(n_1528)
);

OAI21xp5_ASAP7_75t_L g1529 ( 
.A1(n_1369),
.A2(n_992),
.B(n_1044),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1230),
.Y(n_1530)
);

AND2x4_ASAP7_75t_L g1531 ( 
.A(n_1332),
.B(n_1242),
.Y(n_1531)
);

OAI21x1_ASAP7_75t_L g1532 ( 
.A1(n_1223),
.A2(n_1367),
.B(n_1258),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1394),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1534)
);

BUFx12f_ASAP7_75t_L g1535 ( 
.A(n_1491),
.Y(n_1535)
);

O2A1O1Ixp5_ASAP7_75t_L g1536 ( 
.A1(n_1466),
.A2(n_1480),
.B(n_1529),
.C(n_1519),
.Y(n_1536)
);

AND2x2_ASAP7_75t_L g1537 ( 
.A(n_1453),
.B(n_1500),
.Y(n_1537)
);

AND2x4_ASAP7_75t_L g1538 ( 
.A(n_1387),
.B(n_1478),
.Y(n_1538)
);

OAI22xp5_ASAP7_75t_L g1539 ( 
.A1(n_1479),
.A2(n_1493),
.B1(n_1481),
.B2(n_1415),
.Y(n_1539)
);

AND2x2_ASAP7_75t_L g1540 ( 
.A(n_1453),
.B(n_1504),
.Y(n_1540)
);

O2A1O1Ixp33_ASAP7_75t_L g1541 ( 
.A1(n_1512),
.A2(n_1528),
.B(n_1499),
.C(n_1427),
.Y(n_1541)
);

O2A1O1Ixp33_ASAP7_75t_L g1542 ( 
.A1(n_1512),
.A2(n_1528),
.B(n_1499),
.C(n_1427),
.Y(n_1542)
);

HB1xp67_ASAP7_75t_L g1543 ( 
.A(n_1454),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1505),
.B(n_1428),
.Y(n_1544)
);

AND2x4_ASAP7_75t_L g1545 ( 
.A(n_1387),
.B(n_1478),
.Y(n_1545)
);

BUFx6f_ASAP7_75t_L g1546 ( 
.A(n_1426),
.Y(n_1546)
);

OA21x2_ASAP7_75t_L g1547 ( 
.A1(n_1421),
.A2(n_1431),
.B(n_1410),
.Y(n_1547)
);

O2A1O1Ixp5_ASAP7_75t_L g1548 ( 
.A1(n_1402),
.A2(n_1490),
.B(n_1471),
.C(n_1518),
.Y(n_1548)
);

INVx4_ASAP7_75t_L g1549 ( 
.A(n_1391),
.Y(n_1549)
);

INVx1_ASAP7_75t_SL g1550 ( 
.A(n_1517),
.Y(n_1550)
);

BUFx6f_ASAP7_75t_L g1551 ( 
.A(n_1426),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_L g1552 ( 
.A(n_1392),
.B(n_1467),
.Y(n_1552)
);

INVx1_ASAP7_75t_SL g1553 ( 
.A(n_1378),
.Y(n_1553)
);

OA21x2_ASAP7_75t_L g1554 ( 
.A1(n_1460),
.A2(n_1463),
.B(n_1402),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1403),
.Y(n_1555)
);

O2A1O1Ixp33_ASAP7_75t_L g1556 ( 
.A1(n_1469),
.A2(n_1496),
.B(n_1400),
.C(n_1383),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1483),
.B(n_1412),
.Y(n_1557)
);

BUFx3_ASAP7_75t_L g1558 ( 
.A(n_1391),
.Y(n_1558)
);

OAI22xp5_ASAP7_75t_L g1559 ( 
.A1(n_1493),
.A2(n_1507),
.B1(n_1516),
.B2(n_1474),
.Y(n_1559)
);

A2O1A1Ixp33_ASAP7_75t_L g1560 ( 
.A1(n_1496),
.A2(n_1401),
.B(n_1423),
.C(n_1442),
.Y(n_1560)
);

OAI22x1_ASAP7_75t_L g1561 ( 
.A1(n_1438),
.A2(n_1387),
.B1(n_1531),
.B2(n_1478),
.Y(n_1561)
);

HB1xp67_ASAP7_75t_L g1562 ( 
.A(n_1411),
.Y(n_1562)
);

INVx4_ASAP7_75t_L g1563 ( 
.A(n_1391),
.Y(n_1563)
);

OAI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1423),
.A2(n_1422),
.B1(n_1448),
.B2(n_1444),
.Y(n_1564)
);

AOI21xp5_ASAP7_75t_L g1565 ( 
.A1(n_1484),
.A2(n_1489),
.B(n_1487),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1420),
.B(n_1464),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_L g1567 ( 
.A1(n_1484),
.A2(n_1489),
.B(n_1487),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1409),
.A2(n_1389),
.B1(n_1395),
.B2(n_1445),
.Y(n_1568)
);

OR2x2_ASAP7_75t_L g1569 ( 
.A(n_1380),
.B(n_1385),
.Y(n_1569)
);

OA21x2_ASAP7_75t_L g1570 ( 
.A1(n_1425),
.A2(n_1396),
.B(n_1424),
.Y(n_1570)
);

INVx5_ASAP7_75t_L g1571 ( 
.A(n_1459),
.Y(n_1571)
);

AOI21xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1443),
.A2(n_1447),
.B(n_1459),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1390),
.B(n_1473),
.Y(n_1573)
);

AND2x2_ASAP7_75t_L g1574 ( 
.A(n_1390),
.B(n_1473),
.Y(n_1574)
);

AND2x4_ASAP7_75t_L g1575 ( 
.A(n_1459),
.B(n_1475),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1399),
.Y(n_1576)
);

AOI21xp5_ASAP7_75t_L g1577 ( 
.A1(n_1469),
.A2(n_1429),
.B(n_1414),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1411),
.Y(n_1578)
);

O2A1O1Ixp5_ASAP7_75t_L g1579 ( 
.A1(n_1445),
.A2(n_1440),
.B(n_1446),
.C(n_1494),
.Y(n_1579)
);

OAI22xp5_ASAP7_75t_L g1580 ( 
.A1(n_1456),
.A2(n_1451),
.B1(n_1458),
.B2(n_1439),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1386),
.A2(n_1407),
.B(n_1498),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1485),
.B(n_1492),
.Y(n_1582)
);

AOI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1502),
.A2(n_1441),
.B1(n_1486),
.B2(n_1398),
.Y(n_1583)
);

OR2x2_ASAP7_75t_L g1584 ( 
.A(n_1521),
.B(n_1530),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1411),
.Y(n_1585)
);

HB1xp67_ASAP7_75t_L g1586 ( 
.A(n_1432),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1521),
.B(n_1530),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1465),
.B(n_1482),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1436),
.B(n_1495),
.Y(n_1589)
);

BUFx6f_ASAP7_75t_L g1590 ( 
.A(n_1426),
.Y(n_1590)
);

AND2x2_ASAP7_75t_L g1591 ( 
.A(n_1501),
.B(n_1503),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1508),
.B(n_1520),
.Y(n_1592)
);

O2A1O1Ixp33_ASAP7_75t_L g1593 ( 
.A1(n_1416),
.A2(n_1419),
.B(n_1430),
.C(n_1418),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1523),
.B(n_1527),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1435),
.B(n_1413),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1526),
.B(n_1377),
.Y(n_1596)
);

HB1xp67_ASAP7_75t_L g1597 ( 
.A(n_1455),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1386),
.A2(n_1407),
.B(n_1498),
.Y(n_1598)
);

AND2x4_ASAP7_75t_L g1599 ( 
.A(n_1452),
.B(n_1377),
.Y(n_1599)
);

INVxp67_ASAP7_75t_SL g1600 ( 
.A(n_1455),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1455),
.Y(n_1601)
);

BUFx3_ASAP7_75t_L g1602 ( 
.A(n_1524),
.Y(n_1602)
);

A2O1A1Ixp33_ASAP7_75t_L g1603 ( 
.A1(n_1452),
.A2(n_1425),
.B(n_1404),
.C(n_1417),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1382),
.B(n_1461),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1470),
.B(n_1404),
.Y(n_1605)
);

OAI22xp5_ASAP7_75t_L g1606 ( 
.A1(n_1457),
.A2(n_1441),
.B1(n_1524),
.B2(n_1509),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1461),
.B(n_1462),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1437),
.B(n_1524),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1470),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1513),
.Y(n_1610)
);

AOI221x1_ASAP7_75t_SL g1611 ( 
.A1(n_1381),
.A2(n_1509),
.B1(n_1406),
.B2(n_1491),
.C(n_1398),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1510),
.B(n_1450),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1388),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1510),
.B(n_1449),
.Y(n_1614)
);

OAI22xp5_ASAP7_75t_L g1615 ( 
.A1(n_1406),
.A2(n_1434),
.B1(n_1388),
.B2(n_1488),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1449),
.B(n_1522),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1525),
.B(n_1434),
.Y(n_1617)
);

HB1xp67_ASAP7_75t_L g1618 ( 
.A(n_1525),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1408),
.B(n_1405),
.Y(n_1619)
);

OAI211xp5_ASAP7_75t_L g1620 ( 
.A1(n_1488),
.A2(n_1511),
.B(n_1506),
.C(n_1417),
.Y(n_1620)
);

AND2x4_ASAP7_75t_L g1621 ( 
.A(n_1379),
.B(n_1468),
.Y(n_1621)
);

INVx2_ASAP7_75t_L g1622 ( 
.A(n_1472),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1472),
.B(n_1476),
.Y(n_1623)
);

AOI21x1_ASAP7_75t_SL g1624 ( 
.A1(n_1477),
.A2(n_1497),
.B(n_1514),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1497),
.B(n_1532),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1514),
.A2(n_1515),
.B(n_1532),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1515),
.Y(n_1627)
);

AOI21x1_ASAP7_75t_SL g1628 ( 
.A1(n_1384),
.A2(n_1311),
.B(n_1314),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1629)
);

O2A1O1Ixp33_ASAP7_75t_L g1630 ( 
.A1(n_1466),
.A2(n_1480),
.B(n_1529),
.C(n_1519),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1631)
);

OA21x2_ASAP7_75t_L g1632 ( 
.A1(n_1421),
.A2(n_1431),
.B(n_1410),
.Y(n_1632)
);

AOI21x1_ASAP7_75t_SL g1633 ( 
.A1(n_1384),
.A2(n_1311),
.B(n_1314),
.Y(n_1633)
);

OAI22xp5_ASAP7_75t_L g1634 ( 
.A1(n_1479),
.A2(n_1493),
.B1(n_918),
.B2(n_1481),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1393),
.B(n_1397),
.Y(n_1636)
);

OA21x2_ASAP7_75t_L g1637 ( 
.A1(n_1421),
.A2(n_1431),
.B(n_1410),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1638)
);

CKINVDCx16_ASAP7_75t_R g1639 ( 
.A(n_1398),
.Y(n_1639)
);

AOI21x1_ASAP7_75t_SL g1640 ( 
.A1(n_1384),
.A2(n_1311),
.B(n_1314),
.Y(n_1640)
);

AND2x4_ASAP7_75t_L g1641 ( 
.A(n_1387),
.B(n_1478),
.Y(n_1641)
);

AND2x2_ASAP7_75t_L g1642 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1642)
);

AND2x4_ASAP7_75t_L g1643 ( 
.A(n_1387),
.B(n_1478),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1479),
.A2(n_1493),
.B1(n_918),
.B2(n_1481),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1471),
.A2(n_1518),
.B(n_1490),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1433),
.B(n_1453),
.Y(n_1648)
);

OAI22x1_ASAP7_75t_L g1649 ( 
.A1(n_1479),
.A2(n_1415),
.B1(n_1512),
.B2(n_1384),
.Y(n_1649)
);

OAI22xp5_ASAP7_75t_L g1650 ( 
.A1(n_1479),
.A2(n_1493),
.B1(n_918),
.B2(n_1481),
.Y(n_1650)
);

OAI31xp33_ASAP7_75t_SL g1651 ( 
.A1(n_1481),
.A2(n_1480),
.A3(n_1519),
.B(n_1466),
.Y(n_1651)
);

INVxp67_ASAP7_75t_L g1652 ( 
.A(n_1544),
.Y(n_1652)
);

AND2x2_ASAP7_75t_L g1653 ( 
.A(n_1617),
.B(n_1562),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1601),
.Y(n_1654)
);

OAI21xp5_ASAP7_75t_L g1655 ( 
.A1(n_1536),
.A2(n_1630),
.B(n_1634),
.Y(n_1655)
);

OR2x6_ASAP7_75t_L g1656 ( 
.A(n_1577),
.B(n_1572),
.Y(n_1656)
);

INVx2_ASAP7_75t_L g1657 ( 
.A(n_1533),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1636),
.B(n_1566),
.Y(n_1658)
);

NAND2xp5_ASAP7_75t_L g1659 ( 
.A(n_1552),
.B(n_1557),
.Y(n_1659)
);

OA21x2_ASAP7_75t_L g1660 ( 
.A1(n_1579),
.A2(n_1548),
.B(n_1647),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1624),
.A2(n_1567),
.B(n_1565),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1597),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1608),
.B(n_1599),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1578),
.B(n_1585),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1559),
.B(n_1651),
.Y(n_1665)
);

OA21x2_ASAP7_75t_L g1666 ( 
.A1(n_1579),
.A2(n_1548),
.B(n_1603),
.Y(n_1666)
);

NOR2xp67_ASAP7_75t_L g1667 ( 
.A(n_1571),
.B(n_1620),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1649),
.B(n_1537),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1595),
.Y(n_1669)
);

AND2x2_ASAP7_75t_L g1670 ( 
.A(n_1585),
.B(n_1540),
.Y(n_1670)
);

OAI21xp5_ASAP7_75t_L g1671 ( 
.A1(n_1536),
.A2(n_1650),
.B(n_1645),
.Y(n_1671)
);

OR2x6_ASAP7_75t_L g1672 ( 
.A(n_1561),
.B(n_1541),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1576),
.Y(n_1673)
);

AOI21xp5_ASAP7_75t_SL g1674 ( 
.A1(n_1556),
.A2(n_1542),
.B(n_1560),
.Y(n_1674)
);

INVx3_ASAP7_75t_L g1675 ( 
.A(n_1599),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1569),
.Y(n_1676)
);

INVx5_ASAP7_75t_L g1677 ( 
.A(n_1619),
.Y(n_1677)
);

NAND2xp5_ASAP7_75t_L g1678 ( 
.A(n_1573),
.B(n_1574),
.Y(n_1678)
);

AND2x4_ASAP7_75t_L g1679 ( 
.A(n_1599),
.B(n_1612),
.Y(n_1679)
);

OR2x6_ASAP7_75t_L g1680 ( 
.A(n_1581),
.B(n_1598),
.Y(n_1680)
);

AND2x4_ASAP7_75t_L g1681 ( 
.A(n_1538),
.B(n_1545),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1600),
.Y(n_1682)
);

AO21x2_ASAP7_75t_L g1683 ( 
.A1(n_1622),
.A2(n_1627),
.B(n_1609),
.Y(n_1683)
);

AOI21x1_ASAP7_75t_L g1684 ( 
.A1(n_1555),
.A2(n_1610),
.B(n_1618),
.Y(n_1684)
);

NAND2x1_ASAP7_75t_L g1685 ( 
.A(n_1619),
.B(n_1621),
.Y(n_1685)
);

HB1xp67_ASAP7_75t_L g1686 ( 
.A(n_1582),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1584),
.Y(n_1687)
);

INVxp33_ASAP7_75t_SL g1688 ( 
.A(n_1583),
.Y(n_1688)
);

INVx2_ASAP7_75t_L g1689 ( 
.A(n_1616),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1555),
.B(n_1547),
.Y(n_1690)
);

OAI21xp5_ASAP7_75t_L g1691 ( 
.A1(n_1539),
.A2(n_1564),
.B(n_1580),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1586),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1605),
.B(n_1547),
.Y(n_1693)
);

NAND4xp25_ASAP7_75t_L g1694 ( 
.A(n_1611),
.B(n_1593),
.C(n_1553),
.D(n_1550),
.Y(n_1694)
);

OR2x6_ASAP7_75t_L g1695 ( 
.A(n_1619),
.B(n_1554),
.Y(n_1695)
);

BUFx2_ASAP7_75t_L g1696 ( 
.A(n_1614),
.Y(n_1696)
);

AND2x2_ASAP7_75t_L g1697 ( 
.A(n_1547),
.B(n_1637),
.Y(n_1697)
);

BUFx2_ASAP7_75t_L g1698 ( 
.A(n_1543),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1543),
.Y(n_1699)
);

BUFx6f_ASAP7_75t_L g1700 ( 
.A(n_1571),
.Y(n_1700)
);

AO21x1_ASAP7_75t_SL g1701 ( 
.A1(n_1610),
.A2(n_1618),
.B(n_1604),
.Y(n_1701)
);

OR2x2_ASAP7_75t_L g1702 ( 
.A(n_1632),
.B(n_1637),
.Y(n_1702)
);

AO21x2_ASAP7_75t_L g1703 ( 
.A1(n_1623),
.A2(n_1625),
.B(n_1621),
.Y(n_1703)
);

BUFx2_ASAP7_75t_L g1704 ( 
.A(n_1632),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1554),
.B(n_1568),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1587),
.Y(n_1706)
);

NOR2xp33_ASAP7_75t_L g1707 ( 
.A(n_1534),
.B(n_1648),
.Y(n_1707)
);

AO21x2_ASAP7_75t_L g1708 ( 
.A1(n_1592),
.A2(n_1589),
.B(n_1596),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1570),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1709),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1708),
.B(n_1637),
.Y(n_1711)
);

INVx3_ASAP7_75t_L g1712 ( 
.A(n_1685),
.Y(n_1712)
);

INVx2_ASAP7_75t_SL g1713 ( 
.A(n_1677),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1708),
.B(n_1632),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1654),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1709),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1654),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1677),
.B(n_1675),
.Y(n_1718)
);

INVx1_ASAP7_75t_SL g1719 ( 
.A(n_1696),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1708),
.B(n_1594),
.Y(n_1720)
);

OR2x2_ASAP7_75t_L g1721 ( 
.A(n_1689),
.B(n_1570),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1683),
.Y(n_1722)
);

INVx2_ASAP7_75t_L g1723 ( 
.A(n_1683),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1689),
.B(n_1626),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1677),
.B(n_1641),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1683),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1703),
.B(n_1626),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1657),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1703),
.B(n_1626),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1693),
.B(n_1607),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1665),
.A2(n_1535),
.B1(n_1646),
.B2(n_1644),
.Y(n_1731)
);

AND2x2_ASAP7_75t_L g1732 ( 
.A(n_1703),
.B(n_1629),
.Y(n_1732)
);

INVxp67_ASAP7_75t_SL g1733 ( 
.A(n_1682),
.Y(n_1733)
);

AOI22xp33_ASAP7_75t_L g1734 ( 
.A1(n_1691),
.A2(n_1535),
.B1(n_1631),
.B2(n_1642),
.Y(n_1734)
);

NOR4xp25_ASAP7_75t_SL g1735 ( 
.A(n_1704),
.B(n_1633),
.C(n_1640),
.D(n_1628),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_L g1736 ( 
.A(n_1687),
.B(n_1588),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1662),
.Y(n_1737)
);

BUFx2_ASAP7_75t_L g1738 ( 
.A(n_1695),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1697),
.B(n_1690),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1671),
.A2(n_1635),
.B1(n_1638),
.B2(n_1606),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1697),
.B(n_1643),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1687),
.B(n_1591),
.Y(n_1742)
);

INVx1_ASAP7_75t_SL g1743 ( 
.A(n_1696),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1690),
.B(n_1643),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1695),
.Y(n_1745)
);

HB1xp67_ASAP7_75t_SL g1746 ( 
.A(n_1681),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1739),
.B(n_1679),
.Y(n_1747)
);

INVx2_ASAP7_75t_L g1748 ( 
.A(n_1710),
.Y(n_1748)
);

BUFx2_ASAP7_75t_L g1749 ( 
.A(n_1712),
.Y(n_1749)
);

HB1xp67_ASAP7_75t_L g1750 ( 
.A(n_1719),
.Y(n_1750)
);

OAI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1740),
.A2(n_1655),
.B1(n_1674),
.B2(n_1668),
.C(n_1694),
.Y(n_1751)
);

NOR2x1_ASAP7_75t_SL g1752 ( 
.A(n_1713),
.B(n_1701),
.Y(n_1752)
);

INVx2_ASAP7_75t_L g1753 ( 
.A(n_1710),
.Y(n_1753)
);

AND2x4_ASAP7_75t_L g1754 ( 
.A(n_1718),
.B(n_1679),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1737),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1730),
.B(n_1693),
.Y(n_1756)
);

OAI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1740),
.A2(n_1674),
.B1(n_1656),
.B2(n_1672),
.C(n_1659),
.Y(n_1757)
);

OR2x2_ASAP7_75t_L g1758 ( 
.A(n_1730),
.B(n_1739),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1730),
.B(n_1692),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1737),
.Y(n_1760)
);

BUFx2_ASAP7_75t_L g1761 ( 
.A(n_1712),
.Y(n_1761)
);

NOR4xp25_ASAP7_75t_SL g1762 ( 
.A(n_1738),
.B(n_1704),
.C(n_1698),
.D(n_1699),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1715),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1739),
.B(n_1653),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1711),
.A2(n_1714),
.B(n_1722),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1725),
.B(n_1681),
.Y(n_1766)
);

HB1xp67_ASAP7_75t_L g1767 ( 
.A(n_1719),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1715),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1736),
.B(n_1669),
.Y(n_1769)
);

INVxp67_ASAP7_75t_L g1770 ( 
.A(n_1736),
.Y(n_1770)
);

OAI211xp5_ASAP7_75t_SL g1771 ( 
.A1(n_1734),
.A2(n_1652),
.B(n_1658),
.C(n_1673),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1715),
.Y(n_1772)
);

OAI31xp33_ASAP7_75t_L g1773 ( 
.A1(n_1734),
.A2(n_1688),
.A3(n_1575),
.B(n_1545),
.Y(n_1773)
);

HB1xp67_ASAP7_75t_L g1774 ( 
.A(n_1743),
.Y(n_1774)
);

HB1xp67_ASAP7_75t_L g1775 ( 
.A(n_1743),
.Y(n_1775)
);

AOI221xp5_ASAP7_75t_L g1776 ( 
.A1(n_1720),
.A2(n_1688),
.B1(n_1707),
.B2(n_1706),
.C(n_1653),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1732),
.B(n_1663),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1710),
.Y(n_1778)
);

AOI21xp5_ASAP7_75t_L g1779 ( 
.A1(n_1735),
.A2(n_1656),
.B(n_1680),
.Y(n_1779)
);

OR2x6_ASAP7_75t_L g1780 ( 
.A(n_1713),
.B(n_1656),
.Y(n_1780)
);

AO21x2_ASAP7_75t_L g1781 ( 
.A1(n_1722),
.A2(n_1684),
.B(n_1661),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1742),
.B(n_1676),
.Y(n_1782)
);

OAI211xp5_ASAP7_75t_SL g1783 ( 
.A1(n_1731),
.A2(n_1706),
.B(n_1613),
.C(n_1678),
.Y(n_1783)
);

OAI221xp5_ASAP7_75t_L g1784 ( 
.A1(n_1731),
.A2(n_1672),
.B1(n_1667),
.B2(n_1680),
.C(n_1705),
.Y(n_1784)
);

OAI211xp5_ASAP7_75t_L g1785 ( 
.A1(n_1735),
.A2(n_1666),
.B(n_1660),
.C(n_1702),
.Y(n_1785)
);

INVxp67_ASAP7_75t_SL g1786 ( 
.A(n_1720),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1732),
.B(n_1663),
.Y(n_1787)
);

OR2x6_ASAP7_75t_L g1788 ( 
.A(n_1713),
.B(n_1680),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1717),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1746),
.A2(n_1672),
.B1(n_1680),
.B2(n_1571),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1742),
.B(n_1686),
.Y(n_1791)
);

INVx2_ASAP7_75t_SL g1792 ( 
.A(n_1712),
.Y(n_1792)
);

AOI222xp33_ASAP7_75t_L g1793 ( 
.A1(n_1732),
.A2(n_1633),
.B1(n_1640),
.B2(n_1628),
.C1(n_1670),
.C2(n_1664),
.Y(n_1793)
);

INVx2_ASAP7_75t_L g1794 ( 
.A(n_1716),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1721),
.B(n_1692),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1721),
.B(n_1728),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1741),
.B(n_1663),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1738),
.A2(n_1672),
.B1(n_1705),
.B2(n_1666),
.C(n_1660),
.Y(n_1798)
);

INVx2_ASAP7_75t_L g1799 ( 
.A(n_1748),
.Y(n_1799)
);

HB1xp67_ASAP7_75t_L g1800 ( 
.A(n_1763),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1763),
.Y(n_1801)
);

NOR2xp33_ASAP7_75t_L g1802 ( 
.A(n_1751),
.B(n_1639),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1768),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1777),
.B(n_1738),
.Y(n_1804)
);

HB1xp67_ASAP7_75t_L g1805 ( 
.A(n_1768),
.Y(n_1805)
);

INVx2_ASAP7_75t_L g1806 ( 
.A(n_1753),
.Y(n_1806)
);

AND2x2_ASAP7_75t_L g1807 ( 
.A(n_1777),
.B(n_1745),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1786),
.B(n_1724),
.Y(n_1808)
);

INVx2_ASAP7_75t_L g1809 ( 
.A(n_1753),
.Y(n_1809)
);

NOR2x1p5_ASAP7_75t_L g1810 ( 
.A(n_1754),
.B(n_1745),
.Y(n_1810)
);

NAND2xp5_ASAP7_75t_L g1811 ( 
.A(n_1755),
.B(n_1724),
.Y(n_1811)
);

NAND2x1_ASAP7_75t_L g1812 ( 
.A(n_1749),
.B(n_1712),
.Y(n_1812)
);

INVx2_ASAP7_75t_L g1813 ( 
.A(n_1778),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1772),
.Y(n_1814)
);

INVx2_ASAP7_75t_L g1815 ( 
.A(n_1794),
.Y(n_1815)
);

INVx1_ASAP7_75t_L g1816 ( 
.A(n_1789),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1755),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1750),
.Y(n_1818)
);

INVxp67_ASAP7_75t_SL g1819 ( 
.A(n_1765),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1796),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1760),
.Y(n_1821)
);

INVx2_ASAP7_75t_SL g1822 ( 
.A(n_1749),
.Y(n_1822)
);

INVx1_ASAP7_75t_SL g1823 ( 
.A(n_1767),
.Y(n_1823)
);

HB1xp67_ASAP7_75t_L g1824 ( 
.A(n_1760),
.Y(n_1824)
);

NOR2x1p5_ASAP7_75t_L g1825 ( 
.A(n_1754),
.B(n_1745),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1796),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1781),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1759),
.Y(n_1828)
);

NAND3xp33_ASAP7_75t_SL g1829 ( 
.A(n_1762),
.B(n_1714),
.C(n_1729),
.Y(n_1829)
);

INVx4_ASAP7_75t_SL g1830 ( 
.A(n_1788),
.Y(n_1830)
);

OA21x2_ASAP7_75t_L g1831 ( 
.A1(n_1785),
.A2(n_1723),
.B(n_1722),
.Y(n_1831)
);

OA21x2_ASAP7_75t_L g1832 ( 
.A1(n_1798),
.A2(n_1726),
.B(n_1723),
.Y(n_1832)
);

AOI21x1_ASAP7_75t_L g1833 ( 
.A1(n_1779),
.A2(n_1729),
.B(n_1727),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1759),
.Y(n_1834)
);

INVx1_ASAP7_75t_SL g1835 ( 
.A(n_1774),
.Y(n_1835)
);

OR2x2_ASAP7_75t_L g1836 ( 
.A(n_1828),
.B(n_1756),
.Y(n_1836)
);

OR2x2_ASAP7_75t_L g1837 ( 
.A(n_1828),
.B(n_1756),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1814),
.Y(n_1838)
);

NAND4xp25_ASAP7_75t_SL g1839 ( 
.A(n_1818),
.B(n_1776),
.C(n_1793),
.D(n_1784),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1818),
.B(n_1770),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1823),
.B(n_1835),
.Y(n_1841)
);

AND2x2_ASAP7_75t_L g1842 ( 
.A(n_1810),
.B(n_1754),
.Y(n_1842)
);

NOR2xp33_ASAP7_75t_L g1843 ( 
.A(n_1802),
.B(n_1615),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1810),
.B(n_1787),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1825),
.B(n_1787),
.Y(n_1845)
);

OR2x2_ASAP7_75t_L g1846 ( 
.A(n_1834),
.B(n_1823),
.Y(n_1846)
);

AOI221xp5_ASAP7_75t_L g1847 ( 
.A1(n_1829),
.A2(n_1802),
.B1(n_1757),
.B2(n_1819),
.C(n_1835),
.Y(n_1847)
);

INVxp67_ASAP7_75t_L g1848 ( 
.A(n_1824),
.Y(n_1848)
);

NAND3xp33_ASAP7_75t_L g1849 ( 
.A(n_1832),
.B(n_1771),
.C(n_1783),
.Y(n_1849)
);

NOR2xp67_ASAP7_75t_L g1850 ( 
.A(n_1822),
.B(n_1766),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1800),
.Y(n_1851)
);

AND2x2_ASAP7_75t_L g1852 ( 
.A(n_1825),
.B(n_1804),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1814),
.Y(n_1853)
);

NAND4xp25_ASAP7_75t_L g1854 ( 
.A(n_1829),
.B(n_1773),
.C(n_1790),
.D(n_1769),
.Y(n_1854)
);

INVx2_ASAP7_75t_L g1855 ( 
.A(n_1822),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1834),
.B(n_1775),
.Y(n_1856)
);

OR2x2_ASAP7_75t_L g1857 ( 
.A(n_1811),
.B(n_1758),
.Y(n_1857)
);

NAND2xp5_ASAP7_75t_L g1858 ( 
.A(n_1808),
.B(n_1747),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1816),
.Y(n_1859)
);

AND2x2_ASAP7_75t_L g1860 ( 
.A(n_1804),
.B(n_1752),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1808),
.B(n_1747),
.Y(n_1861)
);

INVx2_ASAP7_75t_L g1862 ( 
.A(n_1822),
.Y(n_1862)
);

HB1xp67_ASAP7_75t_L g1863 ( 
.A(n_1824),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1804),
.B(n_1758),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1830),
.B(n_1752),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1800),
.Y(n_1866)
);

OR2x2_ASAP7_75t_L g1867 ( 
.A(n_1811),
.B(n_1795),
.Y(n_1867)
);

INVx1_ASAP7_75t_SL g1868 ( 
.A(n_1830),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1816),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1820),
.B(n_1764),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1817),
.B(n_1795),
.Y(n_1871)
);

AOI322xp5_ASAP7_75t_L g1872 ( 
.A1(n_1819),
.A2(n_1764),
.A3(n_1729),
.B1(n_1727),
.B2(n_1733),
.C1(n_1791),
.C2(n_1782),
.Y(n_1872)
);

NAND4xp25_ASAP7_75t_L g1873 ( 
.A(n_1817),
.B(n_1699),
.C(n_1745),
.D(n_1702),
.Y(n_1873)
);

NOR2xp33_ASAP7_75t_L g1874 ( 
.A(n_1807),
.B(n_1797),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1830),
.Y(n_1875)
);

NOR2x1_ASAP7_75t_L g1876 ( 
.A(n_1812),
.B(n_1761),
.Y(n_1876)
);

AND2x2_ASAP7_75t_L g1877 ( 
.A(n_1830),
.B(n_1807),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1820),
.B(n_1797),
.Y(n_1878)
);

INVxp67_ASAP7_75t_L g1879 ( 
.A(n_1821),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1805),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1830),
.B(n_1761),
.Y(n_1881)
);

A2O1A1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1847),
.A2(n_1812),
.B(n_1745),
.C(n_1727),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1841),
.B(n_1821),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1866),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1840),
.B(n_1820),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1863),
.Y(n_1886)
);

NAND2xp5_ASAP7_75t_L g1887 ( 
.A(n_1872),
.B(n_1820),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1838),
.Y(n_1888)
);

OR2x2_ASAP7_75t_L g1889 ( 
.A(n_1846),
.B(n_1826),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1853),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1859),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_SL g1892 ( 
.A(n_1875),
.B(n_1868),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1846),
.B(n_1826),
.Y(n_1893)
);

INVx2_ASAP7_75t_L g1894 ( 
.A(n_1855),
.Y(n_1894)
);

INVx1_ASAP7_75t_SL g1895 ( 
.A(n_1875),
.Y(n_1895)
);

NOR2xp67_ASAP7_75t_SL g1896 ( 
.A(n_1849),
.B(n_1700),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1843),
.B(n_1874),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1878),
.B(n_1826),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1855),
.Y(n_1899)
);

INVx2_ASAP7_75t_SL g1900 ( 
.A(n_1876),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1869),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1858),
.B(n_1826),
.Y(n_1902)
);

OR2x2_ASAP7_75t_L g1903 ( 
.A(n_1864),
.B(n_1801),
.Y(n_1903)
);

OR2x2_ASAP7_75t_L g1904 ( 
.A(n_1870),
.B(n_1801),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1860),
.B(n_1830),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1860),
.B(n_1807),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1877),
.Y(n_1907)
);

NAND2xp5_ASAP7_75t_L g1908 ( 
.A(n_1861),
.B(n_1856),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1880),
.Y(n_1909)
);

AND2x2_ASAP7_75t_L g1910 ( 
.A(n_1865),
.B(n_1805),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1848),
.B(n_1744),
.Y(n_1911)
);

INVx1_ASAP7_75t_L g1912 ( 
.A(n_1851),
.Y(n_1912)
);

INVx1_ASAP7_75t_L g1913 ( 
.A(n_1851),
.Y(n_1913)
);

AOI21xp33_ASAP7_75t_SL g1914 ( 
.A1(n_1865),
.A2(n_1832),
.B(n_1788),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1879),
.B(n_1744),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1871),
.Y(n_1916)
);

NOR2x1_ASAP7_75t_L g1917 ( 
.A(n_1850),
.B(n_1803),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1852),
.B(n_1833),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1912),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1905),
.B(n_1917),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1906),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1913),
.Y(n_1922)
);

OR2x2_ASAP7_75t_L g1923 ( 
.A(n_1889),
.B(n_1836),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1884),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1905),
.B(n_1852),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1907),
.B(n_1844),
.Y(n_1926)
);

INVx1_ASAP7_75t_L g1927 ( 
.A(n_1884),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_L g1928 ( 
.A(n_1895),
.B(n_1844),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1888),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1886),
.B(n_1845),
.Y(n_1930)
);

AND2x4_ASAP7_75t_L g1931 ( 
.A(n_1900),
.B(n_1842),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1890),
.Y(n_1932)
);

AND2x4_ASAP7_75t_L g1933 ( 
.A(n_1900),
.B(n_1842),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1909),
.B(n_1845),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1906),
.Y(n_1935)
);

AOI22xp5_ASAP7_75t_L g1936 ( 
.A1(n_1896),
.A2(n_1839),
.B1(n_1854),
.B2(n_1877),
.Y(n_1936)
);

HB1xp67_ASAP7_75t_L g1937 ( 
.A(n_1894),
.Y(n_1937)
);

OR2x2_ASAP7_75t_L g1938 ( 
.A(n_1889),
.B(n_1836),
.Y(n_1938)
);

INVx1_ASAP7_75t_SL g1939 ( 
.A(n_1892),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1896),
.B(n_1862),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1891),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1910),
.B(n_1881),
.Y(n_1942)
);

INVx1_ASAP7_75t_L g1943 ( 
.A(n_1901),
.Y(n_1943)
);

INVx1_ASAP7_75t_L g1944 ( 
.A(n_1916),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1910),
.B(n_1881),
.Y(n_1945)
);

O2A1O1Ixp33_ASAP7_75t_L g1946 ( 
.A1(n_1939),
.A2(n_1882),
.B(n_1887),
.C(n_1897),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1926),
.B(n_1908),
.Y(n_1947)
);

OAI21xp5_ASAP7_75t_SL g1948 ( 
.A1(n_1936),
.A2(n_1882),
.B(n_1914),
.Y(n_1948)
);

NOR2xp33_ASAP7_75t_L g1949 ( 
.A(n_1930),
.B(n_1883),
.Y(n_1949)
);

INVxp67_ASAP7_75t_L g1950 ( 
.A(n_1920),
.Y(n_1950)
);

AOI222xp33_ASAP7_75t_L g1951 ( 
.A1(n_1924),
.A2(n_1918),
.B1(n_1885),
.B2(n_1893),
.C1(n_1898),
.C2(n_1902),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_L g1952 ( 
.A(n_1926),
.B(n_1894),
.Y(n_1952)
);

AOI21xp5_ASAP7_75t_L g1953 ( 
.A1(n_1940),
.A2(n_1918),
.B(n_1899),
.Y(n_1953)
);

NAND2x1p5_ASAP7_75t_L g1954 ( 
.A(n_1920),
.B(n_1899),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1937),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1924),
.Y(n_1956)
);

AOI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1928),
.A2(n_1862),
.B(n_1911),
.Y(n_1957)
);

OAI31xp33_ASAP7_75t_L g1958 ( 
.A1(n_1925),
.A2(n_1873),
.A3(n_1903),
.B(n_1904),
.Y(n_1958)
);

O2A1O1Ixp33_ASAP7_75t_L g1959 ( 
.A1(n_1927),
.A2(n_1903),
.B(n_1904),
.C(n_1915),
.Y(n_1959)
);

AOI22xp5_ASAP7_75t_L g1960 ( 
.A1(n_1925),
.A2(n_1788),
.B1(n_1832),
.B2(n_1780),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1927),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1934),
.A2(n_1833),
.B(n_1832),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_L g1963 ( 
.A(n_1945),
.B(n_1942),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1945),
.B(n_1837),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1923),
.Y(n_1965)
);

INVx1_ASAP7_75t_L g1966 ( 
.A(n_1923),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1950),
.B(n_1942),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1965),
.B(n_1944),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1966),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1954),
.Y(n_1970)
);

INVx1_ASAP7_75t_SL g1971 ( 
.A(n_1963),
.Y(n_1971)
);

XNOR2xp5_ASAP7_75t_L g1972 ( 
.A(n_1947),
.B(n_1931),
.Y(n_1972)
);

OR2x2_ASAP7_75t_L g1973 ( 
.A(n_1964),
.B(n_1938),
.Y(n_1973)
);

OAI221xp5_ASAP7_75t_L g1974 ( 
.A1(n_1948),
.A2(n_1944),
.B1(n_1921),
.B2(n_1935),
.C(n_1938),
.Y(n_1974)
);

INVx2_ASAP7_75t_SL g1975 ( 
.A(n_1954),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1952),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_L g1977 ( 
.A(n_1955),
.B(n_1921),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1953),
.B(n_1931),
.Y(n_1978)
);

AND2x2_ASAP7_75t_L g1979 ( 
.A(n_1949),
.B(n_1931),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_L g1980 ( 
.A1(n_1974),
.A2(n_1946),
.B(n_1959),
.Y(n_1980)
);

NAND4xp25_ASAP7_75t_L g1981 ( 
.A(n_1971),
.B(n_1958),
.C(n_1951),
.D(n_1957),
.Y(n_1981)
);

OAI21xp33_ASAP7_75t_L g1982 ( 
.A1(n_1972),
.A2(n_1935),
.B(n_1933),
.Y(n_1982)
);

O2A1O1Ixp5_ASAP7_75t_L g1983 ( 
.A1(n_1970),
.A2(n_1962),
.B(n_1933),
.C(n_1922),
.Y(n_1983)
);

OAI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1973),
.A2(n_1960),
.B1(n_1932),
.B2(n_1943),
.C(n_1941),
.Y(n_1984)
);

AOI211xp5_ASAP7_75t_L g1985 ( 
.A1(n_1978),
.A2(n_1961),
.B(n_1956),
.C(n_1919),
.Y(n_1985)
);

AOI21xp5_ASAP7_75t_L g1986 ( 
.A1(n_1975),
.A2(n_1933),
.B(n_1929),
.Y(n_1986)
);

AOI221xp5_ASAP7_75t_L g1987 ( 
.A1(n_1978),
.A2(n_1929),
.B1(n_1827),
.B2(n_1837),
.C(n_1857),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1967),
.B(n_1979),
.Y(n_1988)
);

AOI21xp5_ASAP7_75t_L g1989 ( 
.A1(n_1975),
.A2(n_1827),
.B(n_1832),
.Y(n_1989)
);

INVx2_ASAP7_75t_L g1990 ( 
.A(n_1988),
.Y(n_1990)
);

INVx1_ASAP7_75t_L g1991 ( 
.A(n_1982),
.Y(n_1991)
);

AOI22xp5_ASAP7_75t_L g1992 ( 
.A1(n_1981),
.A2(n_1979),
.B1(n_1967),
.B2(n_1976),
.Y(n_1992)
);

OAI21xp33_ASAP7_75t_L g1993 ( 
.A1(n_1980),
.A2(n_1973),
.B(n_1977),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1986),
.Y(n_1994)
);

HB1xp67_ASAP7_75t_L g1995 ( 
.A(n_1985),
.Y(n_1995)
);

INVx2_ASAP7_75t_SL g1996 ( 
.A(n_1994),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1993),
.B(n_1969),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_L g1998 ( 
.A(n_1992),
.B(n_1968),
.Y(n_1998)
);

INVx1_ASAP7_75t_L g1999 ( 
.A(n_1990),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1995),
.Y(n_2000)
);

INVx2_ASAP7_75t_SL g2001 ( 
.A(n_1991),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1995),
.B(n_1983),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_2001),
.Y(n_2003)
);

OAI22xp33_ASAP7_75t_L g2004 ( 
.A1(n_2000),
.A2(n_1984),
.B1(n_1987),
.B2(n_1989),
.Y(n_2004)
);

INVx1_ASAP7_75t_L g2005 ( 
.A(n_1996),
.Y(n_2005)
);

NAND4xp25_ASAP7_75t_SL g2006 ( 
.A(n_2000),
.B(n_1827),
.C(n_1857),
.D(n_1867),
.Y(n_2006)
);

NAND3xp33_ASAP7_75t_L g2007 ( 
.A(n_2002),
.B(n_1832),
.C(n_1827),
.Y(n_2007)
);

BUFx2_ASAP7_75t_L g2008 ( 
.A(n_2003),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_2005),
.Y(n_2009)
);

NOR4xp25_ASAP7_75t_L g2010 ( 
.A(n_2004),
.B(n_1998),
.C(n_1999),
.D(n_1997),
.Y(n_2010)
);

NOR3xp33_ASAP7_75t_SL g2011 ( 
.A(n_2010),
.B(n_2006),
.C(n_2007),
.Y(n_2011)
);

AOI22xp33_ASAP7_75t_L g2012 ( 
.A1(n_2011),
.A2(n_2008),
.B1(n_2009),
.B2(n_1831),
.Y(n_2012)
);

AO21x2_ASAP7_75t_L g2013 ( 
.A1(n_2012),
.A2(n_1833),
.B(n_1799),
.Y(n_2013)
);

NAND4xp75_ASAP7_75t_L g2014 ( 
.A(n_2012),
.B(n_1831),
.C(n_1792),
.D(n_1765),
.Y(n_2014)
);

AO22x2_ASAP7_75t_L g2015 ( 
.A1(n_2014),
.A2(n_1809),
.B1(n_1799),
.B2(n_1815),
.Y(n_2015)
);

INVxp67_ASAP7_75t_L g2016 ( 
.A(n_2013),
.Y(n_2016)
);

OAI22xp5_ASAP7_75t_SL g2017 ( 
.A1(n_2016),
.A2(n_1563),
.B1(n_1549),
.B2(n_1602),
.Y(n_2017)
);

XNOR2xp5_ASAP7_75t_L g2018 ( 
.A(n_2015),
.B(n_1558),
.Y(n_2018)
);

OAI221xp5_ASAP7_75t_L g2019 ( 
.A1(n_2018),
.A2(n_1871),
.B1(n_1867),
.B2(n_1563),
.C(n_1549),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_2019),
.B(n_2017),
.Y(n_2020)
);

AO22x2_ASAP7_75t_L g2021 ( 
.A1(n_2020),
.A2(n_1809),
.B1(n_1815),
.B2(n_1806),
.Y(n_2021)
);

OAI21xp5_ASAP7_75t_L g2022 ( 
.A1(n_2021),
.A2(n_1813),
.B(n_1799),
.Y(n_2022)
);

OAI221xp5_ASAP7_75t_L g2023 ( 
.A1(n_2022),
.A2(n_1602),
.B1(n_1558),
.B2(n_1809),
.C(n_1799),
.Y(n_2023)
);

AOI211xp5_ASAP7_75t_L g2024 ( 
.A1(n_2023),
.A2(n_1590),
.B(n_1546),
.C(n_1551),
.Y(n_2024)
);


endmodule