module fake_jpeg_12798_n_429 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_429);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_429;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_0),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_3),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_17),
.Y(n_42)
);

BUFx6f_ASAP7_75t_SL g43 ( 
.A(n_17),
.Y(n_43)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_44),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_45),
.Y(n_107)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_46),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_48),
.Y(n_103)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_23),
.Y(n_49)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_19),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_51),
.Y(n_96)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_31),
.Y(n_52)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_53),
.B(n_1),
.Y(n_134)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_54),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g55 ( 
.A(n_31),
.B(n_16),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_55),
.B(n_62),
.Y(n_125)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_25),
.Y(n_57)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_57),
.Y(n_108)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_58),
.Y(n_97)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_59),
.Y(n_89)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_61),
.Y(n_124)
);

HAxp5_ASAP7_75t_SL g62 ( 
.A(n_41),
.B(n_0),
.CON(n_62),
.SN(n_62)
);

BUFx12_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_63),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_21),
.Y(n_65)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_65),
.Y(n_119)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_66),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_21),
.Y(n_68)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g69 ( 
.A1(n_43),
.A2(n_16),
.B(n_15),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_69),
.B(n_80),
.Y(n_102)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_16),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_86),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_29),
.Y(n_73)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_74),
.Y(n_116)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_35),
.Y(n_75)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx4_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_37),
.Y(n_77)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx4_ASAP7_75t_SL g78 ( 
.A(n_41),
.Y(n_78)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_78),
.Y(n_115)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_37),
.Y(n_79)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_79),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_42),
.B(n_15),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_84),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_82),
.Y(n_122)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_83),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g84 ( 
.A(n_18),
.B(n_0),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_85),
.Y(n_132)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_23),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_87),
.A2(n_61),
.B1(n_83),
.B2(n_71),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_91),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_18),
.B1(n_38),
.B2(n_40),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_93),
.A2(n_99),
.B1(n_104),
.B2(n_111),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_62),
.A2(n_20),
.B1(n_39),
.B2(n_24),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_53),
.A2(n_40),
.B1(n_38),
.B2(n_32),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_45),
.A2(n_57),
.B1(n_54),
.B2(n_47),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_65),
.A2(n_39),
.B1(n_22),
.B2(n_34),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_117),
.A2(n_121),
.B1(n_131),
.B2(n_28),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_67),
.A2(n_30),
.B1(n_36),
.B2(n_26),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_68),
.A2(n_30),
.B1(n_36),
.B2(n_26),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_78),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_117),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_142),
.Y(n_180)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_113),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_136),
.Y(n_193)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_101),
.Y(n_137)
);

HB1xp67_ASAP7_75t_L g199 ( 
.A(n_137),
.Y(n_199)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_138),
.Y(n_177)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_140),
.Y(n_194)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_113),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_143),
.B(n_145),
.Y(n_183)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_95),
.Y(n_145)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_146),
.B(n_147),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_130),
.B(n_64),
.Y(n_147)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_123),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_148),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_97),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

INVx3_ASAP7_75t_L g150 ( 
.A(n_133),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g151 ( 
.A(n_115),
.Y(n_151)
);

OAI31xp33_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_172),
.A3(n_30),
.B(n_32),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_152),
.A2(n_158),
.B1(n_161),
.B2(n_173),
.Y(n_202)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_118),
.Y(n_153)
);

NAND2xp33_ASAP7_75t_SL g200 ( 
.A(n_153),
.B(n_155),
.Y(n_200)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_132),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_154),
.B(n_156),
.Y(n_175)
);

INVx1_ASAP7_75t_SL g155 ( 
.A(n_112),
.Y(n_155)
);

BUFx2_ASAP7_75t_L g156 ( 
.A(n_89),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_157),
.B(n_165),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_102),
.A2(n_82),
.B1(n_77),
.B2(n_73),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_125),
.A2(n_24),
.B(n_39),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g197 ( 
.A1(n_159),
.A2(n_171),
.B(n_28),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_162),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_106),
.A2(n_44),
.B1(n_85),
.B2(n_59),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_90),
.Y(n_162)
);

BUFx2_ASAP7_75t_L g163 ( 
.A(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_163),
.B(n_164),
.Y(n_201)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_91),
.Y(n_165)
);

INVx1_ASAP7_75t_SL g166 ( 
.A(n_96),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_166),
.B(n_167),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_125),
.B(n_36),
.Y(n_167)
);

INVx6_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_168),
.B(n_170),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_105),
.B(n_50),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_96),
.C(n_120),
.Y(n_178)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g171 ( 
.A1(n_99),
.A2(n_22),
.B(n_24),
.Y(n_171)
);

INVx11_ASAP7_75t_L g172 ( 
.A(n_103),
.Y(n_172)
);

AO22x1_ASAP7_75t_L g188 ( 
.A1(n_172),
.A2(n_98),
.B1(n_126),
.B2(n_116),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_111),
.A2(n_32),
.B1(n_26),
.B2(n_28),
.Y(n_173)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_179),
.Y(n_206)
);

AND2x4_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_100),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_144),
.A2(n_108),
.B1(n_114),
.B2(n_110),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_168),
.B1(n_156),
.B2(n_110),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_167),
.B(n_34),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_182),
.B(n_186),
.C(n_169),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_139),
.B(n_127),
.C(n_88),
.Y(n_186)
);

BUFx8_ASAP7_75t_L g221 ( 
.A(n_188),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_173),
.A2(n_108),
.B1(n_126),
.B2(n_116),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_166),
.B1(n_155),
.B2(n_162),
.Y(n_215)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_144),
.A2(n_50),
.A3(n_128),
.B1(n_109),
.B2(n_98),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_190),
.B(n_158),
.Y(n_203)
);

CKINVDCx14_ASAP7_75t_R g228 ( 
.A(n_195),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_197),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_203),
.A2(n_213),
.B1(n_220),
.B2(n_179),
.Y(n_236)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_200),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_204),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_191),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_216),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_207),
.A2(n_180),
.B1(n_198),
.B2(n_193),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_179),
.B(n_169),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_208),
.B(n_215),
.Y(n_238)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_209),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_190),
.A2(n_152),
.B1(n_138),
.B2(n_143),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_210),
.A2(n_222),
.B(n_200),
.Y(n_249)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_201),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_226),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_202),
.A2(n_171),
.B1(n_94),
.B2(n_92),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_SL g214 ( 
.A(n_182),
.B(n_151),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_214),
.B(n_192),
.Y(n_232)
);

NAND3xp33_ASAP7_75t_L g216 ( 
.A(n_174),
.B(n_159),
.C(n_164),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_140),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_218),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_185),
.B(n_182),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_202),
.A2(n_107),
.B1(n_114),
.B2(n_92),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g222 ( 
.A1(n_201),
.A2(n_100),
.B1(n_137),
.B2(n_141),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_177),
.Y(n_224)
);

INVx5_ASAP7_75t_L g233 ( 
.A(n_224),
.Y(n_233)
);

XNOR2x1_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_186),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g226 ( 
.A(n_174),
.B(n_163),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_196),
.B(n_148),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_227),
.B(n_183),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_229),
.B(n_184),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_214),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_211),
.A2(n_197),
.B(n_180),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_235),
.A2(n_216),
.B(n_247),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_236),
.A2(n_221),
.B1(n_215),
.B2(n_187),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_254),
.B1(n_213),
.B2(n_208),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_196),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_241),
.B(n_242),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_219),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g243 ( 
.A(n_208),
.B(n_179),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_243),
.Y(n_276)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_245),
.Y(n_267)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_246),
.Y(n_259)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_223),
.Y(n_248)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_248),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_249),
.A2(n_226),
.B(n_207),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_250),
.B(n_212),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.C(n_253),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_206),
.B(n_192),
.C(n_178),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_206),
.B(n_179),
.C(n_199),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_203),
.A2(n_179),
.B1(n_181),
.B2(n_198),
.Y(n_254)
);

OAI32xp33_ASAP7_75t_L g255 ( 
.A1(n_228),
.A2(n_195),
.A3(n_177),
.B1(n_193),
.B2(n_188),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_221),
.Y(n_281)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_227),
.Y(n_256)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_256),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_258),
.A2(n_239),
.B1(n_233),
.B2(n_187),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_260),
.B(n_188),
.Y(n_301)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_261),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_232),
.B(n_251),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_264),
.C(n_269),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_241),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_263),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_252),
.B(n_218),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_254),
.A2(n_220),
.B1(n_206),
.B2(n_228),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_268),
.A2(n_270),
.B1(n_282),
.B2(n_236),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_225),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_238),
.A2(n_206),
.B1(n_208),
.B2(n_229),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g307 ( 
.A1(n_271),
.A2(n_272),
.B(n_281),
.Y(n_307)
);

MAJx2_ASAP7_75t_L g274 ( 
.A(n_240),
.B(n_214),
.C(n_204),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_274),
.B(n_170),
.C(n_194),
.Y(n_312)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_246),
.Y(n_275)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

FAx1_ASAP7_75t_SL g277 ( 
.A(n_242),
.B(n_204),
.CI(n_221),
.CON(n_277),
.SN(n_277)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_287),
.Y(n_288)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_234),
.Y(n_278)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_278),
.Y(n_298)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_233),
.Y(n_279)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_279),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_238),
.B1(n_231),
.B2(n_243),
.Y(n_296)
);

AOI22x1_ASAP7_75t_L g282 ( 
.A1(n_237),
.A2(n_238),
.B1(n_255),
.B2(n_243),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_235),
.A2(n_221),
.B(n_184),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_283),
.B(n_284),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_249),
.A2(n_221),
.B(n_176),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_234),
.Y(n_285)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_285),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_230),
.B(n_176),
.Y(n_286)
);

INVxp33_ASAP7_75t_SL g305 ( 
.A(n_286),
.Y(n_305)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_244),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_290),
.A2(n_300),
.B1(n_303),
.B2(n_308),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_273),
.B(n_248),
.Y(n_293)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_293),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_267),
.A2(n_231),
.B1(n_256),
.B2(n_245),
.Y(n_294)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_294),
.Y(n_330)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_262),
.B(n_253),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_297),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_296),
.A2(n_306),
.B1(n_272),
.B2(n_277),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_257),
.B(n_239),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g334 ( 
.A(n_301),
.B(n_312),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_269),
.B(n_199),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_310),
.Y(n_331)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_258),
.A2(n_224),
.B1(n_193),
.B2(n_150),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g306 ( 
.A1(n_268),
.A2(n_224),
.B1(n_194),
.B2(n_33),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_281),
.A2(n_142),
.B1(n_136),
.B2(n_94),
.Y(n_308)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_257),
.B(n_188),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_284),
.A2(n_146),
.B1(n_128),
.B2(n_153),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_277),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_309),
.B(n_302),
.C(n_297),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_316),
.B(n_319),
.C(n_326),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g317 ( 
.A(n_293),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_322),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_309),
.B(n_264),
.C(n_270),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_289),
.B(n_271),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_321),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_311),
.B(n_259),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_283),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_304),
.Y(n_324)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_324),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_295),
.B(n_276),
.C(n_260),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_305),
.B(n_265),
.Y(n_327)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_327),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_310),
.B(n_276),
.C(n_274),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_328),
.B(n_333),
.C(n_337),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_292),
.B(n_279),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_329),
.Y(n_349)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_282),
.C(n_280),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_335),
.A2(n_336),
.B1(n_299),
.B2(n_298),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_34),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_301),
.B(n_296),
.C(n_313),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_330),
.A2(n_288),
.B1(n_291),
.B2(n_282),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g375 ( 
.A1(n_339),
.A2(n_350),
.B1(n_354),
.B2(n_6),
.Y(n_375)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_333),
.A2(n_308),
.B1(n_300),
.B2(n_313),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_340),
.A2(n_335),
.B1(n_337),
.B2(n_318),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_316),
.B(n_307),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_341),
.B(n_357),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g342 ( 
.A1(n_322),
.A2(n_307),
.B(n_304),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_342),
.A2(n_6),
.B(n_8),
.Y(n_374)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_345),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_319),
.B(n_303),
.C(n_314),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_347),
.B(n_351),
.C(n_352),
.Y(n_365)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_323),
.A2(n_33),
.B1(n_22),
.B2(n_103),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_325),
.B(n_33),
.C(n_63),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_325),
.B(n_1),
.C(n_2),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_331),
.B(n_1),
.C(n_4),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_353),
.B(n_322),
.C(n_334),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_323),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_SL g356 ( 
.A(n_326),
.B(n_4),
.C(n_5),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_6),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g357 ( 
.A(n_331),
.B(n_4),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_SL g380 ( 
.A(n_360),
.B(n_374),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_349),
.B(n_315),
.Y(n_361)
);

OAI321xp33_ASAP7_75t_L g385 ( 
.A1(n_361),
.A2(n_370),
.A3(n_352),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_385)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_355),
.Y(n_362)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_362),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_348),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_363),
.B(n_367),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_SL g364 ( 
.A(n_341),
.B(n_328),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_SL g377 ( 
.A(n_364),
.B(n_338),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_366),
.A2(n_373),
.B1(n_358),
.B2(n_350),
.Y(n_384)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_344),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_368),
.B(n_369),
.Y(n_387)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_339),
.Y(n_369)
);

O2A1O1Ixp33_ASAP7_75t_L g370 ( 
.A1(n_342),
.A2(n_334),
.B(n_7),
.C(n_8),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_338),
.B(n_6),
.C(n_7),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_371),
.B(n_376),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_340),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g390 ( 
.A1(n_374),
.A2(n_9),
.B(n_11),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_375),
.A2(n_347),
.B1(n_351),
.B2(n_353),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_354),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g395 ( 
.A(n_377),
.B(n_380),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_362),
.B(n_346),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_378),
.B(n_386),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g379 ( 
.A1(n_369),
.A2(n_358),
.B(n_343),
.Y(n_379)
);

OR2x2_ASAP7_75t_L g402 ( 
.A(n_379),
.B(n_385),
.Y(n_402)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_381),
.Y(n_396)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_384),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_364),
.B(n_343),
.C(n_357),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_359),
.B(n_14),
.C(n_11),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_389),
.B(n_390),
.Y(n_401)
);

AOI21xp5_ASAP7_75t_L g391 ( 
.A1(n_387),
.A2(n_361),
.B(n_372),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_391),
.A2(n_394),
.B(n_399),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_384),
.A2(n_375),
.B1(n_366),
.B2(n_367),
.Y(n_392)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_392),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_SL g393 ( 
.A(n_383),
.B(n_371),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g408 ( 
.A(n_393),
.B(n_389),
.Y(n_408)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_379),
.A2(n_365),
.B(n_359),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_388),
.B(n_368),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_398),
.B(n_382),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_386),
.A2(n_365),
.B(n_370),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g403 ( 
.A(n_392),
.B(n_397),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g418 ( 
.A(n_403),
.B(n_410),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_391),
.B(n_377),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_404),
.B(n_407),
.Y(n_419)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_406),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_381),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_408),
.B(n_9),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_402),
.B(n_400),
.Y(n_410)
);

OAI21xp5_ASAP7_75t_SL g411 ( 
.A1(n_395),
.A2(n_373),
.B(n_390),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_L g416 ( 
.A1(n_411),
.A2(n_12),
.B(n_13),
.Y(n_416)
);

NOR2xp67_ASAP7_75t_SL g412 ( 
.A(n_396),
.B(n_9),
.Y(n_412)
);

OAI21x1_ASAP7_75t_SL g413 ( 
.A1(n_412),
.A2(n_401),
.B(n_11),
.Y(n_413)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_413),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_417),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_SL g417 ( 
.A1(n_409),
.A2(n_13),
.B(n_405),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_419),
.B(n_403),
.C(n_409),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_420),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_415),
.Y(n_422)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_422),
.Y(n_425)
);

AO21x1_ASAP7_75t_L g426 ( 
.A1(n_425),
.A2(n_423),
.B(n_422),
.Y(n_426)
);

BUFx24_ASAP7_75t_SL g427 ( 
.A(n_426),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_427),
.A2(n_424),
.B(n_414),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_428),
.B(n_421),
.Y(n_429)
);


endmodule