module real_jpeg_3259_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_293, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_293;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_288;
wire n_166;
wire n_249;
wire n_221;
wire n_176;
wire n_215;
wire n_286;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_255;
wire n_105;
wire n_40;
wire n_173;
wire n_197;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_155;
wire n_113;
wire n_199;
wire n_251;
wire n_93;
wire n_141;
wire n_95;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_285;
wire n_172;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_193;
wire n_99;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_70;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_209;
wire n_55;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_202;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_181;
wire n_85;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_269;
wire n_273;
wire n_89;

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

OAI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

OAI22xp33_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_50),
.B1(n_56),
.B2(n_57),
.Y(n_65)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_1),
.A2(n_26),
.B1(n_31),
.B2(n_50),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_1),
.A2(n_42),
.B1(n_44),
.B2(n_50),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_2),
.A2(n_56),
.B1(n_57),
.B2(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_2),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_2),
.A2(n_42),
.B1(n_44),
.B2(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_2),
.A2(n_26),
.B1(n_31),
.B2(n_63),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_141),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_3),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_141),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_3),
.A2(n_26),
.B1(n_31),
.B2(n_141),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_141),
.Y(n_241)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_104),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_5),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_104),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_5),
.A2(n_26),
.B1(n_31),
.B2(n_104),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_5),
.A2(n_56),
.B1(n_57),
.B2(n_104),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_6),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_6),
.A2(n_56),
.B1(n_57),
.B2(n_162),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_6),
.A2(n_26),
.B1(n_31),
.B2(n_162),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_6),
.A2(n_42),
.B1(n_44),
.B2(n_162),
.Y(n_229)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_7),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_10),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_11),
.A2(n_26),
.B1(n_31),
.B2(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_11),
.A2(n_32),
.B1(n_37),
.B2(n_38),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_11),
.A2(n_32),
.B1(n_56),
.B2(n_57),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_11),
.A2(n_32),
.B1(n_42),
.B2(n_44),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g151 ( 
.A(n_12),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_26),
.C(n_59),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_12),
.A2(n_56),
.B1(n_57),
.B2(n_151),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_12),
.B(n_29),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_12),
.B(n_66),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_12),
.B(n_44),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_12),
.A2(n_44),
.B(n_220),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_12),
.B(n_48),
.Y(n_244)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_12),
.A2(n_37),
.B(n_256),
.Y(n_255)
);

BUFx10_ASAP7_75t_L g39 ( 
.A(n_13),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_14),
.A2(n_42),
.B1(n_44),
.B2(n_76),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_14),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_14),
.A2(n_56),
.B1(n_57),
.B2(n_76),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_14),
.A2(n_37),
.B1(n_38),
.B2(n_76),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_14),
.A2(n_26),
.B1(n_31),
.B2(n_76),
.Y(n_155)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_125),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_123),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_106),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_19),
.B(n_106),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.C(n_87),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_20),
.B(n_67),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_51),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_33),
.B2(n_34),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_22),
.A2(n_23),
.B1(n_52),
.B2(n_168),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_52),
.Y(n_51)
);

AOI21xp33_ASAP7_75t_L g107 ( 
.A1(n_23),
.A2(n_33),
.B(n_51),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_28),
.B(n_30),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_24),
.A2(n_133),
.B(n_135),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g207 ( 
.A1(n_24),
.A2(n_28),
.B1(n_208),
.B2(n_209),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_24),
.A2(n_30),
.B(n_135),
.Y(n_222)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_25),
.B(n_96),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_25),
.A2(n_29),
.B1(n_134),
.B2(n_154),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_25),
.A2(n_93),
.B(n_181),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_25),
.A2(n_29),
.B1(n_151),
.B2(n_200),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_25),
.A2(n_29),
.B1(n_200),
.B2(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

OA22x2_ASAP7_75t_L g61 ( 
.A1(n_26),
.A2(n_31),
.B1(n_59),
.B2(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_26),
.B(n_198),
.Y(n_197)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_28),
.B(n_30),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_28),
.A2(n_95),
.B(n_155),
.Y(n_246)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_29),
.B(n_96),
.Y(n_135)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_45),
.B(n_47),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_35),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_35),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_35),
.A2(n_41),
.B1(n_103),
.B2(n_140),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_35),
.A2(n_41),
.B1(n_140),
.B2(n_161),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_35),
.A2(n_41),
.B1(n_161),
.B2(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_41),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_38),
.B(n_151),
.Y(n_150)
);

NAND3xp33_ASAP7_75t_L g152 ( 
.A(n_38),
.B(n_40),
.C(n_44),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

OA22x2_ASAP7_75t_L g41 ( 
.A1(n_39),
.A2(n_40),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

A2O1A1Ixp33_ASAP7_75t_L g149 ( 
.A1(n_39),
.A2(n_42),
.B(n_150),
.C(n_152),
.Y(n_149)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_41),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

CKINVDCx6p67_ASAP7_75t_R g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_42),
.A2(n_44),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

OAI32xp33_ASAP7_75t_L g218 ( 
.A1(n_44),
.A2(n_57),
.A3(n_80),
.B1(n_219),
.B2(n_221),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_46),
.B(n_48),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_49),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_49),
.B(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_52),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g52 ( 
.A1(n_53),
.A2(n_62),
.B(n_64),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_53),
.A2(n_61),
.B1(n_62),
.B2(n_98),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_53),
.A2(n_61),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_53),
.A2(n_64),
.B(n_70),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_65),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_54),
.A2(n_66),
.B(n_116),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_54),
.A2(n_66),
.B1(n_185),
.B2(n_186),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_54),
.A2(n_66),
.B1(n_185),
.B2(n_193),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_54),
.A2(n_69),
.B(n_235),
.Y(n_234)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_61),
.Y(n_54)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_55)
);

OA22x2_ASAP7_75t_SL g83 ( 
.A1(n_56),
.A2(n_57),
.B1(n_80),
.B2(n_82),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_56),
.B(n_82),
.Y(n_221)
);

CKINVDCx6p67_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_57),
.B(n_190),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx13_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_61),
.B(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_61),
.A2(n_72),
.B(n_98),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_65),
.B(n_66),
.Y(n_64)
);

OAI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_68),
.A2(n_73),
.B(n_86),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_68),
.B(n_73),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

INVxp33_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_77),
.B1(n_84),
.B2(n_85),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_83),
.B(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_101),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g111 ( 
.A1(n_77),
.A2(n_85),
.B(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_77),
.A2(n_84),
.B1(n_239),
.B2(n_240),
.Y(n_238)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_78),
.A2(n_113),
.B(n_143),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g156 ( 
.A1(n_78),
.A2(n_157),
.B(n_158),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_78),
.A2(n_83),
.B1(n_228),
.B2(n_229),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_78),
.A2(n_83),
.B1(n_157),
.B2(n_241),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_83),
.Y(n_78)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_80),
.Y(n_82)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_83),
.B(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_84),
.B(n_101),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_84),
.B(n_159),
.Y(n_158)
);

FAx1_ASAP7_75t_SL g106 ( 
.A(n_86),
.B(n_107),
.CI(n_108),
.CON(n_106),
.SN(n_106)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_87),
.A2(n_88),
.B1(n_287),
.B2(n_288),
.Y(n_286)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_99),
.C(n_102),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_89),
.A2(n_90),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_92),
.B1(n_97),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVxp33_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_99),
.B(n_102),
.Y(n_171)
);

BUFx24_ASAP7_75t_SL g291 ( 
.A(n_106),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_109),
.A2(n_110),
.B1(n_118),
.B2(n_122),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_111),
.A2(n_114),
.B1(n_115),
.B2(n_117),
.Y(n_110)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_111),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_118),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_285),
.B(n_290),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_173),
.B(n_284),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_163),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_128),
.B(n_163),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_144),
.C(n_146),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_129),
.B(n_144),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_130),
.A2(n_131),
.B1(n_137),
.B2(n_138),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_130),
.B(n_139),
.C(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_136),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g275 ( 
.A(n_132),
.B(n_136),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_142),
.Y(n_138)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_143),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_146),
.B(n_268),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_156),
.C(n_160),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g271 ( 
.A(n_147),
.B(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_153),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_148),
.A2(n_149),
.B1(n_153),
.B2(n_264),
.Y(n_263)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_150),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_153),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_156),
.B(n_160),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_172),
.Y(n_163)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_167),
.B(n_169),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_167),
.B(n_169),
.C(n_172),
.Y(n_289)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI321xp33_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_266),
.A3(n_276),
.B1(n_282),
.B2(n_283),
.C(n_293),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_249),
.B(n_265),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_231),
.B(n_248),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_213),
.B(n_230),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_194),
.B(n_212),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_187),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_187),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_182),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_180),
.B(n_184),
.C(n_215),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_181),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_183),
.Y(n_215)
);

INVxp67_ASAP7_75t_L g225 ( 
.A(n_186),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_191),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_188),
.A2(n_189),
.B1(n_191),
.B2(n_192),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_206),
.B(n_211),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_196),
.A2(n_201),
.B(n_205),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_202),
.B(n_204),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g208 ( 
.A(n_203),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_210),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_207),
.B(n_210),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_216),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_223),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_217),
.B(n_224),
.C(n_227),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_222),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_218),
.B(n_222),
.Y(n_236)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_227),
.Y(n_223)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_226),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_229),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_247),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_232),
.B(n_247),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_236),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_236),
.C(n_237),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_238),
.B(n_242),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_238),
.B(n_244),
.C(n_245),
.Y(n_262)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_251),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_260),
.B2(n_261),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_252),
.B(n_262),
.C(n_263),
.Y(n_277)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_257),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_254),
.B(n_258),
.C(n_259),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_267),
.B(n_269),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_267),
.B(n_269),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_273),
.C(n_275),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_270),
.A2(n_271),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_273),
.A2(n_274),
.B1(n_275),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_275),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_289),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_286),
.B(n_289),
.Y(n_290)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);


endmodule