module fake_jpeg_3852_n_315 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_315);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_315;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_15),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx16_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_4),
.B(n_9),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_8),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_37),
.Y(n_45)
);

BUFx12f_ASAP7_75t_SL g36 ( 
.A(n_33),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_36),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_8),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_39),
.Y(n_66)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_0),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_18),
.Y(n_48)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_17),
.B(n_8),
.Y(n_42)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_36),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_46),
.B(n_50),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_48),
.B(n_62),
.Y(n_92)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_41),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_53),
.A2(n_58),
.B1(n_60),
.B2(n_67),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_41),
.A2(n_28),
.B1(n_27),
.B2(n_19),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_54),
.A2(n_59),
.B1(n_22),
.B2(n_42),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_44),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_40),
.A2(n_28),
.B1(n_27),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_25),
.B1(n_20),
.B2(n_23),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_39),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_40),
.B(n_18),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_18),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_59),
.Y(n_81)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_44),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_69),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g67 ( 
.A1(n_40),
.A2(n_32),
.B1(n_30),
.B2(n_21),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_35),
.A2(n_21),
.B1(n_22),
.B2(n_24),
.Y(n_68)
);

OA22x2_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_71),
.B1(n_12),
.B2(n_14),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_24),
.B1(n_22),
.B2(n_26),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g74 ( 
.A(n_47),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_78),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_45),
.B1(n_66),
.B2(n_54),
.Y(n_107)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

INVx11_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_48),
.A2(n_37),
.B(n_29),
.C(n_43),
.Y(n_78)
);

FAx1_ASAP7_75t_SL g80 ( 
.A(n_62),
.B(n_43),
.CI(n_26),
.CON(n_80),
.SN(n_80)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_80),
.B(n_81),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_63),
.B(n_0),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_14),
.B(n_15),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_52),
.B(n_34),
.Y(n_83)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_83),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_43),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_84),
.B(n_86),
.Y(n_102)
);

INVx4_ASAP7_75t_SL g85 ( 
.A(n_46),
.Y(n_85)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_43),
.Y(n_86)
);

A2O1A1Ixp33_ASAP7_75t_L g87 ( 
.A1(n_49),
.A2(n_26),
.B(n_31),
.C(n_12),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_95),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_56),
.B(n_26),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_88),
.B(n_26),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_93),
.A2(n_50),
.B1(n_52),
.B2(n_64),
.Y(n_98)
);

NOR2x1_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_26),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_31),
.Y(n_109)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_66),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_96),
.Y(n_101)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_95),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_97),
.B(n_103),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_93),
.B1(n_87),
.B2(n_94),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_104),
.B(n_106),
.Y(n_133)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_113),
.B1(n_123),
.B2(n_89),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_108),
.B(n_82),
.Y(n_129)
);

OR2x4_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_85),
.Y(n_150)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_72),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_110),
.B(n_112),
.Y(n_144)
);

INVx13_ASAP7_75t_L g112 ( 
.A(n_91),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_45),
.B1(n_65),
.B2(n_61),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_115),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_76),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_117),
.B(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_86),
.Y(n_118)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_75),
.Y(n_120)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_120),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_SL g121 ( 
.A(n_91),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_121),
.Y(n_126)
);

INVx13_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_81),
.A2(n_55),
.B1(n_65),
.B2(n_61),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_105),
.A2(n_94),
.B(n_96),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g168 ( 
.A1(n_124),
.A2(n_150),
.B(n_147),
.Y(n_168)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_123),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_127),
.B(n_130),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_146),
.B1(n_141),
.B2(n_127),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_129),
.B(n_134),
.Y(n_163)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_105),
.B(n_92),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_135),
.A2(n_149),
.B1(n_145),
.B2(n_125),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_101),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_102),
.B(n_92),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_137),
.B(n_140),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_101),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_139),
.B(n_141),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_102),
.B(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_113),
.Y(n_141)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_80),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_147),
.Y(n_177)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_145),
.B(n_146),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_107),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_111),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g148 ( 
.A(n_99),
.B(n_89),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_148),
.B(n_100),
.C(n_110),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_109),
.B(n_80),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_149),
.A2(n_116),
.B(n_115),
.Y(n_160)
);

OA21x2_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_111),
.B(n_104),
.Y(n_153)
);

AO22x1_ASAP7_75t_SL g151 ( 
.A1(n_109),
.A2(n_93),
.B1(n_78),
.B2(n_90),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_151),
.A2(n_98),
.B1(n_93),
.B2(n_100),
.Y(n_162)
);

AO21x1_ASAP7_75t_L g209 ( 
.A1(n_153),
.A2(n_31),
.B(n_69),
.Y(n_209)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_133),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_154),
.B(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_144),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_152),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_157),
.B(n_166),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_173),
.B1(n_172),
.B2(n_162),
.Y(n_199)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_160),
.A2(n_168),
.B(n_172),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_164),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_134),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_179),
.C(n_122),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_143),
.B(n_137),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_167),
.B(n_171),
.Y(n_186)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_169),
.B(n_170),
.Y(n_201)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_151),
.B(n_117),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_151),
.B(n_83),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_128),
.A2(n_79),
.B1(n_114),
.B2(n_106),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_176),
.A2(n_130),
.B1(n_139),
.B2(n_136),
.Y(n_189)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_149),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_178),
.B(n_182),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_124),
.B(n_114),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_125),
.A2(n_79),
.B(n_97),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_181),
.B(n_122),
.Y(n_198)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_184),
.B(n_188),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_175),
.B(n_138),
.Y(n_187)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_187),
.Y(n_230)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_161),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_189),
.A2(n_153),
.B1(n_119),
.B2(n_159),
.Y(n_215)
);

AND2x2_ASAP7_75t_L g192 ( 
.A(n_179),
.B(n_126),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g217 ( 
.A1(n_192),
.A2(n_153),
.B(n_159),
.Y(n_217)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_163),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_193),
.B(n_196),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_138),
.Y(n_194)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_194),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_181),
.B(n_112),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_195),
.B(n_208),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g196 ( 
.A(n_177),
.Y(n_196)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_198),
.B(n_31),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_199),
.A2(n_73),
.B1(n_132),
.B2(n_142),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_126),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_203),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_205),
.C(n_174),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_163),
.B(n_74),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_119),
.B1(n_73),
.B2(n_77),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_204),
.A2(n_166),
.B1(n_119),
.B2(n_169),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_112),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_69),
.C(n_31),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_SL g227 ( 
.A(n_206),
.B(n_203),
.Y(n_227)
);

OAI21xp33_ASAP7_75t_L g207 ( 
.A1(n_177),
.A2(n_10),
.B(n_16),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_207),
.B(n_160),
.Y(n_212)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_180),
.Y(n_208)
);

OA21x2_ASAP7_75t_L g225 ( 
.A1(n_209),
.A2(n_30),
.B(n_32),
.Y(n_225)
);

AOI22x1_ASAP7_75t_SL g210 ( 
.A1(n_191),
.A2(n_172),
.B1(n_176),
.B2(n_171),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_210),
.A2(n_191),
.B(n_201),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_222),
.B1(n_226),
.B2(n_230),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g247 ( 
.A(n_212),
.B(n_186),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_213),
.B(n_214),
.C(n_224),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_174),
.C(n_167),
.Y(n_214)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_215),
.Y(n_242)
);

INVx4_ASAP7_75t_L g216 ( 
.A(n_197),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_216),
.B(n_218),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_217),
.B(n_220),
.Y(n_248)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_190),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_223),
.B(n_225),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_185),
.B(n_32),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_132),
.B1(n_120),
.B2(n_103),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_227),
.B(n_233),
.C(n_202),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_184),
.A2(n_32),
.B1(n_13),
.B2(n_16),
.Y(n_228)
);

A2O1A1Ixp33_ASAP7_75t_L g249 ( 
.A1(n_228),
.A2(n_13),
.B(n_14),
.C(n_11),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_185),
.B(n_11),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_200),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_234),
.B(n_1),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_235),
.A2(n_237),
.B1(n_249),
.B2(n_250),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_217),
.A2(n_219),
.B1(n_210),
.B2(n_192),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g238 ( 
.A(n_221),
.B(n_183),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_238),
.B(n_245),
.Y(n_267)
);

BUFx2_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_239),
.B(n_251),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_240),
.A2(n_254),
.B(n_225),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_241),
.B(n_225),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_193),
.Y(n_245)
);

AOI31xp67_ASAP7_75t_L g246 ( 
.A1(n_227),
.A2(n_192),
.A3(n_198),
.B(n_209),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_246),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_247),
.B(n_233),
.C(n_224),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_206),
.B1(n_186),
.B2(n_120),
.Y(n_250)
);

BUFx2_ASAP7_75t_L g251 ( 
.A(n_231),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_103),
.C(n_57),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_252),
.B(n_214),
.C(n_220),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_229),
.A2(n_75),
.B1(n_57),
.B2(n_55),
.Y(n_253)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_253),
.Y(n_266)
);

NOR2x1_ASAP7_75t_L g254 ( 
.A(n_215),
.B(n_0),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_255),
.B(n_212),
.Y(n_256)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_256),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_249),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_263),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g260 ( 
.A(n_254),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g281 ( 
.A(n_260),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_262),
.A2(n_271),
.B(n_241),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_239),
.B(n_55),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_251),
.B(n_3),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_237),
.A2(n_1),
.B(n_2),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_270),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_236),
.B(n_3),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_246),
.A2(n_242),
.B(n_235),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_271),
.B(n_236),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_274),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_263),
.B(n_250),
.Y(n_274)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_275),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_262),
.B(n_248),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_276),
.B(n_248),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_277),
.B(n_279),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_278),
.B(n_4),
.C(n_6),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g279 ( 
.A1(n_259),
.A2(n_252),
.B(n_244),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_243),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_282),
.B(n_267),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_257),
.B(n_269),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g303 ( 
.A1(n_286),
.A2(n_10),
.B(n_1),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_284),
.B(n_264),
.Y(n_287)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_287),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_288),
.B(n_291),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_294),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_281),
.B(n_258),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_274),
.A2(n_247),
.B1(n_270),
.B2(n_3),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_292),
.B(n_280),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_280),
.A2(n_273),
.B1(n_272),
.B2(n_276),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_295),
.A2(n_272),
.B1(n_4),
.B2(n_7),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_290),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_293),
.B(n_285),
.Y(n_300)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_300),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_301),
.B(n_303),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_1),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_302),
.Y(n_309)
);

AOI321xp33_ASAP7_75t_L g304 ( 
.A1(n_298),
.A2(n_2),
.A3(n_10),
.B1(n_290),
.B2(n_294),
.C(n_297),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_304),
.B(n_305),
.C(n_297),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g308 ( 
.A(n_299),
.B(n_2),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_308),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_310),
.A2(n_311),
.B(n_306),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_307),
.B(n_303),
.C(n_309),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_306),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);


endmodule