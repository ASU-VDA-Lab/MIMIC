module fake_netlist_6_4939_n_4521 (n_52, n_1, n_91, n_326, n_256, n_209, n_367, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_144, n_365, n_125, n_168, n_384, n_297, n_342, n_77, n_106, n_358, n_160, n_131, n_188, n_310, n_186, n_245, n_0, n_368, n_396, n_350, n_78, n_84, n_392, n_142, n_143, n_382, n_180, n_62, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_67, n_15, n_246, n_38, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_389, n_415, n_65, n_230, n_141, n_383, n_200, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_71, n_74, n_229, n_305, n_72, n_173, n_250, n_372, n_111, n_314, n_378, n_413, n_377, n_35, n_183, n_79, n_375, n_338, n_56, n_360, n_119, n_235, n_147, n_191, n_340, n_387, n_39, n_344, n_73, n_428, n_101, n_167, n_174, n_127, n_153, n_156, n_145, n_42, n_133, n_96, n_8, n_371, n_189, n_405, n_213, n_294, n_302, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_20, n_397, n_155, n_109, n_425, n_122, n_45, n_34, n_218, n_70, n_234, n_37, n_381, n_82, n_27, n_236, n_112, n_172, n_270, n_239, n_126, n_414, n_97, n_58, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_9, n_107, n_6, n_417, n_14, n_89, n_374, n_366, n_407, n_103, n_272, n_185, n_348, n_69, n_376, n_390, n_293, n_31, n_334, n_53, n_370, n_44, n_232, n_16, n_163, n_46, n_330, n_298, n_18, n_281, n_258, n_154, n_98, n_260, n_265, n_313, n_279, n_252, n_228, n_356, n_166, n_184, n_216, n_83, n_363, n_395, n_323, n_393, n_411, n_152, n_92, n_321, n_331, n_105, n_227, n_132, n_406, n_102, n_204, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_164, n_292, n_100, n_121, n_307, n_23, n_2, n_291, n_219, n_357, n_150, n_264, n_263, n_325, n_329, n_33, n_408, n_61, n_237, n_244, n_399, n_76, n_243, n_124, n_94, n_282, n_116, n_211, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_240, n_139, n_319, n_41, n_134, n_273, n_95, n_311, n_10, n_403, n_253, n_123, n_136, n_249, n_201, n_386, n_159, n_157, n_162, n_115, n_128, n_241, n_30, n_275, n_43, n_276, n_221, n_423, n_146, n_318, n_303, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_277, n_418, n_113, n_4, n_199, n_138, n_266, n_296, n_268, n_271, n_404, n_158, n_217, n_49, n_210, n_299, n_206, n_5, n_333, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_90, n_347, n_24, n_54, n_328, n_429, n_373, n_87, n_195, n_285, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_339, n_315, n_64, n_288, n_427, n_422, n_135, n_165, n_351, n_259, n_177, n_391, n_364, n_295, n_385, n_388, n_190, n_262, n_187, n_60, n_361, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_4521);

input n_52;
input n_1;
input n_91;
input n_326;
input n_256;
input n_209;
input n_367;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_131;
input n_188;
input n_310;
input n_186;
input n_245;
input n_0;
input n_368;
input n_396;
input n_350;
input n_78;
input n_84;
input n_392;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_67;
input n_15;
input n_246;
input n_38;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_389;
input n_415;
input n_65;
input n_230;
input n_141;
input n_383;
input n_200;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_71;
input n_74;
input n_229;
input n_305;
input n_72;
input n_173;
input n_250;
input n_372;
input n_111;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_79;
input n_375;
input n_338;
input n_56;
input n_360;
input n_119;
input n_235;
input n_147;
input n_191;
input n_340;
input n_387;
input n_39;
input n_344;
input n_73;
input n_428;
input n_101;
input n_167;
input n_174;
input n_127;
input n_153;
input n_156;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_189;
input n_405;
input n_213;
input n_294;
input n_302;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_20;
input n_397;
input n_155;
input n_109;
input n_425;
input n_122;
input n_45;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_58;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_9;
input n_107;
input n_6;
input n_417;
input n_14;
input n_89;
input n_374;
input n_366;
input n_407;
input n_103;
input n_272;
input n_185;
input n_348;
input n_69;
input n_376;
input n_390;
input n_293;
input n_31;
input n_334;
input n_53;
input n_370;
input n_44;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_298;
input n_18;
input n_281;
input n_258;
input n_154;
input n_98;
input n_260;
input n_265;
input n_313;
input n_279;
input n_252;
input n_228;
input n_356;
input n_166;
input n_184;
input n_216;
input n_83;
input n_363;
input n_395;
input n_323;
input n_393;
input n_411;
input n_152;
input n_92;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_406;
input n_102;
input n_204;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_23;
input n_2;
input n_291;
input n_219;
input n_357;
input n_150;
input n_264;
input n_263;
input n_325;
input n_329;
input n_33;
input n_408;
input n_61;
input n_237;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_94;
input n_282;
input n_116;
input n_211;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_273;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_123;
input n_136;
input n_249;
input n_201;
input n_386;
input n_159;
input n_157;
input n_162;
input n_115;
input n_128;
input n_241;
input n_30;
input n_275;
input n_43;
input n_276;
input n_221;
input n_423;
input n_146;
input n_318;
input n_303;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_277;
input n_418;
input n_113;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_268;
input n_271;
input n_404;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_206;
input n_5;
input n_333;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_90;
input n_347;
input n_24;
input n_54;
input n_328;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_339;
input n_315;
input n_64;
input n_288;
input n_427;
input n_422;
input n_135;
input n_165;
input n_351;
input n_259;
input n_177;
input n_391;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_187;
input n_60;
input n_361;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_4521;

wire n_992;
wire n_2542;
wire n_1671;
wire n_2817;
wire n_3660;
wire n_3813;
wire n_801;
wire n_4452;
wire n_3766;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_3254;
wire n_3684;
wire n_1199;
wire n_1674;
wire n_3392;
wire n_741;
wire n_1027;
wire n_1351;
wire n_3266;
wire n_3574;
wire n_625;
wire n_1189;
wire n_3152;
wire n_4154;
wire n_3579;
wire n_1212;
wire n_4251;
wire n_726;
wire n_2157;
wire n_3335;
wire n_2332;
wire n_3783;
wire n_700;
wire n_3773;
wire n_4177;
wire n_1307;
wire n_3178;
wire n_2003;
wire n_3849;
wire n_4127;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_4504;
wire n_3844;
wire n_4388;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_3089;
wire n_3301;
wire n_4395;
wire n_4099;
wire n_1357;
wire n_4241;
wire n_1853;
wire n_3741;
wire n_4517;
wire n_4168;
wire n_783;
wire n_4372;
wire n_2451;
wire n_1738;
wire n_4490;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_3088;
wire n_3443;
wire n_1923;
wire n_3257;
wire n_509;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_3222;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_2977;
wire n_3952;
wire n_1739;
wire n_2051;
wire n_4370;
wire n_2317;
wire n_1380;
wire n_3911;
wire n_2359;
wire n_442;
wire n_480;
wire n_2847;
wire n_1402;
wire n_2557;
wire n_1688;
wire n_1691;
wire n_3332;
wire n_4285;
wire n_4134;
wire n_3465;
wire n_1975;
wire n_1009;
wire n_1930;
wire n_1743;
wire n_2405;
wire n_3706;
wire n_4050;
wire n_1160;
wire n_883;
wire n_2647;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_2997;
wire n_4092;
wire n_1724;
wire n_1032;
wire n_3708;
wire n_2336;
wire n_1247;
wire n_3668;
wire n_4078;
wire n_1547;
wire n_2521;
wire n_3376;
wire n_3046;
wire n_2956;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_3801;
wire n_4249;
wire n_1264;
wire n_1192;
wire n_471;
wire n_3564;
wire n_1844;
wire n_3619;
wire n_4359;
wire n_4087;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_3487;
wire n_4198;
wire n_2382;
wire n_3754;
wire n_2672;
wire n_3030;
wire n_4302;
wire n_2291;
wire n_830;
wire n_2299;
wire n_3340;
wire n_4179;
wire n_461;
wire n_873;
wire n_1371;
wire n_1285;
wire n_2886;
wire n_2974;
wire n_3946;
wire n_1985;
wire n_4213;
wire n_2989;
wire n_447;
wire n_2838;
wire n_2184;
wire n_3395;
wire n_2982;
wire n_1803;
wire n_3427;
wire n_1172;
wire n_4474;
wire n_852;
wire n_2509;
wire n_4065;
wire n_4026;
wire n_2513;
wire n_3282;
wire n_1590;
wire n_2645;
wire n_1532;
wire n_2313;
wire n_2628;
wire n_3071;
wire n_3626;
wire n_3757;
wire n_3904;
wire n_4178;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_2926;
wire n_1704;
wire n_1078;
wire n_544;
wire n_1711;
wire n_2247;
wire n_3106;
wire n_1140;
wire n_2630;
wire n_4273;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_3275;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_4446;
wire n_1263;
wire n_2019;
wire n_3031;
wire n_4029;
wire n_836;
wire n_3345;
wire n_2074;
wire n_4417;
wire n_2447;
wire n_522;
wire n_2919;
wire n_4501;
wire n_3678;
wire n_3440;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_3879;
wire n_4010;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_3080;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_3979;
wire n_658;
wire n_616;
wire n_4308;
wire n_1874;
wire n_4347;
wire n_3165;
wire n_1119;
wire n_2865;
wire n_2825;
wire n_3463;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_2510;
wire n_1735;
wire n_2739;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_1954;
wire n_3023;
wire n_822;
wire n_3232;
wire n_693;
wire n_1313;
wire n_2791;
wire n_3607;
wire n_3750;
wire n_3251;
wire n_1056;
wire n_3877;
wire n_3316;
wire n_4325;
wire n_2212;
wire n_3929;
wire n_758;
wire n_516;
wire n_3494;
wire n_3063;
wire n_1455;
wire n_2418;
wire n_2864;
wire n_1163;
wire n_2729;
wire n_3048;
wire n_4311;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_4060;
wire n_1550;
wire n_2703;
wire n_491;
wire n_3998;
wire n_2786;
wire n_3371;
wire n_1591;
wire n_772;
wire n_3632;
wire n_3122;
wire n_2806;
wire n_1344;
wire n_3261;
wire n_2730;
wire n_2495;
wire n_666;
wire n_4187;
wire n_940;
wire n_770;
wire n_567;
wire n_1971;
wire n_1781;
wire n_2058;
wire n_2090;
wire n_2603;
wire n_2660;
wire n_3028;
wire n_538;
wire n_3829;
wire n_3662;
wire n_2981;
wire n_3076;
wire n_2173;
wire n_4164;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_3624;
wire n_3077;
wire n_3737;
wire n_1345;
wire n_2873;
wire n_1820;
wire n_3452;
wire n_3655;
wire n_494;
wire n_539;
wire n_493;
wire n_3107;
wire n_3825;
wire n_2880;
wire n_3225;
wire n_2394;
wire n_2108;
wire n_3532;
wire n_4117;
wire n_454;
wire n_3948;
wire n_1421;
wire n_2836;
wire n_3664;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_4327;
wire n_1961;
wire n_3047;
wire n_4414;
wire n_1280;
wire n_3765;
wire n_713;
wire n_2655;
wire n_4125;
wire n_1400;
wire n_2625;
wire n_3296;
wire n_2843;
wire n_4221;
wire n_1467;
wire n_3297;
wire n_4250;
wire n_976;
wire n_3760;
wire n_3067;
wire n_2155;
wire n_3906;
wire n_2686;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_4262;
wire n_4392;
wire n_1894;
wire n_2996;
wire n_1231;
wire n_2599;
wire n_2985;
wire n_1978;
wire n_3803;
wire n_2085;
wire n_3963;
wire n_3368;
wire n_917;
wire n_574;
wire n_3639;
wire n_3347;
wire n_2370;
wire n_2612;
wire n_3792;
wire n_907;
wire n_4202;
wire n_1446;
wire n_3938;
wire n_2591;
wire n_3507;
wire n_4334;
wire n_659;
wire n_1815;
wire n_2214;
wire n_3351;
wire n_4253;
wire n_913;
wire n_4110;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_4255;
wire n_4403;
wire n_4071;
wire n_3506;
wire n_4268;
wire n_3568;
wire n_3269;
wire n_4047;
wire n_3531;
wire n_1230;
wire n_3413;
wire n_3850;
wire n_473;
wire n_1193;
wire n_1967;
wire n_3999;
wire n_1054;
wire n_3928;
wire n_559;
wire n_3412;
wire n_2613;
wire n_3535;
wire n_1333;
wire n_2496;
wire n_2708;
wire n_3313;
wire n_1648;
wire n_3189;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_3791;
wire n_4139;
wire n_2011;
wire n_2725;
wire n_2277;
wire n_3164;
wire n_1558;
wire n_1732;
wire n_551;
wire n_2300;
wire n_699;
wire n_1986;
wire n_3943;
wire n_4320;
wire n_4305;
wire n_564;
wire n_2397;
wire n_3884;
wire n_3931;
wire n_4349;
wire n_451;
wire n_824;
wire n_686;
wire n_4102;
wire n_4297;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_3603;
wire n_3871;
wire n_2907;
wire n_577;
wire n_3438;
wire n_2735;
wire n_4141;
wire n_1843;
wire n_619;
wire n_3959;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_521;
wire n_2778;
wire n_4227;
wire n_2850;
wire n_572;
wire n_4314;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_3822;
wire n_4163;
wire n_606;
wire n_1441;
wire n_818;
wire n_3373;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_513;
wire n_645;
wire n_1381;
wire n_2961;
wire n_3812;
wire n_1699;
wire n_3910;
wire n_916;
wire n_3934;
wire n_2093;
wire n_4033;
wire n_4415;
wire n_4296;
wire n_4009;
wire n_2633;
wire n_483;
wire n_3883;
wire n_2207;
wire n_1970;
wire n_2770;
wire n_608;
wire n_2101;
wire n_2696;
wire n_3482;
wire n_4080;
wire n_630;
wire n_2059;
wire n_4507;
wire n_2198;
wire n_3319;
wire n_541;
wire n_512;
wire n_2669;
wire n_2925;
wire n_3728;
wire n_4094;
wire n_4499;
wire n_2073;
wire n_2273;
wire n_3484;
wire n_433;
wire n_3748;
wire n_2546;
wire n_3272;
wire n_3193;
wire n_792;
wire n_2522;
wire n_476;
wire n_3949;
wire n_4364;
wire n_2792;
wire n_1328;
wire n_3396;
wire n_1957;
wire n_2917;
wire n_4354;
wire n_2616;
wire n_3912;
wire n_3118;
wire n_3315;
wire n_3720;
wire n_1907;
wire n_3923;
wire n_2529;
wire n_3900;
wire n_4393;
wire n_1162;
wire n_860;
wire n_1530;
wire n_3798;
wire n_788;
wire n_939;
wire n_3488;
wire n_1543;
wire n_2811;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_3732;
wire n_982;
wire n_4257;
wire n_4458;
wire n_2674;
wire n_2832;
wire n_4226;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_3980;
wire n_932;
wire n_2831;
wire n_2998;
wire n_4318;
wire n_4377;
wire n_3446;
wire n_4158;
wire n_4366;
wire n_3317;
wire n_3857;
wire n_3978;
wire n_1876;
wire n_4107;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_4074;
wire n_3716;
wire n_1873;
wire n_4294;
wire n_905;
wire n_3630;
wire n_3518;
wire n_4445;
wire n_3824;
wire n_3859;
wire n_1866;
wire n_4013;
wire n_1680;
wire n_2692;
wire n_993;
wire n_3842;
wire n_689;
wire n_3248;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_3714;
wire n_3514;
wire n_2228;
wire n_3914;
wire n_4456;
wire n_3397;
wire n_1988;
wire n_2941;
wire n_1278;
wire n_547;
wire n_3575;
wire n_2455;
wire n_2876;
wire n_558;
wire n_2654;
wire n_3036;
wire n_2469;
wire n_4032;
wire n_1064;
wire n_3099;
wire n_1396;
wire n_634;
wire n_2355;
wire n_3927;
wire n_4147;
wire n_4477;
wire n_966;
wire n_3888;
wire n_4511;
wire n_2908;
wire n_3168;
wire n_764;
wire n_4468;
wire n_2751;
wire n_2764;
wire n_3357;
wire n_1663;
wire n_4130;
wire n_4161;
wire n_4337;
wire n_2895;
wire n_2009;
wire n_4172;
wire n_692;
wire n_3403;
wire n_733;
wire n_1793;
wire n_2922;
wire n_3601;
wire n_3882;
wire n_1233;
wire n_1289;
wire n_2714;
wire n_2245;
wire n_487;
wire n_3055;
wire n_3092;
wire n_3492;
wire n_3895;
wire n_3966;
wire n_4369;
wire n_2068;
wire n_1107;
wire n_2866;
wire n_4454;
wire n_2457;
wire n_3294;
wire n_4119;
wire n_1014;
wire n_3734;
wire n_4331;
wire n_3686;
wire n_4520;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_3455;
wire n_4118;
wire n_4502;
wire n_882;
wire n_4503;
wire n_2176;
wire n_2072;
wire n_3649;
wire n_1354;
wire n_2821;
wire n_586;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_2459;
wire n_3746;
wire n_1111;
wire n_1713;
wire n_2971;
wire n_4375;
wire n_715;
wire n_3599;
wire n_2678;
wire n_1251;
wire n_3384;
wire n_3935;
wire n_1265;
wire n_4277;
wire n_2711;
wire n_3490;
wire n_4291;
wire n_4199;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_4319;
wire n_3369;
wire n_3419;
wire n_4441;
wire n_1982;
wire n_3872;
wire n_2878;
wire n_618;
wire n_3012;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_3772;
wire n_3875;
wire n_4478;
wire n_1167;
wire n_1359;
wire n_2818;
wire n_2428;
wire n_3581;
wire n_3794;
wire n_674;
wire n_3247;
wire n_871;
wire n_3069;
wire n_3921;
wire n_922;
wire n_1760;
wire n_1335;
wire n_1927;
wire n_2028;
wire n_3715;
wire n_1069;
wire n_2664;
wire n_2641;
wire n_1722;
wire n_1664;
wire n_612;
wire n_3022;
wire n_3052;
wire n_3725;
wire n_1165;
wire n_3933;
wire n_702;
wire n_2008;
wire n_2749;
wire n_3298;
wire n_2192;
wire n_3346;
wire n_2254;
wire n_2345;
wire n_3281;
wire n_1926;
wire n_1175;
wire n_3273;
wire n_4467;
wire n_2311;
wire n_1386;
wire n_1896;
wire n_2965;
wire n_1747;
wire n_3058;
wire n_1012;
wire n_3691;
wire n_4427;
wire n_780;
wire n_3861;
wire n_675;
wire n_2624;
wire n_4066;
wire n_903;
wire n_4485;
wire n_4146;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_3549;
wire n_2350;
wire n_2804;
wire n_2453;
wire n_4340;
wire n_3891;
wire n_2193;
wire n_3961;
wire n_2676;
wire n_1655;
wire n_3940;
wire n_4072;
wire n_4220;
wire n_928;
wire n_835;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_4371;
wire n_1157;
wire n_3453;
wire n_1750;
wire n_2994;
wire n_1462;
wire n_3410;
wire n_3153;
wire n_3428;
wire n_1188;
wire n_3689;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_3768;
wire n_2206;
wire n_604;
wire n_4004;
wire n_2810;
wire n_2967;
wire n_2319;
wire n_2519;
wire n_4043;
wire n_825;
wire n_4313;
wire n_728;
wire n_4353;
wire n_2916;
wire n_3415;
wire n_1063;
wire n_4292;
wire n_1588;
wire n_3785;
wire n_3942;
wire n_3997;
wire n_2963;
wire n_4041;
wire n_2947;
wire n_3918;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_3145;
wire n_4381;
wire n_1124;
wire n_1624;
wire n_3873;
wire n_3983;
wire n_515;
wire n_2096;
wire n_2980;
wire n_3968;
wire n_4466;
wire n_4418;
wire n_1965;
wire n_3538;
wire n_2476;
wire n_3280;
wire n_598;
wire n_3434;
wire n_4510;
wire n_696;
wire n_1515;
wire n_4473;
wire n_961;
wire n_4356;
wire n_3510;
wire n_437;
wire n_1082;
wire n_1317;
wire n_3227;
wire n_2733;
wire n_2824;
wire n_3289;
wire n_593;
wire n_4169;
wire n_514;
wire n_4055;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_3271;
wire n_950;
wire n_4362;
wire n_4248;
wire n_2812;
wire n_4518;
wire n_484;
wire n_2644;
wire n_2036;
wire n_3326;
wire n_2976;
wire n_2152;
wire n_1709;
wire n_3009;
wire n_2652;
wire n_4200;
wire n_3460;
wire n_2411;
wire n_3719;
wire n_2525;
wire n_1825;
wire n_4361;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_2657;
wire n_1792;
wire n_3827;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2921;
wire n_2409;
wire n_2082;
wire n_3519;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_3889;
wire n_2687;
wire n_3237;
wire n_949;
wire n_1630;
wire n_678;
wire n_2887;
wire n_3809;
wire n_3500;
wire n_3834;
wire n_4245;
wire n_4136;
wire n_3526;
wire n_3707;
wire n_2075;
wire n_4045;
wire n_2194;
wire n_2972;
wire n_2619;
wire n_3139;
wire n_3542;
wire n_4367;
wire n_2763;
wire n_2762;
wire n_4070;
wire n_1987;
wire n_3545;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_3578;
wire n_3885;
wire n_881;
wire n_2271;
wire n_1008;
wire n_3192;
wire n_760;
wire n_3993;
wire n_1546;
wire n_2583;
wire n_590;
wire n_4394;
wire n_4116;
wire n_2606;
wire n_4031;
wire n_2279;
wire n_1033;
wire n_462;
wire n_1052;
wire n_2794;
wire n_1296;
wire n_2663;
wire n_1990;
wire n_3352;
wire n_2391;
wire n_3805;
wire n_3073;
wire n_2431;
wire n_4018;
wire n_2987;
wire n_694;
wire n_2938;
wire n_2150;
wire n_1294;
wire n_2943;
wire n_1420;
wire n_3780;
wire n_3696;
wire n_4082;
wire n_2078;
wire n_1634;
wire n_3252;
wire n_2932;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_3253;
wire n_3337;
wire n_3450;
wire n_3209;
wire n_4002;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2658;
wire n_4329;
wire n_2665;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_3021;
wire n_1391;
wire n_449;
wire n_1523;
wire n_2558;
wire n_2750;
wire n_2775;
wire n_1208;
wire n_2893;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2954;
wire n_3477;
wire n_4288;
wire n_2728;
wire n_2349;
wire n_3128;
wire n_3763;
wire n_4289;
wire n_2684;
wire n_2712;
wire n_1072;
wire n_3146;
wire n_1527;
wire n_1495;
wire n_3733;
wire n_1438;
wire n_495;
wire n_815;
wire n_3953;
wire n_1100;
wire n_585;
wire n_1487;
wire n_4435;
wire n_2691;
wire n_3421;
wire n_840;
wire n_2913;
wire n_3614;
wire n_874;
wire n_4471;
wire n_1756;
wire n_3183;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_2705;
wire n_1969;
wire n_4019;
wire n_2690;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_3405;
wire n_1968;
wire n_898;
wire n_4385;
wire n_1952;
wire n_865;
wire n_3616;
wire n_4228;
wire n_2573;
wire n_3423;
wire n_2646;
wire n_4044;
wire n_3436;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_2535;
wire n_1880;
wire n_3366;
wire n_3442;
wire n_2631;
wire n_4191;
wire n_1364;
wire n_4322;
wire n_3078;
wire n_3644;
wire n_2436;
wire n_3937;
wire n_615;
wire n_2870;
wire n_1249;
wire n_2706;
wire n_3838;
wire n_4287;
wire n_1293;
wire n_2693;
wire n_4137;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_3159;
wire n_1451;
wire n_3941;
wire n_963;
wire n_639;
wire n_794;
wire n_2767;
wire n_3793;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_3727;
wire n_2707;
wire n_3240;
wire n_3576;
wire n_3789;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_3385;
wire n_4350;
wire n_3747;
wire n_3037;
wire n_1646;
wire n_3293;
wire n_872;
wire n_1139;
wire n_1714;
wire n_3922;
wire n_3179;
wire n_718;
wire n_1018;
wire n_3400;
wire n_3729;
wire n_1521;
wire n_1366;
wire n_4000;
wire n_4330;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2897;
wire n_3970;
wire n_4389;
wire n_4483;
wire n_4345;
wire n_2554;
wire n_996;
wire n_532;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_3522;
wire n_1513;
wire n_2747;
wire n_3924;
wire n_3171;
wire n_791;
wire n_1913;
wire n_4216;
wire n_3608;
wire n_510;
wire n_837;
wire n_4315;
wire n_2097;
wire n_2170;
wire n_3459;
wire n_4156;
wire n_3491;
wire n_4240;
wire n_1488;
wire n_2853;
wire n_1808;
wire n_3053;
wire n_948;
wire n_3358;
wire n_2517;
wire n_2713;
wire n_3499;
wire n_704;
wire n_2148;
wire n_4284;
wire n_4162;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_2765;
wire n_2861;
wire n_536;
wire n_3158;
wire n_1788;
wire n_3426;
wire n_1999;
wire n_2731;
wire n_622;
wire n_2590;
wire n_2643;
wire n_3150;
wire n_3018;
wire n_3353;
wire n_3782;
wire n_3975;
wire n_1469;
wire n_2060;
wire n_4479;
wire n_2608;
wire n_1838;
wire n_2638;
wire n_4011;
wire n_1835;
wire n_3470;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_3133;
wire n_2002;
wire n_581;
wire n_2650;
wire n_2138;
wire n_4098;
wire n_4021;
wire n_4476;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_3700;
wire n_2414;
wire n_1340;
wire n_3014;
wire n_3166;
wire n_1771;
wire n_2316;
wire n_4103;
wire n_4058;
wire n_3104;
wire n_631;
wire n_720;
wire n_3435;
wire n_842;
wire n_3148;
wire n_2262;
wire n_3348;
wire n_3229;
wire n_4022;
wire n_1707;
wire n_2239;
wire n_3082;
wire n_3611;
wire n_4310;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_2816;
wire n_797;
wire n_2689;
wire n_2933;
wire n_1473;
wire n_2717;
wire n_1723;
wire n_2191;
wire n_4481;
wire n_1246;
wire n_3799;
wire n_1878;
wire n_2574;
wire n_4475;
wire n_899;
wire n_738;
wire n_2012;
wire n_3497;
wire n_1304;
wire n_1035;
wire n_2842;
wire n_499;
wire n_2675;
wire n_1426;
wire n_3418;
wire n_705;
wire n_3580;
wire n_3775;
wire n_3537;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_4443;
wire n_3887;
wire n_1022;
wire n_614;
wire n_529;
wire n_2069;
wire n_2307;
wire n_3704;
wire n_2362;
wire n_684;
wire n_2539;
wire n_2667;
wire n_2698;
wire n_4123;
wire n_1431;
wire n_4096;
wire n_1615;
wire n_4114;
wire n_1474;
wire n_3312;
wire n_1571;
wire n_3835;
wire n_4286;
wire n_1809;
wire n_3119;
wire n_4280;
wire n_2948;
wire n_1577;
wire n_2958;
wire n_3735;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_4379;
wire n_3731;
wire n_1822;
wire n_486;
wire n_947;
wire n_2936;
wire n_3224;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_3173;
wire n_1992;
wire n_3677;
wire n_3631;
wire n_648;
wire n_657;
wire n_1049;
wire n_3223;
wire n_3996;
wire n_2771;
wire n_2445;
wire n_3020;
wire n_2057;
wire n_2103;
wire n_3140;
wire n_3185;
wire n_3770;
wire n_2605;
wire n_4097;
wire n_1666;
wire n_2772;
wire n_1505;
wire n_803;
wire n_4218;
wire n_4440;
wire n_4402;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_3557;
wire n_2610;
wire n_3654;
wire n_3129;
wire n_3880;
wire n_1849;
wire n_2848;
wire n_919;
wire n_3685;
wire n_2868;
wire n_3620;
wire n_1698;
wire n_478;
wire n_4100;
wire n_2231;
wire n_3609;
wire n_929;
wire n_3832;
wire n_2520;
wire n_1228;
wire n_4264;
wire n_4484;
wire n_2857;
wire n_446;
wire n_3693;
wire n_4497;
wire n_3788;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_4459;
wire n_1299;
wire n_2896;
wire n_526;
wire n_3837;
wire n_2718;
wire n_3019;
wire n_2639;
wire n_3471;
wire n_1183;
wire n_1436;
wire n_2898;
wire n_2251;
wire n_1384;
wire n_3674;
wire n_2494;
wire n_2959;
wire n_4079;
wire n_2501;
wire n_3325;
wire n_3203;
wire n_2238;
wire n_4085;
wire n_2368;
wire n_4464;
wire n_458;
wire n_1070;
wire n_2403;
wire n_3342;
wire n_2837;
wire n_4175;
wire n_998;
wire n_717;
wire n_3200;
wire n_1665;
wire n_4306;
wire n_3600;
wire n_3259;
wire n_2524;
wire n_3167;
wire n_1383;
wire n_2460;
wire n_4224;
wire n_3390;
wire n_3656;
wire n_4339;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_3324;
wire n_3593;
wire n_3341;
wire n_3867;
wire n_4455;
wire n_4453;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_3559;
wire n_4514;
wire n_3025;
wire n_2137;
wire n_1626;
wire n_3191;
wire n_4005;
wire n_1507;
wire n_2482;
wire n_552;
wire n_3810;
wire n_3546;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_3661;
wire n_3006;
wire n_4140;
wire n_2481;
wire n_3561;
wire n_912;
wire n_1857;
wire n_3987;
wire n_1519;
wire n_2144;
wire n_3056;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2424;
wire n_2296;
wire n_3201;
wire n_3633;
wire n_3447;
wire n_4487;
wire n_3971;
wire n_1142;
wire n_2849;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2682;
wire n_3032;
wire n_3103;
wire n_3638;
wire n_2589;
wire n_1395;
wire n_2199;
wire n_2110;
wire n_2661;
wire n_731;
wire n_2877;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_3393;
wire n_527;
wire n_811;
wire n_474;
wire n_1207;
wire n_2442;
wire n_683;
wire n_3627;
wire n_1791;
wire n_1368;
wire n_3451;
wire n_3480;
wire n_1418;
wire n_958;
wire n_1250;
wire n_3331;
wire n_1137;
wire n_3615;
wire n_1897;
wire n_2064;
wire n_880;
wire n_3087;
wire n_3072;
wire n_2053;
wire n_3612;
wire n_3505;
wire n_2259;
wire n_2121;
wire n_2773;
wire n_4222;
wire n_2545;
wire n_3577;
wire n_3540;
wire n_4401;
wire n_889;
wire n_3509;
wire n_2432;
wire n_2710;
wire n_4368;
wire n_1478;
wire n_589;
wire n_3606;
wire n_1310;
wire n_3142;
wire n_3598;
wire n_819;
wire n_2966;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_3591;
wire n_767;
wire n_3641;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2788;
wire n_2218;
wire n_477;
wire n_3196;
wire n_3590;
wire n_2435;
wire n_954;
wire n_4419;
wire n_864;
wire n_2504;
wire n_2797;
wire n_2623;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2892;
wire n_2132;
wire n_2063;
wire n_4120;
wire n_1382;
wire n_1534;
wire n_3892;
wire n_1564;
wire n_1736;
wire n_4069;
wire n_2748;
wire n_4053;
wire n_1483;
wire n_3848;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2860;
wire n_3327;
wire n_2330;
wire n_3441;
wire n_1457;
wire n_505;
wire n_1719;
wire n_3534;
wire n_3718;
wire n_1339;
wire n_1787;
wire n_2701;
wire n_2511;
wire n_537;
wire n_2475;
wire n_3964;
wire n_1993;
wire n_2281;
wire n_4167;
wire n_1427;
wire n_2416;
wire n_2745;
wire n_2617;
wire n_2776;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_3144;
wire n_3705;
wire n_3211;
wire n_3244;
wire n_596;
wire n_3909;
wire n_3944;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_556;
wire n_2784;
wire n_2209;
wire n_2301;
wire n_3582;
wire n_3605;
wire n_3287;
wire n_4223;
wire n_2387;
wire n_3322;
wire n_1755;
wire n_4431;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_3270;
wire n_4387;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2846;
wire n_2464;
wire n_3265;
wire n_1125;
wire n_3755;
wire n_4042;
wire n_970;
wire n_3306;
wire n_2488;
wire n_3640;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_3481;
wire n_2237;
wire n_3026;
wire n_441;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_3090;
wire n_4299;
wire n_444;
wire n_3033;
wire n_3724;
wire n_1252;
wire n_1784;
wire n_3311;
wire n_3571;
wire n_1223;
wire n_3913;
wire n_4276;
wire n_511;
wire n_2990;
wire n_3847;
wire n_1286;
wire n_1775;
wire n_2115;
wire n_1773;
wire n_4430;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_3302;
wire n_2374;
wire n_1681;
wire n_4348;
wire n_520;
wire n_1093;
wire n_4428;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2929;
wire n_2780;
wire n_3323;
wire n_3364;
wire n_3226;
wire n_4020;
wire n_4176;
wire n_4489;
wire n_2596;
wire n_2274;
wire n_3163;
wire n_775;
wire n_4404;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_3407;
wire n_518;
wire n_1531;
wire n_2828;
wire n_1185;
wire n_3856;
wire n_453;
wire n_4236;
wire n_3425;
wire n_2384;
wire n_3894;
wire n_4261;
wire n_4204;
wire n_1745;
wire n_914;
wire n_759;
wire n_3479;
wire n_3127;
wire n_2724;
wire n_1831;
wire n_4496;
wire n_2585;
wire n_2621;
wire n_3623;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_4063;
wire n_1625;
wire n_3986;
wire n_4237;
wire n_2601;
wire n_2160;
wire n_3454;
wire n_4513;
wire n_1453;
wire n_2146;
wire n_4006;
wire n_2502;
wire n_2131;
wire n_488;
wire n_2226;
wire n_2801;
wire n_3646;
wire n_497;
wire n_2920;
wire n_4015;
wire n_773;
wire n_3547;
wire n_1901;
wire n_3869;
wire n_920;
wire n_1374;
wire n_2556;
wire n_2648;
wire n_3212;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_2754;
wire n_1224;
wire n_2783;
wire n_3753;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_3188;
wire n_3742;
wire n_4410;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_2889;
wire n_3243;
wire n_3683;
wire n_4056;
wire n_1617;
wire n_4034;
wire n_3260;
wire n_3370;
wire n_3386;
wire n_3816;
wire n_3960;
wire n_1470;
wire n_2550;
wire n_463;
wire n_3093;
wire n_3175;
wire n_4411;
wire n_3214;
wire n_1243;
wire n_3736;
wire n_848;
wire n_2732;
wire n_2928;
wire n_4206;
wire n_4448;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_2000;
wire n_1917;
wire n_3862;
wire n_4267;
wire n_1580;
wire n_2227;
wire n_4247;
wire n_2270;
wire n_2822;
wire n_1425;
wire n_3169;
wire n_4180;
wire n_3205;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_3284;
wire n_983;
wire n_3109;
wire n_2023;
wire n_3354;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_496;
wire n_2720;
wire n_3126;
wire n_2159;
wire n_906;
wire n_1390;
wire n_2289;
wire n_2315;
wire n_1077;
wire n_1733;
wire n_688;
wire n_1419;
wire n_2863;
wire n_3299;
wire n_3663;
wire n_4386;
wire n_2955;
wire n_2995;
wire n_1731;
wire n_2158;
wire n_3360;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_3051;
wire n_1437;
wire n_4438;
wire n_2135;
wire n_3956;
wire n_3367;
wire n_1645;
wire n_1832;
wire n_4001;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2859;
wire n_2202;
wire n_858;
wire n_2049;
wire n_4149;
wire n_1331;
wire n_613;
wire n_736;
wire n_2627;
wire n_4355;
wire n_501;
wire n_956;
wire n_960;
wire n_2276;
wire n_3234;
wire n_4422;
wire n_3917;
wire n_663;
wire n_856;
wire n_2803;
wire n_2100;
wire n_3314;
wire n_3525;
wire n_2993;
wire n_778;
wire n_1668;
wire n_2777;
wire n_1134;
wire n_3016;
wire n_3566;
wire n_3688;
wire n_3004;
wire n_3202;
wire n_2830;
wire n_2781;
wire n_3220;
wire n_4003;
wire n_4030;
wire n_1129;
wire n_3870;
wire n_4126;
wire n_554;
wire n_602;
wire n_1696;
wire n_2829;
wire n_2181;
wire n_1594;
wire n_1995;
wire n_3751;
wire n_664;
wire n_1869;
wire n_2911;
wire n_3625;
wire n_3804;
wire n_1764;
wire n_4207;
wire n_1429;
wire n_2826;
wire n_1610;
wire n_3084;
wire n_3429;
wire n_4113;
wire n_1889;
wire n_2379;
wire n_435;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_4470;
wire n_587;
wire n_3466;
wire n_3554;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_3901;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_3749;
wire n_1635;
wire n_2942;
wire n_4014;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_4252;
wire n_4357;
wire n_4067;
wire n_607;
wire n_1551;
wire n_4028;
wire n_4054;
wire n_4509;
wire n_2448;
wire n_1103;
wire n_2875;
wire n_3907;
wire n_2555;
wire n_4048;
wire n_4444;
wire n_3338;
wire n_4217;
wire n_3586;
wire n_3462;
wire n_3756;
wire n_2219;
wire n_1203;
wire n_3653;
wire n_3636;
wire n_2851;
wire n_3406;
wire n_820;
wire n_2327;
wire n_951;
wire n_4374;
wire n_2201;
wire n_725;
wire n_952;
wire n_3919;
wire n_999;
wire n_1254;
wire n_2841;
wire n_3349;
wire n_2420;
wire n_3722;
wire n_4400;
wire n_2984;
wire n_575;
wire n_994;
wire n_2263;
wire n_3539;
wire n_3291;
wire n_4399;
wire n_2304;
wire n_4024;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2983;
wire n_2240;
wire n_2278;
wire n_2656;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_3113;
wire n_3194;
wire n_3276;
wire n_1934;
wire n_3250;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_3981;
wire n_4214;
wire n_1728;
wire n_3973;
wire n_557;
wire n_2756;
wire n_3572;
wire n_1871;
wire n_3448;
wire n_4338;
wire n_617;
wire n_3886;
wire n_845;
wire n_807;
wire n_2924;
wire n_1036;
wire n_3595;
wire n_1138;
wire n_3414;
wire n_1661;
wire n_1275;
wire n_2884;
wire n_485;
wire n_1549;
wire n_4420;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_3637;
wire n_3120;
wire n_1468;
wire n_3991;
wire n_2855;
wire n_3651;
wire n_1859;
wire n_2102;
wire n_3516;
wire n_2563;
wire n_3797;
wire n_3926;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_3449;
wire n_1718;
wire n_1749;
wire n_3474;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_4405;
wire n_610;
wire n_4304;
wire n_4234;
wire n_4413;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_4488;
wire n_4101;
wire n_3548;
wire n_3767;
wire n_1024;
wire n_3864;
wire n_4036;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_3670;
wire n_3550;
wire n_3974;
wire n_2052;
wire n_1847;
wire n_3634;
wire n_2302;
wire n_517;
wire n_4211;
wire n_4182;
wire n_1667;
wire n_667;
wire n_1206;
wire n_3230;
wire n_4016;
wire n_621;
wire n_1037;
wire n_1397;
wire n_3268;
wire n_3236;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_3592;
wire n_468;
wire n_2755;
wire n_3141;
wire n_923;
wire n_504;
wire n_1409;
wire n_4230;
wire n_1841;
wire n_3839;
wire n_2637;
wire n_2823;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_3967;
wire n_1503;
wire n_3112;
wire n_2819;
wire n_4328;
wire n_3195;
wire n_466;
wire n_2526;
wire n_3041;
wire n_4274;
wire n_2423;
wire n_1057;
wire n_3277;
wire n_3108;
wire n_2548;
wire n_603;
wire n_991;
wire n_2785;
wire n_1657;
wire n_4270;
wire n_4189;
wire n_4151;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_3817;
wire n_3417;
wire n_2636;
wire n_3131;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_3730;
wire n_1298;
wire n_4124;
wire n_3659;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_3399;
wire n_4397;
wire n_2088;
wire n_3635;
wire n_1611;
wire n_785;
wire n_4155;
wire n_2740;
wire n_746;
wire n_4238;
wire n_609;
wire n_1601;
wire n_3011;
wire n_1960;
wire n_2694;
wire n_2061;
wire n_3416;
wire n_3648;
wire n_1686;
wire n_3498;
wire n_2757;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_3042;
wire n_3213;
wire n_4333;
wire n_3820;
wire n_2309;
wire n_2900;
wire n_2957;
wire n_2607;
wire n_1740;
wire n_2737;
wire n_3994;
wire n_1497;
wire n_2890;
wire n_1168;
wire n_4472;
wire n_1216;
wire n_1943;
wire n_3228;
wire n_3249;
wire n_1320;
wire n_2716;
wire n_3081;
wire n_3657;
wire n_2452;
wire n_1430;
wire n_3650;
wire n_1316;
wire n_1287;
wire n_2722;
wire n_1452;
wire n_2854;
wire n_3672;
wire n_3010;
wire n_2499;
wire n_4152;
wire n_3533;
wire n_3043;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_3464;
wire n_1694;
wire n_1535;
wire n_3137;
wire n_3382;
wire n_4406;
wire n_2486;
wire n_3132;
wire n_3560;
wire n_3723;
wire n_2571;
wire n_3138;
wire n_1596;
wire n_3177;
wire n_1190;
wire n_1734;
wire n_3172;
wire n_4380;
wire n_2902;
wire n_3217;
wire n_1983;
wire n_1938;
wire n_4398;
wire n_2498;
wire n_4219;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_3238;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_3529;
wire n_2235;
wire n_4193;
wire n_3570;
wire n_3394;
wire n_2988;
wire n_3136;
wire n_1350;
wire n_1673;
wire n_3828;
wire n_2232;
wire n_1715;
wire n_3536;
wire n_4192;
wire n_4109;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2894;
wire n_3424;
wire n_3957;
wire n_4131;
wire n_2790;
wire n_4038;
wire n_2037;
wire n_2808;
wire n_3710;
wire n_4159;
wire n_4195;
wire n_3784;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_490;
wire n_3594;
wire n_809;
wire n_1043;
wire n_3819;
wire n_4090;
wire n_3040;
wire n_1797;
wire n_3279;
wire n_1608;
wire n_4165;
wire n_986;
wire n_2305;
wire n_2373;
wire n_1472;
wire n_2120;
wire n_2050;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_3628;
wire n_4144;
wire n_1870;
wire n_2964;
wire n_4174;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_460;
wire n_2169;
wire n_3485;
wire n_4077;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_3402;
wire n_1491;
wire n_2187;
wire n_3501;
wire n_662;
wire n_3475;
wire n_4442;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_3905;
wire n_4434;
wire n_450;
wire n_3262;
wire n_3544;
wire n_4150;
wire n_2904;
wire n_4008;
wire n_2244;
wire n_4290;
wire n_3013;
wire n_3356;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_2789;
wire n_3105;
wire n_3210;
wire n_2872;
wire n_937;
wire n_2257;
wire n_3692;
wire n_4515;
wire n_3845;
wire n_1682;
wire n_2017;
wire n_4516;
wire n_1828;
wire n_1695;
wire n_2046;
wire n_2272;
wire n_2699;
wire n_2200;
wire n_3029;
wire n_4258;
wire n_650;
wire n_3597;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_2760;
wire n_2704;
wire n_3329;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_2738;
wire n_972;
wire n_1405;
wire n_2376;
wire n_3826;
wire n_1406;
wire n_456;
wire n_3790;
wire n_3878;
wire n_2766;
wire n_1332;
wire n_2670;
wire n_2700;
wire n_4323;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_565;
wire n_3134;
wire n_3647;
wire n_1569;
wire n_3681;
wire n_936;
wire n_3045;
wire n_3115;
wire n_1883;
wire n_3821;
wire n_1288;
wire n_4300;
wire n_3318;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_3278;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2970;
wire n_3676;
wire n_2882;
wire n_3666;
wire n_3675;
wire n_4017;
wire n_4260;
wire n_3320;
wire n_2541;
wire n_654;
wire n_2940;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_3050;
wire n_3350;
wire n_2782;
wire n_3977;
wire n_1974;
wire n_3988;
wire n_4122;
wire n_2673;
wire n_2456;
wire n_1720;
wire n_3476;
wire n_2527;
wire n_934;
wire n_482;
wire n_1637;
wire n_2635;
wire n_3307;
wire n_3439;
wire n_3588;
wire n_1407;
wire n_1795;
wire n_2768;
wire n_4209;
wire n_4279;
wire n_2871;
wire n_4135;
wire n_2688;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_3858;
wire n_4321;
wire n_1489;
wire n_4183;
wire n_4298;
wire n_2314;
wire n_3502;
wire n_942;
wire n_3003;
wire n_2798;
wire n_2852;
wire n_1524;
wire n_4128;
wire n_543;
wire n_2229;
wire n_1964;
wire n_4133;
wire n_2288;
wire n_1920;
wire n_2753;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_3292;
wire n_1545;
wire n_4145;
wire n_2007;
wire n_3121;
wire n_2039;
wire n_3388;
wire n_4271;
wire n_1946;
wire n_1355;
wire n_4181;
wire n_1225;
wire n_3184;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_4040;
wire n_804;
wire n_4461;
wire n_464;
wire n_1846;
wire n_3437;
wire n_3245;
wire n_3075;
wire n_2406;
wire n_4111;
wire n_533;
wire n_2390;
wire n_4007;
wire n_806;
wire n_3712;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_584;
wire n_2141;
wire n_2562;
wire n_2642;
wire n_4312;
wire n_1343;
wire n_1522;
wire n_4239;
wire n_2734;
wire n_548;
wire n_1782;
wire n_2383;
wire n_4184;
wire n_2626;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_4037;
wire n_523;
wire n_1319;
wire n_707;
wire n_2986;
wire n_1900;
wire n_3930;
wire n_3246;
wire n_1548;
wire n_799;
wire n_3381;
wire n_3044;
wire n_3562;
wire n_2973;
wire n_1155;
wire n_2536;
wire n_3915;
wire n_2196;
wire n_2629;
wire n_3665;
wire n_1633;
wire n_2195;
wire n_3208;
wire n_2809;
wire n_3007;
wire n_787;
wire n_2172;
wire n_3528;
wire n_3489;
wire n_4343;
wire n_2835;
wire n_1416;
wire n_1528;
wire n_2820;
wire n_2293;
wire n_1146;
wire n_3698;
wire n_2021;
wire n_3355;
wire n_2454;
wire n_2114;
wire n_3074;
wire n_3174;
wire n_1086;
wire n_1066;
wire n_3102;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_4215;
wire n_1282;
wire n_2561;
wire n_550;
wire n_3321;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_2727;
wire n_2962;
wire n_3377;
wire n_2939;
wire n_560;
wire n_1906;
wire n_1484;
wire n_2992;
wire n_3305;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_2533;
wire n_3157;
wire n_3530;
wire n_4185;
wire n_1758;
wire n_3221;
wire n_3267;
wire n_3752;
wire n_2283;
wire n_2869;
wire n_2422;
wire n_1925;
wire n_4378;
wire n_4407;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_3457;
wire n_1229;
wire n_2759;
wire n_3517;
wire n_2945;
wire n_3061;
wire n_3893;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_3762;
wire n_3469;
wire n_3932;
wire n_2266;
wire n_2960;
wire n_3958;
wire n_3005;
wire n_3985;
wire n_2427;
wire n_3151;
wire n_3411;
wire n_1029;
wire n_4196;
wire n_3779;
wire n_1447;
wire n_4519;
wire n_2388;
wire n_3984;
wire n_2056;
wire n_790;
wire n_2611;
wire n_2901;
wire n_3258;
wire n_4358;
wire n_1706;
wire n_4242;
wire n_3389;
wire n_1498;
wire n_3143;
wire n_2653;
wire n_2417;
wire n_4232;
wire n_4190;
wire n_3000;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2680;
wire n_4052;
wire n_2246;
wire n_1047;
wire n_3149;
wire n_3375;
wire n_3899;
wire n_4469;
wire n_3558;
wire n_4084;
wire n_1984;
wire n_3365;
wire n_2236;
wire n_1385;
wire n_3713;
wire n_431;
wire n_3379;
wire n_4326;
wire n_3156;
wire n_459;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_2834;
wire n_3207;
wire n_502;
wire n_2668;
wire n_672;
wire n_4424;
wire n_2441;
wire n_1257;
wire n_3008;
wire n_1751;
wire n_3401;
wire n_2840;
wire n_3197;
wire n_3242;
wire n_3939;
wire n_1375;
wire n_1941;
wire n_3483;
wire n_3613;
wire n_3972;
wire n_4153;
wire n_2128;
wire n_655;
wire n_706;
wire n_1045;
wire n_1794;
wire n_786;
wire n_1650;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_3743;
wire n_3855;
wire n_1872;
wire n_3091;
wire n_4317;
wire n_834;
wire n_4493;
wire n_2695;
wire n_4035;
wire n_3818;
wire n_4269;
wire n_743;
wire n_766;
wire n_3124;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_4088;
wire n_1949;
wire n_3398;
wire n_3761;
wire n_3759;
wire n_545;
wire n_3524;
wire n_2671;
wire n_489;
wire n_2761;
wire n_2885;
wire n_2888;
wire n_2715;
wire n_2793;
wire n_1804;
wire n_2923;
wire n_3776;
wire n_3711;
wire n_4235;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_4301;
wire n_3511;
wire n_2054;
wire n_4143;
wire n_4170;
wire n_729;
wire n_876;
wire n_774;
wire n_3744;
wire n_3642;
wire n_2845;
wire n_1337;
wire n_3097;
wire n_660;
wire n_2062;
wire n_2041;
wire n_2975;
wire n_438;
wire n_1477;
wire n_4421;
wire n_1360;
wire n_2839;
wire n_1860;
wire n_2856;
wire n_1904;
wire n_2874;
wire n_1200;
wire n_4498;
wire n_2070;
wire n_2588;
wire n_479;
wire n_3814;
wire n_1607;
wire n_3781;
wire n_1353;
wire n_1908;
wire n_1777;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2944;
wire n_2614;
wire n_2126;
wire n_3831;
wire n_869;
wire n_1154;
wire n_4492;
wire n_3308;
wire n_1113;
wire n_1600;
wire n_2833;
wire n_2253;
wire n_2758;
wire n_3843;
wire n_2366;
wire n_646;
wire n_528;
wire n_1098;
wire n_3694;
wire n_2937;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_4423;
wire n_3687;
wire n_2216;
wire n_3589;
wire n_2210;
wire n_3602;
wire n_897;
wire n_846;
wire n_3300;
wire n_2978;
wire n_2066;
wire n_3543;
wire n_841;
wire n_1476;
wire n_3621;
wire n_2516;
wire n_3391;
wire n_4376;
wire n_1001;
wire n_508;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_2903;
wire n_3777;
wire n_2827;
wire n_1177;
wire n_3216;
wire n_3458;
wire n_3515;
wire n_1150;
wire n_4203;
wire n_3808;
wire n_3190;
wire n_4505;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_4365;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_2951;
wire n_1118;
wire n_1076;
wire n_4512;
wire n_2949;
wire n_3726;
wire n_1807;
wire n_1007;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_855;
wire n_1592;
wire n_1759;
wire n_2719;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_3758;
wire n_1879;
wire n_853;
wire n_440;
wire n_695;
wire n_3806;
wire n_4081;
wire n_1542;
wire n_2587;
wire n_3199;
wire n_2931;
wire n_875;
wire n_680;
wire n_4462;
wire n_3339;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_3866;
wire n_3787;
wire n_1256;
wire n_3585;
wire n_671;
wire n_3565;
wire n_1953;
wire n_4450;
wire n_933;
wire n_740;
wire n_703;
wire n_3343;
wire n_3303;
wire n_978;
wire n_4157;
wire n_2752;
wire n_4324;
wire n_3135;
wire n_4173;
wire n_1976;
wire n_4382;
wire n_4229;
wire n_2905;
wire n_1291;
wire n_1217;
wire n_3990;
wire n_751;
wire n_749;
wire n_3865;
wire n_1824;
wire n_3954;
wire n_1628;
wire n_4073;
wire n_1324;
wire n_3890;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_3629;
wire n_1435;
wire n_3920;
wire n_969;
wire n_988;
wire n_2140;
wire n_3503;
wire n_3160;
wire n_1065;
wire n_2796;
wire n_3255;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_568;
wire n_3658;
wire n_1516;
wire n_1536;
wire n_3846;
wire n_2163;
wire n_2186;
wire n_3512;
wire n_2029;
wire n_2815;
wire n_1204;
wire n_3951;
wire n_3034;
wire n_823;
wire n_4408;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_4439;
wire n_3569;
wire n_1327;
wire n_1326;
wire n_739;
wire n_955;
wire n_3874;
wire n_1379;
wire n_2528;
wire n_2814;
wire n_2787;
wire n_1338;
wire n_1097;
wire n_2969;
wire n_2395;
wire n_935;
wire n_3027;
wire n_781;
wire n_789;
wire n_1554;
wire n_3231;
wire n_4083;
wire n_4494;
wire n_1130;
wire n_3083;
wire n_4212;
wire n_2979;
wire n_1810;
wire n_2953;
wire n_573;
wire n_769;
wire n_2380;
wire n_676;
wire n_4295;
wire n_1120;
wire n_832;
wire n_1583;
wire n_4480;
wire n_3049;
wire n_1730;
wire n_2295;
wire n_555;
wire n_814;
wire n_2746;
wire n_2946;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_3430;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_4225;
wire n_4171;
wire n_2048;
wire n_3652;
wire n_3830;
wire n_3679;
wire n_2005;
wire n_747;
wire n_3541;
wire n_2565;
wire n_4023;
wire n_1389;
wire n_1105;
wire n_3117;
wire n_721;
wire n_1461;
wire n_742;
wire n_3432;
wire n_535;
wire n_691;
wire n_3617;
wire n_2076;
wire n_2736;
wire n_2883;
wire n_3583;
wire n_3860;
wire n_1408;
wire n_3851;
wire n_3567;
wire n_1196;
wire n_4282;
wire n_1598;
wire n_3493;
wire n_4344;
wire n_2935;
wire n_4046;
wire n_3807;
wire n_863;
wire n_3015;
wire n_2175;
wire n_601;
wire n_2182;
wire n_3774;
wire n_2910;
wire n_1283;
wire n_2385;
wire n_4112;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1848;
wire n_763;
wire n_1147;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_3057;
wire n_3154;
wire n_3701;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_3473;
wire n_895;
wire n_866;
wire n_1227;
wire n_2485;
wire n_2450;
wire n_3739;
wire n_2284;
wire n_3898;
wire n_4432;
wire n_3520;
wire n_2566;
wire n_2287;
wire n_452;
wire n_4352;
wire n_744;
wire n_971;
wire n_4391;
wire n_4416;
wire n_2702;
wire n_3241;
wire n_946;
wire n_2906;
wire n_761;
wire n_1303;
wire n_2769;
wire n_4342;
wire n_4465;
wire n_3622;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_3778;
wire n_4095;
wire n_2438;
wire n_2914;
wire n_1392;
wire n_4495;
wire n_1173;
wire n_1924;
wire n_525;
wire n_2463;
wire n_3363;
wire n_2881;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1702;
wire n_1570;
wire n_1219;
wire n_3551;
wire n_4436;
wire n_3064;
wire n_1780;
wire n_3100;
wire n_3897;
wire n_3721;
wire n_1689;
wire n_2180;
wire n_3372;
wire n_2858;
wire n_3062;
wire n_2679;
wire n_1174;
wire n_3573;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_4106;
wire n_795;
wire n_1501;
wire n_3604;
wire n_1221;
wire n_3334;
wire n_4373;
wire n_4027;
wire n_1245;
wire n_838;
wire n_3215;
wire n_3969;
wire n_3336;
wire n_647;
wire n_4160;
wire n_4231;
wire n_844;
wire n_448;
wire n_2952;
wire n_1017;
wire n_3068;
wire n_3853;
wire n_2117;
wire n_2234;
wire n_4256;
wire n_2779;
wire n_2685;
wire n_3823;
wire n_1083;
wire n_445;
wire n_3553;
wire n_1561;
wire n_4384;
wire n_2741;
wire n_3114;
wire n_930;
wire n_888;
wire n_2465;
wire n_1112;
wire n_2275;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_3811;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2255;
wire n_2112;
wire n_1464;
wire n_1737;
wire n_653;
wire n_2430;
wire n_1414;
wire n_3486;
wire n_4086;
wire n_752;
wire n_908;
wire n_2721;
wire n_2649;
wire n_944;
wire n_4335;
wire n_3556;
wire n_2034;
wire n_576;
wire n_1028;
wire n_3836;
wire n_2106;
wire n_472;
wire n_2862;
wire n_2265;
wire n_2615;
wire n_2683;
wire n_1922;
wire n_563;
wire n_4068;
wire n_2032;
wire n_4409;
wire n_2744;
wire n_4309;
wire n_4363;
wire n_1011;
wire n_2474;
wire n_3703;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_2437;
wire n_839;
wire n_2743;
wire n_3962;
wire n_1973;
wire n_708;
wire n_3181;
wire n_2267;
wire n_3456;
wire n_3035;
wire n_668;
wire n_4166;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_3699;
wire n_4243;
wire n_3204;
wire n_1104;
wire n_854;
wire n_1058;
wire n_3378;
wire n_4025;
wire n_2312;
wire n_498;
wire n_3404;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_3362;
wire n_3745;
wire n_4059;
wire n_1509;
wire n_4188;
wire n_3328;
wire n_1693;
wire n_2934;
wire n_3667;
wire n_3290;
wire n_4121;
wire n_1109;
wire n_3523;
wire n_2222;
wire n_712;
wire n_3256;
wire n_1276;
wire n_3868;
wire n_3802;
wire n_3176;
wire n_3309;
wire n_3671;
wire n_2015;
wire n_2118;
wire n_4142;
wire n_2466;
wire n_2111;
wire n_3982;
wire n_4266;
wire n_2915;
wire n_2530;
wire n_1148;
wire n_2505;
wire n_2188;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2802;
wire n_3796;
wire n_2999;
wire n_4115;
wire n_3840;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_3643;
wire n_3697;
wire n_771;
wire n_1584;
wire n_2425;
wire n_470;
wire n_475;
wire n_924;
wire n_3461;
wire n_3408;
wire n_1582;
wire n_492;
wire n_3680;
wire n_4265;
wire n_2318;
wire n_3286;
wire n_4012;
wire n_2408;
wire n_4246;
wire n_1149;
wire n_3170;
wire n_3513;
wire n_3468;
wire n_3690;
wire n_1184;
wire n_3645;
wire n_2483;
wire n_2950;
wire n_719;
wire n_1972;
wire n_3060;
wire n_3304;
wire n_3682;
wire n_2592;
wire n_3771;
wire n_1525;
wire n_4383;
wire n_4491;
wire n_3098;
wire n_3995;
wire n_4076;
wire n_2594;
wire n_455;
wire n_2666;
wire n_4105;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_4244;
wire n_4486;
wire n_1816;
wire n_4064;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_4049;
wire n_829;
wire n_1362;
wire n_1156;
wire n_4259;
wire n_3123;
wire n_984;
wire n_2600;
wire n_3380;
wire n_1829;
wire n_503;
wire n_2035;
wire n_3508;
wire n_3024;
wire n_1450;
wire n_1638;
wire n_3422;
wire n_868;
wire n_3038;
wire n_570;
wire n_859;
wire n_2033;
wire n_3086;
wire n_735;
wire n_4104;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_3285;
wire n_519;
wire n_4208;
wire n_2523;
wire n_469;
wire n_1218;
wire n_2413;
wire n_500;
wire n_3769;
wire n_1482;
wire n_3361;
wire n_981;
wire n_3596;
wire n_714;
wire n_3478;
wire n_3936;
wire n_1349;
wire n_4346;
wire n_4351;
wire n_4089;
wire n_1144;
wire n_2071;
wire n_3669;
wire n_3863;
wire n_3219;
wire n_2429;
wire n_3130;
wire n_3702;
wire n_985;
wire n_4316;
wire n_2233;
wire n_2440;
wire n_2723;
wire n_481;
wire n_3521;
wire n_3233;
wire n_997;
wire n_1710;
wire n_2800;
wire n_2161;
wire n_3496;
wire n_4437;
wire n_1301;
wire n_2805;
wire n_802;
wire n_561;
wire n_3310;
wire n_980;
wire n_2681;
wire n_1306;
wire n_3264;
wire n_2010;
wire n_4390;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_3096;
wire n_2360;
wire n_3764;
wire n_2047;
wire n_4061;
wire n_2651;
wire n_2095;
wire n_3239;
wire n_1609;
wire n_2174;
wire n_3161;
wire n_2799;
wire n_436;
wire n_4075;
wire n_3344;
wire n_2334;
wire n_3902;
wire n_4062;
wire n_3881;
wire n_3295;
wire n_3947;
wire n_1244;
wire n_1685;
wire n_4396;
wire n_4508;
wire n_1763;
wire n_1998;
wire n_3066;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_2844;
wire n_3101;
wire n_3989;
wire n_756;
wire n_2478;
wire n_1619;
wire n_2303;
wire n_1981;
wire n_2285;
wire n_4233;
wire n_4451;
wire n_1606;
wire n_4332;
wire n_810;
wire n_4108;
wire n_1133;
wire n_4460;
wire n_635;
wire n_1194;
wire n_3374;
wire n_4429;
wire n_4506;
wire n_3786;
wire n_3841;
wire n_2742;
wire n_2640;
wire n_3695;
wire n_4254;
wire n_1051;
wire n_3976;
wire n_4051;
wire n_1552;
wire n_2918;
wire n_583;
wire n_3288;
wire n_1996;
wire n_3563;
wire n_3992;
wire n_2367;
wire n_4307;
wire n_3876;
wire n_2867;
wire n_3198;
wire n_1039;
wire n_1442;
wire n_3495;
wire n_2726;
wire n_1034;
wire n_2043;
wire n_4303;
wire n_1480;
wire n_3125;
wire n_1158;
wire n_2909;
wire n_2248;
wire n_754;
wire n_4293;
wire n_941;
wire n_3552;
wire n_975;
wire n_3206;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_553;
wire n_849;
wire n_2662;
wire n_3147;
wire n_3116;
wire n_3383;
wire n_3709;
wire n_753;
wire n_3925;
wire n_4091;
wire n_1753;
wire n_3095;
wire n_3180;
wire n_3738;
wire n_3359;
wire n_2795;
wire n_3472;
wire n_2471;
wire n_4186;
wire n_467;
wire n_3187;
wire n_2540;
wire n_4412;
wire n_973;
wire n_2807;
wire n_1921;
wire n_3218;
wire n_3610;
wire n_3618;
wire n_3330;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2217;
wire n_2197;
wire n_582;
wire n_2065;
wire n_2879;
wire n_861;
wire n_3717;
wire n_857;
wire n_967;
wire n_4148;
wire n_571;
wire n_2461;
wire n_2215;
wire n_2001;
wire n_2107;
wire n_4341;
wire n_1884;
wire n_2040;
wire n_679;
wire n_4057;
wire n_2968;
wire n_4336;
wire n_4201;
wire n_633;
wire n_1170;
wire n_1629;
wire n_2221;
wire n_665;
wire n_588;
wire n_4263;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_3555;
wire n_1010;
wire n_3444;
wire n_4210;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_3059;
wire n_1166;
wire n_2038;
wire n_4447;
wire n_812;
wire n_2891;
wire n_1131;
wire n_2634;
wire n_1761;
wire n_2709;
wire n_3155;
wire n_3445;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_3110;
wire n_1890;
wire n_1632;
wire n_3017;
wire n_3955;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_3903;
wire n_730;
wire n_1311;
wire n_4132;
wire n_3945;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2697;
wire n_3235;
wire n_3854;
wire n_2308;
wire n_4205;
wire n_2162;
wire n_3908;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_3467;
wire n_3001;
wire n_3587;
wire n_1089;
wire n_4278;
wire n_1887;
wire n_1587;
wire n_3916;
wire n_3527;
wire n_3795;
wire n_2512;
wire n_3950;
wire n_3433;
wire n_3852;
wire n_1365;
wire n_4138;
wire n_4463;
wire n_1417;
wire n_1242;
wire n_2086;
wire n_2185;
wire n_2927;
wire n_3673;
wire n_1836;
wire n_3833;
wire n_4281;
wire n_3815;
wire n_2774;
wire n_3896;
wire n_3039;
wire n_681;
wire n_1226;
wire n_3740;
wire n_3162;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_3094;
wire n_2899;
wire n_3333;
wire n_3274;
wire n_3186;
wire n_640;
wire n_1322;
wire n_4129;
wire n_4457;
wire n_965;
wire n_1899;
wire n_1428;
wire n_4093;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_434;
wire n_1059;
wire n_1197;
wire n_3065;
wire n_3965;
wire n_2632;
wire n_2579;
wire n_722;
wire n_4500;
wire n_862;
wire n_2105;
wire n_3079;
wire n_4360;
wire n_2098;
wire n_3085;
wire n_4433;
wire n_540;
wire n_1423;
wire n_2813;
wire n_1935;
wire n_3584;
wire n_4039;
wire n_3387;
wire n_2027;
wire n_457;
wire n_3070;
wire n_3800;
wire n_2223;
wire n_2091;
wire n_3263;
wire n_3431;
wire n_4197;
wire n_3420;
wire n_2991;
wire n_1915;
wire n_629;
wire n_1621;
wire n_4275;
wire n_4482;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_4283;
wire n_900;
wire n_3504;
wire n_4194;
wire n_1449;
wire n_4426;
wire n_531;
wire n_827;
wire n_2912;
wire n_4272;
wire n_2659;
wire n_2930;
wire n_4425;
wire n_1025;
wire n_3409;
wire n_2419;
wire n_3111;
wire n_2116;
wire n_4449;
wire n_2320;
wire n_1885;
wire n_2677;
wire n_1013;
wire n_3182;
wire n_1259;
wire n_3054;
wire n_3283;
wire n_2183;
wire n_3002;
wire n_1538;
wire n_649;
wire n_1742;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_360),
.Y(n_430)
);

INVx2_ASAP7_75t_SL g431 ( 
.A(n_202),
.Y(n_431)
);

BUFx2_ASAP7_75t_L g432 ( 
.A(n_151),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_291),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_43),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_290),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_405),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_50),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_92),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_131),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_68),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_249),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_300),
.Y(n_442)
);

BUFx6f_ASAP7_75t_L g443 ( 
.A(n_327),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_366),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g445 ( 
.A(n_319),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_323),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_174),
.Y(n_447)
);

CKINVDCx5p33_ASAP7_75t_R g448 ( 
.A(n_418),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_150),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_18),
.Y(n_450)
);

CKINVDCx16_ASAP7_75t_R g451 ( 
.A(n_20),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_63),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_208),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_343),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_209),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_106),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_386),
.Y(n_457)
);

INVx1_ASAP7_75t_SL g458 ( 
.A(n_280),
.Y(n_458)
);

BUFx5_ASAP7_75t_L g459 ( 
.A(n_391),
.Y(n_459)
);

BUFx3_ASAP7_75t_L g460 ( 
.A(n_326),
.Y(n_460)
);

INVx1_ASAP7_75t_SL g461 ( 
.A(n_127),
.Y(n_461)
);

HB1xp67_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g463 ( 
.A(n_358),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_260),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_231),
.Y(n_465)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_98),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_387),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_104),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_37),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_245),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_281),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_117),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_321),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_392),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_268),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_56),
.Y(n_476)
);

BUFx5_ASAP7_75t_L g477 ( 
.A(n_400),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_226),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_292),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_94),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g481 ( 
.A(n_76),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_47),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_393),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_97),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_126),
.Y(n_485)
);

CKINVDCx5p33_ASAP7_75t_R g486 ( 
.A(n_427),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_395),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_121),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_303),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_89),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_163),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_9),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_420),
.Y(n_493)
);

BUFx2_ASAP7_75t_L g494 ( 
.A(n_381),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_361),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_53),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_385),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g498 ( 
.A(n_419),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_62),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_238),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_345),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_225),
.Y(n_502)
);

INVx3_ASAP7_75t_L g503 ( 
.A(n_295),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_350),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_265),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_259),
.Y(n_506)
);

CKINVDCx20_ASAP7_75t_R g507 ( 
.A(n_311),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_216),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_207),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_317),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_282),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_12),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_84),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_339),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_228),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_64),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_285),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_269),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_144),
.Y(n_520)
);

CKINVDCx5p33_ASAP7_75t_R g521 ( 
.A(n_58),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_164),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_336),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_341),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_69),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_36),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_368),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_271),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_390),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_362),
.Y(n_530)
);

CKINVDCx20_ASAP7_75t_R g531 ( 
.A(n_62),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_374),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_289),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_337),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_55),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_124),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_101),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_156),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_234),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_116),
.Y(n_540)
);

CKINVDCx5p33_ASAP7_75t_R g541 ( 
.A(n_162),
.Y(n_541)
);

BUFx3_ASAP7_75t_L g542 ( 
.A(n_356),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_205),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_86),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_417),
.Y(n_545)
);

BUFx3_ASAP7_75t_L g546 ( 
.A(n_179),
.Y(n_546)
);

INVx2_ASAP7_75t_SL g547 ( 
.A(n_359),
.Y(n_547)
);

INVx1_ASAP7_75t_SL g548 ( 
.A(n_402),
.Y(n_548)
);

CKINVDCx20_ASAP7_75t_R g549 ( 
.A(n_226),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_415),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_149),
.Y(n_551)
);

CKINVDCx5p33_ASAP7_75t_R g552 ( 
.A(n_408),
.Y(n_552)
);

CKINVDCx5p33_ASAP7_75t_R g553 ( 
.A(n_335),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_99),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_79),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_363),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_170),
.Y(n_557)
);

CKINVDCx5p33_ASAP7_75t_R g558 ( 
.A(n_426),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_301),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_344),
.Y(n_560)
);

BUFx6f_ASAP7_75t_L g561 ( 
.A(n_351),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_59),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_377),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_97),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_163),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_247),
.Y(n_566)
);

CKINVDCx5p33_ASAP7_75t_R g567 ( 
.A(n_87),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_78),
.Y(n_568)
);

BUFx6f_ASAP7_75t_L g569 ( 
.A(n_370),
.Y(n_569)
);

CKINVDCx5p33_ASAP7_75t_R g570 ( 
.A(n_152),
.Y(n_570)
);

CKINVDCx5p33_ASAP7_75t_R g571 ( 
.A(n_297),
.Y(n_571)
);

CKINVDCx5p33_ASAP7_75t_R g572 ( 
.A(n_302),
.Y(n_572)
);

CKINVDCx5p33_ASAP7_75t_R g573 ( 
.A(n_134),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_42),
.Y(n_574)
);

CKINVDCx5p33_ASAP7_75t_R g575 ( 
.A(n_346),
.Y(n_575)
);

CKINVDCx5p33_ASAP7_75t_R g576 ( 
.A(n_355),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_181),
.Y(n_577)
);

CKINVDCx5p33_ASAP7_75t_R g578 ( 
.A(n_299),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_63),
.Y(n_579)
);

INVx1_ASAP7_75t_SL g580 ( 
.A(n_191),
.Y(n_580)
);

BUFx2_ASAP7_75t_SL g581 ( 
.A(n_56),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_180),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_229),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_8),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_194),
.Y(n_585)
);

BUFx6f_ASAP7_75t_L g586 ( 
.A(n_86),
.Y(n_586)
);

CKINVDCx20_ASAP7_75t_R g587 ( 
.A(n_20),
.Y(n_587)
);

CKINVDCx5p33_ASAP7_75t_R g588 ( 
.A(n_272),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_147),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_193),
.Y(n_590)
);

CKINVDCx5p33_ASAP7_75t_R g591 ( 
.A(n_10),
.Y(n_591)
);

HB1xp67_ASAP7_75t_L g592 ( 
.A(n_236),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_276),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_12),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_251),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_338),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_179),
.Y(n_597)
);

CKINVDCx5p33_ASAP7_75t_R g598 ( 
.A(n_380),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_325),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_184),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_101),
.Y(n_601)
);

BUFx2_ASAP7_75t_L g602 ( 
.A(n_267),
.Y(n_602)
);

BUFx6f_ASAP7_75t_L g603 ( 
.A(n_243),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_139),
.Y(n_604)
);

INVx2_ASAP7_75t_SL g605 ( 
.A(n_246),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_283),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_266),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_1),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_153),
.Y(n_609)
);

HB1xp67_ASAP7_75t_L g610 ( 
.A(n_221),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_288),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_278),
.Y(n_612)
);

BUFx6f_ASAP7_75t_L g613 ( 
.A(n_71),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_320),
.Y(n_614)
);

CKINVDCx5p33_ASAP7_75t_R g615 ( 
.A(n_365),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_91),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_143),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_107),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_349),
.Y(n_619)
);

CKINVDCx5p33_ASAP7_75t_R g620 ( 
.A(n_353),
.Y(n_620)
);

BUFx10_ASAP7_75t_L g621 ( 
.A(n_369),
.Y(n_621)
);

INVx2_ASAP7_75t_L g622 ( 
.A(n_122),
.Y(n_622)
);

CKINVDCx5p33_ASAP7_75t_R g623 ( 
.A(n_157),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_75),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_307),
.Y(n_625)
);

INVx1_ASAP7_75t_L g626 ( 
.A(n_329),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_115),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_373),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_318),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_286),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_334),
.Y(n_631)
);

INVx1_ASAP7_75t_SL g632 ( 
.A(n_135),
.Y(n_632)
);

CKINVDCx20_ASAP7_75t_R g633 ( 
.A(n_220),
.Y(n_633)
);

CKINVDCx5p33_ASAP7_75t_R g634 ( 
.A(n_429),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_287),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_382),
.Y(n_636)
);

CKINVDCx5p33_ASAP7_75t_R g637 ( 
.A(n_296),
.Y(n_637)
);

INVx2_ASAP7_75t_L g638 ( 
.A(n_22),
.Y(n_638)
);

CKINVDCx5p33_ASAP7_75t_R g639 ( 
.A(n_55),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_37),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_39),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_211),
.Y(n_642)
);

CKINVDCx20_ASAP7_75t_R g643 ( 
.A(n_172),
.Y(n_643)
);

BUFx3_ASAP7_75t_L g644 ( 
.A(n_309),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_200),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_2),
.Y(n_646)
);

CKINVDCx14_ASAP7_75t_R g647 ( 
.A(n_153),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_275),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_316),
.Y(n_649)
);

BUFx6f_ASAP7_75t_L g650 ( 
.A(n_17),
.Y(n_650)
);

CKINVDCx20_ASAP7_75t_R g651 ( 
.A(n_26),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_217),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_354),
.Y(n_653)
);

CKINVDCx20_ASAP7_75t_R g654 ( 
.A(n_210),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_412),
.Y(n_655)
);

INVx2_ASAP7_75t_SL g656 ( 
.A(n_411),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_201),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_422),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_41),
.Y(n_659)
);

CKINVDCx5p33_ASAP7_75t_R g660 ( 
.A(n_423),
.Y(n_660)
);

CKINVDCx5p33_ASAP7_75t_R g661 ( 
.A(n_274),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_277),
.Y(n_662)
);

CKINVDCx20_ASAP7_75t_R g663 ( 
.A(n_310),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_398),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_206),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_308),
.Y(n_666)
);

CKINVDCx5p33_ASAP7_75t_R g667 ( 
.A(n_119),
.Y(n_667)
);

CKINVDCx20_ASAP7_75t_R g668 ( 
.A(n_80),
.Y(n_668)
);

CKINVDCx5p33_ASAP7_75t_R g669 ( 
.A(n_315),
.Y(n_669)
);

CKINVDCx5p33_ASAP7_75t_R g670 ( 
.A(n_357),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_54),
.Y(n_671)
);

CKINVDCx5p33_ASAP7_75t_R g672 ( 
.A(n_191),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_367),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_173),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_30),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_110),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_242),
.Y(n_677)
);

CKINVDCx5p33_ASAP7_75t_R g678 ( 
.A(n_399),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_43),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_324),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_193),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_406),
.Y(n_682)
);

CKINVDCx5p33_ASAP7_75t_R g683 ( 
.A(n_26),
.Y(n_683)
);

INVx3_ASAP7_75t_L g684 ( 
.A(n_375),
.Y(n_684)
);

INVx1_ASAP7_75t_L g685 ( 
.A(n_11),
.Y(n_685)
);

INVxp67_ASAP7_75t_L g686 ( 
.A(n_77),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_428),
.Y(n_687)
);

CKINVDCx5p33_ASAP7_75t_R g688 ( 
.A(n_202),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_13),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_71),
.Y(n_690)
);

CKINVDCx20_ASAP7_75t_R g691 ( 
.A(n_168),
.Y(n_691)
);

INVxp67_ASAP7_75t_L g692 ( 
.A(n_108),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_199),
.Y(n_693)
);

CKINVDCx5p33_ASAP7_75t_R g694 ( 
.A(n_184),
.Y(n_694)
);

CKINVDCx5p33_ASAP7_75t_R g695 ( 
.A(n_364),
.Y(n_695)
);

INVx1_ASAP7_75t_L g696 ( 
.A(n_156),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_54),
.Y(n_697)
);

CKINVDCx20_ASAP7_75t_R g698 ( 
.A(n_174),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_211),
.Y(n_699)
);

BUFx10_ASAP7_75t_L g700 ( 
.A(n_332),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_396),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_416),
.Y(n_702)
);

BUFx8_ASAP7_75t_SL g703 ( 
.A(n_205),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_322),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_24),
.Y(n_705)
);

BUFx2_ASAP7_75t_L g706 ( 
.A(n_167),
.Y(n_706)
);

INVx1_ASAP7_75t_SL g707 ( 
.A(n_165),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_194),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_279),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_78),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_206),
.Y(n_711)
);

CKINVDCx5p33_ASAP7_75t_R g712 ( 
.A(n_397),
.Y(n_712)
);

CKINVDCx5p33_ASAP7_75t_R g713 ( 
.A(n_35),
.Y(n_713)
);

BUFx10_ASAP7_75t_L g714 ( 
.A(n_342),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_340),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_378),
.Y(n_716)
);

CKINVDCx5p33_ASAP7_75t_R g717 ( 
.A(n_39),
.Y(n_717)
);

CKINVDCx16_ASAP7_75t_R g718 ( 
.A(n_379),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_347),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_371),
.Y(n_720)
);

BUFx5_ASAP7_75t_L g721 ( 
.A(n_38),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_190),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_165),
.Y(n_723)
);

CKINVDCx20_ASAP7_75t_R g724 ( 
.A(n_352),
.Y(n_724)
);

CKINVDCx14_ASAP7_75t_R g725 ( 
.A(n_116),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_66),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_333),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_293),
.Y(n_728)
);

INVx1_ASAP7_75t_L g729 ( 
.A(n_312),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_270),
.Y(n_730)
);

BUFx10_ASAP7_75t_L g731 ( 
.A(n_227),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_407),
.Y(n_732)
);

CKINVDCx5p33_ASAP7_75t_R g733 ( 
.A(n_331),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_45),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_73),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_149),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_298),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_197),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_139),
.Y(n_739)
);

BUFx2_ASAP7_75t_L g740 ( 
.A(n_404),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_257),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_409),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_232),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_30),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_74),
.Y(n_745)
);

CKINVDCx5p33_ASAP7_75t_R g746 ( 
.A(n_8),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_212),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_210),
.Y(n_748)
);

CKINVDCx20_ASAP7_75t_R g749 ( 
.A(n_284),
.Y(n_749)
);

CKINVDCx5p33_ASAP7_75t_R g750 ( 
.A(n_188),
.Y(n_750)
);

CKINVDCx5p33_ASAP7_75t_R g751 ( 
.A(n_372),
.Y(n_751)
);

CKINVDCx20_ASAP7_75t_R g752 ( 
.A(n_9),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_50),
.Y(n_753)
);

INVx1_ASAP7_75t_SL g754 ( 
.A(n_414),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_348),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_67),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_90),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_313),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_401),
.Y(n_759)
);

CKINVDCx5p33_ASAP7_75t_R g760 ( 
.A(n_394),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_200),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_721),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_703),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_721),
.Y(n_764)
);

INVx1_ASAP7_75t_SL g765 ( 
.A(n_432),
.Y(n_765)
);

CKINVDCx16_ASAP7_75t_R g766 ( 
.A(n_451),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_721),
.Y(n_767)
);

CKINVDCx20_ASAP7_75t_R g768 ( 
.A(n_438),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_721),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_721),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_721),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_721),
.Y(n_772)
);

BUFx3_ASAP7_75t_L g773 ( 
.A(n_460),
.Y(n_773)
);

CKINVDCx5p33_ASAP7_75t_R g774 ( 
.A(n_436),
.Y(n_774)
);

INVx1_ASAP7_75t_L g775 ( 
.A(n_546),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_647),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_546),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_562),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_441),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_562),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_562),
.Y(n_781)
);

CKINVDCx20_ASAP7_75t_R g782 ( 
.A(n_438),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_562),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_562),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_586),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_586),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_586),
.Y(n_787)
);

CKINVDCx20_ASAP7_75t_R g788 ( 
.A(n_525),
.Y(n_788)
);

INVxp67_ASAP7_75t_L g789 ( 
.A(n_706),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_586),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_586),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_725),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_481),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_443),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_434),
.Y(n_795)
);

INVx2_ASAP7_75t_SL g796 ( 
.A(n_731),
.Y(n_796)
);

CKINVDCx5p33_ASAP7_75t_R g797 ( 
.A(n_437),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_613),
.Y(n_798)
);

INVxp67_ASAP7_75t_L g799 ( 
.A(n_610),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_613),
.Y(n_800)
);

BUFx2_ASAP7_75t_L g801 ( 
.A(n_468),
.Y(n_801)
);

CKINVDCx20_ASAP7_75t_R g802 ( 
.A(n_525),
.Y(n_802)
);

INVxp67_ASAP7_75t_SL g803 ( 
.A(n_462),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_439),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_447),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_613),
.Y(n_806)
);

CKINVDCx5p33_ASAP7_75t_R g807 ( 
.A(n_449),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_450),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_613),
.Y(n_809)
);

CKINVDCx5p33_ASAP7_75t_R g810 ( 
.A(n_453),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_455),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_613),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_650),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_650),
.Y(n_814)
);

CKINVDCx20_ASAP7_75t_R g815 ( 
.A(n_531),
.Y(n_815)
);

CKINVDCx5p33_ASAP7_75t_R g816 ( 
.A(n_456),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_650),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_650),
.Y(n_818)
);

INVx1_ASAP7_75t_SL g819 ( 
.A(n_731),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_650),
.Y(n_820)
);

BUFx6f_ASAP7_75t_L g821 ( 
.A(n_443),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_745),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_490),
.Y(n_823)
);

BUFx2_ASAP7_75t_L g824 ( 
.A(n_468),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_745),
.Y(n_825)
);

CKINVDCx5p33_ASAP7_75t_R g826 ( 
.A(n_491),
.Y(n_826)
);

INVx1_ASAP7_75t_SL g827 ( 
.A(n_731),
.Y(n_827)
);

CKINVDCx5p33_ASAP7_75t_R g828 ( 
.A(n_499),
.Y(n_828)
);

CKINVDCx20_ASAP7_75t_R g829 ( 
.A(n_531),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_476),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_745),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_745),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_745),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_508),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_503),
.B(n_0),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_440),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_466),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_469),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_482),
.Y(n_839)
);

INVx1_ASAP7_75t_L g840 ( 
.A(n_484),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_509),
.Y(n_841)
);

CKINVDCx20_ASAP7_75t_R g842 ( 
.A(n_535),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_535),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_514),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_485),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_488),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_442),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_492),
.Y(n_848)
);

CKINVDCx5p33_ASAP7_75t_R g849 ( 
.A(n_446),
.Y(n_849)
);

INVxp67_ASAP7_75t_L g850 ( 
.A(n_581),
.Y(n_850)
);

CKINVDCx5p33_ASAP7_75t_R g851 ( 
.A(n_448),
.Y(n_851)
);

CKINVDCx16_ASAP7_75t_R g852 ( 
.A(n_463),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_496),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_457),
.Y(n_854)
);

BUFx3_ASAP7_75t_L g855 ( 
.A(n_460),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_502),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_513),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_483),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_538),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_555),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_565),
.Y(n_861)
);

CKINVDCx20_ASAP7_75t_R g862 ( 
.A(n_536),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_486),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_487),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_459),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_459),
.Y(n_866)
);

CKINVDCx20_ASAP7_75t_R g867 ( 
.A(n_536),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_568),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_489),
.Y(n_869)
);

CKINVDCx16_ASAP7_75t_R g870 ( 
.A(n_718),
.Y(n_870)
);

HB1xp67_ASAP7_75t_L g871 ( 
.A(n_476),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_500),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_501),
.Y(n_873)
);

CKINVDCx20_ASAP7_75t_R g874 ( 
.A(n_549),
.Y(n_874)
);

BUFx3_ASAP7_75t_L g875 ( 
.A(n_542),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_459),
.Y(n_876)
);

BUFx6f_ASAP7_75t_L g877 ( 
.A(n_443),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_549),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_579),
.Y(n_879)
);

CKINVDCx5p33_ASAP7_75t_R g880 ( 
.A(n_505),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_506),
.Y(n_881)
);

CKINVDCx5p33_ASAP7_75t_R g882 ( 
.A(n_510),
.Y(n_882)
);

BUFx2_ASAP7_75t_L g883 ( 
.A(n_478),
.Y(n_883)
);

CKINVDCx5p33_ASAP7_75t_R g884 ( 
.A(n_515),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_519),
.Y(n_885)
);

BUFx2_ASAP7_75t_L g886 ( 
.A(n_478),
.Y(n_886)
);

INVxp67_ASAP7_75t_L g887 ( 
.A(n_583),
.Y(n_887)
);

CKINVDCx20_ASAP7_75t_R g888 ( 
.A(n_582),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_542),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_524),
.Y(n_890)
);

CKINVDCx5p33_ASAP7_75t_R g891 ( 
.A(n_528),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_533),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_589),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_534),
.Y(n_894)
);

CKINVDCx5p33_ASAP7_75t_R g895 ( 
.A(n_545),
.Y(n_895)
);

BUFx2_ASAP7_75t_L g896 ( 
.A(n_744),
.Y(n_896)
);

INVx1_ASAP7_75t_SL g897 ( 
.A(n_582),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_550),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_552),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_600),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_601),
.Y(n_901)
);

BUFx2_ASAP7_75t_L g902 ( 
.A(n_744),
.Y(n_902)
);

CKINVDCx5p33_ASAP7_75t_R g903 ( 
.A(n_553),
.Y(n_903)
);

INVxp67_ASAP7_75t_L g904 ( 
.A(n_609),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_459),
.Y(n_905)
);

CKINVDCx5p33_ASAP7_75t_R g906 ( 
.A(n_558),
.Y(n_906)
);

CKINVDCx5p33_ASAP7_75t_R g907 ( 
.A(n_563),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_571),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_659),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_572),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_671),
.Y(n_911)
);

INVx1_ASAP7_75t_L g912 ( 
.A(n_685),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_575),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_689),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_690),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_693),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_459),
.Y(n_917)
);

CKINVDCx5p33_ASAP7_75t_R g918 ( 
.A(n_576),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_696),
.Y(n_919)
);

CKINVDCx5p33_ASAP7_75t_R g920 ( 
.A(n_516),
.Y(n_920)
);

CKINVDCx20_ASAP7_75t_R g921 ( 
.A(n_587),
.Y(n_921)
);

HB1xp67_ASAP7_75t_L g922 ( 
.A(n_746),
.Y(n_922)
);

CKINVDCx5p33_ASAP7_75t_R g923 ( 
.A(n_517),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_452),
.Y(n_924)
);

INVx2_ASAP7_75t_L g925 ( 
.A(n_459),
.Y(n_925)
);

CKINVDCx5p33_ASAP7_75t_R g926 ( 
.A(n_520),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_697),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_710),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_578),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_521),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_723),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_738),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_459),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_739),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_522),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_747),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_477),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_587),
.Y(n_938)
);

INVx1_ASAP7_75t_L g939 ( 
.A(n_748),
.Y(n_939)
);

BUFx2_ASAP7_75t_L g940 ( 
.A(n_746),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_443),
.Y(n_941)
);

INVx1_ASAP7_75t_SL g942 ( 
.A(n_594),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_594),
.Y(n_943)
);

CKINVDCx5p33_ASAP7_75t_R g944 ( 
.A(n_526),
.Y(n_944)
);

INVx1_ASAP7_75t_SL g945 ( 
.A(n_633),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_753),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_560),
.Y(n_947)
);

CKINVDCx16_ASAP7_75t_R g948 ( 
.A(n_507),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_560),
.Y(n_949)
);

INVx1_ASAP7_75t_L g950 ( 
.A(n_644),
.Y(n_950)
);

CKINVDCx16_ASAP7_75t_R g951 ( 
.A(n_507),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_644),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_588),
.Y(n_953)
);

CKINVDCx5p33_ASAP7_75t_R g954 ( 
.A(n_598),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_444),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_599),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_612),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_615),
.Y(n_958)
);

CKINVDCx14_ASAP7_75t_R g959 ( 
.A(n_494),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_454),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_503),
.B(n_230),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_633),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_620),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_467),
.Y(n_964)
);

INVxp67_ASAP7_75t_L g965 ( 
.A(n_750),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_471),
.Y(n_966)
);

CKINVDCx5p33_ASAP7_75t_R g967 ( 
.A(n_631),
.Y(n_967)
);

CKINVDCx20_ASAP7_75t_R g968 ( 
.A(n_643),
.Y(n_968)
);

INVx1_ASAP7_75t_L g969 ( 
.A(n_473),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_634),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_637),
.Y(n_971)
);

CKINVDCx20_ASAP7_75t_R g972 ( 
.A(n_643),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_475),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_503),
.B(n_0),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_648),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_493),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_495),
.Y(n_977)
);

BUFx2_ASAP7_75t_L g978 ( 
.A(n_750),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_511),
.Y(n_979)
);

CKINVDCx5p33_ASAP7_75t_R g980 ( 
.A(n_655),
.Y(n_980)
);

CKINVDCx20_ASAP7_75t_R g981 ( 
.A(n_651),
.Y(n_981)
);

BUFx6f_ASAP7_75t_L g982 ( 
.A(n_443),
.Y(n_982)
);

INVx1_ASAP7_75t_SL g983 ( 
.A(n_651),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_512),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_523),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_477),
.Y(n_986)
);

INVx1_ASAP7_75t_L g987 ( 
.A(n_527),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_530),
.Y(n_988)
);

CKINVDCx5p33_ASAP7_75t_R g989 ( 
.A(n_660),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_661),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_532),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_477),
.Y(n_992)
);

BUFx10_ASAP7_75t_L g993 ( 
.A(n_592),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_662),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_556),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_477),
.Y(n_996)
);

INVxp67_ASAP7_75t_SL g997 ( 
.A(n_602),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_477),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_559),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_664),
.Y(n_1000)
);

OR2x2_ASAP7_75t_L g1001 ( 
.A(n_431),
.B(n_1),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_740),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_654),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_593),
.Y(n_1004)
);

INVx1_ASAP7_75t_L g1005 ( 
.A(n_595),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_606),
.Y(n_1006)
);

CKINVDCx20_ASAP7_75t_R g1007 ( 
.A(n_654),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_619),
.Y(n_1008)
);

INVx1_ASAP7_75t_SL g1009 ( 
.A(n_668),
.Y(n_1009)
);

BUFx8_ASAP7_75t_SL g1010 ( 
.A(n_668),
.Y(n_1010)
);

CKINVDCx20_ASAP7_75t_R g1011 ( 
.A(n_691),
.Y(n_1011)
);

CKINVDCx5p33_ASAP7_75t_R g1012 ( 
.A(n_669),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_670),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_677),
.Y(n_1014)
);

BUFx5_ASAP7_75t_L g1015 ( 
.A(n_626),
.Y(n_1015)
);

CKINVDCx20_ASAP7_75t_R g1016 ( 
.A(n_691),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_628),
.Y(n_1017)
);

CKINVDCx5p33_ASAP7_75t_R g1018 ( 
.A(n_678),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_477),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_629),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_682),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_687),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_537),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_477),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_540),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_452),
.Y(n_1026)
);

NOR2xp67_ASAP7_75t_L g1027 ( 
.A(n_684),
.B(n_2),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_541),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_543),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_630),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_635),
.Y(n_1031)
);

CKINVDCx5p33_ASAP7_75t_R g1032 ( 
.A(n_544),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_636),
.Y(n_1033)
);

CKINVDCx5p33_ASAP7_75t_R g1034 ( 
.A(n_554),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_551),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_649),
.Y(n_1036)
);

CKINVDCx5p33_ASAP7_75t_R g1037 ( 
.A(n_557),
.Y(n_1037)
);

CKINVDCx5p33_ASAP7_75t_R g1038 ( 
.A(n_564),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_653),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_658),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_666),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_673),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_715),
.Y(n_1043)
);

CKINVDCx5p33_ASAP7_75t_R g1044 ( 
.A(n_567),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_570),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_573),
.Y(n_1046)
);

CKINVDCx5p33_ASAP7_75t_R g1047 ( 
.A(n_574),
.Y(n_1047)
);

HB1xp67_ASAP7_75t_L g1048 ( 
.A(n_756),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_551),
.Y(n_1049)
);

INVx1_ASAP7_75t_SL g1050 ( 
.A(n_698),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_716),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_729),
.Y(n_1052)
);

CKINVDCx20_ASAP7_75t_R g1053 ( 
.A(n_698),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_577),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_584),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_585),
.Y(n_1056)
);

CKINVDCx20_ASAP7_75t_R g1057 ( 
.A(n_752),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_730),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_732),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_590),
.Y(n_1060)
);

BUFx3_ASAP7_75t_L g1061 ( 
.A(n_621),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_591),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_741),
.Y(n_1063)
);

INVx1_ASAP7_75t_L g1064 ( 
.A(n_742),
.Y(n_1064)
);

INVx2_ASAP7_75t_L g1065 ( 
.A(n_616),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_759),
.Y(n_1066)
);

BUFx10_ASAP7_75t_L g1067 ( 
.A(n_445),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_435),
.Y(n_1068)
);

CKINVDCx16_ASAP7_75t_R g1069 ( 
.A(n_539),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_752),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_561),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_597),
.Y(n_1072)
);

BUFx3_ASAP7_75t_L g1073 ( 
.A(n_621),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_604),
.Y(n_1074)
);

CKINVDCx14_ASAP7_75t_R g1075 ( 
.A(n_621),
.Y(n_1075)
);

BUFx2_ASAP7_75t_L g1076 ( 
.A(n_756),
.Y(n_1076)
);

CKINVDCx5p33_ASAP7_75t_R g1077 ( 
.A(n_608),
.Y(n_1077)
);

BUFx2_ASAP7_75t_L g1078 ( 
.A(n_757),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_539),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_435),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_617),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_618),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_497),
.Y(n_1083)
);

CKINVDCx20_ASAP7_75t_R g1084 ( 
.A(n_596),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_623),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_624),
.Y(n_1086)
);

CKINVDCx20_ASAP7_75t_R g1087 ( 
.A(n_596),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_627),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_757),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_497),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_611),
.Y(n_1091)
);

INVxp33_ASAP7_75t_L g1092 ( 
.A(n_616),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_695),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_518),
.Y(n_1094)
);

CKINVDCx5p33_ASAP7_75t_R g1095 ( 
.A(n_701),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_702),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_704),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_709),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_518),
.Y(n_1099)
);

INVx2_ASAP7_75t_SL g1100 ( 
.A(n_622),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_712),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_719),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_720),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_622),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_727),
.Y(n_1105)
);

INVx1_ASAP7_75t_SL g1106 ( 
.A(n_461),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_529),
.Y(n_1107)
);

CKINVDCx20_ASAP7_75t_R g1108 ( 
.A(n_611),
.Y(n_1108)
);

INVxp67_ASAP7_75t_SL g1109 ( 
.A(n_684),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_529),
.Y(n_1110)
);

CKINVDCx16_ASAP7_75t_R g1111 ( 
.A(n_663),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_607),
.Y(n_1112)
);

CKINVDCx16_ASAP7_75t_R g1113 ( 
.A(n_663),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_607),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_728),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_614),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_614),
.Y(n_1117)
);

BUFx5_ASAP7_75t_L g1118 ( 
.A(n_700),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_680),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_680),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_638),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_638),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_640),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_640),
.Y(n_1124)
);

HB1xp67_ASAP7_75t_L g1125 ( 
.A(n_761),
.Y(n_1125)
);

NOR2xp33_ASAP7_75t_L g1126 ( 
.A(n_959),
.B(n_445),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_773),
.Y(n_1127)
);

CKINVDCx5p33_ASAP7_75t_R g1128 ( 
.A(n_774),
.Y(n_1128)
);

CKINVDCx5p33_ASAP7_75t_R g1129 ( 
.A(n_779),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_847),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_778),
.Y(n_1131)
);

INVx2_ASAP7_75t_L g1132 ( 
.A(n_780),
.Y(n_1132)
);

INVx2_ASAP7_75t_L g1133 ( 
.A(n_780),
.Y(n_1133)
);

INVx1_ASAP7_75t_L g1134 ( 
.A(n_781),
.Y(n_1134)
);

BUFx6f_ASAP7_75t_SL g1135 ( 
.A(n_1061),
.Y(n_1135)
);

CKINVDCx14_ASAP7_75t_R g1136 ( 
.A(n_1075),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_849),
.Y(n_1137)
);

CKINVDCx5p33_ASAP7_75t_R g1138 ( 
.A(n_851),
.Y(n_1138)
);

CKINVDCx20_ASAP7_75t_R g1139 ( 
.A(n_1079),
.Y(n_1139)
);

CKINVDCx5p33_ASAP7_75t_R g1140 ( 
.A(n_854),
.Y(n_1140)
);

NOR2xp67_ASAP7_75t_L g1141 ( 
.A(n_965),
.B(n_684),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_858),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_863),
.B(n_504),
.Y(n_1143)
);

BUFx2_ASAP7_75t_L g1144 ( 
.A(n_793),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_864),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_783),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_784),
.Y(n_1147)
);

CKINVDCx20_ASAP7_75t_R g1148 ( 
.A(n_1079),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_869),
.B(n_504),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_785),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_786),
.Y(n_1151)
);

INVxp67_ASAP7_75t_SL g1152 ( 
.A(n_850),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_787),
.Y(n_1153)
);

CKINVDCx20_ASAP7_75t_R g1154 ( 
.A(n_1084),
.Y(n_1154)
);

CKINVDCx20_ASAP7_75t_R g1155 ( 
.A(n_1084),
.Y(n_1155)
);

CKINVDCx20_ASAP7_75t_R g1156 ( 
.A(n_1087),
.Y(n_1156)
);

NOR2xp67_ASAP7_75t_L g1157 ( 
.A(n_872),
.B(n_547),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_790),
.Y(n_1158)
);

CKINVDCx5p33_ASAP7_75t_R g1159 ( 
.A(n_873),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_791),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_798),
.Y(n_1161)
);

CKINVDCx20_ASAP7_75t_R g1162 ( 
.A(n_1087),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_1108),
.Y(n_1163)
);

CKINVDCx20_ASAP7_75t_R g1164 ( 
.A(n_1108),
.Y(n_1164)
);

INVxp33_ASAP7_75t_SL g1165 ( 
.A(n_763),
.Y(n_1165)
);

HB1xp67_ASAP7_75t_L g1166 ( 
.A(n_793),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_800),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_806),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_809),
.Y(n_1169)
);

INVxp67_ASAP7_75t_SL g1170 ( 
.A(n_773),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_812),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_813),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_814),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_817),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_818),
.Y(n_1175)
);

CKINVDCx20_ASAP7_75t_R g1176 ( 
.A(n_768),
.Y(n_1176)
);

CKINVDCx5p33_ASAP7_75t_R g1177 ( 
.A(n_880),
.Y(n_1177)
);

CKINVDCx20_ASAP7_75t_R g1178 ( 
.A(n_768),
.Y(n_1178)
);

CKINVDCx5p33_ASAP7_75t_R g1179 ( 
.A(n_881),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_882),
.B(n_547),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_884),
.Y(n_1181)
);

INVx1_ASAP7_75t_L g1182 ( 
.A(n_820),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_885),
.B(n_566),
.Y(n_1183)
);

CKINVDCx16_ASAP7_75t_R g1184 ( 
.A(n_948),
.Y(n_1184)
);

CKINVDCx5p33_ASAP7_75t_R g1185 ( 
.A(n_890),
.Y(n_1185)
);

CKINVDCx20_ASAP7_75t_R g1186 ( 
.A(n_782),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_782),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_822),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_891),
.Y(n_1189)
);

CKINVDCx5p33_ASAP7_75t_R g1190 ( 
.A(n_892),
.Y(n_1190)
);

CKINVDCx20_ASAP7_75t_R g1191 ( 
.A(n_788),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_825),
.Y(n_1192)
);

INVxp67_ASAP7_75t_SL g1193 ( 
.A(n_855),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_894),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_895),
.B(n_566),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_898),
.Y(n_1196)
);

INVxp67_ASAP7_75t_L g1197 ( 
.A(n_1106),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_831),
.Y(n_1198)
);

NOR2xp67_ASAP7_75t_L g1199 ( 
.A(n_899),
.B(n_605),
.Y(n_1199)
);

CKINVDCx20_ASAP7_75t_R g1200 ( 
.A(n_788),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_903),
.Y(n_1201)
);

CKINVDCx20_ASAP7_75t_R g1202 ( 
.A(n_802),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_832),
.Y(n_1203)
);

CKINVDCx20_ASAP7_75t_R g1204 ( 
.A(n_802),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_795),
.Y(n_1205)
);

INVxp67_ASAP7_75t_L g1206 ( 
.A(n_830),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_906),
.Y(n_1207)
);

CKINVDCx5p33_ASAP7_75t_R g1208 ( 
.A(n_907),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_855),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_833),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_955),
.Y(n_1211)
);

BUFx2_ASAP7_75t_SL g1212 ( 
.A(n_1118),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_960),
.Y(n_1213)
);

CKINVDCx20_ASAP7_75t_R g1214 ( 
.A(n_815),
.Y(n_1214)
);

XNOR2xp5_ASAP7_75t_L g1215 ( 
.A(n_815),
.B(n_724),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_964),
.Y(n_1216)
);

CKINVDCx5p33_ASAP7_75t_R g1217 ( 
.A(n_908),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_910),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_913),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_918),
.Y(n_1220)
);

CKINVDCx14_ASAP7_75t_R g1221 ( 
.A(n_776),
.Y(n_1221)
);

CKINVDCx5p33_ASAP7_75t_R g1222 ( 
.A(n_929),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_953),
.Y(n_1223)
);

CKINVDCx16_ASAP7_75t_R g1224 ( 
.A(n_951),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_966),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_969),
.Y(n_1226)
);

CKINVDCx20_ASAP7_75t_R g1227 ( 
.A(n_829),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_954),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_956),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_973),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_957),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_976),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_958),
.Y(n_1233)
);

INVxp33_ASAP7_75t_SL g1234 ( 
.A(n_763),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_963),
.Y(n_1235)
);

INVxp67_ASAP7_75t_SL g1236 ( 
.A(n_875),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_967),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_794),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_970),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_977),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_979),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_984),
.Y(n_1242)
);

NAND2xp5_ASAP7_75t_L g1243 ( 
.A(n_971),
.B(n_605),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_985),
.Y(n_1244)
);

INVxp67_ASAP7_75t_SL g1245 ( 
.A(n_875),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_975),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_987),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_795),
.Y(n_1248)
);

CKINVDCx20_ASAP7_75t_R g1249 ( 
.A(n_829),
.Y(n_1249)
);

CKINVDCx20_ASAP7_75t_R g1250 ( 
.A(n_842),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_988),
.Y(n_1251)
);

CKINVDCx20_ASAP7_75t_R g1252 ( 
.A(n_842),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_991),
.Y(n_1253)
);

INVx1_ASAP7_75t_SL g1254 ( 
.A(n_1010),
.Y(n_1254)
);

CKINVDCx20_ASAP7_75t_R g1255 ( 
.A(n_843),
.Y(n_1255)
);

CKINVDCx5p33_ASAP7_75t_R g1256 ( 
.A(n_980),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_995),
.Y(n_1257)
);

INVxp67_ASAP7_75t_L g1258 ( 
.A(n_871),
.Y(n_1258)
);

INVxp33_ASAP7_75t_SL g1259 ( 
.A(n_989),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_990),
.B(n_656),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_999),
.Y(n_1261)
);

NOR2xp33_ASAP7_75t_L g1262 ( 
.A(n_994),
.B(n_656),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1004),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1005),
.Y(n_1264)
);

CKINVDCx5p33_ASAP7_75t_R g1265 ( 
.A(n_1000),
.Y(n_1265)
);

CKINVDCx16_ASAP7_75t_R g1266 ( 
.A(n_1069),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1006),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1008),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1017),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1020),
.Y(n_1270)
);

CKINVDCx5p33_ASAP7_75t_R g1271 ( 
.A(n_1012),
.Y(n_1271)
);

CKINVDCx5p33_ASAP7_75t_R g1272 ( 
.A(n_1013),
.Y(n_1272)
);

INVxp67_ASAP7_75t_SL g1273 ( 
.A(n_889),
.Y(n_1273)
);

CKINVDCx5p33_ASAP7_75t_R g1274 ( 
.A(n_1014),
.Y(n_1274)
);

CKINVDCx5p33_ASAP7_75t_R g1275 ( 
.A(n_1018),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1030),
.Y(n_1276)
);

CKINVDCx20_ASAP7_75t_R g1277 ( 
.A(n_843),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1031),
.Y(n_1278)
);

CKINVDCx14_ASAP7_75t_R g1279 ( 
.A(n_776),
.Y(n_1279)
);

INVx1_ASAP7_75t_L g1280 ( 
.A(n_1033),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1036),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1021),
.B(n_733),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_794),
.Y(n_1283)
);

CKINVDCx20_ASAP7_75t_R g1284 ( 
.A(n_862),
.Y(n_1284)
);

INVxp33_ASAP7_75t_L g1285 ( 
.A(n_922),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_1022),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_1093),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1039),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_1095),
.Y(n_1289)
);

CKINVDCx16_ASAP7_75t_R g1290 ( 
.A(n_1091),
.Y(n_1290)
);

CKINVDCx5p33_ASAP7_75t_R g1291 ( 
.A(n_1096),
.Y(n_1291)
);

CKINVDCx20_ASAP7_75t_R g1292 ( 
.A(n_862),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1040),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_1097),
.Y(n_1294)
);

INVxp67_ASAP7_75t_L g1295 ( 
.A(n_1048),
.Y(n_1295)
);

INVxp67_ASAP7_75t_L g1296 ( 
.A(n_1125),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1041),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1098),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1042),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_794),
.Y(n_1300)
);

CKINVDCx20_ASAP7_75t_R g1301 ( 
.A(n_867),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_1101),
.Y(n_1302)
);

INVx1_ASAP7_75t_L g1303 ( 
.A(n_1043),
.Y(n_1303)
);

INVxp67_ASAP7_75t_SL g1304 ( 
.A(n_889),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_867),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1051),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1052),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_874),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1058),
.Y(n_1309)
);

CKINVDCx20_ASAP7_75t_R g1310 ( 
.A(n_874),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1059),
.Y(n_1311)
);

CKINVDCx20_ASAP7_75t_R g1312 ( 
.A(n_878),
.Y(n_1312)
);

NOR2xp33_ASAP7_75t_L g1313 ( 
.A(n_1102),
.B(n_458),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1063),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1064),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_1066),
.Y(n_1316)
);

CKINVDCx20_ASAP7_75t_R g1317 ( 
.A(n_878),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1103),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_836),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_797),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_888),
.Y(n_1321)
);

CKINVDCx5p33_ASAP7_75t_R g1322 ( 
.A(n_1105),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_837),
.Y(n_1323)
);

BUFx3_ASAP7_75t_L g1324 ( 
.A(n_961),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_838),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_839),
.Y(n_1326)
);

CKINVDCx20_ASAP7_75t_R g1327 ( 
.A(n_888),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_1115),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_797),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_840),
.Y(n_1330)
);

INVx1_ASAP7_75t_SL g1331 ( 
.A(n_897),
.Y(n_1331)
);

CKINVDCx20_ASAP7_75t_R g1332 ( 
.A(n_921),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_845),
.Y(n_1333)
);

CKINVDCx20_ASAP7_75t_R g1334 ( 
.A(n_921),
.Y(n_1334)
);

CKINVDCx20_ASAP7_75t_R g1335 ( 
.A(n_938),
.Y(n_1335)
);

CKINVDCx20_ASAP7_75t_R g1336 ( 
.A(n_938),
.Y(n_1336)
);

CKINVDCx5p33_ASAP7_75t_R g1337 ( 
.A(n_804),
.Y(n_1337)
);

CKINVDCx20_ASAP7_75t_R g1338 ( 
.A(n_943),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_804),
.Y(n_1339)
);

INVxp67_ASAP7_75t_L g1340 ( 
.A(n_801),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_846),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_997),
.B(n_498),
.Y(n_1342)
);

NOR2xp33_ASAP7_75t_L g1343 ( 
.A(n_1002),
.B(n_548),
.Y(n_1343)
);

CKINVDCx20_ASAP7_75t_R g1344 ( 
.A(n_943),
.Y(n_1344)
);

CKINVDCx16_ASAP7_75t_R g1345 ( 
.A(n_1111),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_805),
.Y(n_1346)
);

CKINVDCx20_ASAP7_75t_R g1347 ( 
.A(n_968),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_805),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_R g1349 ( 
.A(n_807),
.B(n_724),
.Y(n_1349)
);

CKINVDCx5p33_ASAP7_75t_R g1350 ( 
.A(n_807),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_848),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_968),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_853),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_808),
.Y(n_1354)
);

CKINVDCx20_ASAP7_75t_R g1355 ( 
.A(n_972),
.Y(n_1355)
);

INVxp67_ASAP7_75t_SL g1356 ( 
.A(n_1109),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_856),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_857),
.Y(n_1358)
);

CKINVDCx5p33_ASAP7_75t_R g1359 ( 
.A(n_808),
.Y(n_1359)
);

INVxp33_ASAP7_75t_SL g1360 ( 
.A(n_792),
.Y(n_1360)
);

CKINVDCx16_ASAP7_75t_R g1361 ( 
.A(n_1113),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_859),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_810),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_810),
.Y(n_1364)
);

CKINVDCx20_ASAP7_75t_R g1365 ( 
.A(n_972),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_860),
.Y(n_1366)
);

CKINVDCx16_ASAP7_75t_R g1367 ( 
.A(n_766),
.Y(n_1367)
);

INVxp67_ASAP7_75t_L g1368 ( 
.A(n_824),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_861),
.Y(n_1369)
);

CKINVDCx5p33_ASAP7_75t_R g1370 ( 
.A(n_811),
.Y(n_1370)
);

NOR2xp33_ASAP7_75t_L g1371 ( 
.A(n_792),
.B(n_625),
.Y(n_1371)
);

NOR2xp33_ASAP7_75t_L g1372 ( 
.A(n_803),
.B(n_754),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_868),
.Y(n_1373)
);

CKINVDCx20_ASAP7_75t_R g1374 ( 
.A(n_981),
.Y(n_1374)
);

BUFx2_ASAP7_75t_L g1375 ( 
.A(n_811),
.Y(n_1375)
);

CKINVDCx5p33_ASAP7_75t_R g1376 ( 
.A(n_816),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_879),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_816),
.Y(n_1378)
);

INVxp67_ASAP7_75t_SL g1379 ( 
.A(n_947),
.Y(n_1379)
);

INVxp67_ASAP7_75t_SL g1380 ( 
.A(n_949),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_893),
.Y(n_1381)
);

INVx1_ASAP7_75t_L g1382 ( 
.A(n_900),
.Y(n_1382)
);

BUFx3_ASAP7_75t_L g1383 ( 
.A(n_961),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_901),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_823),
.Y(n_1385)
);

CKINVDCx20_ASAP7_75t_R g1386 ( 
.A(n_981),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_909),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_911),
.Y(n_1388)
);

CKINVDCx20_ASAP7_75t_R g1389 ( 
.A(n_1003),
.Y(n_1389)
);

INVxp67_ASAP7_75t_L g1390 ( 
.A(n_883),
.Y(n_1390)
);

NOR2xp33_ASAP7_75t_L g1391 ( 
.A(n_1061),
.B(n_430),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_823),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_912),
.Y(n_1393)
);

CKINVDCx20_ASAP7_75t_R g1394 ( 
.A(n_1003),
.Y(n_1394)
);

BUFx2_ASAP7_75t_SL g1395 ( 
.A(n_1118),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_914),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_826),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_826),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_828),
.Y(n_1399)
);

BUFx2_ASAP7_75t_L g1400 ( 
.A(n_828),
.Y(n_1400)
);

CKINVDCx5p33_ASAP7_75t_R g1401 ( 
.A(n_834),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_915),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_916),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1007),
.Y(n_1404)
);

CKINVDCx5p33_ASAP7_75t_R g1405 ( 
.A(n_834),
.Y(n_1405)
);

CKINVDCx20_ASAP7_75t_R g1406 ( 
.A(n_1007),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_919),
.Y(n_1407)
);

HB1xp67_ASAP7_75t_L g1408 ( 
.A(n_841),
.Y(n_1408)
);

CKINVDCx16_ASAP7_75t_R g1409 ( 
.A(n_852),
.Y(n_1409)
);

NOR2xp33_ASAP7_75t_L g1410 ( 
.A(n_1073),
.B(n_430),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_927),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_928),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_R g1413 ( 
.A(n_841),
.B(n_749),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_931),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1118),
.B(n_737),
.Y(n_1415)
);

CKINVDCx20_ASAP7_75t_R g1416 ( 
.A(n_1011),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_932),
.Y(n_1417)
);

NOR2xp33_ASAP7_75t_L g1418 ( 
.A(n_1073),
.B(n_433),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_R g1419 ( 
.A(n_844),
.B(n_749),
.Y(n_1419)
);

INVxp33_ASAP7_75t_SL g1420 ( 
.A(n_844),
.Y(n_1420)
);

INVxp67_ASAP7_75t_SL g1421 ( 
.A(n_950),
.Y(n_1421)
);

CKINVDCx20_ASAP7_75t_R g1422 ( 
.A(n_1011),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_934),
.Y(n_1423)
);

HB1xp67_ASAP7_75t_L g1424 ( 
.A(n_920),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_936),
.Y(n_1425)
);

NOR2xp33_ASAP7_75t_L g1426 ( 
.A(n_1067),
.B(n_433),
.Y(n_1426)
);

CKINVDCx20_ASAP7_75t_R g1427 ( 
.A(n_1016),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_SL g1428 ( 
.A(n_961),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_939),
.Y(n_1429)
);

CKINVDCx20_ASAP7_75t_R g1430 ( 
.A(n_1016),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_946),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1132),
.Y(n_1432)
);

INVx2_ASAP7_75t_L g1433 ( 
.A(n_1132),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1319),
.Y(n_1434)
);

BUFx6f_ASAP7_75t_L g1435 ( 
.A(n_1238),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1127),
.B(n_775),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1356),
.B(n_1324),
.Y(n_1437)
);

BUFx12f_ASAP7_75t_L g1438 ( 
.A(n_1128),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1323),
.Y(n_1439)
);

INVx3_ASAP7_75t_L g1440 ( 
.A(n_1238),
.Y(n_1440)
);

BUFx6f_ASAP7_75t_L g1441 ( 
.A(n_1283),
.Y(n_1441)
);

AND2x4_ASAP7_75t_L g1442 ( 
.A(n_1127),
.B(n_777),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1324),
.Y(n_1443)
);

BUFx6f_ASAP7_75t_L g1444 ( 
.A(n_1283),
.Y(n_1444)
);

NAND2xp5_ASAP7_75t_L g1445 ( 
.A(n_1383),
.B(n_1118),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1383),
.B(n_1143),
.Y(n_1446)
);

BUFx3_ASAP7_75t_L g1447 ( 
.A(n_1211),
.Y(n_1447)
);

NOR2xp33_ASAP7_75t_L g1448 ( 
.A(n_1170),
.B(n_920),
.Y(n_1448)
);

INVxp67_ASAP7_75t_L g1449 ( 
.A(n_1197),
.Y(n_1449)
);

BUFx6f_ASAP7_75t_L g1450 ( 
.A(n_1300),
.Y(n_1450)
);

AND2x4_ASAP7_75t_L g1451 ( 
.A(n_1193),
.B(n_952),
.Y(n_1451)
);

AND2x6_ASAP7_75t_L g1452 ( 
.A(n_1149),
.B(n_561),
.Y(n_1452)
);

INVx3_ASAP7_75t_L g1453 ( 
.A(n_1300),
.Y(n_1453)
);

AND2x2_ASAP7_75t_L g1454 ( 
.A(n_1136),
.B(n_1152),
.Y(n_1454)
);

INVxp33_ASAP7_75t_SL g1455 ( 
.A(n_1349),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1372),
.B(n_765),
.Y(n_1456)
);

AND2x2_ASAP7_75t_SL g1457 ( 
.A(n_1313),
.B(n_1001),
.Y(n_1457)
);

INVx3_ASAP7_75t_L g1458 ( 
.A(n_1133),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1415),
.A2(n_771),
.B(n_764),
.Y(n_1459)
);

BUFx6f_ASAP7_75t_L g1460 ( 
.A(n_1213),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1325),
.Y(n_1461)
);

CKINVDCx20_ASAP7_75t_R g1462 ( 
.A(n_1176),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1216),
.Y(n_1463)
);

BUFx6f_ASAP7_75t_L g1464 ( 
.A(n_1225),
.Y(n_1464)
);

BUFx3_ASAP7_75t_L g1465 ( 
.A(n_1226),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1326),
.Y(n_1466)
);

AND2x6_ASAP7_75t_L g1467 ( 
.A(n_1195),
.B(n_561),
.Y(n_1467)
);

AOI22xp5_ASAP7_75t_L g1468 ( 
.A1(n_1342),
.A2(n_870),
.B1(n_926),
.B2(n_923),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_L g1469 ( 
.A(n_1260),
.B(n_1118),
.Y(n_1469)
);

INVx2_ASAP7_75t_L g1470 ( 
.A(n_1133),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1330),
.Y(n_1471)
);

OAI22xp5_ASAP7_75t_SL g1472 ( 
.A1(n_1215),
.A2(n_1057),
.B1(n_1070),
.B2(n_1053),
.Y(n_1472)
);

AOI22xp5_ASAP7_75t_L g1473 ( 
.A1(n_1343),
.A2(n_1371),
.B1(n_1206),
.B2(n_1295),
.Y(n_1473)
);

AOI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1258),
.A2(n_923),
.B1(n_930),
.B2(n_926),
.Y(n_1474)
);

INVx3_ASAP7_75t_L g1475 ( 
.A(n_1150),
.Y(n_1475)
);

CKINVDCx5p33_ASAP7_75t_R g1476 ( 
.A(n_1413),
.Y(n_1476)
);

NOR2xp33_ASAP7_75t_L g1477 ( 
.A(n_1209),
.B(n_930),
.Y(n_1477)
);

CKINVDCx5p33_ASAP7_75t_R g1478 ( 
.A(n_1419),
.Y(n_1478)
);

INVx1_ASAP7_75t_L g1479 ( 
.A(n_1333),
.Y(n_1479)
);

NOR2x1_ASAP7_75t_L g1480 ( 
.A(n_1157),
.B(n_835),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1341),
.Y(n_1481)
);

BUFx6f_ASAP7_75t_L g1482 ( 
.A(n_1230),
.Y(n_1482)
);

NAND2xp33_ASAP7_75t_L g1483 ( 
.A(n_1183),
.B(n_1118),
.Y(n_1483)
);

INVx3_ASAP7_75t_L g1484 ( 
.A(n_1150),
.Y(n_1484)
);

OAI21x1_ASAP7_75t_L g1485 ( 
.A1(n_1243),
.A2(n_771),
.B(n_764),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_R g1486 ( 
.A(n_1221),
.B(n_935),
.Y(n_1486)
);

BUFx6f_ASAP7_75t_L g1487 ( 
.A(n_1232),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1331),
.Y(n_1488)
);

OAI22xp5_ASAP7_75t_L g1489 ( 
.A1(n_1296),
.A2(n_974),
.B1(n_1027),
.B2(n_789),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1351),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_L g1491 ( 
.A(n_1240),
.Y(n_1491)
);

BUFx6f_ASAP7_75t_L g1492 ( 
.A(n_1241),
.Y(n_1492)
);

NAND2xp33_ASAP7_75t_L g1493 ( 
.A(n_1242),
.B(n_1118),
.Y(n_1493)
);

AND2x2_ASAP7_75t_L g1494 ( 
.A(n_1285),
.B(n_819),
.Y(n_1494)
);

BUFx6f_ASAP7_75t_L g1495 ( 
.A(n_1244),
.Y(n_1495)
);

AND2x2_ASAP7_75t_L g1496 ( 
.A(n_1236),
.B(n_827),
.Y(n_1496)
);

AND2x2_ASAP7_75t_L g1497 ( 
.A(n_1245),
.B(n_796),
.Y(n_1497)
);

AND2x6_ASAP7_75t_L g1498 ( 
.A(n_1262),
.B(n_561),
.Y(n_1498)
);

INVx2_ASAP7_75t_L g1499 ( 
.A(n_1169),
.Y(n_1499)
);

NAND2xp5_ASAP7_75t_L g1500 ( 
.A(n_1273),
.B(n_1015),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1340),
.A2(n_944),
.B1(n_1023),
.B2(n_935),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1169),
.Y(n_1502)
);

INVx2_ASAP7_75t_L g1503 ( 
.A(n_1171),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1353),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1304),
.B(n_1180),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1379),
.B(n_1380),
.Y(n_1506)
);

AND2x4_ASAP7_75t_L g1507 ( 
.A(n_1421),
.B(n_887),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1171),
.Y(n_1508)
);

NOR2xp33_ASAP7_75t_SL g1509 ( 
.A(n_1259),
.B(n_942),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1426),
.B(n_796),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1357),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1358),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1362),
.Y(n_1513)
);

BUFx6f_ASAP7_75t_L g1514 ( 
.A(n_1247),
.Y(n_1514)
);

NOR2xp33_ASAP7_75t_L g1515 ( 
.A(n_1282),
.B(n_944),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1366),
.Y(n_1516)
);

INVx4_ASAP7_75t_L g1517 ( 
.A(n_1129),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1279),
.Y(n_1518)
);

OR2x6_ASAP7_75t_L g1519 ( 
.A(n_1144),
.B(n_886),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1391),
.B(n_1023),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_1175),
.Y(n_1521)
);

OAI21x1_ASAP7_75t_L g1522 ( 
.A1(n_1175),
.A2(n_767),
.B(n_762),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1199),
.B(n_1015),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1369),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_L g1525 ( 
.A(n_1251),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1141),
.B(n_904),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1212),
.B(n_1015),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1373),
.Y(n_1528)
);

AND2x4_ASAP7_75t_L g1529 ( 
.A(n_1377),
.B(n_1026),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1381),
.B(n_1026),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1382),
.Y(n_1531)
);

BUFx12f_ASAP7_75t_L g1532 ( 
.A(n_1130),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1198),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1395),
.B(n_1015),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1126),
.B(n_1015),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1410),
.B(n_1025),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1198),
.Y(n_1537)
);

BUFx6f_ASAP7_75t_L g1538 ( 
.A(n_1253),
.Y(n_1538)
);

INVx2_ASAP7_75t_L g1539 ( 
.A(n_1131),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1367),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1384),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1134),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1418),
.B(n_1146),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1387),
.Y(n_1544)
);

INVx3_ASAP7_75t_L g1545 ( 
.A(n_1147),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1151),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_L g1547 ( 
.A(n_1257),
.B(n_561),
.Y(n_1547)
);

INVx6_ASAP7_75t_L g1548 ( 
.A(n_1409),
.Y(n_1548)
);

CKINVDCx5p33_ASAP7_75t_R g1549 ( 
.A(n_1137),
.Y(n_1549)
);

INVx2_ASAP7_75t_L g1550 ( 
.A(n_1153),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1388),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1158),
.A2(n_770),
.B(n_769),
.Y(n_1552)
);

AOI22x1_ASAP7_75t_SL g1553 ( 
.A1(n_1176),
.A2(n_1053),
.B1(n_1070),
.B2(n_1057),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_1184),
.Y(n_1554)
);

INVx6_ASAP7_75t_L g1555 ( 
.A(n_1224),
.Y(n_1555)
);

BUFx6f_ASAP7_75t_L g1556 ( 
.A(n_1261),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1393),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1396),
.B(n_1402),
.Y(n_1558)
);

AND2x4_ASAP7_75t_L g1559 ( 
.A(n_1403),
.B(n_1035),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_L g1560 ( 
.A(n_1263),
.Y(n_1560)
);

INVx5_ASAP7_75t_L g1561 ( 
.A(n_1428),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1368),
.B(n_1025),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_L g1563 ( 
.A(n_1160),
.B(n_1015),
.Y(n_1563)
);

NOR2xp33_ASAP7_75t_L g1564 ( 
.A(n_1390),
.B(n_1028),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1407),
.Y(n_1565)
);

INVx2_ASAP7_75t_L g1566 ( 
.A(n_1161),
.Y(n_1566)
);

INVx3_ASAP7_75t_L g1567 ( 
.A(n_1167),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1138),
.B(n_569),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1168),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1205),
.B(n_1028),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1266),
.B(n_945),
.Y(n_1571)
);

AND2x4_ASAP7_75t_L g1572 ( 
.A(n_1411),
.B(n_1035),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1412),
.Y(n_1573)
);

BUFx6f_ASAP7_75t_L g1574 ( 
.A(n_1264),
.Y(n_1574)
);

INVx3_ASAP7_75t_L g1575 ( 
.A(n_1172),
.Y(n_1575)
);

CKINVDCx5p33_ASAP7_75t_R g1576 ( 
.A(n_1290),
.Y(n_1576)
);

AND2x4_ASAP7_75t_L g1577 ( 
.A(n_1414),
.B(n_1049),
.Y(n_1577)
);

INVx1_ASAP7_75t_L g1578 ( 
.A(n_1417),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1423),
.Y(n_1579)
);

NOR2xp33_ASAP7_75t_L g1580 ( 
.A(n_1267),
.B(n_1029),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1248),
.B(n_1029),
.Y(n_1581)
);

HB1xp67_ASAP7_75t_L g1582 ( 
.A(n_1268),
.Y(n_1582)
);

CKINVDCx20_ASAP7_75t_R g1583 ( 
.A(n_1178),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1425),
.B(n_1049),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1173),
.Y(n_1585)
);

AND2x2_ASAP7_75t_L g1586 ( 
.A(n_1375),
.B(n_1032),
.Y(n_1586)
);

HB1xp67_ASAP7_75t_L g1587 ( 
.A(n_1269),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1429),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1345),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1431),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1270),
.Y(n_1591)
);

INVx2_ASAP7_75t_L g1592 ( 
.A(n_1174),
.Y(n_1592)
);

OAI22x1_ASAP7_75t_SL g1593 ( 
.A1(n_1178),
.A2(n_962),
.B1(n_1009),
.B2(n_983),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1276),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1278),
.Y(n_1595)
);

HB1xp67_ASAP7_75t_L g1596 ( 
.A(n_1280),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1182),
.Y(n_1597)
);

INVx2_ASAP7_75t_L g1598 ( 
.A(n_1188),
.Y(n_1598)
);

INVx5_ASAP7_75t_L g1599 ( 
.A(n_1428),
.Y(n_1599)
);

INVx2_ASAP7_75t_L g1600 ( 
.A(n_1192),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1400),
.B(n_1032),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1281),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1203),
.B(n_1015),
.Y(n_1603)
);

INVx1_ASAP7_75t_L g1604 ( 
.A(n_1288),
.Y(n_1604)
);

NAND2x1p5_ASAP7_75t_L g1605 ( 
.A(n_1293),
.B(n_569),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1210),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1297),
.Y(n_1607)
);

INVx3_ASAP7_75t_L g1608 ( 
.A(n_1299),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1303),
.B(n_1034),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1306),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1307),
.Y(n_1611)
);

BUFx6f_ASAP7_75t_L g1612 ( 
.A(n_1309),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_SL g1613 ( 
.A(n_1140),
.B(n_569),
.Y(n_1613)
);

AND2x4_ASAP7_75t_L g1614 ( 
.A(n_1311),
.B(n_1065),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1314),
.B(n_772),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1315),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1316),
.B(n_1034),
.Y(n_1617)
);

INVx4_ASAP7_75t_L g1618 ( 
.A(n_1142),
.Y(n_1618)
);

BUFx6f_ASAP7_75t_L g1619 ( 
.A(n_1145),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1428),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1135),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_SL g1622 ( 
.A(n_1159),
.B(n_569),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1135),
.Y(n_1623)
);

CKINVDCx6p67_ASAP7_75t_R g1624 ( 
.A(n_1361),
.Y(n_1624)
);

AND2x6_ASAP7_75t_L g1625 ( 
.A(n_1254),
.B(n_569),
.Y(n_1625)
);

BUFx6f_ASAP7_75t_L g1626 ( 
.A(n_1177),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1135),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1179),
.B(n_1037),
.Y(n_1628)
);

OA21x2_ASAP7_75t_L g1629 ( 
.A1(n_1181),
.A2(n_1080),
.B(n_1068),
.Y(n_1629)
);

INVx2_ASAP7_75t_L g1630 ( 
.A(n_1320),
.Y(n_1630)
);

AND2x4_ASAP7_75t_L g1631 ( 
.A(n_1408),
.B(n_1065),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1185),
.Y(n_1632)
);

OA21x2_ASAP7_75t_L g1633 ( 
.A1(n_1189),
.A2(n_1090),
.B(n_1083),
.Y(n_1633)
);

CKINVDCx16_ASAP7_75t_R g1634 ( 
.A(n_1139),
.Y(n_1634)
);

AND2x4_ASAP7_75t_L g1635 ( 
.A(n_1424),
.B(n_1104),
.Y(n_1635)
);

AND2x4_ASAP7_75t_L g1636 ( 
.A(n_1166),
.B(n_1104),
.Y(n_1636)
);

NOR2xp33_ASAP7_75t_R g1637 ( 
.A(n_1329),
.B(n_1337),
.Y(n_1637)
);

AND2x4_ASAP7_75t_L g1638 ( 
.A(n_1190),
.B(n_1121),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1194),
.B(n_1121),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1196),
.B(n_1037),
.Y(n_1640)
);

OAI22xp5_ASAP7_75t_L g1641 ( 
.A1(n_1201),
.A2(n_1044),
.B1(n_1045),
.B2(n_1038),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1207),
.B(n_1038),
.Y(n_1642)
);

BUFx3_ASAP7_75t_L g1643 ( 
.A(n_1339),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1208),
.Y(n_1644)
);

OAI22xp5_ASAP7_75t_L g1645 ( 
.A1(n_1217),
.A2(n_1045),
.B1(n_1046),
.B2(n_1044),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_SL g1646 ( 
.A(n_1218),
.B(n_603),
.Y(n_1646)
);

BUFx3_ASAP7_75t_L g1647 ( 
.A(n_1346),
.Y(n_1647)
);

OAI22x1_ASAP7_75t_R g1648 ( 
.A1(n_1186),
.A2(n_1050),
.B1(n_761),
.B2(n_1047),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1219),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1348),
.Y(n_1650)
);

BUFx3_ASAP7_75t_L g1651 ( 
.A(n_1350),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1220),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1222),
.B(n_924),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1223),
.Y(n_1654)
);

OAI22xp5_ASAP7_75t_L g1655 ( 
.A1(n_1228),
.A2(n_1047),
.B1(n_1054),
.B2(n_1046),
.Y(n_1655)
);

AND3x1_ASAP7_75t_L g1656 ( 
.A(n_1420),
.B(n_657),
.C(n_431),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1229),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1231),
.Y(n_1658)
);

INVx3_ASAP7_75t_L g1659 ( 
.A(n_1233),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1235),
.Y(n_1660)
);

AND2x2_ASAP7_75t_L g1661 ( 
.A(n_1237),
.B(n_1054),
.Y(n_1661)
);

INVx1_ASAP7_75t_L g1662 ( 
.A(n_1239),
.Y(n_1662)
);

CKINVDCx20_ASAP7_75t_R g1663 ( 
.A(n_1186),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1246),
.Y(n_1664)
);

AOI22x1_ASAP7_75t_SL g1665 ( 
.A1(n_1187),
.A2(n_641),
.B1(n_642),
.B2(n_639),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1256),
.B(n_1055),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1265),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1271),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1272),
.B(n_1055),
.Y(n_1669)
);

AND2x4_ASAP7_75t_L g1670 ( 
.A(n_1274),
.B(n_924),
.Y(n_1670)
);

INVx2_ASAP7_75t_L g1671 ( 
.A(n_1275),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1286),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1287),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1289),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1291),
.B(n_1056),
.Y(n_1675)
);

BUFx2_ASAP7_75t_L g1676 ( 
.A(n_1187),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1294),
.Y(n_1677)
);

AND2x2_ASAP7_75t_L g1678 ( 
.A(n_1298),
.B(n_1056),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1302),
.Y(n_1679)
);

OAI22xp5_ASAP7_75t_L g1680 ( 
.A1(n_1318),
.A2(n_1062),
.B1(n_1072),
.B2(n_1060),
.Y(n_1680)
);

BUFx6f_ASAP7_75t_L g1681 ( 
.A(n_1322),
.Y(n_1681)
);

OA21x2_ASAP7_75t_L g1682 ( 
.A1(n_1328),
.A2(n_1099),
.B(n_1094),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1354),
.Y(n_1683)
);

BUFx12f_ASAP7_75t_L g1684 ( 
.A(n_1359),
.Y(n_1684)
);

INVx3_ASAP7_75t_L g1685 ( 
.A(n_1363),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1364),
.Y(n_1686)
);

INVx2_ASAP7_75t_L g1687 ( 
.A(n_1370),
.Y(n_1687)
);

BUFx6f_ASAP7_75t_L g1688 ( 
.A(n_1376),
.Y(n_1688)
);

BUFx6f_ASAP7_75t_L g1689 ( 
.A(n_1378),
.Y(n_1689)
);

OA21x2_ASAP7_75t_L g1690 ( 
.A1(n_1385),
.A2(n_1110),
.B(n_1107),
.Y(n_1690)
);

INVx1_ASAP7_75t_L g1691 ( 
.A(n_1392),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1397),
.B(n_1060),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1398),
.B(n_896),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1399),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1401),
.Y(n_1695)
);

INVx3_ASAP7_75t_L g1696 ( 
.A(n_1405),
.Y(n_1696)
);

OAI21x1_ASAP7_75t_L g1697 ( 
.A1(n_1360),
.A2(n_866),
.B(n_865),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1165),
.B(n_1062),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1234),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1139),
.Y(n_1700)
);

INVx1_ASAP7_75t_L g1701 ( 
.A(n_1148),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1148),
.B(n_1072),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1154),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1154),
.Y(n_1704)
);

BUFx6f_ASAP7_75t_L g1705 ( 
.A(n_1155),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1155),
.B(n_1074),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1156),
.Y(n_1707)
);

OA21x2_ASAP7_75t_L g1708 ( 
.A1(n_1156),
.A2(n_1114),
.B(n_1112),
.Y(n_1708)
);

BUFx6f_ASAP7_75t_L g1709 ( 
.A(n_1162),
.Y(n_1709)
);

AND2x2_ASAP7_75t_L g1710 ( 
.A(n_1162),
.B(n_1074),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1163),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1163),
.B(n_1077),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1164),
.Y(n_1713)
);

NAND2xp33_ASAP7_75t_L g1714 ( 
.A(n_1164),
.B(n_603),
.Y(n_1714)
);

BUFx6f_ASAP7_75t_L g1715 ( 
.A(n_1191),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1430),
.Y(n_1716)
);

BUFx6f_ASAP7_75t_L g1717 ( 
.A(n_1191),
.Y(n_1717)
);

BUFx8_ASAP7_75t_L g1718 ( 
.A(n_1200),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1200),
.B(n_1077),
.Y(n_1719)
);

OA21x2_ASAP7_75t_L g1720 ( 
.A1(n_1202),
.A2(n_1117),
.B(n_1116),
.Y(n_1720)
);

INVx3_ASAP7_75t_L g1721 ( 
.A(n_1522),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1529),
.Y(n_1722)
);

BUFx6f_ASAP7_75t_L g1723 ( 
.A(n_1443),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1488),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1529),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1432),
.Y(n_1726)
);

NAND2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1456),
.B(n_657),
.Y(n_1727)
);

INVx3_ASAP7_75t_L g1728 ( 
.A(n_1552),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1432),
.Y(n_1729)
);

INVx3_ASAP7_75t_L g1730 ( 
.A(n_1552),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1433),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1530),
.Y(n_1732)
);

OAI21x1_ASAP7_75t_L g1733 ( 
.A1(n_1485),
.A2(n_866),
.B(n_865),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1449),
.B(n_902),
.Y(n_1734)
);

INVx2_ASAP7_75t_L g1735 ( 
.A(n_1433),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1530),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1488),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1559),
.Y(n_1738)
);

INVx3_ASAP7_75t_L g1739 ( 
.A(n_1552),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1446),
.B(n_1081),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1437),
.B(n_1081),
.Y(n_1741)
);

AND2x6_ASAP7_75t_L g1742 ( 
.A(n_1621),
.B(n_603),
.Y(n_1742)
);

INVx3_ASAP7_75t_L g1743 ( 
.A(n_1697),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1470),
.Y(n_1744)
);

INVx3_ASAP7_75t_L g1745 ( 
.A(n_1435),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1470),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1449),
.B(n_940),
.Y(n_1747)
);

BUFx2_ASAP7_75t_L g1748 ( 
.A(n_1494),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1457),
.B(n_1082),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1559),
.Y(n_1750)
);

INVx2_ASAP7_75t_L g1751 ( 
.A(n_1499),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1499),
.Y(n_1752)
);

AND2x4_ASAP7_75t_L g1753 ( 
.A(n_1443),
.B(n_1122),
.Y(n_1753)
);

HB1xp67_ASAP7_75t_L g1754 ( 
.A(n_1705),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1502),
.Y(n_1755)
);

AND2x2_ASAP7_75t_SL g1756 ( 
.A(n_1457),
.B(n_603),
.Y(n_1756)
);

INVx2_ASAP7_75t_L g1757 ( 
.A(n_1502),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1572),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1572),
.Y(n_1759)
);

AND2x2_ASAP7_75t_L g1760 ( 
.A(n_1510),
.B(n_978),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1577),
.Y(n_1761)
);

BUFx6f_ASAP7_75t_L g1762 ( 
.A(n_1460),
.Y(n_1762)
);

BUFx6f_ASAP7_75t_L g1763 ( 
.A(n_1460),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1577),
.Y(n_1764)
);

BUFx6f_ASAP7_75t_L g1765 ( 
.A(n_1460),
.Y(n_1765)
);

OA21x2_ASAP7_75t_L g1766 ( 
.A1(n_1563),
.A2(n_905),
.B(n_876),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1548),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1584),
.Y(n_1768)
);

BUFx6f_ASAP7_75t_L g1769 ( 
.A(n_1460),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1584),
.Y(n_1770)
);

OR2x2_ASAP7_75t_L g1771 ( 
.A(n_1571),
.B(n_1076),
.Y(n_1771)
);

BUFx2_ASAP7_75t_L g1772 ( 
.A(n_1707),
.Y(n_1772)
);

INVx3_ASAP7_75t_L g1773 ( 
.A(n_1435),
.Y(n_1773)
);

NAND2xp5_ASAP7_75t_L g1774 ( 
.A(n_1515),
.B(n_1082),
.Y(n_1774)
);

INVx2_ASAP7_75t_L g1775 ( 
.A(n_1503),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1515),
.B(n_1085),
.Y(n_1776)
);

INVx1_ASAP7_75t_SL g1777 ( 
.A(n_1462),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1503),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1614),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1508),
.Y(n_1780)
);

INVx3_ASAP7_75t_L g1781 ( 
.A(n_1435),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1508),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1521),
.Y(n_1783)
);

AND2x4_ASAP7_75t_L g1784 ( 
.A(n_1447),
.B(n_1123),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1614),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1616),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1616),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1463),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1521),
.Y(n_1789)
);

NOR2xp33_ASAP7_75t_SL g1790 ( 
.A(n_1455),
.B(n_1085),
.Y(n_1790)
);

BUFx6f_ASAP7_75t_L g1791 ( 
.A(n_1463),
.Y(n_1791)
);

INVx2_ASAP7_75t_L g1792 ( 
.A(n_1533),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1533),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1434),
.Y(n_1794)
);

CKINVDCx16_ASAP7_75t_R g1795 ( 
.A(n_1634),
.Y(n_1795)
);

INVx3_ASAP7_75t_L g1796 ( 
.A(n_1435),
.Y(n_1796)
);

OR2x2_ASAP7_75t_L g1797 ( 
.A(n_1707),
.B(n_1078),
.Y(n_1797)
);

INVx4_ASAP7_75t_L g1798 ( 
.A(n_1441),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1506),
.B(n_1086),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1537),
.Y(n_1800)
);

BUFx6f_ASAP7_75t_L g1801 ( 
.A(n_1463),
.Y(n_1801)
);

AND2x2_ASAP7_75t_L g1802 ( 
.A(n_1497),
.B(n_1089),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1537),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1439),
.Y(n_1804)
);

AND2x2_ASAP7_75t_L g1805 ( 
.A(n_1496),
.B(n_1092),
.Y(n_1805)
);

BUFx6f_ASAP7_75t_L g1806 ( 
.A(n_1463),
.Y(n_1806)
);

INVx2_ASAP7_75t_L g1807 ( 
.A(n_1458),
.Y(n_1807)
);

NAND2xp5_ASAP7_75t_L g1808 ( 
.A(n_1506),
.B(n_1086),
.Y(n_1808)
);

INVxp67_ASAP7_75t_L g1809 ( 
.A(n_1564),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1461),
.Y(n_1810)
);

HB1xp67_ASAP7_75t_L g1811 ( 
.A(n_1705),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1458),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1466),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1471),
.Y(n_1814)
);

OA21x2_ASAP7_75t_L g1815 ( 
.A1(n_1603),
.A2(n_905),
.B(n_876),
.Y(n_1815)
);

CKINVDCx5p33_ASAP7_75t_R g1816 ( 
.A(n_1476),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1440),
.Y(n_1817)
);

INVx1_ASAP7_75t_SL g1818 ( 
.A(n_1462),
.Y(n_1818)
);

NAND2xp5_ASAP7_75t_SL g1819 ( 
.A(n_1469),
.B(n_603),
.Y(n_1819)
);

INVx3_ASAP7_75t_L g1820 ( 
.A(n_1441),
.Y(n_1820)
);

HB1xp67_ASAP7_75t_L g1821 ( 
.A(n_1705),
.Y(n_1821)
);

BUFx6f_ASAP7_75t_L g1822 ( 
.A(n_1464),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1479),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1481),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1440),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1535),
.B(n_1088),
.Y(n_1826)
);

BUFx2_ASAP7_75t_L g1827 ( 
.A(n_1711),
.Y(n_1827)
);

NOR2xp33_ASAP7_75t_L g1828 ( 
.A(n_1473),
.B(n_1088),
.Y(n_1828)
);

AND2x4_ASAP7_75t_L g1829 ( 
.A(n_1447),
.B(n_1124),
.Y(n_1829)
);

HB1xp67_ASAP7_75t_L g1830 ( 
.A(n_1705),
.Y(n_1830)
);

AND2x2_ASAP7_75t_L g1831 ( 
.A(n_1526),
.B(n_799),
.Y(n_1831)
);

INVx2_ASAP7_75t_L g1832 ( 
.A(n_1453),
.Y(n_1832)
);

HB1xp67_ASAP7_75t_L g1833 ( 
.A(n_1709),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1490),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1526),
.B(n_993),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1453),
.Y(n_1836)
);

AND2x4_ASAP7_75t_L g1837 ( 
.A(n_1465),
.B(n_711),
.Y(n_1837)
);

BUFx6f_ASAP7_75t_L g1838 ( 
.A(n_1464),
.Y(n_1838)
);

BUFx6f_ASAP7_75t_L g1839 ( 
.A(n_1464),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1504),
.Y(n_1840)
);

AND2x4_ASAP7_75t_L g1841 ( 
.A(n_1465),
.B(n_711),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1511),
.Y(n_1842)
);

INVx2_ASAP7_75t_L g1843 ( 
.A(n_1475),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1451),
.B(n_993),
.Y(n_1844)
);

NOR2xp33_ASAP7_75t_SL g1845 ( 
.A(n_1455),
.B(n_700),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1543),
.B(n_1119),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_SL g1847 ( 
.A(n_1653),
.B(n_743),
.Y(n_1847)
);

INVx1_ASAP7_75t_L g1848 ( 
.A(n_1512),
.Y(n_1848)
);

OAI22xp5_ASAP7_75t_SL g1849 ( 
.A1(n_1472),
.A2(n_1204),
.B1(n_1214),
.B2(n_1202),
.Y(n_1849)
);

AND2x4_ASAP7_75t_L g1850 ( 
.A(n_1558),
.B(n_1100),
.Y(n_1850)
);

BUFx8_ASAP7_75t_L g1851 ( 
.A(n_1676),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1513),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1475),
.Y(n_1853)
);

INVxp67_ASAP7_75t_L g1854 ( 
.A(n_1564),
.Y(n_1854)
);

INVx1_ASAP7_75t_L g1855 ( 
.A(n_1516),
.Y(n_1855)
);

INVx3_ASAP7_75t_L g1856 ( 
.A(n_1441),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_SL g1857 ( 
.A(n_1653),
.B(n_464),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1524),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1528),
.Y(n_1859)
);

INVx2_ASAP7_75t_L g1860 ( 
.A(n_1484),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1709),
.Y(n_1861)
);

XOR2x2_ASAP7_75t_L g1862 ( 
.A(n_1656),
.B(n_1468),
.Y(n_1862)
);

OAI22xp5_ASAP7_75t_SL g1863 ( 
.A1(n_1583),
.A2(n_1430),
.B1(n_1214),
.B2(n_1227),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1531),
.Y(n_1864)
);

BUFx6f_ASAP7_75t_L g1865 ( 
.A(n_1464),
.Y(n_1865)
);

INVx2_ASAP7_75t_L g1866 ( 
.A(n_1484),
.Y(n_1866)
);

NAND2xp33_ASAP7_75t_R g1867 ( 
.A(n_1708),
.B(n_645),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1541),
.Y(n_1868)
);

INVx4_ASAP7_75t_L g1869 ( 
.A(n_1441),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1539),
.Y(n_1870)
);

INVx2_ASAP7_75t_L g1871 ( 
.A(n_1539),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1544),
.Y(n_1872)
);

INVx3_ASAP7_75t_L g1873 ( 
.A(n_1444),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1551),
.Y(n_1874)
);

BUFx6f_ASAP7_75t_L g1875 ( 
.A(n_1482),
.Y(n_1875)
);

NOR2xp33_ASAP7_75t_L g1876 ( 
.A(n_1617),
.B(n_993),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1608),
.B(n_1119),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1557),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1608),
.B(n_1119),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1565),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1573),
.Y(n_1881)
);

BUFx6f_ASAP7_75t_L g1882 ( 
.A(n_1482),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1545),
.B(n_1067),
.Y(n_1883)
);

NAND2xp5_ASAP7_75t_SL g1884 ( 
.A(n_1670),
.B(n_464),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1545),
.B(n_1067),
.Y(n_1885)
);

AOI22xp5_ASAP7_75t_L g1886 ( 
.A1(n_1448),
.A2(n_470),
.B1(n_474),
.B2(n_465),
.Y(n_1886)
);

INVx2_ASAP7_75t_L g1887 ( 
.A(n_1542),
.Y(n_1887)
);

INVx2_ASAP7_75t_L g1888 ( 
.A(n_1542),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1546),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1546),
.Y(n_1890)
);

CKINVDCx5p33_ASAP7_75t_R g1891 ( 
.A(n_1476),
.Y(n_1891)
);

NOR2xp33_ASAP7_75t_L g1892 ( 
.A(n_1582),
.B(n_472),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1550),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1567),
.B(n_1120),
.Y(n_1894)
);

INVx1_ASAP7_75t_L g1895 ( 
.A(n_1578),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1579),
.Y(n_1896)
);

NAND2xp5_ASAP7_75t_L g1897 ( 
.A(n_1567),
.B(n_1575),
.Y(n_1897)
);

HB1xp67_ASAP7_75t_L g1898 ( 
.A(n_1709),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1451),
.B(n_1100),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1507),
.B(n_917),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1588),
.Y(n_1901)
);

AND2x4_ASAP7_75t_L g1902 ( 
.A(n_1558),
.B(n_233),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1550),
.Y(n_1903)
);

BUFx6f_ASAP7_75t_L g1904 ( 
.A(n_1482),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1507),
.B(n_1631),
.Y(n_1905)
);

INVx2_ASAP7_75t_L g1906 ( 
.A(n_1566),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1590),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_SL g1908 ( 
.A(n_1478),
.B(n_700),
.Y(n_1908)
);

INVx2_ASAP7_75t_L g1909 ( 
.A(n_1566),
.Y(n_1909)
);

INVx2_ASAP7_75t_L g1910 ( 
.A(n_1569),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1591),
.Y(n_1911)
);

BUFx6f_ASAP7_75t_L g1912 ( 
.A(n_1482),
.Y(n_1912)
);

BUFx2_ASAP7_75t_L g1913 ( 
.A(n_1711),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1594),
.Y(n_1914)
);

AND2x6_ASAP7_75t_L g1915 ( 
.A(n_1621),
.B(n_917),
.Y(n_1915)
);

CKINVDCx16_ASAP7_75t_R g1916 ( 
.A(n_1486),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1595),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1569),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1585),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1602),
.Y(n_1920)
);

BUFx2_ASAP7_75t_L g1921 ( 
.A(n_1716),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1604),
.B(n_235),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1607),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1610),
.Y(n_1924)
);

AND2x2_ASAP7_75t_L g1925 ( 
.A(n_1631),
.B(n_925),
.Y(n_1925)
);

CKINVDCx5p33_ASAP7_75t_R g1926 ( 
.A(n_1478),
.Y(n_1926)
);

OA21x2_ASAP7_75t_L g1927 ( 
.A1(n_1459),
.A2(n_933),
.B(n_925),
.Y(n_1927)
);

CKINVDCx20_ASAP7_75t_R g1928 ( 
.A(n_1583),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1582),
.Y(n_1929)
);

BUFx6f_ASAP7_75t_SL g1930 ( 
.A(n_1619),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1587),
.Y(n_1931)
);

INVx2_ASAP7_75t_L g1932 ( 
.A(n_1585),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1587),
.Y(n_1933)
);

OA21x2_ASAP7_75t_L g1934 ( 
.A1(n_1500),
.A2(n_1615),
.B(n_1445),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1596),
.Y(n_1935)
);

INVxp67_ASAP7_75t_L g1936 ( 
.A(n_1509),
.Y(n_1936)
);

INVx2_ASAP7_75t_L g1937 ( 
.A(n_1592),
.Y(n_1937)
);

XOR2xp5_ASAP7_75t_L g1938 ( 
.A(n_1553),
.B(n_1204),
.Y(n_1938)
);

BUFx6f_ASAP7_75t_L g1939 ( 
.A(n_1487),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1596),
.Y(n_1940)
);

INVx3_ASAP7_75t_L g1941 ( 
.A(n_1444),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1592),
.Y(n_1942)
);

INVxp33_ASAP7_75t_SL g1943 ( 
.A(n_1637),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1562),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1597),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1575),
.B(n_465),
.Y(n_1946)
);

INVx4_ASAP7_75t_L g1947 ( 
.A(n_1444),
.Y(n_1947)
);

BUFx2_ASAP7_75t_L g1948 ( 
.A(n_1716),
.Y(n_1948)
);

INVxp67_ASAP7_75t_L g1949 ( 
.A(n_1580),
.Y(n_1949)
);

AND2x4_ASAP7_75t_L g1950 ( 
.A(n_1436),
.B(n_237),
.Y(n_1950)
);

INVx1_ASAP7_75t_L g1951 ( 
.A(n_1597),
.Y(n_1951)
);

INVx2_ASAP7_75t_L g1952 ( 
.A(n_1598),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1635),
.B(n_1670),
.Y(n_1953)
);

INVx3_ASAP7_75t_L g1954 ( 
.A(n_1444),
.Y(n_1954)
);

INVx3_ASAP7_75t_L g1955 ( 
.A(n_1450),
.Y(n_1955)
);

INVx2_ASAP7_75t_L g1956 ( 
.A(n_1598),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1505),
.B(n_1448),
.Y(n_1957)
);

INVx3_ASAP7_75t_L g1958 ( 
.A(n_1450),
.Y(n_1958)
);

OR2x2_ASAP7_75t_L g1959 ( 
.A(n_1702),
.B(n_580),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1600),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1635),
.B(n_933),
.Y(n_1961)
);

BUFx6f_ASAP7_75t_L g1962 ( 
.A(n_1487),
.Y(n_1962)
);

OAI21x1_ASAP7_75t_L g1963 ( 
.A1(n_1527),
.A2(n_986),
.B(n_937),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1600),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1477),
.B(n_470),
.Y(n_1965)
);

BUFx6f_ASAP7_75t_L g1966 ( 
.A(n_1487),
.Y(n_1966)
);

BUFx6f_ASAP7_75t_L g1967 ( 
.A(n_1487),
.Y(n_1967)
);

INVx1_ASAP7_75t_L g1968 ( 
.A(n_1606),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1606),
.Y(n_1969)
);

OAI21x1_ASAP7_75t_L g1970 ( 
.A1(n_1534),
.A2(n_986),
.B(n_937),
.Y(n_1970)
);

AND2x4_ASAP7_75t_L g1971 ( 
.A(n_1436),
.B(n_239),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1638),
.B(n_992),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1477),
.B(n_474),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1450),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1442),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1442),
.Y(n_1976)
);

INVxp33_ASAP7_75t_L g1977 ( 
.A(n_1648),
.Y(n_1977)
);

BUFx6f_ASAP7_75t_L g1978 ( 
.A(n_1491),
.Y(n_1978)
);

INVx1_ASAP7_75t_L g1979 ( 
.A(n_1636),
.Y(n_1979)
);

OA21x2_ASAP7_75t_L g1980 ( 
.A1(n_1523),
.A2(n_996),
.B(n_992),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1580),
.A2(n_751),
.B1(n_755),
.B2(n_479),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1636),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1491),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1491),
.B(n_479),
.Y(n_1984)
);

BUFx6f_ASAP7_75t_L g1985 ( 
.A(n_1491),
.Y(n_1985)
);

INVx2_ASAP7_75t_L g1986 ( 
.A(n_1450),
.Y(n_1986)
);

INVx1_ASAP7_75t_L g1987 ( 
.A(n_1492),
.Y(n_1987)
);

INVxp67_ASAP7_75t_L g1988 ( 
.A(n_1609),
.Y(n_1988)
);

AND2x4_ASAP7_75t_L g1989 ( 
.A(n_1620),
.B(n_240),
.Y(n_1989)
);

BUFx6f_ASAP7_75t_L g1990 ( 
.A(n_1492),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1609),
.B(n_632),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1492),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1638),
.B(n_996),
.Y(n_1993)
);

OA21x2_ASAP7_75t_L g1994 ( 
.A1(n_1568),
.A2(n_1019),
.B(n_998),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1492),
.Y(n_1995)
);

INVx1_ASAP7_75t_SL g1996 ( 
.A(n_1663),
.Y(n_1996)
);

INVx3_ASAP7_75t_L g1997 ( 
.A(n_1495),
.Y(n_1997)
);

AND2x4_ASAP7_75t_L g1998 ( 
.A(n_1639),
.B(n_241),
.Y(n_1998)
);

BUFx2_ASAP7_75t_L g1999 ( 
.A(n_1519),
.Y(n_1999)
);

CKINVDCx5p33_ASAP7_75t_R g2000 ( 
.A(n_1486),
.Y(n_2000)
);

AND2x4_ASAP7_75t_L g2001 ( 
.A(n_1639),
.B(n_244),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1495),
.Y(n_2002)
);

BUFx2_ASAP7_75t_L g2003 ( 
.A(n_1519),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1495),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1519),
.Y(n_2005)
);

OAI22xp5_ASAP7_75t_SL g2006 ( 
.A1(n_1663),
.A2(n_1427),
.B1(n_1249),
.B2(n_1250),
.Y(n_2006)
);

INVx1_ASAP7_75t_L g2007 ( 
.A(n_1495),
.Y(n_2007)
);

AND2x4_ASAP7_75t_L g2008 ( 
.A(n_1514),
.B(n_248),
.Y(n_2008)
);

INVx2_ASAP7_75t_L g2009 ( 
.A(n_1514),
.Y(n_2009)
);

NAND2xp5_ASAP7_75t_L g2010 ( 
.A(n_1514),
.B(n_751),
.Y(n_2010)
);

BUFx6f_ASAP7_75t_L g2011 ( 
.A(n_1514),
.Y(n_2011)
);

INVx1_ASAP7_75t_L g2012 ( 
.A(n_1525),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1525),
.B(n_755),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1525),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1525),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1538),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1538),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1538),
.Y(n_2018)
);

INVx1_ASAP7_75t_L g2019 ( 
.A(n_1538),
.Y(n_2019)
);

INVx1_ASAP7_75t_L g2020 ( 
.A(n_1556),
.Y(n_2020)
);

INVx2_ASAP7_75t_L g2021 ( 
.A(n_1726),
.Y(n_2021)
);

INVx2_ASAP7_75t_SL g2022 ( 
.A(n_1737),
.Y(n_2022)
);

INVx1_ASAP7_75t_SL g2023 ( 
.A(n_1748),
.Y(n_2023)
);

NAND2xp33_ASAP7_75t_L g2024 ( 
.A(n_1762),
.B(n_1619),
.Y(n_2024)
);

INVx1_ASAP7_75t_L g2025 ( 
.A(n_1870),
.Y(n_2025)
);

INVx1_ASAP7_75t_L g2026 ( 
.A(n_1870),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1871),
.Y(n_2027)
);

INVx1_ASAP7_75t_SL g2028 ( 
.A(n_1748),
.Y(n_2028)
);

AOI22xp33_ASAP7_75t_L g2029 ( 
.A1(n_1756),
.A2(n_1467),
.B1(n_1498),
.B2(n_1452),
.Y(n_2029)
);

NOR2x1p5_ASAP7_75t_L g2030 ( 
.A(n_1767),
.B(n_1624),
.Y(n_2030)
);

NOR2xp33_ASAP7_75t_SL g2031 ( 
.A(n_1943),
.B(n_1549),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1871),
.Y(n_2032)
);

NAND2xp5_ASAP7_75t_L g2033 ( 
.A(n_1957),
.B(n_1520),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1900),
.B(n_1536),
.Y(n_2034)
);

INVx2_ASAP7_75t_SL g2035 ( 
.A(n_1850),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1900),
.B(n_1690),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1805),
.B(n_1570),
.Y(n_2037)
);

INVx2_ASAP7_75t_L g2038 ( 
.A(n_1726),
.Y(n_2038)
);

INVx1_ASAP7_75t_L g2039 ( 
.A(n_1887),
.Y(n_2039)
);

INVx1_ASAP7_75t_L g2040 ( 
.A(n_1887),
.Y(n_2040)
);

INVx1_ASAP7_75t_L g2041 ( 
.A(n_1888),
.Y(n_2041)
);

INVx3_ASAP7_75t_L g2042 ( 
.A(n_1762),
.Y(n_2042)
);

INVx2_ASAP7_75t_SL g2043 ( 
.A(n_1850),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1972),
.B(n_1690),
.Y(n_2044)
);

AOI22xp5_ASAP7_75t_L g2045 ( 
.A1(n_1756),
.A2(n_1483),
.B1(n_1633),
.B2(n_1629),
.Y(n_2045)
);

HB1xp67_ASAP7_75t_L g2046 ( 
.A(n_1772),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1972),
.B(n_1690),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1888),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_L g2049 ( 
.A(n_1993),
.B(n_1949),
.Y(n_2049)
);

INVx3_ASAP7_75t_L g2050 ( 
.A(n_1762),
.Y(n_2050)
);

NOR3xp33_ASAP7_75t_L g2051 ( 
.A(n_1991),
.B(n_1749),
.C(n_1828),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1805),
.B(n_1581),
.Y(n_2052)
);

OAI21xp33_ASAP7_75t_L g2053 ( 
.A1(n_1991),
.A2(n_1474),
.B(n_1501),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1993),
.B(n_1629),
.Y(n_2054)
);

INVx2_ASAP7_75t_L g2055 ( 
.A(n_1729),
.Y(n_2055)
);

BUFx2_ASAP7_75t_L g2056 ( 
.A(n_1724),
.Y(n_2056)
);

AND2x6_ASAP7_75t_L g2057 ( 
.A(n_1728),
.B(n_1623),
.Y(n_2057)
);

NAND3xp33_ASAP7_75t_L g2058 ( 
.A(n_1828),
.B(n_1645),
.C(n_1641),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1889),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_L g2060 ( 
.A1(n_1728),
.A2(n_1467),
.B1(n_1498),
.B2(n_1452),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1998),
.B(n_2001),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_1889),
.Y(n_2062)
);

INVx1_ASAP7_75t_L g2063 ( 
.A(n_1890),
.Y(n_2063)
);

NOR2xp33_ASAP7_75t_L g2064 ( 
.A(n_1809),
.B(n_1692),
.Y(n_2064)
);

AO22x2_ASAP7_75t_L g2065 ( 
.A1(n_1988),
.A2(n_1854),
.B1(n_1774),
.B2(n_1776),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1998),
.B(n_1619),
.Y(n_2066)
);

OR2x6_ASAP7_75t_L g2067 ( 
.A(n_1767),
.B(n_1548),
.Y(n_2067)
);

AOI22xp33_ASAP7_75t_L g2068 ( 
.A1(n_1728),
.A2(n_1467),
.B1(n_1498),
.B2(n_1452),
.Y(n_2068)
);

INVx2_ASAP7_75t_SL g2069 ( 
.A(n_1850),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_L g2070 ( 
.A(n_1925),
.B(n_1629),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1890),
.Y(n_2071)
);

INVx2_ASAP7_75t_L g2072 ( 
.A(n_1729),
.Y(n_2072)
);

OAI22xp33_ASAP7_75t_L g2073 ( 
.A1(n_1799),
.A2(n_1630),
.B1(n_1695),
.B2(n_1687),
.Y(n_2073)
);

INVx1_ASAP7_75t_L g2074 ( 
.A(n_1893),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1731),
.Y(n_2075)
);

NOR2xp33_ASAP7_75t_L g2076 ( 
.A(n_1944),
.B(n_1628),
.Y(n_2076)
);

INVx2_ASAP7_75t_L g2077 ( 
.A(n_1731),
.Y(n_2077)
);

INVxp67_ASAP7_75t_SL g2078 ( 
.A(n_1762),
.Y(n_2078)
);

INVx2_ASAP7_75t_SL g2079 ( 
.A(n_1837),
.Y(n_2079)
);

INVx3_ASAP7_75t_L g2080 ( 
.A(n_1763),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_1925),
.B(n_1633),
.Y(n_2081)
);

INVx3_ASAP7_75t_L g2082 ( 
.A(n_1763),
.Y(n_2082)
);

INVx4_ASAP7_75t_L g2083 ( 
.A(n_1723),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1893),
.Y(n_2084)
);

AND2x2_ASAP7_75t_SL g2085 ( 
.A(n_2008),
.B(n_1714),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1735),
.Y(n_2086)
);

INVx2_ASAP7_75t_SL g2087 ( 
.A(n_1837),
.Y(n_2087)
);

AND2x2_ASAP7_75t_SL g2088 ( 
.A(n_2008),
.B(n_1714),
.Y(n_2088)
);

AND2x6_ASAP7_75t_L g2089 ( 
.A(n_1730),
.B(n_1623),
.Y(n_2089)
);

BUFx3_ASAP7_75t_L g2090 ( 
.A(n_1723),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1763),
.Y(n_2091)
);

BUFx2_ASAP7_75t_L g2092 ( 
.A(n_1928),
.Y(n_2092)
);

INVx2_ASAP7_75t_SL g2093 ( 
.A(n_1837),
.Y(n_2093)
);

INVx1_ASAP7_75t_L g2094 ( 
.A(n_1903),
.Y(n_2094)
);

BUFx10_ASAP7_75t_L g2095 ( 
.A(n_1930),
.Y(n_2095)
);

AOI22xp33_ASAP7_75t_L g2096 ( 
.A1(n_1730),
.A2(n_1467),
.B1(n_1498),
.B2(n_1452),
.Y(n_2096)
);

INVx2_ASAP7_75t_L g2097 ( 
.A(n_1735),
.Y(n_2097)
);

NOR2xp33_ASAP7_75t_L g2098 ( 
.A(n_1808),
.B(n_1642),
.Y(n_2098)
);

INVx2_ASAP7_75t_L g2099 ( 
.A(n_1744),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1998),
.B(n_2001),
.Y(n_2100)
);

INVx5_ASAP7_75t_L g2101 ( 
.A(n_1763),
.Y(n_2101)
);

AOI22xp33_ASAP7_75t_SL g2102 ( 
.A1(n_1845),
.A2(n_1619),
.B1(n_1632),
.B2(n_1626),
.Y(n_2102)
);

INVx2_ASAP7_75t_L g2103 ( 
.A(n_1744),
.Y(n_2103)
);

INVx3_ASAP7_75t_L g2104 ( 
.A(n_1765),
.Y(n_2104)
);

NAND2xp33_ASAP7_75t_L g2105 ( 
.A(n_1765),
.B(n_1626),
.Y(n_2105)
);

NOR2xp33_ASAP7_75t_L g2106 ( 
.A(n_1740),
.B(n_1669),
.Y(n_2106)
);

INVx2_ASAP7_75t_L g2107 ( 
.A(n_1746),
.Y(n_2107)
);

INVx2_ASAP7_75t_L g2108 ( 
.A(n_1746),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_2001),
.B(n_1626),
.Y(n_2109)
);

AOI22xp5_ASAP7_75t_L g2110 ( 
.A1(n_1826),
.A2(n_1483),
.B1(n_1682),
.B2(n_1633),
.Y(n_2110)
);

INVx3_ASAP7_75t_L g2111 ( 
.A(n_1765),
.Y(n_2111)
);

BUFx3_ASAP7_75t_L g2112 ( 
.A(n_1723),
.Y(n_2112)
);

AND2x6_ASAP7_75t_L g2113 ( 
.A(n_1730),
.B(n_1627),
.Y(n_2113)
);

NAND2xp33_ASAP7_75t_SL g2114 ( 
.A(n_1930),
.B(n_1686),
.Y(n_2114)
);

INVx3_ASAP7_75t_L g2115 ( 
.A(n_1765),
.Y(n_2115)
);

INVx1_ASAP7_75t_L g2116 ( 
.A(n_1903),
.Y(n_2116)
);

AND2x6_ASAP7_75t_L g2117 ( 
.A(n_1739),
.B(n_1627),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_1751),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_L g2119 ( 
.A1(n_1739),
.A2(n_1467),
.B1(n_1498),
.B2(n_1452),
.Y(n_2119)
);

BUFx3_ASAP7_75t_L g2120 ( 
.A(n_1723),
.Y(n_2120)
);

AND2x4_ASAP7_75t_L g2121 ( 
.A(n_1905),
.B(n_1626),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1906),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1751),
.Y(n_2123)
);

INVx1_ASAP7_75t_L g2124 ( 
.A(n_1906),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_1752),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_1752),
.Y(n_2126)
);

NOR2xp33_ASAP7_75t_L g2127 ( 
.A(n_1959),
.B(n_1675),
.Y(n_2127)
);

NAND2xp5_ASAP7_75t_L g2128 ( 
.A(n_1961),
.B(n_1682),
.Y(n_2128)
);

INVx2_ASAP7_75t_L g2129 ( 
.A(n_1755),
.Y(n_2129)
);

INVx2_ASAP7_75t_L g2130 ( 
.A(n_1755),
.Y(n_2130)
);

BUFx3_ASAP7_75t_L g2131 ( 
.A(n_1772),
.Y(n_2131)
);

INVx3_ASAP7_75t_L g2132 ( 
.A(n_1769),
.Y(n_2132)
);

INVx2_ASAP7_75t_SL g2133 ( 
.A(n_1841),
.Y(n_2133)
);

AO21x2_ASAP7_75t_L g2134 ( 
.A1(n_1733),
.A2(n_1493),
.B(n_1568),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1961),
.B(n_1682),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_SL g2136 ( 
.A(n_1769),
.B(n_1632),
.Y(n_2136)
);

BUFx3_ASAP7_75t_L g2137 ( 
.A(n_1827),
.Y(n_2137)
);

NAND2xp5_ASAP7_75t_L g2138 ( 
.A(n_1846),
.B(n_1708),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_1757),
.Y(n_2139)
);

INVx3_ASAP7_75t_L g2140 ( 
.A(n_1769),
.Y(n_2140)
);

BUFx3_ASAP7_75t_L g2141 ( 
.A(n_1827),
.Y(n_2141)
);

AND2x6_ASAP7_75t_L g2142 ( 
.A(n_1739),
.B(n_1632),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1757),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_1909),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1741),
.B(n_1708),
.Y(n_2145)
);

NAND2xp5_ASAP7_75t_L g2146 ( 
.A(n_1897),
.B(n_1720),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1909),
.Y(n_2147)
);

INVx2_ASAP7_75t_SL g2148 ( 
.A(n_1841),
.Y(n_2148)
);

NOR2xp33_ASAP7_75t_L g2149 ( 
.A(n_1959),
.B(n_1630),
.Y(n_2149)
);

INVx4_ASAP7_75t_L g2150 ( 
.A(n_1930),
.Y(n_2150)
);

INVx5_ASAP7_75t_L g2151 ( 
.A(n_1769),
.Y(n_2151)
);

INVx3_ASAP7_75t_L g2152 ( 
.A(n_1788),
.Y(n_2152)
);

OAI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_1965),
.A2(n_1671),
.B1(n_1644),
.B2(n_1687),
.Y(n_2153)
);

CKINVDCx11_ASAP7_75t_R g2154 ( 
.A(n_1928),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1973),
.B(n_1720),
.Y(n_2155)
);

XNOR2xp5_ASAP7_75t_L g2156 ( 
.A(n_1863),
.B(n_1540),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_1775),
.A2(n_1720),
.B1(n_1493),
.B2(n_707),
.Y(n_2157)
);

INVx4_ASAP7_75t_L g2158 ( 
.A(n_1788),
.Y(n_2158)
);

INVx1_ASAP7_75t_L g2159 ( 
.A(n_1910),
.Y(n_2159)
);

NAND2xp5_ASAP7_75t_L g2160 ( 
.A(n_1802),
.B(n_1556),
.Y(n_2160)
);

NOR3xp33_ASAP7_75t_L g2161 ( 
.A(n_1936),
.B(n_1680),
.C(n_1655),
.Y(n_2161)
);

BUFx6f_ASAP7_75t_L g2162 ( 
.A(n_1788),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_1910),
.Y(n_2163)
);

NAND2xp5_ASAP7_75t_SL g2164 ( 
.A(n_1788),
.B(n_1632),
.Y(n_2164)
);

INVx1_ASAP7_75t_L g2165 ( 
.A(n_1918),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1802),
.B(n_1556),
.Y(n_2166)
);

BUFx6f_ASAP7_75t_L g2167 ( 
.A(n_1791),
.Y(n_2167)
);

INVx2_ASAP7_75t_L g2168 ( 
.A(n_1775),
.Y(n_2168)
);

NOR2xp33_ASAP7_75t_L g2169 ( 
.A(n_1760),
.B(n_1517),
.Y(n_2169)
);

INVx4_ASAP7_75t_L g2170 ( 
.A(n_1791),
.Y(n_2170)
);

INVx4_ASAP7_75t_L g2171 ( 
.A(n_1791),
.Y(n_2171)
);

NAND2xp5_ASAP7_75t_SL g2172 ( 
.A(n_1791),
.B(n_1674),
.Y(n_2172)
);

INVx1_ASAP7_75t_SL g2173 ( 
.A(n_1771),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1899),
.B(n_1556),
.Y(n_2174)
);

NAND2xp5_ASAP7_75t_L g2175 ( 
.A(n_1899),
.B(n_1560),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_1918),
.Y(n_2176)
);

HB1xp67_ASAP7_75t_SL g2177 ( 
.A(n_1851),
.Y(n_2177)
);

NAND2xp33_ASAP7_75t_L g2178 ( 
.A(n_1801),
.B(n_1674),
.Y(n_2178)
);

BUFx4f_ASAP7_75t_L g2179 ( 
.A(n_1989),
.Y(n_2179)
);

AND2x2_ASAP7_75t_L g2180 ( 
.A(n_1760),
.B(n_1586),
.Y(n_2180)
);

OR2x6_ASAP7_75t_L g2181 ( 
.A(n_1999),
.B(n_1548),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1919),
.Y(n_2182)
);

HB1xp67_ASAP7_75t_L g2183 ( 
.A(n_1913),
.Y(n_2183)
);

AND2x4_ASAP7_75t_L g2184 ( 
.A(n_1905),
.B(n_1674),
.Y(n_2184)
);

OAI22xp5_ASAP7_75t_L g2185 ( 
.A1(n_1929),
.A2(n_1931),
.B1(n_1935),
.B2(n_1933),
.Y(n_2185)
);

NAND2xp5_ASAP7_75t_SL g2186 ( 
.A(n_1801),
.B(n_1674),
.Y(n_2186)
);

INVx1_ASAP7_75t_L g2187 ( 
.A(n_1919),
.Y(n_2187)
);

INVx2_ASAP7_75t_SL g2188 ( 
.A(n_1841),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1932),
.Y(n_2189)
);

INVxp33_ASAP7_75t_L g2190 ( 
.A(n_1892),
.Y(n_2190)
);

INVx3_ASAP7_75t_L g2191 ( 
.A(n_1801),
.Y(n_2191)
);

BUFx2_ASAP7_75t_L g2192 ( 
.A(n_1754),
.Y(n_2192)
);

INVx2_ASAP7_75t_L g2193 ( 
.A(n_1778),
.Y(n_2193)
);

NOR2xp33_ASAP7_75t_L g2194 ( 
.A(n_1892),
.B(n_1517),
.Y(n_2194)
);

INVx2_ASAP7_75t_SL g2195 ( 
.A(n_1797),
.Y(n_2195)
);

INVxp33_ASAP7_75t_L g2196 ( 
.A(n_1734),
.Y(n_2196)
);

OAI22xp5_ASAP7_75t_L g2197 ( 
.A1(n_1940),
.A2(n_1671),
.B1(n_1644),
.B2(n_1695),
.Y(n_2197)
);

NOR2xp33_ASAP7_75t_L g2198 ( 
.A(n_1734),
.B(n_1618),
.Y(n_2198)
);

OR2x6_ASAP7_75t_L g2199 ( 
.A(n_1999),
.B(n_1555),
.Y(n_2199)
);

OAI22xp33_ASAP7_75t_L g2200 ( 
.A1(n_1908),
.A2(n_1681),
.B1(n_1688),
.B2(n_1686),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1932),
.Y(n_2201)
);

INVx2_ASAP7_75t_L g2202 ( 
.A(n_1778),
.Y(n_2202)
);

INVx2_ASAP7_75t_SL g2203 ( 
.A(n_1797),
.Y(n_2203)
);

INVx4_ASAP7_75t_L g2204 ( 
.A(n_1801),
.Y(n_2204)
);

INVx2_ASAP7_75t_L g2205 ( 
.A(n_1780),
.Y(n_2205)
);

INVx2_ASAP7_75t_L g2206 ( 
.A(n_1780),
.Y(n_2206)
);

INVx2_ASAP7_75t_L g2207 ( 
.A(n_1782),
.Y(n_2207)
);

BUFx10_ASAP7_75t_L g2208 ( 
.A(n_1876),
.Y(n_2208)
);

NAND3xp33_ASAP7_75t_L g2209 ( 
.A(n_1876),
.B(n_1886),
.C(n_1981),
.Y(n_2209)
);

INVx3_ASAP7_75t_L g2210 ( 
.A(n_1806),
.Y(n_2210)
);

INVx3_ASAP7_75t_L g2211 ( 
.A(n_1806),
.Y(n_2211)
);

NAND2xp5_ASAP7_75t_L g2212 ( 
.A(n_1937),
.B(n_1560),
.Y(n_2212)
);

BUFx6f_ASAP7_75t_L g2213 ( 
.A(n_1806),
.Y(n_2213)
);

CKINVDCx5p33_ASAP7_75t_R g2214 ( 
.A(n_1943),
.Y(n_2214)
);

INVx3_ASAP7_75t_L g2215 ( 
.A(n_1806),
.Y(n_2215)
);

INVx2_ASAP7_75t_L g2216 ( 
.A(n_1782),
.Y(n_2216)
);

NOR2xp33_ASAP7_75t_L g2217 ( 
.A(n_1747),
.B(n_1618),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_1783),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_1937),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_1945),
.Y(n_2220)
);

AOI22xp33_ASAP7_75t_L g2221 ( 
.A1(n_1783),
.A2(n_705),
.B1(n_1622),
.B2(n_1613),
.Y(n_2221)
);

NAND2xp33_ASAP7_75t_L g2222 ( 
.A(n_1822),
.B(n_1681),
.Y(n_2222)
);

INVx2_ASAP7_75t_SL g2223 ( 
.A(n_1953),
.Y(n_2223)
);

AND2x6_ASAP7_75t_L g2224 ( 
.A(n_1902),
.B(n_1681),
.Y(n_2224)
);

INVx1_ASAP7_75t_L g2225 ( 
.A(n_1945),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1822),
.Y(n_2226)
);

INVx2_ASAP7_75t_L g2227 ( 
.A(n_1789),
.Y(n_2227)
);

NAND2xp33_ASAP7_75t_L g2228 ( 
.A(n_1822),
.B(n_1681),
.Y(n_2228)
);

AOI22xp5_ASAP7_75t_L g2229 ( 
.A1(n_1953),
.A2(n_1601),
.B1(n_1661),
.B2(n_1640),
.Y(n_2229)
);

INVx1_ASAP7_75t_L g2230 ( 
.A(n_1952),
.Y(n_2230)
);

INVx3_ASAP7_75t_L g2231 ( 
.A(n_1822),
.Y(n_2231)
);

INVx2_ASAP7_75t_L g2232 ( 
.A(n_1789),
.Y(n_2232)
);

INVx2_ASAP7_75t_L g2233 ( 
.A(n_1792),
.Y(n_2233)
);

XNOR2xp5_ASAP7_75t_L g2234 ( 
.A(n_2006),
.B(n_1540),
.Y(n_2234)
);

INVx2_ASAP7_75t_L g2235 ( 
.A(n_1792),
.Y(n_2235)
);

NAND2xp5_ASAP7_75t_L g2236 ( 
.A(n_1952),
.B(n_1560),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1956),
.Y(n_2237)
);

INVx1_ASAP7_75t_L g2238 ( 
.A(n_1956),
.Y(n_2238)
);

INVx4_ASAP7_75t_L g2239 ( 
.A(n_1838),
.Y(n_2239)
);

INVx2_ASAP7_75t_L g2240 ( 
.A(n_1793),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1960),
.Y(n_2241)
);

CKINVDCx20_ASAP7_75t_R g2242 ( 
.A(n_1795),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1793),
.Y(n_2243)
);

XNOR2xp5_ASAP7_75t_L g2244 ( 
.A(n_1938),
.B(n_1554),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_1960),
.Y(n_2245)
);

AOI22xp5_ASAP7_75t_L g2246 ( 
.A1(n_1902),
.A2(n_1678),
.B1(n_1666),
.B2(n_1560),
.Y(n_2246)
);

NAND2xp5_ASAP7_75t_L g2247 ( 
.A(n_1969),
.B(n_1574),
.Y(n_2247)
);

INVxp33_ASAP7_75t_L g2248 ( 
.A(n_1747),
.Y(n_2248)
);

INVx2_ASAP7_75t_L g2249 ( 
.A(n_1800),
.Y(n_2249)
);

OAI22xp5_ASAP7_75t_L g2250 ( 
.A1(n_1902),
.A2(n_1691),
.B1(n_1694),
.B2(n_1683),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_SL g2251 ( 
.A(n_1838),
.B(n_1686),
.Y(n_2251)
);

AOI22xp33_ASAP7_75t_L g2252 ( 
.A1(n_1800),
.A2(n_1803),
.B1(n_2008),
.B2(n_1969),
.Y(n_2252)
);

OR2x2_ASAP7_75t_L g2253 ( 
.A(n_1771),
.B(n_1706),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_1913),
.B(n_1659),
.Y(n_2254)
);

INVx1_ASAP7_75t_L g2255 ( 
.A(n_1803),
.Y(n_2255)
);

NOR2xp33_ASAP7_75t_L g2256 ( 
.A(n_1921),
.B(n_1659),
.Y(n_2256)
);

AND2x2_ASAP7_75t_SL g2257 ( 
.A(n_1922),
.B(n_1709),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_SL g2258 ( 
.A(n_1838),
.B(n_1686),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1786),
.B(n_1787),
.Y(n_2259)
);

INVx2_ASAP7_75t_L g2260 ( 
.A(n_1807),
.Y(n_2260)
);

NOR2xp33_ASAP7_75t_L g2261 ( 
.A(n_1921),
.B(n_1685),
.Y(n_2261)
);

NAND2xp5_ASAP7_75t_SL g2262 ( 
.A(n_1838),
.B(n_1688),
.Y(n_2262)
);

OR2x6_ASAP7_75t_L g2263 ( 
.A(n_2003),
.B(n_1555),
.Y(n_2263)
);

INVx2_ASAP7_75t_L g2264 ( 
.A(n_1807),
.Y(n_2264)
);

OR2x6_ASAP7_75t_L g2265 ( 
.A(n_2003),
.B(n_1555),
.Y(n_2265)
);

BUFx2_ASAP7_75t_L g2266 ( 
.A(n_1811),
.Y(n_2266)
);

AND2x6_ASAP7_75t_L g2267 ( 
.A(n_1743),
.B(n_1688),
.Y(n_2267)
);

INVx5_ASAP7_75t_L g2268 ( 
.A(n_1839),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_L g2269 ( 
.A(n_1839),
.B(n_1688),
.Y(n_2269)
);

INVx1_ASAP7_75t_L g2270 ( 
.A(n_1942),
.Y(n_2270)
);

INVx1_ASAP7_75t_L g2271 ( 
.A(n_1951),
.Y(n_2271)
);

NAND2xp5_ASAP7_75t_SL g2272 ( 
.A(n_1839),
.B(n_1689),
.Y(n_2272)
);

OR2x2_ASAP7_75t_L g2273 ( 
.A(n_1777),
.B(n_1719),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_1812),
.Y(n_2274)
);

BUFx6f_ASAP7_75t_L g2275 ( 
.A(n_1839),
.Y(n_2275)
);

INVx1_ASAP7_75t_L g2276 ( 
.A(n_1964),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_1968),
.B(n_1574),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_1722),
.Y(n_2278)
);

INVx3_ASAP7_75t_L g2279 ( 
.A(n_1865),
.Y(n_2279)
);

INVx3_ASAP7_75t_L g2280 ( 
.A(n_1865),
.Y(n_2280)
);

NAND2xp5_ASAP7_75t_SL g2281 ( 
.A(n_1865),
.B(n_1689),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_1725),
.Y(n_2282)
);

NOR2xp33_ASAP7_75t_L g2283 ( 
.A(n_1948),
.B(n_1685),
.Y(n_2283)
);

BUFx3_ASAP7_75t_L g2284 ( 
.A(n_1948),
.Y(n_2284)
);

INVx1_ASAP7_75t_L g2285 ( 
.A(n_1732),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_1794),
.B(n_1574),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1812),
.Y(n_2287)
);

XNOR2xp5_ASAP7_75t_L g2288 ( 
.A(n_1938),
.B(n_1554),
.Y(n_2288)
);

INVx1_ASAP7_75t_SL g2289 ( 
.A(n_1818),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_1736),
.Y(n_2290)
);

NAND2xp5_ASAP7_75t_L g2291 ( 
.A(n_1804),
.B(n_1574),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_1738),
.Y(n_2292)
);

AND2x2_ASAP7_75t_L g2293 ( 
.A(n_1844),
.B(n_1696),
.Y(n_2293)
);

AND2x2_ASAP7_75t_L g2294 ( 
.A(n_1844),
.B(n_1696),
.Y(n_2294)
);

INVx1_ASAP7_75t_SL g2295 ( 
.A(n_1996),
.Y(n_2295)
);

INVx2_ASAP7_75t_L g2296 ( 
.A(n_1843),
.Y(n_2296)
);

INVx4_ASAP7_75t_L g2297 ( 
.A(n_1865),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_1810),
.B(n_1611),
.Y(n_2298)
);

AOI22xp33_ASAP7_75t_L g2299 ( 
.A1(n_1727),
.A2(n_1862),
.B1(n_1994),
.B2(n_1922),
.Y(n_2299)
);

INVx2_ASAP7_75t_L g2300 ( 
.A(n_1843),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_1750),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1853),
.Y(n_2302)
);

INVx2_ASAP7_75t_L g2303 ( 
.A(n_1853),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1758),
.Y(n_2304)
);

NAND2xp5_ASAP7_75t_SL g2305 ( 
.A(n_1875),
.B(n_1689),
.Y(n_2305)
);

NAND2xp5_ASAP7_75t_L g2306 ( 
.A(n_1813),
.B(n_1611),
.Y(n_2306)
);

NAND2xp5_ASAP7_75t_L g2307 ( 
.A(n_1814),
.B(n_1611),
.Y(n_2307)
);

CKINVDCx5p33_ASAP7_75t_R g2308 ( 
.A(n_2000),
.Y(n_2308)
);

INVx8_ASAP7_75t_L g2309 ( 
.A(n_1915),
.Y(n_2309)
);

INVx1_ASAP7_75t_SL g2310 ( 
.A(n_1821),
.Y(n_2310)
);

CKINVDCx5p33_ASAP7_75t_R g2311 ( 
.A(n_2000),
.Y(n_2311)
);

INVx1_ASAP7_75t_L g2312 ( 
.A(n_1759),
.Y(n_2312)
);

INVx1_ASAP7_75t_SL g2313 ( 
.A(n_1830),
.Y(n_2313)
);

AOI21x1_ASAP7_75t_L g2314 ( 
.A1(n_1819),
.A2(n_1622),
.B(n_1613),
.Y(n_2314)
);

INVx5_ASAP7_75t_L g2315 ( 
.A(n_1875),
.Y(n_2315)
);

NOR2xp33_ASAP7_75t_L g2316 ( 
.A(n_1790),
.B(n_1650),
.Y(n_2316)
);

INVx1_ASAP7_75t_L g2317 ( 
.A(n_1761),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1860),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_1823),
.B(n_1611),
.Y(n_2319)
);

INVx2_ASAP7_75t_SL g2320 ( 
.A(n_1831),
.Y(n_2320)
);

NOR2xp33_ASAP7_75t_L g2321 ( 
.A(n_1831),
.B(n_1857),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_1727),
.A2(n_1646),
.B1(n_686),
.B2(n_692),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_1824),
.B(n_1612),
.Y(n_2323)
);

NAND2xp5_ASAP7_75t_L g2324 ( 
.A(n_1834),
.B(n_1612),
.Y(n_2324)
);

AND2x2_ASAP7_75t_L g2325 ( 
.A(n_2180),
.B(n_1835),
.Y(n_2325)
);

BUFx6f_ASAP7_75t_SL g2326 ( 
.A(n_2181),
.Y(n_2326)
);

INVx1_ASAP7_75t_L g2327 ( 
.A(n_2025),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2033),
.B(n_2098),
.Y(n_2328)
);

INVx2_ASAP7_75t_L g2329 ( 
.A(n_2021),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_SL g2330 ( 
.A(n_2200),
.B(n_1689),
.Y(n_2330)
);

NAND2xp5_ASAP7_75t_L g2331 ( 
.A(n_2098),
.B(n_2106),
.Y(n_2331)
);

INVx2_ASAP7_75t_SL g2332 ( 
.A(n_2022),
.Y(n_2332)
);

INVx1_ASAP7_75t_L g2333 ( 
.A(n_2026),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_2027),
.Y(n_2334)
);

NOR2xp67_ASAP7_75t_L g2335 ( 
.A(n_2150),
.B(n_1438),
.Y(n_2335)
);

NAND2xp5_ASAP7_75t_SL g2336 ( 
.A(n_2200),
.B(n_1643),
.Y(n_2336)
);

INVx1_ASAP7_75t_L g2337 ( 
.A(n_2032),
.Y(n_2337)
);

OR2x2_ASAP7_75t_L g2338 ( 
.A(n_2173),
.B(n_1700),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_SL g2339 ( 
.A(n_2169),
.B(n_1643),
.Y(n_2339)
);

INVx2_ASAP7_75t_L g2340 ( 
.A(n_2021),
.Y(n_2340)
);

NAND2xp5_ASAP7_75t_SL g2341 ( 
.A(n_2169),
.B(n_1647),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_2190),
.B(n_2064),
.Y(n_2342)
);

NOR2xp33_ASAP7_75t_L g2343 ( 
.A(n_2190),
.B(n_1816),
.Y(n_2343)
);

INVx4_ASAP7_75t_SL g2344 ( 
.A(n_2224),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2106),
.B(n_1922),
.Y(n_2345)
);

INVx2_ASAP7_75t_L g2346 ( 
.A(n_2038),
.Y(n_2346)
);

AND2x2_ASAP7_75t_L g2347 ( 
.A(n_2037),
.B(n_1835),
.Y(n_2347)
);

NAND2xp5_ASAP7_75t_L g2348 ( 
.A(n_2127),
.B(n_1840),
.Y(n_2348)
);

INVx2_ASAP7_75t_SL g2349 ( 
.A(n_2131),
.Y(n_2349)
);

NOR2xp33_ASAP7_75t_L g2350 ( 
.A(n_2064),
.B(n_1816),
.Y(n_2350)
);

AND2x2_ASAP7_75t_L g2351 ( 
.A(n_2052),
.B(n_1833),
.Y(n_2351)
);

INVx2_ASAP7_75t_L g2352 ( 
.A(n_2038),
.Y(n_2352)
);

NOR2xp33_ASAP7_75t_L g2353 ( 
.A(n_2194),
.B(n_1891),
.Y(n_2353)
);

XOR2xp5_ASAP7_75t_L g2354 ( 
.A(n_2242),
.B(n_1576),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2055),
.Y(n_2355)
);

NAND2xp5_ASAP7_75t_SL g2356 ( 
.A(n_2198),
.B(n_1647),
.Y(n_2356)
);

BUFx6f_ASAP7_75t_L g2357 ( 
.A(n_2162),
.Y(n_2357)
);

INVx2_ASAP7_75t_SL g2358 ( 
.A(n_2131),
.Y(n_2358)
);

NOR2xp33_ASAP7_75t_L g2359 ( 
.A(n_2194),
.B(n_1891),
.Y(n_2359)
);

NAND2xp5_ASAP7_75t_L g2360 ( 
.A(n_2127),
.B(n_1842),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2039),
.Y(n_2361)
);

BUFx6f_ASAP7_75t_L g2362 ( 
.A(n_2162),
.Y(n_2362)
);

NAND2xp5_ASAP7_75t_L g2363 ( 
.A(n_2034),
.B(n_1848),
.Y(n_2363)
);

NAND2xp5_ASAP7_75t_SL g2364 ( 
.A(n_2198),
.B(n_1651),
.Y(n_2364)
);

AO221x1_ASAP7_75t_L g2365 ( 
.A1(n_2073),
.A2(n_1717),
.B1(n_1715),
.B2(n_1849),
.C(n_1489),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_SL g2366 ( 
.A(n_2217),
.B(n_1651),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2076),
.B(n_1926),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_2040),
.Y(n_2368)
);

INVx2_ASAP7_75t_L g2369 ( 
.A(n_2055),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_SL g2370 ( 
.A(n_2217),
.B(n_1649),
.Y(n_2370)
);

NOR2xp33_ASAP7_75t_L g2371 ( 
.A(n_2076),
.B(n_1926),
.Y(n_2371)
);

NAND2xp5_ASAP7_75t_SL g2372 ( 
.A(n_2254),
.B(n_1652),
.Y(n_2372)
);

INVx1_ASAP7_75t_L g2373 ( 
.A(n_2041),
.Y(n_2373)
);

INVx1_ASAP7_75t_L g2374 ( 
.A(n_2048),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2059),
.Y(n_2375)
);

BUFx6f_ASAP7_75t_L g2376 ( 
.A(n_2162),
.Y(n_2376)
);

INVx1_ASAP7_75t_L g2377 ( 
.A(n_2062),
.Y(n_2377)
);

INVx4_ASAP7_75t_L g2378 ( 
.A(n_2067),
.Y(n_2378)
);

INVxp67_ASAP7_75t_SL g2379 ( 
.A(n_2252),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2051),
.B(n_1852),
.Y(n_2380)
);

NAND2xp5_ASAP7_75t_L g2381 ( 
.A(n_2051),
.B(n_1855),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_2063),
.Y(n_2382)
);

INVx2_ASAP7_75t_L g2383 ( 
.A(n_2086),
.Y(n_2383)
);

NAND2xp5_ASAP7_75t_L g2384 ( 
.A(n_2049),
.B(n_1858),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2071),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_SL g2386 ( 
.A(n_2254),
.B(n_1654),
.Y(n_2386)
);

NOR3xp33_ASAP7_75t_L g2387 ( 
.A(n_2053),
.B(n_1712),
.C(n_1710),
.Y(n_2387)
);

NAND2xp5_ASAP7_75t_SL g2388 ( 
.A(n_2256),
.B(n_1657),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_2160),
.B(n_1859),
.Y(n_2389)
);

INVxp67_ASAP7_75t_L g2390 ( 
.A(n_2056),
.Y(n_2390)
);

INVx1_ASAP7_75t_SL g2391 ( 
.A(n_2023),
.Y(n_2391)
);

NAND3xp33_ASAP7_75t_L g2392 ( 
.A(n_2209),
.B(n_1693),
.C(n_1701),
.Y(n_2392)
);

AND2x2_ASAP7_75t_L g2393 ( 
.A(n_2149),
.B(n_1861),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2074),
.Y(n_2394)
);

INVx1_ASAP7_75t_L g2395 ( 
.A(n_2084),
.Y(n_2395)
);

NOR2xp33_ASAP7_75t_SL g2396 ( 
.A(n_2085),
.B(n_1438),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_2085),
.B(n_1864),
.Y(n_2397)
);

INVx2_ASAP7_75t_SL g2398 ( 
.A(n_2137),
.Y(n_2398)
);

INVx1_ASAP7_75t_L g2399 ( 
.A(n_2094),
.Y(n_2399)
);

BUFx6f_ASAP7_75t_L g2400 ( 
.A(n_2162),
.Y(n_2400)
);

OR2x6_ASAP7_75t_L g2401 ( 
.A(n_2067),
.B(n_1715),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_2116),
.Y(n_2402)
);

NOR2xp67_ASAP7_75t_L g2403 ( 
.A(n_2150),
.B(n_1532),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_2122),
.Y(n_2404)
);

NOR2xp67_ASAP7_75t_L g2405 ( 
.A(n_2308),
.B(n_1532),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2124),
.Y(n_2406)
);

INVx1_ASAP7_75t_L g2407 ( 
.A(n_2144),
.Y(n_2407)
);

NAND2xp5_ASAP7_75t_L g2408 ( 
.A(n_2088),
.B(n_1868),
.Y(n_2408)
);

INVx2_ASAP7_75t_SL g2409 ( 
.A(n_2137),
.Y(n_2409)
);

INVxp33_ASAP7_75t_L g2410 ( 
.A(n_2253),
.Y(n_2410)
);

NAND2xp5_ASAP7_75t_L g2411 ( 
.A(n_2166),
.B(n_2149),
.Y(n_2411)
);

NOR2xp67_ASAP7_75t_SL g2412 ( 
.A(n_2101),
.B(n_1561),
.Y(n_2412)
);

NAND2xp5_ASAP7_75t_SL g2413 ( 
.A(n_2256),
.B(n_1658),
.Y(n_2413)
);

BUFx3_ASAP7_75t_L g2414 ( 
.A(n_2141),
.Y(n_2414)
);

INVx1_ASAP7_75t_L g2415 ( 
.A(n_2147),
.Y(n_2415)
);

NOR2xp33_ASAP7_75t_L g2416 ( 
.A(n_2196),
.B(n_1660),
.Y(n_2416)
);

NAND2xp5_ASAP7_75t_L g2417 ( 
.A(n_2088),
.B(n_1872),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2086),
.Y(n_2418)
);

AOI22xp33_ASAP7_75t_L g2419 ( 
.A1(n_2058),
.A2(n_1950),
.B1(n_1971),
.B2(n_1862),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2061),
.B(n_1874),
.Y(n_2420)
);

NAND2xp5_ASAP7_75t_L g2421 ( 
.A(n_2061),
.B(n_1878),
.Y(n_2421)
);

NOR2xp33_ASAP7_75t_L g2422 ( 
.A(n_2196),
.B(n_2248),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2195),
.Y(n_2423)
);

NAND2xp5_ASAP7_75t_SL g2424 ( 
.A(n_2121),
.B(n_1662),
.Y(n_2424)
);

INVx2_ASAP7_75t_L g2425 ( 
.A(n_2097),
.Y(n_2425)
);

NOR2xp33_ASAP7_75t_L g2426 ( 
.A(n_2248),
.B(n_1664),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2100),
.B(n_1880),
.Y(n_2427)
);

NOR2xp33_ASAP7_75t_L g2428 ( 
.A(n_2028),
.B(n_1667),
.Y(n_2428)
);

NAND2xp5_ASAP7_75t_SL g2429 ( 
.A(n_2121),
.B(n_1668),
.Y(n_2429)
);

NOR2xp33_ASAP7_75t_L g2430 ( 
.A(n_2273),
.B(n_2261),
.Y(n_2430)
);

AND3x4_ASAP7_75t_L g2431 ( 
.A(n_2161),
.B(n_1989),
.C(n_1977),
.Y(n_2431)
);

INVx2_ASAP7_75t_L g2432 ( 
.A(n_2097),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_2159),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2100),
.B(n_1881),
.Y(n_2434)
);

NAND2xp5_ASAP7_75t_SL g2435 ( 
.A(n_2184),
.B(n_1672),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_2261),
.B(n_1673),
.Y(n_2436)
);

OR2x6_ASAP7_75t_L g2437 ( 
.A(n_2067),
.B(n_1715),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2099),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2099),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_SL g2440 ( 
.A(n_2184),
.B(n_1677),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_L g2441 ( 
.A(n_2145),
.B(n_1895),
.Y(n_2441)
);

A2O1A1Ixp33_ASAP7_75t_L g2442 ( 
.A1(n_2321),
.A2(n_1901),
.B(n_1907),
.C(n_1896),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2174),
.B(n_1911),
.Y(n_2443)
);

CKINVDCx20_ASAP7_75t_R g2444 ( 
.A(n_2242),
.Y(n_2444)
);

AO221x1_ASAP7_75t_L g2445 ( 
.A1(n_2073),
.A2(n_1717),
.B1(n_1715),
.B2(n_1704),
.C(n_1713),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2103),
.Y(n_2446)
);

AND2x2_ASAP7_75t_L g2447 ( 
.A(n_2203),
.B(n_1898),
.Y(n_2447)
);

INVxp67_ASAP7_75t_SL g2448 ( 
.A(n_2252),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2163),
.Y(n_2449)
);

NOR2xp67_ASAP7_75t_L g2450 ( 
.A(n_2311),
.B(n_1684),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2175),
.B(n_1914),
.Y(n_2451)
);

INVx8_ASAP7_75t_L g2452 ( 
.A(n_2181),
.Y(n_2452)
);

AND2x2_ASAP7_75t_L g2453 ( 
.A(n_2141),
.B(n_1979),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_SL g2454 ( 
.A(n_2102),
.B(n_1679),
.Y(n_2454)
);

INVx2_ASAP7_75t_L g2455 ( 
.A(n_2103),
.Y(n_2455)
);

NOR2xp33_ASAP7_75t_L g2456 ( 
.A(n_2283),
.B(n_1703),
.Y(n_2456)
);

INVx2_ASAP7_75t_SL g2457 ( 
.A(n_2284),
.Y(n_2457)
);

NAND2xp33_ASAP7_75t_L g2458 ( 
.A(n_2224),
.B(n_1915),
.Y(n_2458)
);

BUFx6f_ASAP7_75t_L g2459 ( 
.A(n_2167),
.Y(n_2459)
);

HB1xp67_ASAP7_75t_L g2460 ( 
.A(n_2284),
.Y(n_2460)
);

BUFx2_ASAP7_75t_L g2461 ( 
.A(n_2046),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2165),
.Y(n_2462)
);

NOR2xp33_ASAP7_75t_L g2463 ( 
.A(n_2283),
.B(n_1227),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_SL g2464 ( 
.A(n_2102),
.B(n_1637),
.Y(n_2464)
);

NOR2xp33_ASAP7_75t_L g2465 ( 
.A(n_2208),
.B(n_1249),
.Y(n_2465)
);

NAND3xp33_ASAP7_75t_L g2466 ( 
.A(n_2321),
.B(n_1867),
.C(n_1857),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2107),
.Y(n_2467)
);

NOR2xp33_ASAP7_75t_L g2468 ( 
.A(n_2208),
.B(n_2289),
.Y(n_2468)
);

AND2x2_ASAP7_75t_L g2469 ( 
.A(n_2046),
.B(n_1982),
.Y(n_2469)
);

NAND2xp5_ASAP7_75t_L g2470 ( 
.A(n_2155),
.B(n_1917),
.Y(n_2470)
);

AND2x2_ASAP7_75t_L g2471 ( 
.A(n_2183),
.B(n_2293),
.Y(n_2471)
);

OR2x2_ASAP7_75t_L g2472 ( 
.A(n_2295),
.B(n_1717),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2176),
.Y(n_2473)
);

NOR2xp33_ASAP7_75t_L g2474 ( 
.A(n_2316),
.B(n_1250),
.Y(n_2474)
);

NAND2xp33_ASAP7_75t_L g2475 ( 
.A(n_2224),
.B(n_1915),
.Y(n_2475)
);

INVx1_ASAP7_75t_L g2476 ( 
.A(n_2182),
.Y(n_2476)
);

INVx1_ASAP7_75t_L g2477 ( 
.A(n_2187),
.Y(n_2477)
);

NAND2xp5_ASAP7_75t_L g2478 ( 
.A(n_2044),
.B(n_1920),
.Y(n_2478)
);

NOR2xp33_ASAP7_75t_L g2479 ( 
.A(n_2316),
.B(n_1252),
.Y(n_2479)
);

INVx2_ASAP7_75t_L g2480 ( 
.A(n_2107),
.Y(n_2480)
);

NOR2xp33_ASAP7_75t_L g2481 ( 
.A(n_2183),
.B(n_2229),
.Y(n_2481)
);

BUFx5_ASAP7_75t_L g2482 ( 
.A(n_2057),
.Y(n_2482)
);

AND2x2_ASAP7_75t_L g2483 ( 
.A(n_2294),
.B(n_1454),
.Y(n_2483)
);

INVx2_ASAP7_75t_L g2484 ( 
.A(n_2108),
.Y(n_2484)
);

NAND2xp5_ASAP7_75t_L g2485 ( 
.A(n_2047),
.B(n_1923),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2320),
.B(n_1252),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2031),
.B(n_1255),
.Y(n_2487)
);

INVx2_ASAP7_75t_L g2488 ( 
.A(n_2108),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2189),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2310),
.B(n_1784),
.Y(n_2490)
);

INVxp33_ASAP7_75t_L g2491 ( 
.A(n_2092),
.Y(n_2491)
);

NAND2xp5_ASAP7_75t_L g2492 ( 
.A(n_2257),
.B(n_1924),
.Y(n_2492)
);

NOR2xp67_ASAP7_75t_L g2493 ( 
.A(n_2214),
.B(n_1684),
.Y(n_2493)
);

NAND2xp5_ASAP7_75t_L g2494 ( 
.A(n_2257),
.B(n_1950),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2201),
.Y(n_2495)
);

NAND2xp5_ASAP7_75t_L g2496 ( 
.A(n_2224),
.B(n_1950),
.Y(n_2496)
);

CKINVDCx20_ASAP7_75t_R g2497 ( 
.A(n_2154),
.Y(n_2497)
);

NAND2xp5_ASAP7_75t_L g2498 ( 
.A(n_2224),
.B(n_1971),
.Y(n_2498)
);

NAND2xp5_ASAP7_75t_SL g2499 ( 
.A(n_2246),
.B(n_1916),
.Y(n_2499)
);

NAND2xp5_ASAP7_75t_L g2500 ( 
.A(n_2153),
.B(n_1971),
.Y(n_2500)
);

INVx2_ASAP7_75t_L g2501 ( 
.A(n_2168),
.Y(n_2501)
);

HB1xp67_ASAP7_75t_L g2502 ( 
.A(n_2181),
.Y(n_2502)
);

BUFx5_ASAP7_75t_L g2503 ( 
.A(n_2057),
.Y(n_2503)
);

INVx2_ASAP7_75t_L g2504 ( 
.A(n_2168),
.Y(n_2504)
);

AOI221xp5_ASAP7_75t_L g2505 ( 
.A1(n_2322),
.A2(n_1977),
.B1(n_1593),
.B2(n_1884),
.C(n_480),
.Y(n_2505)
);

INVx1_ASAP7_75t_L g2506 ( 
.A(n_2219),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2220),
.Y(n_2507)
);

HB1xp67_ASAP7_75t_L g2508 ( 
.A(n_2199),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2167),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2225),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2079),
.B(n_1784),
.Y(n_2511)
);

INVx3_ASAP7_75t_L g2512 ( 
.A(n_2167),
.Y(n_2512)
);

NAND2xp5_ASAP7_75t_L g2513 ( 
.A(n_2036),
.B(n_2002),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2054),
.B(n_2002),
.Y(n_2514)
);

INVx2_ASAP7_75t_L g2515 ( 
.A(n_2205),
.Y(n_2515)
);

INVx3_ASAP7_75t_L g2516 ( 
.A(n_2167),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2299),
.B(n_2009),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_2230),
.Y(n_2518)
);

INVxp67_ASAP7_75t_L g2519 ( 
.A(n_2192),
.Y(n_2519)
);

AND2x2_ASAP7_75t_L g2520 ( 
.A(n_2313),
.B(n_1784),
.Y(n_2520)
);

BUFx3_ASAP7_75t_L g2521 ( 
.A(n_2199),
.Y(n_2521)
);

NAND2xp33_ASAP7_75t_L g2522 ( 
.A(n_2267),
.B(n_1915),
.Y(n_2522)
);

INVx3_ASAP7_75t_L g2523 ( 
.A(n_2213),
.Y(n_2523)
);

NOR2xp33_ASAP7_75t_L g2524 ( 
.A(n_2223),
.B(n_1255),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2213),
.Y(n_2525)
);

BUFx6f_ASAP7_75t_L g2526 ( 
.A(n_2213),
.Y(n_2526)
);

NAND2xp5_ASAP7_75t_L g2527 ( 
.A(n_2299),
.B(n_2009),
.Y(n_2527)
);

NAND2xp5_ASAP7_75t_L g2528 ( 
.A(n_2138),
.B(n_2014),
.Y(n_2528)
);

INVxp67_ASAP7_75t_L g2529 ( 
.A(n_2266),
.Y(n_2529)
);

INVx1_ASAP7_75t_L g2530 ( 
.A(n_2237),
.Y(n_2530)
);

NAND2xp33_ASAP7_75t_L g2531 ( 
.A(n_2267),
.B(n_1915),
.Y(n_2531)
);

NAND2xp5_ASAP7_75t_L g2532 ( 
.A(n_2146),
.B(n_2065),
.Y(n_2532)
);

INVxp67_ASAP7_75t_L g2533 ( 
.A(n_2185),
.Y(n_2533)
);

INVx1_ASAP7_75t_L g2534 ( 
.A(n_2238),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2205),
.Y(n_2535)
);

NAND2xp33_ASAP7_75t_L g2536 ( 
.A(n_2267),
.B(n_1915),
.Y(n_2536)
);

HB1xp67_ASAP7_75t_L g2537 ( 
.A(n_2199),
.Y(n_2537)
);

BUFx6f_ASAP7_75t_SL g2538 ( 
.A(n_2263),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_2241),
.Y(n_2539)
);

NOR2xp33_ASAP7_75t_L g2540 ( 
.A(n_2197),
.B(n_1277),
.Y(n_2540)
);

INVx2_ASAP7_75t_L g2541 ( 
.A(n_2206),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2245),
.Y(n_2542)
);

AOI221xp5_ASAP7_75t_L g2543 ( 
.A1(n_2322),
.A2(n_1884),
.B1(n_2005),
.B2(n_1847),
.C(n_1646),
.Y(n_2543)
);

INVx1_ASAP7_75t_L g2544 ( 
.A(n_2255),
.Y(n_2544)
);

BUFx8_ASAP7_75t_L g2545 ( 
.A(n_2035),
.Y(n_2545)
);

INVx1_ASAP7_75t_L g2546 ( 
.A(n_2206),
.Y(n_2546)
);

NAND3xp33_ASAP7_75t_L g2547 ( 
.A(n_2161),
.B(n_1867),
.C(n_1698),
.Y(n_2547)
);

BUFx6f_ASAP7_75t_L g2548 ( 
.A(n_2213),
.Y(n_2548)
);

NOR2xp33_ASAP7_75t_L g2549 ( 
.A(n_2250),
.B(n_1277),
.Y(n_2549)
);

NOR2x1p5_ASAP7_75t_L g2550 ( 
.A(n_2278),
.B(n_1576),
.Y(n_2550)
);

AOI22xp5_ASAP7_75t_L g2551 ( 
.A1(n_2179),
.A2(n_1847),
.B1(n_1885),
.B2(n_1883),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2207),
.Y(n_2552)
);

NAND2xp5_ASAP7_75t_SL g2553 ( 
.A(n_2179),
.B(n_1717),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_2065),
.B(n_2014),
.Y(n_2554)
);

NOR2xp33_ASAP7_75t_L g2555 ( 
.A(n_2066),
.B(n_1284),
.Y(n_2555)
);

NAND2xp5_ASAP7_75t_L g2556 ( 
.A(n_2065),
.B(n_2018),
.Y(n_2556)
);

NAND2xp5_ASAP7_75t_L g2557 ( 
.A(n_2070),
.B(n_2018),
.Y(n_2557)
);

INVx1_ASAP7_75t_L g2558 ( 
.A(n_2207),
.Y(n_2558)
);

NAND2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2043),
.B(n_1561),
.Y(n_2559)
);

NAND2xp5_ASAP7_75t_SL g2560 ( 
.A(n_2069),
.B(n_1561),
.Y(n_2560)
);

NAND2xp33_ASAP7_75t_SL g2561 ( 
.A(n_2030),
.B(n_2066),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2233),
.Y(n_2562)
);

NOR2xp33_ASAP7_75t_L g2563 ( 
.A(n_2109),
.B(n_1284),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2233),
.Y(n_2564)
);

INVx2_ASAP7_75t_SL g2565 ( 
.A(n_2263),
.Y(n_2565)
);

INVx1_ASAP7_75t_L g2566 ( 
.A(n_2235),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2235),
.Y(n_2567)
);

NAND2xp5_ASAP7_75t_L g2568 ( 
.A(n_2081),
.B(n_1997),
.Y(n_2568)
);

OR2x2_ASAP7_75t_L g2569 ( 
.A(n_2087),
.B(n_1589),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_SL g2570 ( 
.A(n_2114),
.B(n_1561),
.Y(n_2570)
);

AOI21xp5_ASAP7_75t_L g2571 ( 
.A1(n_2345),
.A2(n_2105),
.B(n_2024),
.Y(n_2571)
);

AOI22xp33_ASAP7_75t_SL g2572 ( 
.A1(n_2331),
.A2(n_1301),
.B1(n_1305),
.B2(n_1292),
.Y(n_2572)
);

NAND2xp5_ASAP7_75t_L g2573 ( 
.A(n_2331),
.B(n_2093),
.Y(n_2573)
);

OR2x2_ASAP7_75t_L g2574 ( 
.A(n_2328),
.B(n_2005),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2342),
.B(n_2393),
.Y(n_2575)
);

AND2x2_ASAP7_75t_L g2576 ( 
.A(n_2430),
.B(n_1753),
.Y(n_2576)
);

INVx3_ASAP7_75t_L g2577 ( 
.A(n_2357),
.Y(n_2577)
);

NOR2xp33_ASAP7_75t_L g2578 ( 
.A(n_2350),
.B(n_2367),
.Y(n_2578)
);

NAND2xp5_ASAP7_75t_L g2579 ( 
.A(n_2328),
.B(n_2188),
.Y(n_2579)
);

BUFx6f_ASAP7_75t_SL g2580 ( 
.A(n_2414),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2411),
.B(n_2133),
.Y(n_2581)
);

NAND2xp5_ASAP7_75t_L g2582 ( 
.A(n_2360),
.B(n_2148),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2327),
.Y(n_2583)
);

NAND2xp5_ASAP7_75t_L g2584 ( 
.A(n_2348),
.B(n_2282),
.Y(n_2584)
);

NAND2xp5_ASAP7_75t_L g2585 ( 
.A(n_2348),
.B(n_2285),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2329),
.Y(n_2586)
);

INVx2_ASAP7_75t_SL g2587 ( 
.A(n_2332),
.Y(n_2587)
);

NOR2xp33_ASAP7_75t_L g2588 ( 
.A(n_2371),
.B(n_1292),
.Y(n_2588)
);

NAND2xp5_ASAP7_75t_L g2589 ( 
.A(n_2345),
.B(n_2290),
.Y(n_2589)
);

NOR2xp33_ASAP7_75t_L g2590 ( 
.A(n_2353),
.B(n_1301),
.Y(n_2590)
);

NOR2xp33_ASAP7_75t_L g2591 ( 
.A(n_2359),
.B(n_1305),
.Y(n_2591)
);

NAND2xp5_ASAP7_75t_L g2592 ( 
.A(n_2436),
.B(n_2292),
.Y(n_2592)
);

A2O1A1Ixp33_ASAP7_75t_L g2593 ( 
.A1(n_2547),
.A2(n_2110),
.B(n_2109),
.C(n_2045),
.Y(n_2593)
);

OR2x6_ASAP7_75t_L g2594 ( 
.A(n_2452),
.B(n_2263),
.Y(n_2594)
);

AOI22xp33_ASAP7_75t_L g2595 ( 
.A1(n_2387),
.A2(n_1975),
.B1(n_1976),
.B2(n_2301),
.Y(n_2595)
);

O2A1O1Ixp33_ASAP7_75t_L g2596 ( 
.A1(n_2336),
.A2(n_1984),
.B(n_2269),
.C(n_1946),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2333),
.Y(n_2597)
);

INVx2_ASAP7_75t_L g2598 ( 
.A(n_2340),
.Y(n_2598)
);

CKINVDCx5p33_ASAP7_75t_R g2599 ( 
.A(n_2444),
.Y(n_2599)
);

HB1xp67_ASAP7_75t_L g2600 ( 
.A(n_2461),
.Y(n_2600)
);

NAND2xp5_ASAP7_75t_L g2601 ( 
.A(n_2384),
.B(n_2304),
.Y(n_2601)
);

AOI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2419),
.A2(n_2365),
.B1(n_2466),
.B2(n_2481),
.Y(n_2602)
);

NAND2xp5_ASAP7_75t_L g2603 ( 
.A(n_2363),
.B(n_2312),
.Y(n_2603)
);

BUFx6f_ASAP7_75t_L g2604 ( 
.A(n_2452),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2533),
.B(n_2317),
.Y(n_2605)
);

AND2x4_ASAP7_75t_L g2606 ( 
.A(n_2378),
.B(n_2090),
.Y(n_2606)
);

INVx4_ASAP7_75t_L g2607 ( 
.A(n_2452),
.Y(n_2607)
);

NAND2xp5_ASAP7_75t_SL g2608 ( 
.A(n_2428),
.B(n_2114),
.Y(n_2608)
);

CKINVDCx5p33_ASAP7_75t_R g2609 ( 
.A(n_2497),
.Y(n_2609)
);

BUFx6f_ASAP7_75t_L g2610 ( 
.A(n_2357),
.Y(n_2610)
);

NAND2xp5_ASAP7_75t_L g2611 ( 
.A(n_2483),
.B(n_2221),
.Y(n_2611)
);

INVx3_ASAP7_75t_L g2612 ( 
.A(n_2357),
.Y(n_2612)
);

AND2x2_ASAP7_75t_L g2613 ( 
.A(n_2471),
.B(n_1753),
.Y(n_2613)
);

CKINVDCx5p33_ASAP7_75t_R g2614 ( 
.A(n_2326),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2351),
.B(n_1753),
.Y(n_2615)
);

INVx1_ASAP7_75t_L g2616 ( 
.A(n_2334),
.Y(n_2616)
);

AND2x2_ASAP7_75t_L g2617 ( 
.A(n_2325),
.B(n_1829),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2337),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2410),
.B(n_1308),
.Y(n_2619)
);

AOI22xp5_ASAP7_75t_L g2620 ( 
.A1(n_2463),
.A2(n_1589),
.B1(n_1699),
.B2(n_1310),
.Y(n_2620)
);

INVx2_ASAP7_75t_L g2621 ( 
.A(n_2346),
.Y(n_2621)
);

HB1xp67_ASAP7_75t_L g2622 ( 
.A(n_2391),
.Y(n_2622)
);

NAND2xp5_ASAP7_75t_L g2623 ( 
.A(n_2389),
.B(n_2221),
.Y(n_2623)
);

CKINVDCx5p33_ASAP7_75t_R g2624 ( 
.A(n_2326),
.Y(n_2624)
);

NOR2xp33_ASAP7_75t_L g2625 ( 
.A(n_2343),
.B(n_1308),
.Y(n_2625)
);

AOI22xp33_ASAP7_75t_L g2626 ( 
.A1(n_2431),
.A2(n_2271),
.B1(n_2276),
.B2(n_2270),
.Y(n_2626)
);

NAND2xp5_ASAP7_75t_L g2627 ( 
.A(n_2347),
.B(n_1829),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2380),
.B(n_1829),
.Y(n_2628)
);

NAND2xp5_ASAP7_75t_SL g2629 ( 
.A(n_2391),
.B(n_2095),
.Y(n_2629)
);

NAND2xp5_ASAP7_75t_L g2630 ( 
.A(n_2380),
.B(n_2128),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2330),
.A2(n_2543),
.B1(n_2464),
.B2(n_2454),
.Y(n_2631)
);

NAND2xp5_ASAP7_75t_SL g2632 ( 
.A(n_2416),
.B(n_2095),
.Y(n_2632)
);

INVx5_ASAP7_75t_L g2633 ( 
.A(n_2362),
.Y(n_2633)
);

NOR2xp33_ASAP7_75t_SL g2634 ( 
.A(n_2405),
.B(n_1310),
.Y(n_2634)
);

INVx8_ASAP7_75t_L g2635 ( 
.A(n_2401),
.Y(n_2635)
);

NAND2xp5_ASAP7_75t_SL g2636 ( 
.A(n_2426),
.B(n_2156),
.Y(n_2636)
);

AND2x2_ASAP7_75t_L g2637 ( 
.A(n_2469),
.B(n_2265),
.Y(n_2637)
);

AND2x6_ASAP7_75t_SL g2638 ( 
.A(n_2465),
.B(n_2265),
.Y(n_2638)
);

NAND2xp5_ASAP7_75t_L g2639 ( 
.A(n_2381),
.B(n_2135),
.Y(n_2639)
);

CKINVDCx5p33_ASAP7_75t_R g2640 ( 
.A(n_2538),
.Y(n_2640)
);

AOI22xp33_ASAP7_75t_L g2641 ( 
.A1(n_2381),
.A2(n_2259),
.B1(n_2157),
.B2(n_1989),
.Y(n_2641)
);

NAND2xp5_ASAP7_75t_L g2642 ( 
.A(n_2456),
.B(n_1764),
.Y(n_2642)
);

NAND2xp5_ASAP7_75t_L g2643 ( 
.A(n_2443),
.B(n_1768),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2361),
.Y(n_2644)
);

NAND2xp5_ASAP7_75t_L g2645 ( 
.A(n_2451),
.B(n_1770),
.Y(n_2645)
);

INVx3_ASAP7_75t_L g2646 ( 
.A(n_2362),
.Y(n_2646)
);

NAND2xp33_ASAP7_75t_SL g2647 ( 
.A(n_2378),
.B(n_2275),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2490),
.B(n_2265),
.Y(n_2648)
);

INVx2_ASAP7_75t_SL g2649 ( 
.A(n_2472),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2368),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2352),
.Y(n_2651)
);

AND2x2_ASAP7_75t_L g2652 ( 
.A(n_2520),
.B(n_1779),
.Y(n_2652)
);

INVx2_ASAP7_75t_L g2653 ( 
.A(n_2355),
.Y(n_2653)
);

NAND2xp5_ASAP7_75t_L g2654 ( 
.A(n_2397),
.B(n_1785),
.Y(n_2654)
);

INVx1_ASAP7_75t_SL g2655 ( 
.A(n_2338),
.Y(n_2655)
);

NOR3xp33_ASAP7_75t_L g2656 ( 
.A(n_2392),
.B(n_1480),
.C(n_1984),
.Y(n_2656)
);

NOR2xp33_ASAP7_75t_L g2657 ( 
.A(n_2540),
.B(n_1312),
.Y(n_2657)
);

NAND2xp5_ASAP7_75t_L g2658 ( 
.A(n_2397),
.B(n_2157),
.Y(n_2658)
);

NOR2xp33_ASAP7_75t_L g2659 ( 
.A(n_2390),
.B(n_1312),
.Y(n_2659)
);

AOI22xp33_ASAP7_75t_L g2660 ( 
.A1(n_2555),
.A2(n_1625),
.B1(n_2112),
.B2(n_2090),
.Y(n_2660)
);

INVx1_ASAP7_75t_L g2661 ( 
.A(n_2373),
.Y(n_2661)
);

AND2x6_ASAP7_75t_SL g2662 ( 
.A(n_2486),
.B(n_1718),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_SL g2663 ( 
.A(n_2487),
.B(n_2234),
.Y(n_2663)
);

NAND2xp5_ASAP7_75t_L g2664 ( 
.A(n_2408),
.B(n_2286),
.Y(n_2664)
);

AOI22xp33_ASAP7_75t_SL g2665 ( 
.A1(n_2549),
.A2(n_1321),
.B1(n_1327),
.B2(n_1317),
.Y(n_2665)
);

NAND2xp5_ASAP7_75t_SL g2666 ( 
.A(n_2524),
.B(n_2291),
.Y(n_2666)
);

NAND2xp5_ASAP7_75t_L g2667 ( 
.A(n_2408),
.B(n_2298),
.Y(n_2667)
);

NAND2xp5_ASAP7_75t_SL g2668 ( 
.A(n_2339),
.B(n_2306),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2374),
.Y(n_2669)
);

CKINVDCx5p33_ASAP7_75t_R g2670 ( 
.A(n_2538),
.Y(n_2670)
);

NOR2xp33_ASAP7_75t_L g2671 ( 
.A(n_2474),
.B(n_1317),
.Y(n_2671)
);

INVx2_ASAP7_75t_L g2672 ( 
.A(n_2369),
.Y(n_2672)
);

NAND2xp5_ASAP7_75t_SL g2673 ( 
.A(n_2341),
.B(n_2307),
.Y(n_2673)
);

NAND2xp5_ASAP7_75t_L g2674 ( 
.A(n_2417),
.B(n_2319),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2375),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2417),
.B(n_2323),
.Y(n_2676)
);

NAND2xp5_ASAP7_75t_L g2677 ( 
.A(n_2478),
.B(n_2324),
.Y(n_2677)
);

NOR2xp33_ASAP7_75t_L g2678 ( 
.A(n_2479),
.B(n_1321),
.Y(n_2678)
);

INVx3_ASAP7_75t_L g2679 ( 
.A(n_2362),
.Y(n_2679)
);

INVx2_ASAP7_75t_L g2680 ( 
.A(n_2383),
.Y(n_2680)
);

NOR2xp33_ASAP7_75t_L g2681 ( 
.A(n_2370),
.B(n_1327),
.Y(n_2681)
);

NAND2xp5_ASAP7_75t_SL g2682 ( 
.A(n_2396),
.B(n_1851),
.Y(n_2682)
);

INVx1_ASAP7_75t_L g2683 ( 
.A(n_2377),
.Y(n_2683)
);

NAND2xp5_ASAP7_75t_L g2684 ( 
.A(n_2478),
.B(n_2112),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2382),
.Y(n_2685)
);

INVx2_ASAP7_75t_SL g2686 ( 
.A(n_2545),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2385),
.Y(n_2687)
);

INVx4_ASAP7_75t_L g2688 ( 
.A(n_2344),
.Y(n_2688)
);

HB1xp67_ASAP7_75t_L g2689 ( 
.A(n_2460),
.Y(n_2689)
);

INVx2_ASAP7_75t_L g2690 ( 
.A(n_2418),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2394),
.Y(n_2691)
);

NAND2xp5_ASAP7_75t_SL g2692 ( 
.A(n_2396),
.B(n_2349),
.Y(n_2692)
);

O2A1O1Ixp33_ASAP7_75t_L g2693 ( 
.A1(n_2442),
.A2(n_2364),
.B(n_2366),
.C(n_2356),
.Y(n_2693)
);

AOI21xp5_ASAP7_75t_L g2694 ( 
.A1(n_2500),
.A2(n_2222),
.B(n_2178),
.Y(n_2694)
);

NAND2xp5_ASAP7_75t_L g2695 ( 
.A(n_2485),
.B(n_2120),
.Y(n_2695)
);

NAND2xp5_ASAP7_75t_L g2696 ( 
.A(n_2485),
.B(n_2120),
.Y(n_2696)
);

NAND2xp5_ASAP7_75t_L g2697 ( 
.A(n_2422),
.B(n_2010),
.Y(n_2697)
);

NAND2xp5_ASAP7_75t_SL g2698 ( 
.A(n_2358),
.B(n_1851),
.Y(n_2698)
);

BUFx3_ASAP7_75t_L g2699 ( 
.A(n_2545),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2395),
.Y(n_2700)
);

AOI21xp5_ASAP7_75t_L g2701 ( 
.A1(n_2441),
.A2(n_2228),
.B(n_2029),
.Y(n_2701)
);

BUFx2_ASAP7_75t_L g2702 ( 
.A(n_2401),
.Y(n_2702)
);

INVx2_ASAP7_75t_L g2703 ( 
.A(n_2425),
.Y(n_2703)
);

NAND3xp33_ASAP7_75t_L g2704 ( 
.A(n_2505),
.B(n_1718),
.C(n_1334),
.Y(n_2704)
);

AOI22xp33_ASAP7_75t_L g2705 ( 
.A1(n_2445),
.A2(n_2258),
.B1(n_2262),
.B2(n_2251),
.Y(n_2705)
);

NAND2xp5_ASAP7_75t_SL g2706 ( 
.A(n_2398),
.B(n_2083),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2441),
.B(n_2013),
.Y(n_2707)
);

INVx2_ASAP7_75t_L g2708 ( 
.A(n_2432),
.Y(n_2708)
);

NOR2xp33_ASAP7_75t_SL g2709 ( 
.A(n_2450),
.B(n_1332),
.Y(n_2709)
);

NAND2xp5_ASAP7_75t_L g2710 ( 
.A(n_2470),
.B(n_2251),
.Y(n_2710)
);

NAND2xp5_ASAP7_75t_L g2711 ( 
.A(n_2470),
.B(n_2258),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2399),
.Y(n_2712)
);

CKINVDCx20_ASAP7_75t_R g2713 ( 
.A(n_2354),
.Y(n_2713)
);

NAND2xp5_ASAP7_75t_L g2714 ( 
.A(n_2379),
.B(n_2262),
.Y(n_2714)
);

INVx2_ASAP7_75t_SL g2715 ( 
.A(n_2550),
.Y(n_2715)
);

O2A1O1Ixp33_ASAP7_75t_L g2716 ( 
.A1(n_2554),
.A2(n_2272),
.B(n_2305),
.C(n_2281),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2453),
.B(n_2260),
.Y(n_2717)
);

BUFx8_ASAP7_75t_L g2718 ( 
.A(n_2409),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_SL g2719 ( 
.A(n_2457),
.B(n_2083),
.Y(n_2719)
);

AND2x6_ASAP7_75t_SL g2720 ( 
.A(n_2468),
.B(n_2563),
.Y(n_2720)
);

AOI22xp5_ASAP7_75t_L g2721 ( 
.A1(n_2499),
.A2(n_2429),
.B1(n_2435),
.B2(n_2424),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_SL g2722 ( 
.A(n_2447),
.B(n_2101),
.Y(n_2722)
);

INVx1_ASAP7_75t_L g2723 ( 
.A(n_2402),
.Y(n_2723)
);

NOR2xp33_ASAP7_75t_L g2724 ( 
.A(n_2372),
.B(n_1332),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2448),
.B(n_2272),
.Y(n_2725)
);

NAND2x1p5_ASAP7_75t_L g2726 ( 
.A(n_2412),
.B(n_2158),
.Y(n_2726)
);

NOR2xp33_ASAP7_75t_L g2727 ( 
.A(n_2386),
.B(n_1334),
.Y(n_2727)
);

NOR2xp33_ASAP7_75t_L g2728 ( 
.A(n_2388),
.B(n_1335),
.Y(n_2728)
);

AOI22xp33_ASAP7_75t_L g2729 ( 
.A1(n_2532),
.A2(n_2305),
.B1(n_2281),
.B2(n_2164),
.Y(n_2729)
);

NAND2xp5_ASAP7_75t_SL g2730 ( 
.A(n_2519),
.B(n_2529),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2532),
.A2(n_2164),
.B1(n_2172),
.B2(n_2136),
.Y(n_2731)
);

AOI22xp5_ASAP7_75t_L g2732 ( 
.A1(n_2440),
.A2(n_1336),
.B1(n_1338),
.B2(n_1335),
.Y(n_2732)
);

OAI22xp5_ASAP7_75t_SL g2733 ( 
.A1(n_2437),
.A2(n_1338),
.B1(n_1344),
.B2(n_1336),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_SL g2734 ( 
.A(n_2493),
.B(n_2101),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2404),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2406),
.Y(n_2736)
);

NOR2xp33_ASAP7_75t_L g2737 ( 
.A(n_2413),
.B(n_1344),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2407),
.Y(n_2738)
);

NAND2xp5_ASAP7_75t_L g2739 ( 
.A(n_2492),
.B(n_2136),
.Y(n_2739)
);

AOI221xp5_ASAP7_75t_L g2740 ( 
.A1(n_2561),
.A2(n_665),
.B1(n_667),
.B2(n_652),
.C(n_646),
.Y(n_2740)
);

NAND2xp5_ASAP7_75t_L g2741 ( 
.A(n_2420),
.B(n_2172),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2420),
.B(n_2186),
.Y(n_2742)
);

NOR2xp33_ASAP7_75t_L g2743 ( 
.A(n_2491),
.B(n_1347),
.Y(n_2743)
);

NOR2xp33_ASAP7_75t_L g2744 ( 
.A(n_2423),
.B(n_1347),
.Y(n_2744)
);

OAI22xp5_ASAP7_75t_L g2745 ( 
.A1(n_2494),
.A2(n_2498),
.B1(n_2496),
.B2(n_2517),
.Y(n_2745)
);

NAND2xp5_ASAP7_75t_SL g2746 ( 
.A(n_2569),
.B(n_2101),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_SL g2747 ( 
.A(n_2335),
.B(n_2151),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2421),
.B(n_2427),
.Y(n_2748)
);

OR2x6_ASAP7_75t_L g2749 ( 
.A(n_2437),
.B(n_2309),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2421),
.B(n_2186),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_SL g2751 ( 
.A(n_2403),
.B(n_2151),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2502),
.B(n_2264),
.Y(n_2752)
);

NAND2xp5_ASAP7_75t_L g2753 ( 
.A(n_2427),
.B(n_2142),
.Y(n_2753)
);

NAND2xp5_ASAP7_75t_SL g2754 ( 
.A(n_2551),
.B(n_2151),
.Y(n_2754)
);

INVx1_ASAP7_75t_L g2755 ( 
.A(n_2415),
.Y(n_2755)
);

NOR2xp33_ASAP7_75t_L g2756 ( 
.A(n_2434),
.B(n_1352),
.Y(n_2756)
);

NAND2xp5_ASAP7_75t_L g2757 ( 
.A(n_2434),
.B(n_2142),
.Y(n_2757)
);

NOR2xp33_ASAP7_75t_L g2758 ( 
.A(n_2511),
.B(n_1352),
.Y(n_2758)
);

NAND2xp5_ASAP7_75t_L g2759 ( 
.A(n_2517),
.B(n_2142),
.Y(n_2759)
);

NAND2xp5_ASAP7_75t_L g2760 ( 
.A(n_2527),
.B(n_2142),
.Y(n_2760)
);

OR2x2_ASAP7_75t_L g2761 ( 
.A(n_2508),
.B(n_2244),
.Y(n_2761)
);

NAND2xp5_ASAP7_75t_L g2762 ( 
.A(n_2527),
.B(n_2142),
.Y(n_2762)
);

AOI22xp33_ASAP7_75t_L g2763 ( 
.A1(n_2565),
.A2(n_1625),
.B1(n_1612),
.B2(n_2057),
.Y(n_2763)
);

OAI22xp5_ASAP7_75t_L g2764 ( 
.A1(n_2437),
.A2(n_2029),
.B1(n_2078),
.B2(n_2554),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2528),
.B(n_1894),
.Y(n_2765)
);

AOI22xp33_ASAP7_75t_L g2766 ( 
.A1(n_2556),
.A2(n_2302),
.B1(n_2303),
.B2(n_2296),
.Y(n_2766)
);

OAI21xp5_ASAP7_75t_L g2767 ( 
.A1(n_2693),
.A2(n_2556),
.B(n_2553),
.Y(n_2767)
);

AND2x2_ASAP7_75t_L g2768 ( 
.A(n_2575),
.B(n_2537),
.Y(n_2768)
);

BUFx8_ASAP7_75t_SL g2769 ( 
.A(n_2599),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2583),
.Y(n_2770)
);

NAND2xp5_ASAP7_75t_L g2771 ( 
.A(n_2578),
.B(n_2521),
.Y(n_2771)
);

OAI21x1_ASAP7_75t_L g2772 ( 
.A1(n_2694),
.A2(n_1733),
.B(n_1963),
.Y(n_2772)
);

INVx11_ASAP7_75t_L g2773 ( 
.A(n_2718),
.Y(n_2773)
);

NOR2xp67_ASAP7_75t_L g2774 ( 
.A(n_2587),
.B(n_1518),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2576),
.B(n_2433),
.Y(n_2775)
);

AO21x1_ASAP7_75t_L g2776 ( 
.A1(n_2693),
.A2(n_2568),
.B(n_2514),
.Y(n_2776)
);

NAND2xp5_ASAP7_75t_L g2777 ( 
.A(n_2592),
.B(n_2449),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2597),
.Y(n_2778)
);

O2A1O1Ixp33_ASAP7_75t_L g2779 ( 
.A1(n_2608),
.A2(n_2560),
.B(n_2559),
.C(n_2570),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_SL g2780 ( 
.A(n_2642),
.B(n_2655),
.Y(n_2780)
);

NAND2xp5_ASAP7_75t_L g2781 ( 
.A(n_2603),
.B(n_2462),
.Y(n_2781)
);

NAND2xp5_ASAP7_75t_SL g2782 ( 
.A(n_2636),
.B(n_1355),
.Y(n_2782)
);

AO21x1_ASAP7_75t_L g2783 ( 
.A1(n_2596),
.A2(n_2568),
.B(n_2514),
.Y(n_2783)
);

A2O1A1Ixp33_ASAP7_75t_L g2784 ( 
.A1(n_2631),
.A2(n_2458),
.B(n_2475),
.C(n_2473),
.Y(n_2784)
);

AOI21xp5_ASAP7_75t_L g2785 ( 
.A1(n_2694),
.A2(n_2531),
.B(n_2522),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2601),
.B(n_2476),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2697),
.B(n_2477),
.Y(n_2787)
);

NAND2xp5_ASAP7_75t_L g2788 ( 
.A(n_2756),
.B(n_2489),
.Y(n_2788)
);

AOI21xp5_ASAP7_75t_L g2789 ( 
.A1(n_2571),
.A2(n_2536),
.B(n_2528),
.Y(n_2789)
);

INVx2_ASAP7_75t_SL g2790 ( 
.A(n_2718),
.Y(n_2790)
);

AOI21xp5_ASAP7_75t_L g2791 ( 
.A1(n_2571),
.A2(n_2557),
.B(n_2513),
.Y(n_2791)
);

AOI21xp5_ASAP7_75t_L g2792 ( 
.A1(n_2707),
.A2(n_2557),
.B(n_2513),
.Y(n_2792)
);

NOR2xp33_ASAP7_75t_L g2793 ( 
.A(n_2588),
.B(n_1355),
.Y(n_2793)
);

AOI21xp5_ASAP7_75t_L g2794 ( 
.A1(n_2701),
.A2(n_2268),
.B(n_2151),
.Y(n_2794)
);

AOI21xp5_ASAP7_75t_L g2795 ( 
.A1(n_2701),
.A2(n_2677),
.B(n_2639),
.Y(n_2795)
);

OAI21xp5_ASAP7_75t_L g2796 ( 
.A1(n_2596),
.A2(n_2314),
.B(n_2277),
.Y(n_2796)
);

INVx2_ASAP7_75t_SL g2797 ( 
.A(n_2622),
.Y(n_2797)
);

BUFx6f_ASAP7_75t_L g2798 ( 
.A(n_2604),
.Y(n_2798)
);

INVx2_ASAP7_75t_L g2799 ( 
.A(n_2586),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2616),
.Y(n_2800)
);

NOR3xp33_ASAP7_75t_L g2801 ( 
.A(n_2704),
.B(n_2663),
.C(n_2657),
.Y(n_2801)
);

OAI22xp5_ASAP7_75t_L g2802 ( 
.A1(n_2626),
.A2(n_2177),
.B1(n_1374),
.B2(n_1386),
.Y(n_2802)
);

NAND2xp5_ASAP7_75t_SL g2803 ( 
.A(n_2721),
.B(n_1365),
.Y(n_2803)
);

NAND2xp5_ASAP7_75t_L g2804 ( 
.A(n_2573),
.B(n_2495),
.Y(n_2804)
);

INVx3_ASAP7_75t_L g2805 ( 
.A(n_2688),
.Y(n_2805)
);

NOR2x1_ASAP7_75t_R g2806 ( 
.A(n_2609),
.B(n_2154),
.Y(n_2806)
);

OAI21xp5_ASAP7_75t_L g2807 ( 
.A1(n_2623),
.A2(n_1879),
.B(n_1877),
.Y(n_2807)
);

O2A1O1Ixp33_ASAP7_75t_L g2808 ( 
.A1(n_2692),
.A2(n_1374),
.B(n_1386),
.C(n_1365),
.Y(n_2808)
);

OAI21xp5_ASAP7_75t_L g2809 ( 
.A1(n_2656),
.A2(n_2236),
.B(n_2212),
.Y(n_2809)
);

NAND2x1p5_ASAP7_75t_L g2810 ( 
.A(n_2688),
.B(n_2268),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2584),
.B(n_2506),
.Y(n_2811)
);

BUFx3_ASAP7_75t_L g2812 ( 
.A(n_2622),
.Y(n_2812)
);

AOI21xp5_ASAP7_75t_L g2813 ( 
.A1(n_2630),
.A2(n_2315),
.B(n_2268),
.Y(n_2813)
);

A2O1A1Ixp33_ASAP7_75t_L g2814 ( 
.A1(n_2631),
.A2(n_2507),
.B(n_2518),
.C(n_2510),
.Y(n_2814)
);

NOR2xp33_ASAP7_75t_SL g2815 ( 
.A(n_2634),
.B(n_2267),
.Y(n_2815)
);

AOI21xp5_ASAP7_75t_L g2816 ( 
.A1(n_2593),
.A2(n_2315),
.B(n_2268),
.Y(n_2816)
);

AOI21xp5_ASAP7_75t_L g2817 ( 
.A1(n_2765),
.A2(n_2315),
.B(n_2068),
.Y(n_2817)
);

NAND2xp5_ASAP7_75t_L g2818 ( 
.A(n_2585),
.B(n_2530),
.Y(n_2818)
);

AOI22xp5_ASAP7_75t_L g2819 ( 
.A1(n_2671),
.A2(n_1394),
.B1(n_1404),
.B2(n_1389),
.Y(n_2819)
);

HB1xp67_ASAP7_75t_L g2820 ( 
.A(n_2600),
.Y(n_2820)
);

OAI21xp5_ASAP7_75t_L g2821 ( 
.A1(n_2759),
.A2(n_1819),
.B(n_2247),
.Y(n_2821)
);

AOI21xp5_ASAP7_75t_L g2822 ( 
.A1(n_2754),
.A2(n_2315),
.B(n_2068),
.Y(n_2822)
);

BUFx6f_ASAP7_75t_L g2823 ( 
.A(n_2604),
.Y(n_2823)
);

INVx11_ASAP7_75t_L g2824 ( 
.A(n_2580),
.Y(n_2824)
);

AOI21xp5_ASAP7_75t_L g2825 ( 
.A1(n_2710),
.A2(n_2096),
.B(n_2060),
.Y(n_2825)
);

AOI21xp5_ASAP7_75t_L g2826 ( 
.A1(n_2711),
.A2(n_2096),
.B(n_2060),
.Y(n_2826)
);

NOR2xp67_ASAP7_75t_L g2827 ( 
.A(n_2607),
.B(n_1518),
.Y(n_2827)
);

AOI21xp5_ASAP7_75t_L g2828 ( 
.A1(n_2589),
.A2(n_2119),
.B(n_2078),
.Y(n_2828)
);

NAND2xp5_ASAP7_75t_SL g2829 ( 
.A(n_2681),
.B(n_1389),
.Y(n_2829)
);

AO21x1_ASAP7_75t_L g2830 ( 
.A1(n_2764),
.A2(n_2539),
.B(n_2534),
.Y(n_2830)
);

BUFx3_ASAP7_75t_L g2831 ( 
.A(n_2699),
.Y(n_2831)
);

AOI21xp5_ASAP7_75t_L g2832 ( 
.A1(n_2641),
.A2(n_2119),
.B(n_2134),
.Y(n_2832)
);

AOI21xp5_ASAP7_75t_L g2833 ( 
.A1(n_2641),
.A2(n_2134),
.B(n_1882),
.Y(n_2833)
);

INVx1_ASAP7_75t_L g2834 ( 
.A(n_2618),
.Y(n_2834)
);

AOI21xp5_ASAP7_75t_L g2835 ( 
.A1(n_2748),
.A2(n_1882),
.B(n_1875),
.Y(n_2835)
);

AOI21xp5_ASAP7_75t_L g2836 ( 
.A1(n_2628),
.A2(n_1882),
.B(n_1875),
.Y(n_2836)
);

NAND2xp5_ASAP7_75t_L g2837 ( 
.A(n_2579),
.B(n_2582),
.Y(n_2837)
);

AOI21xp33_ASAP7_75t_L g2838 ( 
.A1(n_2602),
.A2(n_2544),
.B(n_2542),
.Y(n_2838)
);

INVx2_ASAP7_75t_L g2839 ( 
.A(n_2598),
.Y(n_2839)
);

OAI22xp5_ASAP7_75t_L g2840 ( 
.A1(n_2626),
.A2(n_1404),
.B1(n_1406),
.B2(n_1394),
.Y(n_2840)
);

OAI22xp5_ASAP7_75t_L g2841 ( 
.A1(n_2665),
.A2(n_1416),
.B1(n_1422),
.B2(n_1406),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2749),
.Y(n_2842)
);

INVx3_ASAP7_75t_L g2843 ( 
.A(n_2749),
.Y(n_2843)
);

INVx1_ASAP7_75t_L g2844 ( 
.A(n_2644),
.Y(n_2844)
);

AOI21xp5_ASAP7_75t_L g2845 ( 
.A1(n_2684),
.A2(n_1904),
.B(n_1882),
.Y(n_2845)
);

AOI21xp5_ASAP7_75t_L g2846 ( 
.A1(n_2695),
.A2(n_1912),
.B(n_1904),
.Y(n_2846)
);

NAND2xp5_ASAP7_75t_L g2847 ( 
.A(n_2574),
.B(n_1625),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2650),
.Y(n_2848)
);

NAND2xp5_ASAP7_75t_L g2849 ( 
.A(n_2605),
.B(n_1625),
.Y(n_2849)
);

O2A1O1Ixp33_ASAP7_75t_L g2850 ( 
.A1(n_2666),
.A2(n_1422),
.B(n_1427),
.C(n_1416),
.Y(n_2850)
);

BUFx6f_ASAP7_75t_L g2851 ( 
.A(n_2604),
.Y(n_2851)
);

INVx1_ASAP7_75t_L g2852 ( 
.A(n_2661),
.Y(n_2852)
);

OAI22xp5_ASAP7_75t_L g2853 ( 
.A1(n_2665),
.A2(n_2288),
.B1(n_2558),
.B2(n_2546),
.Y(n_2853)
);

AOI21xp5_ASAP7_75t_L g2854 ( 
.A1(n_2696),
.A2(n_1912),
.B(n_1904),
.Y(n_2854)
);

OAI21xp33_ASAP7_75t_L g2855 ( 
.A1(n_2590),
.A2(n_674),
.B(n_672),
.Y(n_2855)
);

AOI22xp5_ASAP7_75t_L g2856 ( 
.A1(n_2678),
.A2(n_1625),
.B1(n_1665),
.B2(n_1612),
.Y(n_2856)
);

AND2x2_ASAP7_75t_L g2857 ( 
.A(n_2613),
.B(n_2318),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2669),
.Y(n_2858)
);

NAND2xp5_ASAP7_75t_L g2859 ( 
.A(n_2717),
.B(n_2438),
.Y(n_2859)
);

AOI21xp5_ASAP7_75t_L g2860 ( 
.A1(n_2668),
.A2(n_1912),
.B(n_1904),
.Y(n_2860)
);

INVx3_ASAP7_75t_L g2861 ( 
.A(n_2749),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2675),
.Y(n_2862)
);

NOR3xp33_ASAP7_75t_L g2863 ( 
.A(n_2591),
.B(n_676),
.C(n_675),
.Y(n_2863)
);

NOR2xp33_ASAP7_75t_L g2864 ( 
.A(n_2625),
.B(n_2512),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2683),
.Y(n_2865)
);

AOI21xp5_ASAP7_75t_L g2866 ( 
.A1(n_2673),
.A2(n_1939),
.B(n_1912),
.Y(n_2866)
);

NAND2xp5_ASAP7_75t_SL g2867 ( 
.A(n_2724),
.B(n_2344),
.Y(n_2867)
);

AOI21xp33_ASAP7_75t_L g2868 ( 
.A1(n_2611),
.A2(n_1934),
.B(n_2562),
.Y(n_2868)
);

INVx1_ASAP7_75t_L g2869 ( 
.A(n_2685),
.Y(n_2869)
);

NOR2xp33_ASAP7_75t_L g2870 ( 
.A(n_2619),
.B(n_2512),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2615),
.B(n_2439),
.Y(n_2871)
);

INVx3_ASAP7_75t_L g2872 ( 
.A(n_2607),
.Y(n_2872)
);

O2A1O1Ixp33_ASAP7_75t_L g2873 ( 
.A1(n_2632),
.A2(n_1547),
.B(n_1987),
.C(n_1983),
.Y(n_2873)
);

AOI21xp5_ASAP7_75t_L g2874 ( 
.A1(n_2741),
.A2(n_1962),
.B(n_1939),
.Y(n_2874)
);

AOI21xp5_ASAP7_75t_L g2875 ( 
.A1(n_2742),
.A2(n_1962),
.B(n_1939),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2581),
.B(n_2446),
.Y(n_2876)
);

NAND2xp5_ASAP7_75t_L g2877 ( 
.A(n_2643),
.B(n_2455),
.Y(n_2877)
);

AOI21xp5_ASAP7_75t_L g2878 ( 
.A1(n_2750),
.A2(n_1962),
.B(n_1939),
.Y(n_2878)
);

AOI21xp5_ASAP7_75t_L g2879 ( 
.A1(n_2658),
.A2(n_1966),
.B(n_1962),
.Y(n_2879)
);

AOI21xp33_ASAP7_75t_L g2880 ( 
.A1(n_2745),
.A2(n_1934),
.B(n_2564),
.Y(n_2880)
);

NAND2xp5_ASAP7_75t_L g2881 ( 
.A(n_2645),
.B(n_2467),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2652),
.B(n_2480),
.Y(n_2882)
);

OAI22xp5_ASAP7_75t_L g2883 ( 
.A1(n_2620),
.A2(n_2567),
.B1(n_2566),
.B2(n_2158),
.Y(n_2883)
);

OAI21x1_ASAP7_75t_L g2884 ( 
.A1(n_2716),
.A2(n_1970),
.B(n_1963),
.Y(n_2884)
);

BUFx6f_ASAP7_75t_L g2885 ( 
.A(n_2610),
.Y(n_2885)
);

NAND2xp5_ASAP7_75t_L g2886 ( 
.A(n_2654),
.B(n_2484),
.Y(n_2886)
);

BUFx3_ASAP7_75t_L g2887 ( 
.A(n_2600),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2617),
.B(n_2488),
.Y(n_2888)
);

AOI21xp5_ASAP7_75t_L g2889 ( 
.A1(n_2664),
.A2(n_1967),
.B(n_1966),
.Y(n_2889)
);

INVx2_ASAP7_75t_L g2890 ( 
.A(n_2621),
.Y(n_2890)
);

O2A1O1Ixp5_ASAP7_75t_L g2891 ( 
.A1(n_2682),
.A2(n_2504),
.B(n_2515),
.C(n_2501),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_SL g2892 ( 
.A(n_2727),
.B(n_2344),
.Y(n_2892)
);

O2A1O1Ixp33_ASAP7_75t_SL g2893 ( 
.A1(n_2747),
.A2(n_1995),
.B(n_2004),
.C(n_1992),
.Y(n_2893)
);

AOI21xp5_ASAP7_75t_L g2894 ( 
.A1(n_2667),
.A2(n_2676),
.B(n_2674),
.Y(n_2894)
);

NAND2xp5_ASAP7_75t_L g2895 ( 
.A(n_2758),
.B(n_2535),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2728),
.B(n_2541),
.Y(n_2896)
);

OAI21xp5_ASAP7_75t_L g2897 ( 
.A1(n_2656),
.A2(n_2012),
.B(n_2007),
.Y(n_2897)
);

NOR2xp33_ASAP7_75t_L g2898 ( 
.A(n_2659),
.B(n_2743),
.Y(n_2898)
);

AOI21xp5_ASAP7_75t_L g2899 ( 
.A1(n_2714),
.A2(n_1967),
.B(n_1966),
.Y(n_2899)
);

AOI21x1_ASAP7_75t_L g2900 ( 
.A1(n_2760),
.A2(n_1970),
.B(n_1927),
.Y(n_2900)
);

A2O1A1Ixp33_ASAP7_75t_L g2901 ( 
.A1(n_2737),
.A2(n_2015),
.B(n_2017),
.C(n_2016),
.Y(n_2901)
);

AOI21xp5_ASAP7_75t_L g2902 ( 
.A1(n_2725),
.A2(n_1967),
.B(n_1966),
.Y(n_2902)
);

INVx1_ASAP7_75t_SL g2903 ( 
.A(n_2689),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2627),
.B(n_2552),
.Y(n_2904)
);

INVx3_ASAP7_75t_L g2905 ( 
.A(n_2606),
.Y(n_2905)
);

NOR2xp33_ASAP7_75t_L g2906 ( 
.A(n_2744),
.B(n_2516),
.Y(n_2906)
);

AOI22xp5_ASAP7_75t_L g2907 ( 
.A1(n_2709),
.A2(n_2267),
.B1(n_2019),
.B2(n_2020),
.Y(n_2907)
);

AOI21xp5_ASAP7_75t_L g2908 ( 
.A1(n_2753),
.A2(n_1978),
.B(n_1967),
.Y(n_2908)
);

INVx1_ASAP7_75t_L g2909 ( 
.A(n_2687),
.Y(n_2909)
);

NOR3xp33_ASAP7_75t_L g2910 ( 
.A(n_2740),
.B(n_681),
.C(n_679),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2691),
.Y(n_2911)
);

AND2x2_ASAP7_75t_SL g2912 ( 
.A(n_2660),
.B(n_2376),
.Y(n_2912)
);

OAI22xp5_ASAP7_75t_L g2913 ( 
.A1(n_2572),
.A2(n_2170),
.B1(n_2204),
.B2(n_2171),
.Y(n_2913)
);

AOI21xp5_ASAP7_75t_L g2914 ( 
.A1(n_2757),
.A2(n_1985),
.B(n_1978),
.Y(n_2914)
);

AND2x2_ASAP7_75t_L g2915 ( 
.A(n_2637),
.B(n_714),
.Y(n_2915)
);

OAI21xp5_ASAP7_75t_L g2916 ( 
.A1(n_2595),
.A2(n_1866),
.B(n_1860),
.Y(n_2916)
);

OAI22xp5_ASAP7_75t_L g2917 ( 
.A1(n_2572),
.A2(n_2170),
.B1(n_2204),
.B2(n_2171),
.Y(n_2917)
);

AOI21xp5_ASAP7_75t_L g2918 ( 
.A1(n_2762),
.A2(n_1985),
.B(n_1978),
.Y(n_2918)
);

HB1xp67_ASAP7_75t_L g2919 ( 
.A(n_2689),
.Y(n_2919)
);

OAI21xp5_ASAP7_75t_L g2920 ( 
.A1(n_2716),
.A2(n_1866),
.B(n_2274),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2649),
.B(n_2739),
.Y(n_2921)
);

INVx1_ASAP7_75t_SL g2922 ( 
.A(n_2648),
.Y(n_2922)
);

NOR2xp67_ASAP7_75t_L g2923 ( 
.A(n_2715),
.B(n_2516),
.Y(n_2923)
);

NOR2xp33_ASAP7_75t_L g2924 ( 
.A(n_2732),
.B(n_2523),
.Y(n_2924)
);

AOI21xp5_ASAP7_75t_L g2925 ( 
.A1(n_2647),
.A2(n_1985),
.B(n_1978),
.Y(n_2925)
);

O2A1O1Ixp33_ASAP7_75t_L g2926 ( 
.A1(n_2730),
.A2(n_1547),
.B(n_1605),
.C(n_1997),
.Y(n_2926)
);

NAND2xp5_ASAP7_75t_L g2927 ( 
.A(n_2752),
.B(n_2720),
.Y(n_2927)
);

NAND2xp5_ASAP7_75t_L g2928 ( 
.A(n_2700),
.B(n_2274),
.Y(n_2928)
);

OAI22xp5_ASAP7_75t_L g2929 ( 
.A1(n_2733),
.A2(n_2239),
.B1(n_2297),
.B2(n_2275),
.Y(n_2929)
);

NAND2xp5_ASAP7_75t_L g2930 ( 
.A(n_2712),
.B(n_2287),
.Y(n_2930)
);

OAI21xp5_ASAP7_75t_L g2931 ( 
.A1(n_2740),
.A2(n_2300),
.B(n_2287),
.Y(n_2931)
);

AO21x1_ASAP7_75t_L g2932 ( 
.A1(n_2722),
.A2(n_1605),
.B(n_2239),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2723),
.Y(n_2933)
);

O2A1O1Ixp33_ASAP7_75t_L g2934 ( 
.A1(n_2746),
.A2(n_2629),
.B(n_2698),
.C(n_2734),
.Y(n_2934)
);

BUFx6f_ASAP7_75t_L g2935 ( 
.A(n_2610),
.Y(n_2935)
);

OAI21xp5_ASAP7_75t_L g2936 ( 
.A1(n_2729),
.A2(n_2300),
.B(n_1934),
.Y(n_2936)
);

NAND2xp5_ASAP7_75t_L g2937 ( 
.A(n_2735),
.B(n_2072),
.Y(n_2937)
);

AOI21xp5_ASAP7_75t_L g2938 ( 
.A1(n_2726),
.A2(n_1990),
.B(n_1985),
.Y(n_2938)
);

INVx2_ASAP7_75t_L g2939 ( 
.A(n_2651),
.Y(n_2939)
);

NOR2xp67_ASAP7_75t_L g2940 ( 
.A(n_2761),
.B(n_2523),
.Y(n_2940)
);

AOI21xp5_ASAP7_75t_L g2941 ( 
.A1(n_2726),
.A2(n_2011),
.B(n_1990),
.Y(n_2941)
);

OAI21xp5_ASAP7_75t_L g2942 ( 
.A1(n_2729),
.A2(n_1994),
.B(n_2240),
.Y(n_2942)
);

AOI21x1_ASAP7_75t_L g2943 ( 
.A1(n_2706),
.A2(n_1927),
.B(n_1974),
.Y(n_2943)
);

OAI21xp5_ASAP7_75t_L g2944 ( 
.A1(n_2731),
.A2(n_2705),
.B(n_2766),
.Y(n_2944)
);

OAI21xp33_ASAP7_75t_L g2945 ( 
.A1(n_2731),
.A2(n_688),
.B(n_683),
.Y(n_2945)
);

OAI21xp5_ASAP7_75t_L g2946 ( 
.A1(n_2705),
.A2(n_2077),
.B(n_2075),
.Y(n_2946)
);

NOR2xp33_ASAP7_75t_L g2947 ( 
.A(n_2713),
.B(n_2525),
.Y(n_2947)
);

BUFx6f_ASAP7_75t_L g2948 ( 
.A(n_2610),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_2702),
.Y(n_2949)
);

NAND2x1p5_ASAP7_75t_L g2950 ( 
.A(n_2633),
.B(n_2297),
.Y(n_2950)
);

INVx3_ASAP7_75t_L g2951 ( 
.A(n_2606),
.Y(n_2951)
);

O2A1O1Ixp33_ASAP7_75t_L g2952 ( 
.A1(n_2751),
.A2(n_1997),
.B(n_2123),
.C(n_2118),
.Y(n_2952)
);

NOR2x1p5_ASAP7_75t_SL g2953 ( 
.A(n_2653),
.B(n_2482),
.Y(n_2953)
);

AOI21xp5_ASAP7_75t_L g2954 ( 
.A1(n_2763),
.A2(n_2011),
.B(n_1990),
.Y(n_2954)
);

AOI21xp5_ASAP7_75t_L g2955 ( 
.A1(n_2766),
.A2(n_2011),
.B(n_1990),
.Y(n_2955)
);

O2A1O1Ixp33_ASAP7_75t_L g2956 ( 
.A1(n_2736),
.A2(n_2126),
.B(n_2129),
.C(n_2125),
.Y(n_2956)
);

OR2x2_ASAP7_75t_L g2957 ( 
.A(n_2738),
.B(n_2525),
.Y(n_2957)
);

AOI21xp5_ASAP7_75t_L g2958 ( 
.A1(n_2635),
.A2(n_2011),
.B(n_2309),
.Y(n_2958)
);

BUFx2_ASAP7_75t_L g2959 ( 
.A(n_2812),
.Y(n_2959)
);

OR2x6_ASAP7_75t_L g2960 ( 
.A(n_2944),
.B(n_2635),
.Y(n_2960)
);

INVx2_ASAP7_75t_L g2961 ( 
.A(n_2799),
.Y(n_2961)
);

OR2x2_ASAP7_75t_L g2962 ( 
.A(n_2922),
.B(n_2903),
.Y(n_2962)
);

BUFx2_ASAP7_75t_L g2963 ( 
.A(n_2887),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2837),
.B(n_2755),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_SL g2965 ( 
.A(n_2801),
.B(n_2614),
.Y(n_2965)
);

INVx2_ASAP7_75t_SL g2966 ( 
.A(n_2824),
.Y(n_2966)
);

BUFx4f_ASAP7_75t_L g2967 ( 
.A(n_2798),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2894),
.B(n_2672),
.Y(n_2968)
);

INVx2_ASAP7_75t_L g2969 ( 
.A(n_2839),
.Y(n_2969)
);

INVx1_ASAP7_75t_L g2970 ( 
.A(n_2770),
.Y(n_2970)
);

NOR2xp33_ASAP7_75t_R g2971 ( 
.A(n_2905),
.B(n_2624),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2795),
.B(n_2811),
.Y(n_2972)
);

BUFx3_ASAP7_75t_L g2973 ( 
.A(n_2831),
.Y(n_2973)
);

INVx2_ASAP7_75t_L g2974 ( 
.A(n_2890),
.Y(n_2974)
);

AND2x4_ASAP7_75t_L g2975 ( 
.A(n_2842),
.B(n_2594),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2778),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2805),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2800),
.Y(n_2978)
);

INVx2_ASAP7_75t_L g2979 ( 
.A(n_2939),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2780),
.B(n_2680),
.Y(n_2980)
);

OR2x6_ASAP7_75t_L g2981 ( 
.A(n_2785),
.B(n_2635),
.Y(n_2981)
);

INVx2_ASAP7_75t_L g2982 ( 
.A(n_2957),
.Y(n_2982)
);

NAND2xp5_ASAP7_75t_L g2983 ( 
.A(n_2777),
.B(n_2690),
.Y(n_2983)
);

INVx1_ASAP7_75t_L g2984 ( 
.A(n_2834),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2844),
.Y(n_2985)
);

AND2x4_ASAP7_75t_L g2986 ( 
.A(n_2842),
.B(n_2594),
.Y(n_2986)
);

BUFx6f_ASAP7_75t_L g2987 ( 
.A(n_2885),
.Y(n_2987)
);

BUFx6f_ASAP7_75t_L g2988 ( 
.A(n_2885),
.Y(n_2988)
);

NAND2xp5_ASAP7_75t_L g2989 ( 
.A(n_2788),
.B(n_2703),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2848),
.Y(n_2990)
);

AND2x2_ASAP7_75t_L g2991 ( 
.A(n_2768),
.B(n_2594),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2852),
.Y(n_2992)
);

AOI22xp33_ASAP7_75t_L g2993 ( 
.A1(n_2910),
.A2(n_2863),
.B1(n_2803),
.B2(n_2898),
.Y(n_2993)
);

NAND2xp5_ASAP7_75t_L g2994 ( 
.A(n_2787),
.B(n_2708),
.Y(n_2994)
);

INVx1_ASAP7_75t_L g2995 ( 
.A(n_2858),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2922),
.B(n_2775),
.Y(n_2996)
);

BUFx6f_ASAP7_75t_L g2997 ( 
.A(n_2885),
.Y(n_2997)
);

NAND2xp5_ASAP7_75t_SL g2998 ( 
.A(n_2940),
.B(n_2640),
.Y(n_2998)
);

CKINVDCx20_ASAP7_75t_R g2999 ( 
.A(n_2769),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_L g3000 ( 
.A(n_2921),
.B(n_2638),
.Y(n_3000)
);

NAND2xp5_ASAP7_75t_L g3001 ( 
.A(n_2804),
.B(n_2577),
.Y(n_3001)
);

INVx3_ASAP7_75t_L g3002 ( 
.A(n_2805),
.Y(n_3002)
);

NAND2xp5_ASAP7_75t_SL g3003 ( 
.A(n_2927),
.B(n_2670),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2781),
.B(n_2577),
.Y(n_3004)
);

A2O1A1Ixp33_ASAP7_75t_L g3005 ( 
.A1(n_2945),
.A2(n_2719),
.B(n_2686),
.C(n_2646),
.Y(n_3005)
);

BUFx6f_ASAP7_75t_L g3006 ( 
.A(n_2935),
.Y(n_3006)
);

INVx2_ASAP7_75t_SL g3007 ( 
.A(n_2773),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2862),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2786),
.B(n_2612),
.Y(n_3009)
);

BUFx6f_ASAP7_75t_L g3010 ( 
.A(n_2935),
.Y(n_3010)
);

INVx1_ASAP7_75t_SL g3011 ( 
.A(n_2903),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2896),
.B(n_2612),
.Y(n_3012)
);

BUFx2_ASAP7_75t_L g3013 ( 
.A(n_2949),
.Y(n_3013)
);

NAND2xp5_ASAP7_75t_SL g3014 ( 
.A(n_2934),
.B(n_2633),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2818),
.B(n_2646),
.Y(n_3015)
);

CKINVDCx20_ASAP7_75t_R g3016 ( 
.A(n_2771),
.Y(n_3016)
);

BUFx2_ASAP7_75t_L g3017 ( 
.A(n_2820),
.Y(n_3017)
);

BUFx3_ASAP7_75t_L g3018 ( 
.A(n_2798),
.Y(n_3018)
);

INVx3_ASAP7_75t_L g3019 ( 
.A(n_2905),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2870),
.B(n_2679),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2865),
.Y(n_3021)
);

INVx1_ASAP7_75t_L g3022 ( 
.A(n_2869),
.Y(n_3022)
);

BUFx6f_ASAP7_75t_L g3023 ( 
.A(n_2935),
.Y(n_3023)
);

NAND2xp5_ASAP7_75t_L g3024 ( 
.A(n_2792),
.B(n_2679),
.Y(n_3024)
);

BUFx12f_ASAP7_75t_L g3025 ( 
.A(n_2798),
.Y(n_3025)
);

AOI22xp33_ASAP7_75t_L g3026 ( 
.A1(n_2841),
.A2(n_714),
.B1(n_2580),
.B2(n_2089),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2909),
.Y(n_3027)
);

INVx3_ASAP7_75t_L g3028 ( 
.A(n_2951),
.Y(n_3028)
);

BUFx8_ASAP7_75t_L g3029 ( 
.A(n_2790),
.Y(n_3029)
);

NAND2xp5_ASAP7_75t_SL g3030 ( 
.A(n_2808),
.B(n_2633),
.Y(n_3030)
);

INVx1_ASAP7_75t_L g3031 ( 
.A(n_2911),
.Y(n_3031)
);

INVxp67_ASAP7_75t_SL g3032 ( 
.A(n_2919),
.Y(n_3032)
);

NAND2xp5_ASAP7_75t_L g3033 ( 
.A(n_2886),
.B(n_2633),
.Y(n_3033)
);

OR2x2_ASAP7_75t_L g3034 ( 
.A(n_2797),
.B(n_1994),
.Y(n_3034)
);

INVx3_ASAP7_75t_L g3035 ( 
.A(n_2951),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2933),
.Y(n_3036)
);

INVx2_ASAP7_75t_L g3037 ( 
.A(n_2857),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2928),
.Y(n_3038)
);

INVx3_ASAP7_75t_L g3039 ( 
.A(n_2823),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_SL g3040 ( 
.A(n_2856),
.B(n_2482),
.Y(n_3040)
);

BUFx4f_ASAP7_75t_L g3041 ( 
.A(n_2823),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2930),
.Y(n_3042)
);

HB1xp67_ASAP7_75t_L g3043 ( 
.A(n_2859),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2937),
.Y(n_3044)
);

BUFx4f_ASAP7_75t_L g3045 ( 
.A(n_2823),
.Y(n_3045)
);

AO221x1_ASAP7_75t_L g3046 ( 
.A1(n_2843),
.A2(n_2400),
.B1(n_2509),
.B2(n_2459),
.C(n_2376),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2876),
.Y(n_3047)
);

BUFx6f_ASAP7_75t_L g3048 ( 
.A(n_2948),
.Y(n_3048)
);

AND3x1_ASAP7_75t_SL g3049 ( 
.A(n_2850),
.B(n_2662),
.C(n_699),
.Y(n_3049)
);

AOI21xp5_ASAP7_75t_L g3050 ( 
.A1(n_2791),
.A2(n_2309),
.B(n_2275),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2882),
.Y(n_3051)
);

NAND2xp5_ASAP7_75t_L g3052 ( 
.A(n_2895),
.B(n_694),
.Y(n_3052)
);

AOI22xp33_ASAP7_75t_L g3053 ( 
.A1(n_2840),
.A2(n_714),
.B1(n_2089),
.B2(n_2057),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_SL g3054 ( 
.A(n_2815),
.B(n_2482),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2871),
.Y(n_3055)
);

INVx2_ASAP7_75t_L g3056 ( 
.A(n_2888),
.Y(n_3056)
);

AND2x6_ASAP7_75t_L g3057 ( 
.A(n_2843),
.B(n_2376),
.Y(n_3057)
);

BUFx12f_ASAP7_75t_SL g3058 ( 
.A(n_2851),
.Y(n_3058)
);

INVx1_ASAP7_75t_SL g3059 ( 
.A(n_2906),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2948),
.Y(n_3060)
);

NAND2xp5_ASAP7_75t_L g3061 ( 
.A(n_2864),
.B(n_708),
.Y(n_3061)
);

NAND2xp5_ASAP7_75t_SL g3062 ( 
.A(n_2815),
.B(n_2482),
.Y(n_3062)
);

INVx1_ASAP7_75t_SL g3063 ( 
.A(n_2912),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2830),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2924),
.B(n_758),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2776),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2877),
.B(n_713),
.Y(n_3067)
);

NOR2xp33_ASAP7_75t_L g3068 ( 
.A(n_2793),
.B(n_758),
.Y(n_3068)
);

NAND2xp5_ASAP7_75t_SL g3069 ( 
.A(n_2838),
.B(n_2802),
.Y(n_3069)
);

NOR2xp33_ASAP7_75t_L g3070 ( 
.A(n_2819),
.B(n_2829),
.Y(n_3070)
);

AND2x4_ASAP7_75t_L g3071 ( 
.A(n_2861),
.B(n_2400),
.Y(n_3071)
);

BUFx6f_ASAP7_75t_L g3072 ( 
.A(n_2948),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2851),
.Y(n_3073)
);

NOR2xp33_ASAP7_75t_L g3074 ( 
.A(n_2782),
.B(n_760),
.Y(n_3074)
);

NAND2xp5_ASAP7_75t_SL g3075 ( 
.A(n_2853),
.B(n_2482),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2915),
.B(n_760),
.Y(n_3076)
);

BUFx6f_ASAP7_75t_L g3077 ( 
.A(n_2851),
.Y(n_3077)
);

AND2x4_ASAP7_75t_L g3078 ( 
.A(n_2861),
.B(n_2400),
.Y(n_3078)
);

OAI22xp5_ASAP7_75t_L g3079 ( 
.A1(n_2814),
.A2(n_722),
.B1(n_726),
.B2(n_717),
.Y(n_3079)
);

INVx2_ASAP7_75t_L g3080 ( 
.A(n_2904),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2881),
.B(n_734),
.Y(n_3081)
);

AOI21xp5_ASAP7_75t_L g3082 ( 
.A1(n_2832),
.A2(n_2275),
.B(n_1743),
.Y(n_3082)
);

NAND2xp5_ASAP7_75t_SL g3083 ( 
.A(n_2779),
.B(n_2503),
.Y(n_3083)
);

BUFx6f_ASAP7_75t_L g3084 ( 
.A(n_2872),
.Y(n_3084)
);

NAND2xp5_ASAP7_75t_L g3085 ( 
.A(n_2867),
.B(n_735),
.Y(n_3085)
);

INVx2_ASAP7_75t_L g3086 ( 
.A(n_2891),
.Y(n_3086)
);

AOI22xp33_ASAP7_75t_L g3087 ( 
.A1(n_2855),
.A2(n_2089),
.B1(n_2113),
.B2(n_2057),
.Y(n_3087)
);

BUFx2_ASAP7_75t_L g3088 ( 
.A(n_2872),
.Y(n_3088)
);

BUFx6f_ASAP7_75t_L g3089 ( 
.A(n_2950),
.Y(n_3089)
);

INVx1_ASAP7_75t_L g3090 ( 
.A(n_2783),
.Y(n_3090)
);

NOR2x1p5_ASAP7_75t_L g3091 ( 
.A(n_2847),
.B(n_2548),
.Y(n_3091)
);

AND3x2_ASAP7_75t_SL g3092 ( 
.A(n_2806),
.B(n_1019),
.C(n_998),
.Y(n_3092)
);

AOI22xp5_ASAP7_75t_L g3093 ( 
.A1(n_2892),
.A2(n_736),
.B1(n_2113),
.B2(n_2089),
.Y(n_3093)
);

BUFx3_ASAP7_75t_L g3094 ( 
.A(n_2947),
.Y(n_3094)
);

BUFx2_ASAP7_75t_L g3095 ( 
.A(n_2950),
.Y(n_3095)
);

OAI22xp5_ASAP7_75t_L g3096 ( 
.A1(n_2784),
.A2(n_2243),
.B1(n_2249),
.B2(n_2240),
.Y(n_3096)
);

INVx1_ASAP7_75t_L g3097 ( 
.A(n_2767),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2953),
.Y(n_3098)
);

AND2x2_ASAP7_75t_L g3099 ( 
.A(n_2897),
.B(n_2459),
.Y(n_3099)
);

INVx1_ASAP7_75t_L g3100 ( 
.A(n_2956),
.Y(n_3100)
);

INVx3_ASAP7_75t_L g3101 ( 
.A(n_2810),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2920),
.Y(n_3102)
);

AND2x4_ASAP7_75t_L g3103 ( 
.A(n_2923),
.B(n_2459),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2936),
.Y(n_3104)
);

NAND2xp5_ASAP7_75t_L g3105 ( 
.A(n_2809),
.B(n_2243),
.Y(n_3105)
);

NAND2xp5_ASAP7_75t_SL g3106 ( 
.A(n_2907),
.B(n_2503),
.Y(n_3106)
);

INVx2_ASAP7_75t_L g3107 ( 
.A(n_2943),
.Y(n_3107)
);

BUFx4f_ASAP7_75t_L g3108 ( 
.A(n_2810),
.Y(n_3108)
);

INVx2_ASAP7_75t_SL g3109 ( 
.A(n_2929),
.Y(n_3109)
);

INVx3_ASAP7_75t_L g3110 ( 
.A(n_2900),
.Y(n_3110)
);

INVxp67_ASAP7_75t_L g3111 ( 
.A(n_2774),
.Y(n_3111)
);

INVx2_ASAP7_75t_L g3112 ( 
.A(n_2884),
.Y(n_3112)
);

AND2x2_ASAP7_75t_L g3113 ( 
.A(n_2883),
.B(n_2509),
.Y(n_3113)
);

INVx1_ASAP7_75t_L g3114 ( 
.A(n_2936),
.Y(n_3114)
);

AND2x6_ASAP7_75t_L g3115 ( 
.A(n_2849),
.B(n_2509),
.Y(n_3115)
);

BUFx6f_ASAP7_75t_L g3116 ( 
.A(n_2772),
.Y(n_3116)
);

INVx3_ASAP7_75t_SL g3117 ( 
.A(n_2827),
.Y(n_3117)
);

AND2x2_ASAP7_75t_L g3118 ( 
.A(n_2807),
.B(n_2931),
.Y(n_3118)
);

BUFx3_ASAP7_75t_L g3119 ( 
.A(n_2913),
.Y(n_3119)
);

INVx2_ASAP7_75t_L g3120 ( 
.A(n_2946),
.Y(n_3120)
);

INVx2_ASAP7_75t_L g3121 ( 
.A(n_2916),
.Y(n_3121)
);

NAND2xp5_ASAP7_75t_L g3122 ( 
.A(n_2789),
.B(n_2249),
.Y(n_3122)
);

INVx5_ASAP7_75t_L g3123 ( 
.A(n_2932),
.Y(n_3123)
);

NAND2xp5_ASAP7_75t_L g3124 ( 
.A(n_2828),
.B(n_2130),
.Y(n_3124)
);

BUFx6f_ASAP7_75t_L g3125 ( 
.A(n_2958),
.Y(n_3125)
);

CKINVDCx11_ASAP7_75t_R g3126 ( 
.A(n_2917),
.Y(n_3126)
);

NOR2xp33_ASAP7_75t_L g3127 ( 
.A(n_2901),
.B(n_2526),
.Y(n_3127)
);

AND2x2_ASAP7_75t_L g3128 ( 
.A(n_2821),
.B(n_2526),
.Y(n_3128)
);

AOI22xp5_ASAP7_75t_L g3129 ( 
.A1(n_2821),
.A2(n_2089),
.B1(n_2117),
.B2(n_2113),
.Y(n_3129)
);

A2O1A1Ixp33_ASAP7_75t_L g3130 ( 
.A1(n_2833),
.A2(n_2926),
.B(n_2816),
.C(n_2817),
.Y(n_3130)
);

AOI22xp33_ASAP7_75t_L g3131 ( 
.A1(n_2796),
.A2(n_2113),
.B1(n_2117),
.B2(n_1742),
.Y(n_3131)
);

CKINVDCx5p33_ASAP7_75t_R g3132 ( 
.A(n_2813),
.Y(n_3132)
);

INVx1_ASAP7_75t_L g3133 ( 
.A(n_2942),
.Y(n_3133)
);

INVx2_ASAP7_75t_SL g3134 ( 
.A(n_2893),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2942),
.Y(n_3135)
);

NAND2xp5_ASAP7_75t_L g3136 ( 
.A(n_2825),
.B(n_2139),
.Y(n_3136)
);

CKINVDCx5p33_ASAP7_75t_R g3137 ( 
.A(n_2938),
.Y(n_3137)
);

NAND2xp5_ASAP7_75t_L g3138 ( 
.A(n_2826),
.B(n_2143),
.Y(n_3138)
);

INVx3_ASAP7_75t_SL g3139 ( 
.A(n_2908),
.Y(n_3139)
);

CKINVDCx5p33_ASAP7_75t_R g3140 ( 
.A(n_2941),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2918),
.B(n_2193),
.Y(n_3141)
);

AO22x1_ASAP7_75t_L g3142 ( 
.A1(n_2873),
.A2(n_2113),
.B1(n_2117),
.B2(n_1742),
.Y(n_3142)
);

CKINVDCx14_ASAP7_75t_R g3143 ( 
.A(n_2925),
.Y(n_3143)
);

NAND2xp5_ASAP7_75t_L g3144 ( 
.A(n_2879),
.B(n_2202),
.Y(n_3144)
);

BUFx3_ASAP7_75t_L g3145 ( 
.A(n_2952),
.Y(n_3145)
);

HB1xp67_ASAP7_75t_L g3146 ( 
.A(n_2955),
.Y(n_3146)
);

NOR2xp33_ASAP7_75t_L g3147 ( 
.A(n_2914),
.B(n_2526),
.Y(n_3147)
);

NAND2xp5_ASAP7_75t_L g3148 ( 
.A(n_2836),
.B(n_2216),
.Y(n_3148)
);

NAND2xp5_ASAP7_75t_L g3149 ( 
.A(n_2845),
.B(n_2218),
.Y(n_3149)
);

INVx2_ASAP7_75t_L g3150 ( 
.A(n_2860),
.Y(n_3150)
);

AND2x4_ASAP7_75t_L g3151 ( 
.A(n_2866),
.B(n_2548),
.Y(n_3151)
);

NAND2xp5_ASAP7_75t_L g3152 ( 
.A(n_2846),
.B(n_2227),
.Y(n_3152)
);

INVx4_ASAP7_75t_L g3153 ( 
.A(n_2822),
.Y(n_3153)
);

BUFx6f_ASAP7_75t_L g3154 ( 
.A(n_2854),
.Y(n_3154)
);

INVx1_ASAP7_75t_L g3155 ( 
.A(n_2899),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_2868),
.B(n_2232),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_2902),
.Y(n_3157)
);

OR2x2_ASAP7_75t_L g3158 ( 
.A(n_2889),
.B(n_2548),
.Y(n_3158)
);

NAND2xp5_ASAP7_75t_L g3159 ( 
.A(n_2874),
.B(n_2117),
.Y(n_3159)
);

NAND2xp5_ASAP7_75t_L g3160 ( 
.A(n_2875),
.B(n_2117),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_3011),
.Y(n_3161)
);

OR2x6_ASAP7_75t_SL g3162 ( 
.A(n_3132),
.B(n_1024),
.Y(n_3162)
);

A2O1A1Ixp33_ASAP7_75t_L g3163 ( 
.A1(n_3070),
.A2(n_2835),
.B(n_2880),
.C(n_2878),
.Y(n_3163)
);

BUFx2_ASAP7_75t_L g3164 ( 
.A(n_2959),
.Y(n_3164)
);

AND2x4_ASAP7_75t_L g3165 ( 
.A(n_3032),
.B(n_2794),
.Y(n_3165)
);

AND2x2_ASAP7_75t_L g3166 ( 
.A(n_2991),
.B(n_3),
.Y(n_3166)
);

AOI22xp33_ASAP7_75t_L g3167 ( 
.A1(n_3069),
.A2(n_1742),
.B1(n_2954),
.B2(n_1024),
.Y(n_3167)
);

INVx2_ASAP7_75t_L g3168 ( 
.A(n_2985),
.Y(n_3168)
);

INVx3_ASAP7_75t_L g3169 ( 
.A(n_3084),
.Y(n_3169)
);

HB1xp67_ASAP7_75t_L g3170 ( 
.A(n_3011),
.Y(n_3170)
);

AOI22xp5_ASAP7_75t_L g3171 ( 
.A1(n_2993),
.A2(n_1742),
.B1(n_2503),
.B2(n_1599),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_2996),
.B(n_3),
.Y(n_3172)
);

O2A1O1Ixp5_ASAP7_75t_SL g3173 ( 
.A1(n_3066),
.A2(n_1743),
.B(n_2050),
.C(n_2042),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2990),
.Y(n_3174)
);

INVx1_ASAP7_75t_SL g3175 ( 
.A(n_3059),
.Y(n_3175)
);

NOR2xp33_ASAP7_75t_L g3176 ( 
.A(n_3094),
.B(n_4),
.Y(n_3176)
);

INVx2_ASAP7_75t_L g3177 ( 
.A(n_3008),
.Y(n_3177)
);

INVx3_ASAP7_75t_L g3178 ( 
.A(n_3084),
.Y(n_3178)
);

AND2x6_ASAP7_75t_L g3179 ( 
.A(n_3097),
.B(n_2042),
.Y(n_3179)
);

AND2x4_ASAP7_75t_L g3180 ( 
.A(n_2975),
.B(n_2050),
.Y(n_3180)
);

INVxp67_ASAP7_75t_L g3181 ( 
.A(n_3013),
.Y(n_3181)
);

OR2x6_ASAP7_75t_SL g3182 ( 
.A(n_3137),
.B(n_1974),
.Y(n_3182)
);

NAND2xp5_ASAP7_75t_L g3183 ( 
.A(n_3043),
.B(n_4),
.Y(n_3183)
);

AOI21x1_ASAP7_75t_L g3184 ( 
.A1(n_3014),
.A2(n_1927),
.B(n_1986),
.Y(n_3184)
);

BUFx2_ASAP7_75t_L g3185 ( 
.A(n_2963),
.Y(n_3185)
);

OAI21x1_ASAP7_75t_L g3186 ( 
.A1(n_3082),
.A2(n_1721),
.B(n_2080),
.Y(n_3186)
);

OAI21xp33_ASAP7_75t_SL g3187 ( 
.A1(n_3063),
.A2(n_2082),
.B(n_2080),
.Y(n_3187)
);

AOI22xp5_ASAP7_75t_L g3188 ( 
.A1(n_2965),
.A2(n_1742),
.B1(n_2503),
.B2(n_1599),
.Y(n_3188)
);

A2O1A1Ixp33_ASAP7_75t_SL g3189 ( 
.A1(n_3143),
.A2(n_2091),
.B(n_2104),
.C(n_2082),
.Y(n_3189)
);

INVxp67_ASAP7_75t_L g3190 ( 
.A(n_3017),
.Y(n_3190)
);

AND2x4_ASAP7_75t_L g3191 ( 
.A(n_2975),
.B(n_2091),
.Y(n_3191)
);

INVx4_ASAP7_75t_L g3192 ( 
.A(n_3084),
.Y(n_3192)
);

AOI21xp5_ASAP7_75t_L g3193 ( 
.A1(n_2972),
.A2(n_1869),
.B(n_1798),
.Y(n_3193)
);

BUFx2_ASAP7_75t_L g3194 ( 
.A(n_2971),
.Y(n_3194)
);

NAND2xp5_ASAP7_75t_SL g3195 ( 
.A(n_3059),
.B(n_2503),
.Y(n_3195)
);

BUFx2_ASAP7_75t_SL g3196 ( 
.A(n_2999),
.Y(n_3196)
);

NAND2xp5_ASAP7_75t_SL g3197 ( 
.A(n_3140),
.B(n_1599),
.Y(n_3197)
);

O2A1O1Ixp33_ASAP7_75t_L g3198 ( 
.A1(n_3030),
.A2(n_2111),
.B(n_2115),
.C(n_2104),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2970),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_3047),
.B(n_5),
.Y(n_3200)
);

BUFx6f_ASAP7_75t_L g3201 ( 
.A(n_2987),
.Y(n_3201)
);

AOI22xp33_ASAP7_75t_L g3202 ( 
.A1(n_3126),
.A2(n_1742),
.B1(n_2115),
.B2(n_2111),
.Y(n_3202)
);

INVx1_ASAP7_75t_SL g3203 ( 
.A(n_3016),
.Y(n_3203)
);

BUFx3_ASAP7_75t_L g3204 ( 
.A(n_2973),
.Y(n_3204)
);

OAI22x1_ASAP7_75t_L g3205 ( 
.A1(n_3063),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_3205)
);

BUFx8_ASAP7_75t_L g3206 ( 
.A(n_3007),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_3020),
.B(n_6),
.Y(n_3207)
);

OAI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_3026),
.A2(n_2280),
.B1(n_2132),
.B2(n_2152),
.Y(n_3208)
);

AOI21xp5_ASAP7_75t_L g3209 ( 
.A1(n_2972),
.A2(n_1869),
.B(n_1798),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_2976),
.Y(n_3210)
);

AO32x1_ASAP7_75t_L g3211 ( 
.A1(n_3109),
.A2(n_1986),
.A3(n_1947),
.B1(n_1869),
.B2(n_1798),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_L g3212 ( 
.A(n_3055),
.B(n_7),
.Y(n_3212)
);

BUFx6f_ASAP7_75t_L g3213 ( 
.A(n_2987),
.Y(n_3213)
);

NAND2xp5_ASAP7_75t_SL g3214 ( 
.A(n_3000),
.B(n_1599),
.Y(n_3214)
);

BUFx6f_ASAP7_75t_L g3215 ( 
.A(n_2987),
.Y(n_3215)
);

INVx3_ASAP7_75t_L g3216 ( 
.A(n_2986),
.Y(n_3216)
);

INVx3_ASAP7_75t_L g3217 ( 
.A(n_2986),
.Y(n_3217)
);

OR2x6_ASAP7_75t_L g3218 ( 
.A(n_2960),
.B(n_2132),
.Y(n_3218)
);

INVx1_ASAP7_75t_L g3219 ( 
.A(n_2978),
.Y(n_3219)
);

BUFx10_ASAP7_75t_L g3220 ( 
.A(n_2966),
.Y(n_3220)
);

BUFx3_ASAP7_75t_L g3221 ( 
.A(n_3029),
.Y(n_3221)
);

INVx4_ASAP7_75t_L g3222 ( 
.A(n_3089),
.Y(n_3222)
);

BUFx6f_ASAP7_75t_L g3223 ( 
.A(n_2988),
.Y(n_3223)
);

O2A1O1Ixp33_ASAP7_75t_L g3224 ( 
.A1(n_3079),
.A2(n_2152),
.B(n_2191),
.C(n_2140),
.Y(n_3224)
);

NAND2xp5_ASAP7_75t_SL g3225 ( 
.A(n_3125),
.B(n_2998),
.Y(n_3225)
);

AOI22xp33_ASAP7_75t_SL g3226 ( 
.A1(n_3119),
.A2(n_2191),
.B1(n_2210),
.B2(n_2140),
.Y(n_3226)
);

OAI22xp33_ASAP7_75t_L g3227 ( 
.A1(n_2960),
.A2(n_2211),
.B1(n_2215),
.B2(n_2210),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_2960),
.A2(n_2215),
.B1(n_2226),
.B2(n_2211),
.Y(n_3228)
);

BUFx6f_ASAP7_75t_L g3229 ( 
.A(n_2988),
.Y(n_3229)
);

BUFx5_ASAP7_75t_L g3230 ( 
.A(n_3155),
.Y(n_3230)
);

NAND2xp5_ASAP7_75t_L g3231 ( 
.A(n_3056),
.B(n_10),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_2984),
.Y(n_3232)
);

AOI21xp5_ASAP7_75t_L g3233 ( 
.A1(n_3130),
.A2(n_1947),
.B(n_2226),
.Y(n_3233)
);

OAI221xp5_ASAP7_75t_L g3234 ( 
.A1(n_3068),
.A2(n_1832),
.B1(n_1836),
.B2(n_1825),
.C(n_1817),
.Y(n_3234)
);

BUFx2_ASAP7_75t_L g3235 ( 
.A(n_2962),
.Y(n_3235)
);

NOR2xp33_ASAP7_75t_L g3236 ( 
.A(n_3003),
.B(n_11),
.Y(n_3236)
);

CKINVDCx6p67_ASAP7_75t_R g3237 ( 
.A(n_3025),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_3089),
.Y(n_3238)
);

AOI22xp33_ASAP7_75t_L g3239 ( 
.A1(n_3040),
.A2(n_2279),
.B1(n_2280),
.B2(n_2231),
.Y(n_3239)
);

BUFx2_ASAP7_75t_L g3240 ( 
.A(n_3088),
.Y(n_3240)
);

NAND2xp5_ASAP7_75t_L g3241 ( 
.A(n_3080),
.B(n_13),
.Y(n_3241)
);

BUFx6f_ASAP7_75t_L g3242 ( 
.A(n_2988),
.Y(n_3242)
);

INVx3_ASAP7_75t_L g3243 ( 
.A(n_3089),
.Y(n_3243)
);

OAI22xp5_ASAP7_75t_L g3244 ( 
.A1(n_3074),
.A2(n_2279),
.B1(n_2231),
.B2(n_1745),
.Y(n_3244)
);

NAND2xp5_ASAP7_75t_L g3245 ( 
.A(n_3051),
.B(n_14),
.Y(n_3245)
);

OAI22xp33_ASAP7_75t_L g3246 ( 
.A1(n_3079),
.A2(n_1745),
.B1(n_1781),
.B2(n_1773),
.Y(n_3246)
);

HB1xp67_ASAP7_75t_L g3247 ( 
.A(n_2982),
.Y(n_3247)
);

AOI22xp5_ASAP7_75t_L g3248 ( 
.A1(n_3049),
.A2(n_1825),
.B1(n_1832),
.B2(n_1817),
.Y(n_3248)
);

AOI21xp5_ASAP7_75t_L g3249 ( 
.A1(n_3050),
.A2(n_1947),
.B(n_1773),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3037),
.B(n_14),
.Y(n_3250)
);

A2O1A1Ixp33_ASAP7_75t_L g3251 ( 
.A1(n_3065),
.A2(n_1745),
.B(n_1781),
.C(n_1773),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3027),
.Y(n_3252)
);

NAND2xp5_ASAP7_75t_L g3253 ( 
.A(n_2964),
.B(n_15),
.Y(n_3253)
);

NAND2xp5_ASAP7_75t_SL g3254 ( 
.A(n_3125),
.B(n_1836),
.Y(n_3254)
);

NAND2xp5_ASAP7_75t_SL g3255 ( 
.A(n_3125),
.B(n_1781),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3036),
.B(n_15),
.Y(n_3256)
);

AND2x4_ASAP7_75t_L g3257 ( 
.A(n_2992),
.B(n_2995),
.Y(n_3257)
);

CKINVDCx5p33_ASAP7_75t_R g3258 ( 
.A(n_3029),
.Y(n_3258)
);

AND2x2_ASAP7_75t_L g3259 ( 
.A(n_3021),
.B(n_16),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_3044),
.B(n_3012),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3022),
.Y(n_3261)
);

AOI21xp5_ASAP7_75t_L g3262 ( 
.A1(n_3118),
.A2(n_1820),
.B(n_1796),
.Y(n_3262)
);

AOI21xp5_ASAP7_75t_L g3263 ( 
.A1(n_2968),
.A2(n_3083),
.B(n_3024),
.Y(n_3263)
);

BUFx2_ASAP7_75t_R g3264 ( 
.A(n_3018),
.Y(n_3264)
);

INVx1_ASAP7_75t_L g3265 ( 
.A(n_3031),
.Y(n_3265)
);

BUFx8_ASAP7_75t_L g3266 ( 
.A(n_3073),
.Y(n_3266)
);

AND2x4_ASAP7_75t_L g3267 ( 
.A(n_2981),
.B(n_1796),
.Y(n_3267)
);

HB1xp67_ASAP7_75t_L g3268 ( 
.A(n_3024),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3064),
.Y(n_3269)
);

O2A1O1Ixp33_ASAP7_75t_L g3270 ( 
.A1(n_3005),
.A2(n_1796),
.B(n_1856),
.C(n_1820),
.Y(n_3270)
);

AOI22xp5_ASAP7_75t_L g3271 ( 
.A1(n_3075),
.A2(n_1820),
.B1(n_1873),
.B2(n_1856),
.Y(n_3271)
);

INVx2_ASAP7_75t_L g3272 ( 
.A(n_2961),
.Y(n_3272)
);

AOI21xp5_ASAP7_75t_L g3273 ( 
.A1(n_2968),
.A2(n_1873),
.B(n_1856),
.Y(n_3273)
);

AOI21xp5_ASAP7_75t_L g3274 ( 
.A1(n_3142),
.A2(n_1941),
.B(n_1873),
.Y(n_3274)
);

OR2x6_ASAP7_75t_L g3275 ( 
.A(n_2981),
.B(n_1941),
.Y(n_3275)
);

NAND2xp5_ASAP7_75t_L g3276 ( 
.A(n_3001),
.B(n_16),
.Y(n_3276)
);

NAND2xp5_ASAP7_75t_SL g3277 ( 
.A(n_3108),
.B(n_2989),
.Y(n_3277)
);

BUFx6f_ASAP7_75t_L g3278 ( 
.A(n_2997),
.Y(n_3278)
);

O2A1O1Ixp33_ASAP7_75t_L g3279 ( 
.A1(n_3085),
.A2(n_3061),
.B(n_3100),
.C(n_3052),
.Y(n_3279)
);

O2A1O1Ixp33_ASAP7_75t_SL g3280 ( 
.A1(n_3111),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_3280)
);

AOI21xp5_ASAP7_75t_L g3281 ( 
.A1(n_3146),
.A2(n_1954),
.B(n_1941),
.Y(n_3281)
);

INVxp67_ASAP7_75t_L g3282 ( 
.A(n_3060),
.Y(n_3282)
);

BUFx2_ASAP7_75t_L g3283 ( 
.A(n_3058),
.Y(n_3283)
);

INVx5_ASAP7_75t_SL g3284 ( 
.A(n_3077),
.Y(n_3284)
);

OAI22xp5_ASAP7_75t_L g3285 ( 
.A1(n_3053),
.A2(n_1955),
.B1(n_1958),
.B2(n_1954),
.Y(n_3285)
);

OAI22xp5_ASAP7_75t_L g3286 ( 
.A1(n_3093),
.A2(n_1955),
.B1(n_1958),
.B2(n_1954),
.Y(n_3286)
);

O2A1O1Ixp5_ASAP7_75t_SL g3287 ( 
.A1(n_3090),
.A2(n_1955),
.B(n_1958),
.C(n_1721),
.Y(n_3287)
);

INVx3_ASAP7_75t_L g3288 ( 
.A(n_2977),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3098),
.Y(n_3289)
);

HB1xp67_ASAP7_75t_L g3290 ( 
.A(n_3128),
.Y(n_3290)
);

BUFx12f_ASAP7_75t_L g3291 ( 
.A(n_3077),
.Y(n_3291)
);

HB1xp67_ASAP7_75t_L g3292 ( 
.A(n_3033),
.Y(n_3292)
);

NAND2xp5_ASAP7_75t_L g3293 ( 
.A(n_3004),
.B(n_19),
.Y(n_3293)
);

AOI21xp5_ASAP7_75t_L g3294 ( 
.A1(n_3122),
.A2(n_1980),
.B(n_1815),
.Y(n_3294)
);

INVx2_ASAP7_75t_L g3295 ( 
.A(n_2969),
.Y(n_3295)
);

INVx2_ASAP7_75t_L g3296 ( 
.A(n_2974),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2979),
.Y(n_3297)
);

O2A1O1Ixp33_ASAP7_75t_L g3298 ( 
.A1(n_3145),
.A2(n_1721),
.B(n_23),
.C(n_21),
.Y(n_3298)
);

INVxp67_ASAP7_75t_L g3299 ( 
.A(n_3076),
.Y(n_3299)
);

BUFx3_ASAP7_75t_L g3300 ( 
.A(n_3077),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_2980),
.Y(n_3301)
);

BUFx6f_ASAP7_75t_L g3302 ( 
.A(n_2997),
.Y(n_3302)
);

BUFx2_ASAP7_75t_L g3303 ( 
.A(n_3095),
.Y(n_3303)
);

NAND2xp5_ASAP7_75t_L g3304 ( 
.A(n_3009),
.B(n_21),
.Y(n_3304)
);

INVx2_ASAP7_75t_L g3305 ( 
.A(n_3038),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3042),
.Y(n_3306)
);

BUFx3_ASAP7_75t_L g3307 ( 
.A(n_2997),
.Y(n_3307)
);

INVx1_ASAP7_75t_L g3308 ( 
.A(n_3157),
.Y(n_3308)
);

AND2x2_ASAP7_75t_L g3309 ( 
.A(n_3099),
.B(n_22),
.Y(n_3309)
);

INVx3_ASAP7_75t_L g3310 ( 
.A(n_2977),
.Y(n_3310)
);

OAI22xp5_ASAP7_75t_L g3311 ( 
.A1(n_3127),
.A2(n_1815),
.B1(n_1766),
.B2(n_1980),
.Y(n_3311)
);

AND2x4_ASAP7_75t_L g3312 ( 
.A(n_2981),
.B(n_250),
.Y(n_3312)
);

INVx3_ASAP7_75t_L g3313 ( 
.A(n_3002),
.Y(n_3313)
);

INVx5_ASAP7_75t_L g3314 ( 
.A(n_3154),
.Y(n_3314)
);

HB1xp67_ASAP7_75t_L g3315 ( 
.A(n_3033),
.Y(n_3315)
);

INVx2_ASAP7_75t_SL g3316 ( 
.A(n_3006),
.Y(n_3316)
);

A2O1A1Ixp33_ASAP7_75t_L g3317 ( 
.A1(n_3108),
.A2(n_25),
.B(n_23),
.C(n_24),
.Y(n_3317)
);

NAND2xp5_ASAP7_75t_L g3318 ( 
.A(n_3015),
.B(n_25),
.Y(n_3318)
);

A2O1A1Ixp33_ASAP7_75t_L g3319 ( 
.A1(n_3102),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_3319)
);

AOI22xp33_ASAP7_75t_L g3320 ( 
.A1(n_3153),
.A2(n_1766),
.B1(n_821),
.B2(n_877),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3105),
.Y(n_3321)
);

OAI21x1_ASAP7_75t_L g3322 ( 
.A1(n_3112),
.A2(n_253),
.B(n_252),
.Y(n_3322)
);

INVx2_ASAP7_75t_L g3323 ( 
.A(n_3034),
.Y(n_3323)
);

BUFx6f_ASAP7_75t_L g3324 ( 
.A(n_3006),
.Y(n_3324)
);

INVx2_ASAP7_75t_L g3325 ( 
.A(n_3158),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_3105),
.Y(n_3326)
);

BUFx2_ASAP7_75t_L g3327 ( 
.A(n_3019),
.Y(n_3327)
);

INVx2_ASAP7_75t_L g3328 ( 
.A(n_3019),
.Y(n_3328)
);

A2O1A1Ixp33_ASAP7_75t_L g3329 ( 
.A1(n_3120),
.A2(n_3106),
.B(n_3114),
.C(n_3104),
.Y(n_3329)
);

O2A1O1Ixp5_ASAP7_75t_L g3330 ( 
.A1(n_3153),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_3330)
);

INVx2_ASAP7_75t_L g3331 ( 
.A(n_3028),
.Y(n_3331)
);

AND2x4_ASAP7_75t_L g3332 ( 
.A(n_3028),
.B(n_254),
.Y(n_3332)
);

NAND2xp5_ASAP7_75t_L g3333 ( 
.A(n_2983),
.B(n_31),
.Y(n_3333)
);

AOI22xp5_ASAP7_75t_L g3334 ( 
.A1(n_3091),
.A2(n_821),
.B1(n_877),
.B2(n_794),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_3086),
.Y(n_3335)
);

NAND2xp5_ASAP7_75t_SL g3336 ( 
.A(n_3035),
.B(n_821),
.Y(n_3336)
);

NAND2x1_ASAP7_75t_SL g3337 ( 
.A(n_3117),
.B(n_31),
.Y(n_3337)
);

CKINVDCx8_ASAP7_75t_R g3338 ( 
.A(n_3006),
.Y(n_3338)
);

O2A1O1Ixp33_ASAP7_75t_L g3339 ( 
.A1(n_3067),
.A2(n_34),
.B(n_32),
.C(n_33),
.Y(n_3339)
);

AND2x2_ASAP7_75t_L g3340 ( 
.A(n_3035),
.B(n_32),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_L g3341 ( 
.A(n_2994),
.B(n_33),
.Y(n_3341)
);

INVx1_ASAP7_75t_L g3342 ( 
.A(n_3144),
.Y(n_3342)
);

NAND2xp5_ASAP7_75t_SL g3343 ( 
.A(n_3101),
.B(n_3002),
.Y(n_3343)
);

NAND2xp5_ASAP7_75t_L g3344 ( 
.A(n_3081),
.B(n_34),
.Y(n_3344)
);

NOR2xp33_ASAP7_75t_L g3345 ( 
.A(n_3039),
.B(n_35),
.Y(n_3345)
);

INVx1_ASAP7_75t_L g3346 ( 
.A(n_3144),
.Y(n_3346)
);

INVx5_ASAP7_75t_L g3347 ( 
.A(n_3154),
.Y(n_3347)
);

AOI21xp5_ASAP7_75t_L g3348 ( 
.A1(n_3122),
.A2(n_877),
.B(n_821),
.Y(n_3348)
);

BUFx2_ASAP7_75t_L g3349 ( 
.A(n_3010),
.Y(n_3349)
);

A2O1A1Ixp33_ASAP7_75t_L g3350 ( 
.A1(n_3133),
.A2(n_40),
.B(n_36),
.C(n_38),
.Y(n_3350)
);

INVx1_ASAP7_75t_L g3351 ( 
.A(n_3141),
.Y(n_3351)
);

HB1xp67_ASAP7_75t_L g3352 ( 
.A(n_3147),
.Y(n_3352)
);

INVx1_ASAP7_75t_L g3353 ( 
.A(n_3141),
.Y(n_3353)
);

INVx3_ASAP7_75t_L g3354 ( 
.A(n_3010),
.Y(n_3354)
);

AOI22xp33_ASAP7_75t_L g3355 ( 
.A1(n_3113),
.A2(n_941),
.B1(n_982),
.B2(n_877),
.Y(n_3355)
);

BUFx2_ASAP7_75t_L g3356 ( 
.A(n_3010),
.Y(n_3356)
);

BUFx6f_ASAP7_75t_L g3357 ( 
.A(n_3023),
.Y(n_3357)
);

NOR2xp33_ASAP7_75t_L g3358 ( 
.A(n_3039),
.B(n_40),
.Y(n_3358)
);

INVx2_ASAP7_75t_L g3359 ( 
.A(n_3150),
.Y(n_3359)
);

INVx5_ASAP7_75t_L g3360 ( 
.A(n_3154),
.Y(n_3360)
);

INVx6_ASAP7_75t_L g3361 ( 
.A(n_3023),
.Y(n_3361)
);

NAND2xp5_ASAP7_75t_L g3362 ( 
.A(n_3121),
.B(n_41),
.Y(n_3362)
);

AOI21xp5_ASAP7_75t_L g3363 ( 
.A1(n_3054),
.A2(n_982),
.B(n_941),
.Y(n_3363)
);

BUFx2_ASAP7_75t_L g3364 ( 
.A(n_3023),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_3124),
.Y(n_3365)
);

NAND2xp5_ASAP7_75t_L g3366 ( 
.A(n_3136),
.B(n_42),
.Y(n_3366)
);

INVx2_ASAP7_75t_L g3367 ( 
.A(n_3048),
.Y(n_3367)
);

HB1xp67_ASAP7_75t_L g3368 ( 
.A(n_3151),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_L g3369 ( 
.A(n_3103),
.B(n_44),
.Y(n_3369)
);

OAI22xp5_ASAP7_75t_L g3370 ( 
.A1(n_3087),
.A2(n_1071),
.B1(n_982),
.B2(n_941),
.Y(n_3370)
);

HB1xp67_ASAP7_75t_L g3371 ( 
.A(n_3151),
.Y(n_3371)
);

INVx3_ASAP7_75t_L g3372 ( 
.A(n_3257),
.Y(n_3372)
);

AND2x2_ASAP7_75t_L g3373 ( 
.A(n_3235),
.B(n_3135),
.Y(n_3373)
);

AOI21xp5_ASAP7_75t_L g3374 ( 
.A1(n_3263),
.A2(n_3062),
.B(n_3124),
.Y(n_3374)
);

AND2x2_ASAP7_75t_SL g3375 ( 
.A(n_3312),
.B(n_2967),
.Y(n_3375)
);

INVx2_ASAP7_75t_L g3376 ( 
.A(n_3257),
.Y(n_3376)
);

NAND2xp5_ASAP7_75t_L g3377 ( 
.A(n_3268),
.B(n_3110),
.Y(n_3377)
);

BUFx3_ASAP7_75t_L g3378 ( 
.A(n_3206),
.Y(n_3378)
);

AO22x1_ASAP7_75t_L g3379 ( 
.A1(n_3194),
.A2(n_3057),
.B1(n_3123),
.B2(n_3101),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3290),
.B(n_3110),
.Y(n_3380)
);

INVx2_ASAP7_75t_L g3381 ( 
.A(n_3325),
.Y(n_3381)
);

INVx3_ASAP7_75t_L g3382 ( 
.A(n_3222),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3214),
.A2(n_3115),
.B1(n_3139),
.B2(n_3134),
.Y(n_3383)
);

AOI22xp33_ASAP7_75t_L g3384 ( 
.A1(n_3236),
.A2(n_3115),
.B1(n_3046),
.B2(n_3138),
.Y(n_3384)
);

OAI22xp5_ASAP7_75t_L g3385 ( 
.A1(n_3350),
.A2(n_3129),
.B1(n_3131),
.B2(n_3123),
.Y(n_3385)
);

INVx4_ASAP7_75t_SL g3386 ( 
.A(n_3221),
.Y(n_3386)
);

NOR2xp67_ASAP7_75t_L g3387 ( 
.A(n_3335),
.B(n_3123),
.Y(n_3387)
);

INVx1_ASAP7_75t_L g3388 ( 
.A(n_3199),
.Y(n_3388)
);

INVx2_ASAP7_75t_L g3389 ( 
.A(n_3168),
.Y(n_3389)
);

AOI22xp5_ASAP7_75t_L g3390 ( 
.A1(n_3317),
.A2(n_3129),
.B1(n_3115),
.B2(n_3096),
.Y(n_3390)
);

OAI22xp5_ASAP7_75t_L g3391 ( 
.A1(n_3319),
.A2(n_3041),
.B1(n_3045),
.B2(n_2967),
.Y(n_3391)
);

OAI21x1_ASAP7_75t_L g3392 ( 
.A1(n_3287),
.A2(n_3348),
.B(n_3173),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3210),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3219),
.Y(n_3394)
);

AOI22xp33_ASAP7_75t_L g3395 ( 
.A1(n_3352),
.A2(n_3115),
.B1(n_3078),
.B2(n_3071),
.Y(n_3395)
);

INVx2_ASAP7_75t_L g3396 ( 
.A(n_3174),
.Y(n_3396)
);

INVx3_ASAP7_75t_L g3397 ( 
.A(n_3222),
.Y(n_3397)
);

NOR2xp33_ASAP7_75t_SL g3398 ( 
.A(n_3264),
.B(n_3041),
.Y(n_3398)
);

OR2x6_ASAP7_75t_L g3399 ( 
.A(n_3218),
.B(n_3116),
.Y(n_3399)
);

O2A1O1Ixp33_ASAP7_75t_L g3400 ( 
.A1(n_3298),
.A2(n_3160),
.B(n_3159),
.C(n_3149),
.Y(n_3400)
);

BUFx6f_ASAP7_75t_L g3401 ( 
.A(n_3201),
.Y(n_3401)
);

A2O1A1Ixp33_ASAP7_75t_L g3402 ( 
.A1(n_3339),
.A2(n_3045),
.B(n_3092),
.C(n_3103),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3232),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3261),
.Y(n_3404)
);

NAND2xp5_ASAP7_75t_L g3405 ( 
.A(n_3292),
.B(n_3156),
.Y(n_3405)
);

OR2x6_ASAP7_75t_L g3406 ( 
.A(n_3218),
.B(n_3116),
.Y(n_3406)
);

CKINVDCx11_ASAP7_75t_R g3407 ( 
.A(n_3220),
.Y(n_3407)
);

AOI22xp33_ASAP7_75t_L g3408 ( 
.A1(n_3312),
.A2(n_3078),
.B1(n_3071),
.B2(n_3057),
.Y(n_3408)
);

INVx5_ASAP7_75t_L g3409 ( 
.A(n_3179),
.Y(n_3409)
);

BUFx8_ASAP7_75t_L g3410 ( 
.A(n_3283),
.Y(n_3410)
);

NAND2xp5_ASAP7_75t_L g3411 ( 
.A(n_3315),
.B(n_3107),
.Y(n_3411)
);

INVx3_ASAP7_75t_L g3412 ( 
.A(n_3238),
.Y(n_3412)
);

AND2x2_ASAP7_75t_L g3413 ( 
.A(n_3164),
.B(n_3185),
.Y(n_3413)
);

CKINVDCx6p67_ASAP7_75t_R g3414 ( 
.A(n_3196),
.Y(n_3414)
);

INVx2_ASAP7_75t_SL g3415 ( 
.A(n_3204),
.Y(n_3415)
);

INVxp67_ASAP7_75t_L g3416 ( 
.A(n_3161),
.Y(n_3416)
);

INVx1_ASAP7_75t_L g3417 ( 
.A(n_3265),
.Y(n_3417)
);

AOI221xp5_ASAP7_75t_L g3418 ( 
.A1(n_3205),
.A2(n_3148),
.B1(n_3152),
.B2(n_3159),
.C(n_3160),
.Y(n_3418)
);

BUFx6f_ASAP7_75t_L g3419 ( 
.A(n_3201),
.Y(n_3419)
);

NOR2xp33_ASAP7_75t_SL g3420 ( 
.A(n_3314),
.B(n_3347),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3342),
.B(n_3116),
.Y(n_3421)
);

NAND2xp33_ASAP7_75t_L g3422 ( 
.A(n_3258),
.B(n_3057),
.Y(n_3422)
);

BUFx2_ASAP7_75t_L g3423 ( 
.A(n_3240),
.Y(n_3423)
);

INVx2_ASAP7_75t_SL g3424 ( 
.A(n_3266),
.Y(n_3424)
);

INVx1_ASAP7_75t_L g3425 ( 
.A(n_3289),
.Y(n_3425)
);

AOI22xp33_ASAP7_75t_L g3426 ( 
.A1(n_3197),
.A2(n_3057),
.B1(n_3072),
.B2(n_3048),
.Y(n_3426)
);

NOR2xp33_ASAP7_75t_L g3427 ( 
.A(n_3299),
.B(n_3072),
.Y(n_3427)
);

AOI22xp33_ASAP7_75t_L g3428 ( 
.A1(n_3225),
.A2(n_3072),
.B1(n_3096),
.B2(n_982),
.Y(n_3428)
);

INVx2_ASAP7_75t_L g3429 ( 
.A(n_3177),
.Y(n_3429)
);

AOI21xp5_ASAP7_75t_L g3430 ( 
.A1(n_3279),
.A2(n_1071),
.B(n_941),
.Y(n_3430)
);

NAND2xp5_ASAP7_75t_L g3431 ( 
.A(n_3247),
.B(n_3170),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3252),
.Y(n_3432)
);

INVx5_ASAP7_75t_L g3433 ( 
.A(n_3179),
.Y(n_3433)
);

INVxp67_ASAP7_75t_SL g3434 ( 
.A(n_3269),
.Y(n_3434)
);

NAND2xp33_ASAP7_75t_L g3435 ( 
.A(n_3179),
.B(n_1071),
.Y(n_3435)
);

INVx3_ASAP7_75t_L g3436 ( 
.A(n_3238),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3346),
.B(n_3351),
.Y(n_3437)
);

AND2x2_ASAP7_75t_SL g3438 ( 
.A(n_3303),
.B(n_1071),
.Y(n_3438)
);

BUFx6f_ASAP7_75t_L g3439 ( 
.A(n_3201),
.Y(n_3439)
);

NAND2xp5_ASAP7_75t_L g3440 ( 
.A(n_3301),
.B(n_44),
.Y(n_3440)
);

BUFx2_ASAP7_75t_L g3441 ( 
.A(n_3368),
.Y(n_3441)
);

AOI21xp5_ASAP7_75t_L g3442 ( 
.A1(n_3163),
.A2(n_45),
.B(n_46),
.Y(n_3442)
);

AOI22xp33_ASAP7_75t_L g3443 ( 
.A1(n_3176),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_3443)
);

AOI21xp5_ASAP7_75t_L g3444 ( 
.A1(n_3193),
.A2(n_48),
.B(n_49),
.Y(n_3444)
);

INVx3_ASAP7_75t_L g3445 ( 
.A(n_3243),
.Y(n_3445)
);

NAND2xp5_ASAP7_75t_L g3446 ( 
.A(n_3260),
.B(n_49),
.Y(n_3446)
);

AOI22xp5_ASAP7_75t_L g3447 ( 
.A1(n_3280),
.A2(n_53),
.B1(n_51),
.B2(n_52),
.Y(n_3447)
);

INVx2_ASAP7_75t_L g3448 ( 
.A(n_3305),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3308),
.Y(n_3449)
);

BUFx2_ASAP7_75t_L g3450 ( 
.A(n_3371),
.Y(n_3450)
);

NAND2xp5_ASAP7_75t_L g3451 ( 
.A(n_3190),
.B(n_51),
.Y(n_3451)
);

HB1xp67_ASAP7_75t_L g3452 ( 
.A(n_3181),
.Y(n_3452)
);

NOR2x1_ASAP7_75t_SL g3453 ( 
.A(n_3275),
.B(n_52),
.Y(n_3453)
);

AOI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3209),
.A2(n_57),
.B(n_58),
.Y(n_3454)
);

CKINVDCx5p33_ASAP7_75t_R g3455 ( 
.A(n_3206),
.Y(n_3455)
);

AO21x1_ASAP7_75t_L g3456 ( 
.A1(n_3183),
.A2(n_57),
.B(n_59),
.Y(n_3456)
);

INVx3_ASAP7_75t_L g3457 ( 
.A(n_3243),
.Y(n_3457)
);

NOR2xp67_ASAP7_75t_L g3458 ( 
.A(n_3314),
.B(n_60),
.Y(n_3458)
);

INVx1_ASAP7_75t_SL g3459 ( 
.A(n_3175),
.Y(n_3459)
);

BUFx3_ASAP7_75t_L g3460 ( 
.A(n_3220),
.Y(n_3460)
);

INVx2_ASAP7_75t_L g3461 ( 
.A(n_3306),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3297),
.Y(n_3462)
);

OAI21xp33_ASAP7_75t_L g3463 ( 
.A1(n_3344),
.A2(n_3366),
.B(n_3253),
.Y(n_3463)
);

AOI222xp33_ASAP7_75t_L g3464 ( 
.A1(n_3333),
.A2(n_60),
.B1(n_61),
.B2(n_64),
.C1(n_65),
.C2(n_66),
.Y(n_3464)
);

INVx4_ASAP7_75t_L g3465 ( 
.A(n_3213),
.Y(n_3465)
);

INVx2_ASAP7_75t_L g3466 ( 
.A(n_3272),
.Y(n_3466)
);

BUFx2_ASAP7_75t_L g3467 ( 
.A(n_3216),
.Y(n_3467)
);

AND2x4_ASAP7_75t_L g3468 ( 
.A(n_3217),
.B(n_3165),
.Y(n_3468)
);

AOI22xp33_ASAP7_75t_L g3469 ( 
.A1(n_3277),
.A2(n_67),
.B1(n_61),
.B2(n_65),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_3314),
.B(n_255),
.Y(n_3470)
);

AND2x2_ASAP7_75t_L g3471 ( 
.A(n_3217),
.B(n_68),
.Y(n_3471)
);

INVx2_ASAP7_75t_SL g3472 ( 
.A(n_3266),
.Y(n_3472)
);

BUFx3_ASAP7_75t_L g3473 ( 
.A(n_3291),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3353),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3295),
.Y(n_3475)
);

BUFx6f_ASAP7_75t_L g3476 ( 
.A(n_3213),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3365),
.B(n_3321),
.Y(n_3477)
);

INVx4_ASAP7_75t_L g3478 ( 
.A(n_3213),
.Y(n_3478)
);

AND2x2_ASAP7_75t_L g3479 ( 
.A(n_3327),
.B(n_69),
.Y(n_3479)
);

BUFx6f_ASAP7_75t_L g3480 ( 
.A(n_3215),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3296),
.Y(n_3481)
);

NOR2xp33_ASAP7_75t_L g3482 ( 
.A(n_3162),
.B(n_70),
.Y(n_3482)
);

AOI22xp33_ASAP7_75t_L g3483 ( 
.A1(n_3166),
.A2(n_73),
.B1(n_70),
.B2(n_72),
.Y(n_3483)
);

BUFx3_ASAP7_75t_L g3484 ( 
.A(n_3300),
.Y(n_3484)
);

BUFx2_ASAP7_75t_L g3485 ( 
.A(n_3349),
.Y(n_3485)
);

AND2x4_ASAP7_75t_L g3486 ( 
.A(n_3165),
.B(n_72),
.Y(n_3486)
);

NAND2xp5_ASAP7_75t_L g3487 ( 
.A(n_3326),
.B(n_74),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_SL g3488 ( 
.A(n_3347),
.B(n_256),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3359),
.Y(n_3489)
);

BUFx6f_ASAP7_75t_L g3490 ( 
.A(n_3215),
.Y(n_3490)
);

BUFx2_ASAP7_75t_L g3491 ( 
.A(n_3356),
.Y(n_3491)
);

NAND2xp5_ASAP7_75t_L g3492 ( 
.A(n_3323),
.B(n_75),
.Y(n_3492)
);

INVx1_ASAP7_75t_L g3493 ( 
.A(n_3328),
.Y(n_3493)
);

BUFx3_ASAP7_75t_L g3494 ( 
.A(n_3307),
.Y(n_3494)
);

AND2x2_ASAP7_75t_L g3495 ( 
.A(n_3282),
.B(n_76),
.Y(n_3495)
);

INVx2_ASAP7_75t_SL g3496 ( 
.A(n_3361),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3329),
.B(n_77),
.Y(n_3497)
);

INVx3_ASAP7_75t_SL g3498 ( 
.A(n_3237),
.Y(n_3498)
);

AOI21xp5_ASAP7_75t_L g3499 ( 
.A1(n_3233),
.A2(n_79),
.B(n_80),
.Y(n_3499)
);

BUFx3_ASAP7_75t_L g3500 ( 
.A(n_3361),
.Y(n_3500)
);

CKINVDCx16_ASAP7_75t_R g3501 ( 
.A(n_3182),
.Y(n_3501)
);

OR2x2_ASAP7_75t_L g3502 ( 
.A(n_3331),
.B(n_81),
.Y(n_3502)
);

AOI21xp5_ASAP7_75t_L g3503 ( 
.A1(n_3270),
.A2(n_81),
.B(n_82),
.Y(n_3503)
);

INVx2_ASAP7_75t_L g3504 ( 
.A(n_3288),
.Y(n_3504)
);

NAND2xp5_ASAP7_75t_L g3505 ( 
.A(n_3230),
.B(n_82),
.Y(n_3505)
);

NAND2xp5_ASAP7_75t_L g3506 ( 
.A(n_3230),
.B(n_83),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3288),
.Y(n_3507)
);

NAND2xp5_ASAP7_75t_L g3508 ( 
.A(n_3230),
.B(n_83),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3310),
.Y(n_3509)
);

INVx2_ASAP7_75t_SL g3510 ( 
.A(n_3215),
.Y(n_3510)
);

AOI22xp33_ASAP7_75t_L g3511 ( 
.A1(n_3309),
.A2(n_87),
.B1(n_84),
.B2(n_85),
.Y(n_3511)
);

BUFx2_ASAP7_75t_L g3512 ( 
.A(n_3364),
.Y(n_3512)
);

INVx5_ASAP7_75t_L g3513 ( 
.A(n_3179),
.Y(n_3513)
);

INVxp67_ASAP7_75t_SL g3514 ( 
.A(n_3310),
.Y(n_3514)
);

NOR2xp33_ASAP7_75t_L g3515 ( 
.A(n_3203),
.B(n_85),
.Y(n_3515)
);

BUFx6f_ASAP7_75t_L g3516 ( 
.A(n_3223),
.Y(n_3516)
);

NAND2xp5_ASAP7_75t_L g3517 ( 
.A(n_3230),
.B(n_88),
.Y(n_3517)
);

INVx3_ASAP7_75t_SL g3518 ( 
.A(n_3207),
.Y(n_3518)
);

AND2x2_ASAP7_75t_L g3519 ( 
.A(n_3172),
.B(n_88),
.Y(n_3519)
);

NOR2x1_ASAP7_75t_L g3520 ( 
.A(n_3313),
.B(n_89),
.Y(n_3520)
);

INVxp67_ASAP7_75t_SL g3521 ( 
.A(n_3313),
.Y(n_3521)
);

NOR2x1_ASAP7_75t_L g3522 ( 
.A(n_3192),
.B(n_91),
.Y(n_3522)
);

INVx3_ASAP7_75t_L g3523 ( 
.A(n_3192),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3367),
.Y(n_3524)
);

NAND2xp5_ASAP7_75t_L g3525 ( 
.A(n_3276),
.B(n_92),
.Y(n_3525)
);

OR2x4_ASAP7_75t_L g3526 ( 
.A(n_3369),
.B(n_93),
.Y(n_3526)
);

INVx2_ASAP7_75t_SL g3527 ( 
.A(n_3223),
.Y(n_3527)
);

INVx1_ASAP7_75t_L g3528 ( 
.A(n_3259),
.Y(n_3528)
);

INVx3_ASAP7_75t_L g3529 ( 
.A(n_3169),
.Y(n_3529)
);

INVxp67_ASAP7_75t_L g3530 ( 
.A(n_3293),
.Y(n_3530)
);

AND2x4_ASAP7_75t_L g3531 ( 
.A(n_3275),
.B(n_93),
.Y(n_3531)
);

BUFx3_ASAP7_75t_L g3532 ( 
.A(n_3223),
.Y(n_3532)
);

INVx2_ASAP7_75t_L g3533 ( 
.A(n_3343),
.Y(n_3533)
);

BUFx3_ASAP7_75t_L g3534 ( 
.A(n_3229),
.Y(n_3534)
);

HB1xp67_ASAP7_75t_L g3535 ( 
.A(n_3195),
.Y(n_3535)
);

NOR2xp33_ASAP7_75t_L g3536 ( 
.A(n_3304),
.B(n_95),
.Y(n_3536)
);

NAND2xp5_ASAP7_75t_L g3537 ( 
.A(n_3318),
.B(n_95),
.Y(n_3537)
);

INVx1_ASAP7_75t_L g3538 ( 
.A(n_3256),
.Y(n_3538)
);

INVx1_ASAP7_75t_L g3539 ( 
.A(n_3241),
.Y(n_3539)
);

NOR2xp33_ASAP7_75t_L g3540 ( 
.A(n_3463),
.B(n_3341),
.Y(n_3540)
);

AOI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3464),
.A2(n_3171),
.B1(n_3187),
.B2(n_3345),
.Y(n_3541)
);

A2O1A1Ixp33_ASAP7_75t_SL g3542 ( 
.A1(n_3442),
.A2(n_3358),
.B(n_3362),
.C(n_3200),
.Y(n_3542)
);

INVx1_ASAP7_75t_L g3543 ( 
.A(n_3425),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3388),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3463),
.B(n_3245),
.Y(n_3545)
);

OAI21x1_ASAP7_75t_L g3546 ( 
.A1(n_3374),
.A2(n_3262),
.B(n_3184),
.Y(n_3546)
);

OR2x6_ASAP7_75t_L g3547 ( 
.A(n_3379),
.B(n_3281),
.Y(n_3547)
);

A2O1A1Ixp33_ASAP7_75t_L g3548 ( 
.A1(n_3447),
.A2(n_3337),
.B(n_3330),
.C(n_3224),
.Y(n_3548)
);

NAND2xp5_ASAP7_75t_L g3549 ( 
.A(n_3474),
.B(n_3212),
.Y(n_3549)
);

INVx2_ASAP7_75t_L g3550 ( 
.A(n_3372),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3423),
.B(n_3178),
.Y(n_3551)
);

INVx2_ASAP7_75t_L g3552 ( 
.A(n_3372),
.Y(n_3552)
);

OAI21x1_ASAP7_75t_L g3553 ( 
.A1(n_3430),
.A2(n_3186),
.B(n_3273),
.Y(n_3553)
);

OAI21x1_ASAP7_75t_L g3554 ( 
.A1(n_3505),
.A2(n_3508),
.B(n_3506),
.Y(n_3554)
);

AND2x2_ASAP7_75t_L g3555 ( 
.A(n_3441),
.B(n_3178),
.Y(n_3555)
);

INVx1_ASAP7_75t_L g3556 ( 
.A(n_3393),
.Y(n_3556)
);

AOI21xp5_ASAP7_75t_L g3557 ( 
.A1(n_3435),
.A2(n_3211),
.B(n_3347),
.Y(n_3557)
);

NAND2xp5_ASAP7_75t_L g3558 ( 
.A(n_3434),
.B(n_3231),
.Y(n_3558)
);

OA21x2_ASAP7_75t_L g3559 ( 
.A1(n_3377),
.A2(n_3294),
.B(n_3363),
.Y(n_3559)
);

AOI22x1_ASAP7_75t_L g3560 ( 
.A1(n_3464),
.A2(n_3340),
.B1(n_3250),
.B2(n_3332),
.Y(n_3560)
);

INVx2_ASAP7_75t_L g3561 ( 
.A(n_3376),
.Y(n_3561)
);

OAI22xp5_ASAP7_75t_L g3562 ( 
.A1(n_3447),
.A2(n_3226),
.B1(n_3228),
.B2(n_3167),
.Y(n_3562)
);

OAI21xp5_ASAP7_75t_L g3563 ( 
.A1(n_3499),
.A2(n_3251),
.B(n_3198),
.Y(n_3563)
);

OAI21x1_ASAP7_75t_L g3564 ( 
.A1(n_3505),
.A2(n_3322),
.B(n_3255),
.Y(n_3564)
);

NAND2x1p5_ASAP7_75t_L g3565 ( 
.A(n_3409),
.B(n_3360),
.Y(n_3565)
);

OAI21x1_ASAP7_75t_L g3566 ( 
.A1(n_3506),
.A2(n_3249),
.B(n_3274),
.Y(n_3566)
);

AND2x2_ASAP7_75t_L g3567 ( 
.A(n_3450),
.B(n_3360),
.Y(n_3567)
);

AO32x2_ASAP7_75t_L g3568 ( 
.A1(n_3510),
.A2(n_3316),
.A3(n_3311),
.B1(n_3244),
.B2(n_3286),
.Y(n_3568)
);

INVxp67_ASAP7_75t_SL g3569 ( 
.A(n_3377),
.Y(n_3569)
);

OA21x2_ASAP7_75t_L g3570 ( 
.A1(n_3387),
.A2(n_3254),
.B(n_3336),
.Y(n_3570)
);

OAI21x1_ASAP7_75t_L g3571 ( 
.A1(n_3517),
.A2(n_3354),
.B(n_3320),
.Y(n_3571)
);

INVx1_ASAP7_75t_L g3572 ( 
.A(n_3394),
.Y(n_3572)
);

OAI21x1_ASAP7_75t_L g3573 ( 
.A1(n_3517),
.A2(n_3355),
.B(n_3334),
.Y(n_3573)
);

INVx1_ASAP7_75t_L g3574 ( 
.A(n_3403),
.Y(n_3574)
);

NAND2xp5_ASAP7_75t_L g3575 ( 
.A(n_3437),
.B(n_3416),
.Y(n_3575)
);

INVx1_ASAP7_75t_L g3576 ( 
.A(n_3404),
.Y(n_3576)
);

INVx2_ASAP7_75t_SL g3577 ( 
.A(n_3410),
.Y(n_3577)
);

O2A1O1Ixp33_ASAP7_75t_L g3578 ( 
.A1(n_3497),
.A2(n_3189),
.B(n_3246),
.C(n_3227),
.Y(n_3578)
);

OAI21x1_ASAP7_75t_L g3579 ( 
.A1(n_3400),
.A2(n_3271),
.B(n_3239),
.Y(n_3579)
);

NOR2xp33_ASAP7_75t_L g3580 ( 
.A(n_3530),
.B(n_3180),
.Y(n_3580)
);

OAI21x1_ASAP7_75t_L g3581 ( 
.A1(n_3392),
.A2(n_3370),
.B(n_3208),
.Y(n_3581)
);

AND2x4_ASAP7_75t_L g3582 ( 
.A(n_3468),
.B(n_3360),
.Y(n_3582)
);

AOI21xp5_ASAP7_75t_L g3583 ( 
.A1(n_3444),
.A2(n_3234),
.B(n_3211),
.Y(n_3583)
);

CKINVDCx20_ASAP7_75t_R g3584 ( 
.A(n_3414),
.Y(n_3584)
);

INVx2_ASAP7_75t_L g3585 ( 
.A(n_3417),
.Y(n_3585)
);

INVx1_ASAP7_75t_L g3586 ( 
.A(n_3462),
.Y(n_3586)
);

OAI21x1_ASAP7_75t_L g3587 ( 
.A1(n_3421),
.A2(n_3188),
.B(n_3285),
.Y(n_3587)
);

O2A1O1Ixp33_ASAP7_75t_SL g3588 ( 
.A1(n_3424),
.A2(n_3338),
.B(n_3248),
.C(n_3284),
.Y(n_3588)
);

AOI21x1_ASAP7_75t_L g3589 ( 
.A1(n_3497),
.A2(n_3267),
.B(n_3191),
.Y(n_3589)
);

OAI21x1_ASAP7_75t_L g3590 ( 
.A1(n_3421),
.A2(n_3202),
.B(n_3267),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3449),
.Y(n_3591)
);

BUFx3_ASAP7_75t_L g3592 ( 
.A(n_3410),
.Y(n_3592)
);

BUFx3_ASAP7_75t_L g3593 ( 
.A(n_3378),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3504),
.Y(n_3594)
);

AOI221xp5_ASAP7_75t_L g3595 ( 
.A1(n_3443),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.C(n_100),
.Y(n_3595)
);

OAI21x1_ASAP7_75t_L g3596 ( 
.A1(n_3387),
.A2(n_3454),
.B(n_3397),
.Y(n_3596)
);

NAND2xp5_ASAP7_75t_L g3597 ( 
.A(n_3437),
.B(n_3229),
.Y(n_3597)
);

OAI21x1_ASAP7_75t_L g3598 ( 
.A1(n_3382),
.A2(n_3284),
.B(n_3242),
.Y(n_3598)
);

OA21x2_ASAP7_75t_L g3599 ( 
.A1(n_3477),
.A2(n_3191),
.B(n_3180),
.Y(n_3599)
);

A2O1A1Ixp33_ASAP7_75t_L g3600 ( 
.A1(n_3482),
.A2(n_3332),
.B(n_3242),
.C(n_3278),
.Y(n_3600)
);

OAI21x1_ASAP7_75t_L g3601 ( 
.A1(n_3382),
.A2(n_3242),
.B(n_3229),
.Y(n_3601)
);

AND2x4_ASAP7_75t_L g3602 ( 
.A(n_3468),
.B(n_3278),
.Y(n_3602)
);

OR2x6_ASAP7_75t_L g3603 ( 
.A(n_3399),
.B(n_3278),
.Y(n_3603)
);

OA21x2_ASAP7_75t_L g3604 ( 
.A1(n_3477),
.A2(n_3324),
.B(n_3302),
.Y(n_3604)
);

AO21x2_ASAP7_75t_L g3605 ( 
.A1(n_3411),
.A2(n_3324),
.B(n_3302),
.Y(n_3605)
);

OAI21x1_ASAP7_75t_L g3606 ( 
.A1(n_3397),
.A2(n_3324),
.B(n_3302),
.Y(n_3606)
);

INVx1_ASAP7_75t_SL g3607 ( 
.A(n_3459),
.Y(n_3607)
);

NAND2x1p5_ASAP7_75t_L g3608 ( 
.A(n_3409),
.B(n_3357),
.Y(n_3608)
);

OAI21x1_ASAP7_75t_L g3609 ( 
.A1(n_3523),
.A2(n_3357),
.B(n_96),
.Y(n_3609)
);

INVx3_ASAP7_75t_L g3610 ( 
.A(n_3412),
.Y(n_3610)
);

NOR2xp33_ASAP7_75t_L g3611 ( 
.A(n_3498),
.B(n_3357),
.Y(n_3611)
);

AOI21xp5_ASAP7_75t_L g3612 ( 
.A1(n_3420),
.A2(n_100),
.B(n_102),
.Y(n_3612)
);

INVxp67_ASAP7_75t_L g3613 ( 
.A(n_3431),
.Y(n_3613)
);

OAI22xp5_ASAP7_75t_L g3614 ( 
.A1(n_3501),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_3614)
);

INVx1_ASAP7_75t_L g3615 ( 
.A(n_3475),
.Y(n_3615)
);

INVx3_ASAP7_75t_L g3616 ( 
.A(n_3412),
.Y(n_3616)
);

INVx4_ASAP7_75t_L g3617 ( 
.A(n_3407),
.Y(n_3617)
);

CKINVDCx20_ASAP7_75t_R g3618 ( 
.A(n_3455),
.Y(n_3618)
);

HB1xp67_ASAP7_75t_L g3619 ( 
.A(n_3535),
.Y(n_3619)
);

AO21x2_ASAP7_75t_L g3620 ( 
.A1(n_3487),
.A2(n_103),
.B(n_105),
.Y(n_3620)
);

OA21x2_ASAP7_75t_L g3621 ( 
.A1(n_3487),
.A2(n_105),
.B(n_106),
.Y(n_3621)
);

OAI21x1_ASAP7_75t_L g3622 ( 
.A1(n_3523),
.A2(n_107),
.B(n_108),
.Y(n_3622)
);

AND2x2_ASAP7_75t_L g3623 ( 
.A(n_3413),
.B(n_109),
.Y(n_3623)
);

OAI21x1_ASAP7_75t_SL g3624 ( 
.A1(n_3456),
.A2(n_109),
.B(n_110),
.Y(n_3624)
);

OAI22xp5_ASAP7_75t_L g3625 ( 
.A1(n_3390),
.A2(n_3469),
.B1(n_3483),
.B2(n_3511),
.Y(n_3625)
);

NAND2xp33_ASAP7_75t_L g3626 ( 
.A(n_3522),
.B(n_111),
.Y(n_3626)
);

BUFx3_ASAP7_75t_L g3627 ( 
.A(n_3460),
.Y(n_3627)
);

BUFx2_ASAP7_75t_SL g3628 ( 
.A(n_3472),
.Y(n_3628)
);

CKINVDCx20_ASAP7_75t_R g3629 ( 
.A(n_3473),
.Y(n_3629)
);

OAI21x1_ASAP7_75t_L g3630 ( 
.A1(n_3384),
.A2(n_111),
.B(n_112),
.Y(n_3630)
);

OAI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_3503),
.A2(n_112),
.B(n_113),
.Y(n_3631)
);

OAI21x1_ASAP7_75t_L g3632 ( 
.A1(n_3383),
.A2(n_113),
.B(n_114),
.Y(n_3632)
);

INVx1_ASAP7_75t_L g3633 ( 
.A(n_3481),
.Y(n_3633)
);

NAND2xp5_ASAP7_75t_L g3634 ( 
.A(n_3373),
.B(n_114),
.Y(n_3634)
);

NOR2xp33_ASAP7_75t_L g3635 ( 
.A(n_3539),
.B(n_115),
.Y(n_3635)
);

OR2x2_ASAP7_75t_L g3636 ( 
.A(n_3405),
.B(n_117),
.Y(n_3636)
);

OAI21xp5_ASAP7_75t_L g3637 ( 
.A1(n_3520),
.A2(n_118),
.B(n_119),
.Y(n_3637)
);

INVx3_ASAP7_75t_L g3638 ( 
.A(n_3436),
.Y(n_3638)
);

OAI222xp33_ASAP7_75t_L g3639 ( 
.A1(n_3390),
.A2(n_118),
.B1(n_120),
.B2(n_121),
.C1(n_122),
.C2(n_123),
.Y(n_3639)
);

OAI21x1_ASAP7_75t_L g3640 ( 
.A1(n_3492),
.A2(n_120),
.B(n_123),
.Y(n_3640)
);

BUFx6f_ASAP7_75t_L g3641 ( 
.A(n_3401),
.Y(n_3641)
);

INVx4_ASAP7_75t_L g3642 ( 
.A(n_3386),
.Y(n_3642)
);

INVx1_ASAP7_75t_L g3643 ( 
.A(n_3448),
.Y(n_3643)
);

OAI21x1_ASAP7_75t_L g3644 ( 
.A1(n_3492),
.A2(n_124),
.B(n_125),
.Y(n_3644)
);

INVx2_ASAP7_75t_L g3645 ( 
.A(n_3507),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3461),
.Y(n_3646)
);

NAND3xp33_ASAP7_75t_SL g3647 ( 
.A(n_3402),
.B(n_125),
.C(n_126),
.Y(n_3647)
);

INVx1_ASAP7_75t_L g3648 ( 
.A(n_3389),
.Y(n_3648)
);

OAI21x1_ASAP7_75t_L g3649 ( 
.A1(n_3436),
.A2(n_127),
.B(n_128),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3420),
.A2(n_128),
.B(n_129),
.Y(n_3650)
);

INVx1_ASAP7_75t_L g3651 ( 
.A(n_3396),
.Y(n_3651)
);

INVx1_ASAP7_75t_L g3652 ( 
.A(n_3429),
.Y(n_3652)
);

NAND2xp5_ASAP7_75t_L g3653 ( 
.A(n_3432),
.B(n_129),
.Y(n_3653)
);

OA21x2_ASAP7_75t_L g3654 ( 
.A1(n_3533),
.A2(n_3418),
.B(n_3509),
.Y(n_3654)
);

AO31x2_ASAP7_75t_L g3655 ( 
.A1(n_3489),
.A2(n_3385),
.A3(n_3478),
.B(n_3465),
.Y(n_3655)
);

AND2x4_ASAP7_75t_L g3656 ( 
.A(n_3514),
.B(n_130),
.Y(n_3656)
);

INVx2_ASAP7_75t_L g3657 ( 
.A(n_3524),
.Y(n_3657)
);

O2A1O1Ixp33_ASAP7_75t_L g3658 ( 
.A1(n_3391),
.A2(n_130),
.B(n_131),
.C(n_132),
.Y(n_3658)
);

INVx1_ASAP7_75t_L g3659 ( 
.A(n_3466),
.Y(n_3659)
);

OAI21x1_ASAP7_75t_L g3660 ( 
.A1(n_3445),
.A2(n_132),
.B(n_133),
.Y(n_3660)
);

INVx1_ASAP7_75t_L g3661 ( 
.A(n_3381),
.Y(n_3661)
);

AOI21xp5_ASAP7_75t_L g3662 ( 
.A1(n_3385),
.A2(n_133),
.B(n_134),
.Y(n_3662)
);

OAI21x1_ASAP7_75t_L g3663 ( 
.A1(n_3457),
.A2(n_3426),
.B(n_3529),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3493),
.Y(n_3664)
);

NAND2x1p5_ASAP7_75t_L g3665 ( 
.A(n_3409),
.B(n_258),
.Y(n_3665)
);

OAI22xp5_ASAP7_75t_SL g3666 ( 
.A1(n_3526),
.A2(n_136),
.B1(n_137),
.B2(n_138),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3467),
.B(n_137),
.Y(n_3667)
);

INVx1_ASAP7_75t_SL g3668 ( 
.A(n_3485),
.Y(n_3668)
);

NAND2xp5_ASAP7_75t_L g3669 ( 
.A(n_3521),
.B(n_138),
.Y(n_3669)
);

INVxp67_ASAP7_75t_L g3670 ( 
.A(n_3452),
.Y(n_3670)
);

INVx2_ASAP7_75t_L g3671 ( 
.A(n_3604),
.Y(n_3671)
);

HB1xp67_ASAP7_75t_L g3672 ( 
.A(n_3619),
.Y(n_3672)
);

INVx5_ASAP7_75t_L g3673 ( 
.A(n_3642),
.Y(n_3673)
);

INVx2_ASAP7_75t_L g3674 ( 
.A(n_3604),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3567),
.B(n_3491),
.Y(n_3675)
);

OAI22xp5_ASAP7_75t_L g3676 ( 
.A1(n_3541),
.A2(n_3375),
.B1(n_3438),
.B2(n_3408),
.Y(n_3676)
);

INVx6_ASAP7_75t_L g3677 ( 
.A(n_3642),
.Y(n_3677)
);

NOR2xp33_ASAP7_75t_L g3678 ( 
.A(n_3617),
.B(n_3518),
.Y(n_3678)
);

AOI21x1_ASAP7_75t_L g3679 ( 
.A1(n_3669),
.A2(n_3440),
.B(n_3451),
.Y(n_3679)
);

AO21x1_ASAP7_75t_L g3680 ( 
.A1(n_3612),
.A2(n_3650),
.B(n_3614),
.Y(n_3680)
);

AOI22xp33_ASAP7_75t_SL g3681 ( 
.A1(n_3560),
.A2(n_3536),
.B1(n_3453),
.B2(n_3515),
.Y(n_3681)
);

OR2x2_ASAP7_75t_L g3682 ( 
.A(n_3569),
.B(n_3380),
.Y(n_3682)
);

INVx3_ASAP7_75t_L g3683 ( 
.A(n_3582),
.Y(n_3683)
);

AOI22xp33_ASAP7_75t_L g3684 ( 
.A1(n_3647),
.A2(n_3486),
.B1(n_3488),
.B2(n_3470),
.Y(n_3684)
);

NAND2x1p5_ASAP7_75t_L g3685 ( 
.A(n_3570),
.B(n_3433),
.Y(n_3685)
);

OAI21x1_ASAP7_75t_SL g3686 ( 
.A1(n_3612),
.A2(n_3415),
.B(n_3446),
.Y(n_3686)
);

INVx2_ASAP7_75t_L g3687 ( 
.A(n_3605),
.Y(n_3687)
);

INVx2_ASAP7_75t_L g3688 ( 
.A(n_3599),
.Y(n_3688)
);

INVx3_ASAP7_75t_L g3689 ( 
.A(n_3582),
.Y(n_3689)
);

INVx2_ASAP7_75t_L g3690 ( 
.A(n_3599),
.Y(n_3690)
);

BUFx2_ASAP7_75t_R g3691 ( 
.A(n_3628),
.Y(n_3691)
);

AOI22xp5_ASAP7_75t_L g3692 ( 
.A1(n_3625),
.A2(n_3391),
.B1(n_3486),
.B2(n_3531),
.Y(n_3692)
);

INVx1_ASAP7_75t_L g3693 ( 
.A(n_3543),
.Y(n_3693)
);

BUFx4f_ASAP7_75t_SL g3694 ( 
.A(n_3618),
.Y(n_3694)
);

INVx1_ASAP7_75t_L g3695 ( 
.A(n_3544),
.Y(n_3695)
);

INVx2_ASAP7_75t_L g3696 ( 
.A(n_3550),
.Y(n_3696)
);

AOI21x1_ASAP7_75t_L g3697 ( 
.A1(n_3669),
.A2(n_3537),
.B(n_3458),
.Y(n_3697)
);

AOI22xp33_ASAP7_75t_L g3698 ( 
.A1(n_3625),
.A2(n_3538),
.B1(n_3528),
.B2(n_3458),
.Y(n_3698)
);

BUFx2_ASAP7_75t_L g3699 ( 
.A(n_3617),
.Y(n_3699)
);

AOI21x1_ASAP7_75t_L g3700 ( 
.A1(n_3653),
.A2(n_3537),
.B(n_3479),
.Y(n_3700)
);

INVx6_ASAP7_75t_L g3701 ( 
.A(n_3592),
.Y(n_3701)
);

AO21x1_ASAP7_75t_L g3702 ( 
.A1(n_3650),
.A2(n_3427),
.B(n_3398),
.Y(n_3702)
);

BUFx12f_ASAP7_75t_L g3703 ( 
.A(n_3577),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3556),
.Y(n_3704)
);

INVx2_ASAP7_75t_L g3705 ( 
.A(n_3552),
.Y(n_3705)
);

AOI22xp33_ASAP7_75t_L g3706 ( 
.A1(n_3662),
.A2(n_3525),
.B1(n_3531),
.B2(n_3519),
.Y(n_3706)
);

HB1xp67_ASAP7_75t_L g3707 ( 
.A(n_3554),
.Y(n_3707)
);

AND2x2_ASAP7_75t_L g3708 ( 
.A(n_3602),
.B(n_3512),
.Y(n_3708)
);

BUFx10_ASAP7_75t_L g3709 ( 
.A(n_3656),
.Y(n_3709)
);

INVx1_ASAP7_75t_L g3710 ( 
.A(n_3572),
.Y(n_3710)
);

BUFx3_ASAP7_75t_L g3711 ( 
.A(n_3629),
.Y(n_3711)
);

AND2x4_ASAP7_75t_L g3712 ( 
.A(n_3655),
.B(n_3529),
.Y(n_3712)
);

CKINVDCx11_ASAP7_75t_R g3713 ( 
.A(n_3584),
.Y(n_3713)
);

INVx1_ASAP7_75t_L g3714 ( 
.A(n_3574),
.Y(n_3714)
);

AND2x2_ASAP7_75t_L g3715 ( 
.A(n_3602),
.B(n_3484),
.Y(n_3715)
);

INVx1_ASAP7_75t_L g3716 ( 
.A(n_3576),
.Y(n_3716)
);

OAI21x1_ASAP7_75t_L g3717 ( 
.A1(n_3663),
.A2(n_3395),
.B(n_3502),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3591),
.Y(n_3718)
);

AOI22xp33_ASAP7_75t_SL g3719 ( 
.A1(n_3666),
.A2(n_3398),
.B1(n_3513),
.B2(n_3433),
.Y(n_3719)
);

OAI22xp5_ASAP7_75t_L g3720 ( 
.A1(n_3541),
.A2(n_3428),
.B1(n_3433),
.B2(n_3513),
.Y(n_3720)
);

OA21x2_ASAP7_75t_L g3721 ( 
.A1(n_3596),
.A2(n_3471),
.B(n_3495),
.Y(n_3721)
);

AOI22xp33_ASAP7_75t_L g3722 ( 
.A1(n_3662),
.A2(n_3422),
.B1(n_3494),
.B2(n_3500),
.Y(n_3722)
);

OAI22xp5_ASAP7_75t_L g3723 ( 
.A1(n_3666),
.A2(n_3513),
.B1(n_3406),
.B2(n_3399),
.Y(n_3723)
);

AOI22xp33_ASAP7_75t_L g3724 ( 
.A1(n_3631),
.A2(n_3399),
.B1(n_3406),
.B2(n_3496),
.Y(n_3724)
);

NAND2x1p5_ASAP7_75t_L g3725 ( 
.A(n_3570),
.B(n_3465),
.Y(n_3725)
);

INVx2_ASAP7_75t_SL g3726 ( 
.A(n_3593),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_3637),
.A2(n_3406),
.B1(n_3478),
.B2(n_3401),
.Y(n_3727)
);

INVx2_ASAP7_75t_L g3728 ( 
.A(n_3610),
.Y(n_3728)
);

BUFx2_ASAP7_75t_L g3729 ( 
.A(n_3655),
.Y(n_3729)
);

INVx1_ASAP7_75t_L g3730 ( 
.A(n_3585),
.Y(n_3730)
);

AND2x2_ASAP7_75t_L g3731 ( 
.A(n_3551),
.B(n_3386),
.Y(n_3731)
);

INVx1_ASAP7_75t_L g3732 ( 
.A(n_3586),
.Y(n_3732)
);

AOI22xp33_ASAP7_75t_L g3733 ( 
.A1(n_3631),
.A2(n_3532),
.B1(n_3534),
.B2(n_3527),
.Y(n_3733)
);

INVx1_ASAP7_75t_SL g3734 ( 
.A(n_3668),
.Y(n_3734)
);

OAI22xp5_ASAP7_75t_L g3735 ( 
.A1(n_3637),
.A2(n_3516),
.B1(n_3490),
.B2(n_3480),
.Y(n_3735)
);

INVx5_ASAP7_75t_L g3736 ( 
.A(n_3547),
.Y(n_3736)
);

AOI22xp33_ASAP7_75t_SL g3737 ( 
.A1(n_3626),
.A2(n_3516),
.B1(n_3490),
.B2(n_3480),
.Y(n_3737)
);

BUFx3_ASAP7_75t_L g3738 ( 
.A(n_3627),
.Y(n_3738)
);

HB1xp67_ASAP7_75t_L g3739 ( 
.A(n_3607),
.Y(n_3739)
);

AOI22xp33_ASAP7_75t_L g3740 ( 
.A1(n_3540),
.A2(n_3516),
.B1(n_3490),
.B2(n_3480),
.Y(n_3740)
);

INVx1_ASAP7_75t_L g3741 ( 
.A(n_3664),
.Y(n_3741)
);

INVx2_ASAP7_75t_L g3742 ( 
.A(n_3610),
.Y(n_3742)
);

INVx1_ASAP7_75t_L g3743 ( 
.A(n_3615),
.Y(n_3743)
);

OR2x2_ASAP7_75t_L g3744 ( 
.A(n_3613),
.B(n_3419),
.Y(n_3744)
);

AOI22xp5_ASAP7_75t_L g3745 ( 
.A1(n_3595),
.A2(n_3476),
.B1(n_3439),
.B2(n_3419),
.Y(n_3745)
);

AO22x1_ASAP7_75t_L g3746 ( 
.A1(n_3545),
.A2(n_3476),
.B1(n_3439),
.B2(n_3419),
.Y(n_3746)
);

INVx1_ASAP7_75t_L g3747 ( 
.A(n_3633),
.Y(n_3747)
);

INVx2_ASAP7_75t_L g3748 ( 
.A(n_3616),
.Y(n_3748)
);

INVx2_ASAP7_75t_SL g3749 ( 
.A(n_3555),
.Y(n_3749)
);

AOI22xp33_ASAP7_75t_L g3750 ( 
.A1(n_3595),
.A2(n_3476),
.B1(n_3439),
.B2(n_142),
.Y(n_3750)
);

AND2x4_ASAP7_75t_L g3751 ( 
.A(n_3655),
.B(n_140),
.Y(n_3751)
);

OAI22xp33_ASAP7_75t_L g3752 ( 
.A1(n_3547),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_3752)
);

BUFx2_ASAP7_75t_R g3753 ( 
.A(n_3620),
.Y(n_3753)
);

INVx8_ASAP7_75t_L g3754 ( 
.A(n_3656),
.Y(n_3754)
);

OR2x2_ASAP7_75t_L g3755 ( 
.A(n_3670),
.B(n_141),
.Y(n_3755)
);

OAI22xp33_ASAP7_75t_L g3756 ( 
.A1(n_3547),
.A2(n_3603),
.B1(n_3607),
.B2(n_3614),
.Y(n_3756)
);

BUFx6f_ASAP7_75t_L g3757 ( 
.A(n_3641),
.Y(n_3757)
);

INVx1_ASAP7_75t_L g3758 ( 
.A(n_3643),
.Y(n_3758)
);

OR2x6_ASAP7_75t_L g3759 ( 
.A(n_3565),
.B(n_143),
.Y(n_3759)
);

AND2x4_ASAP7_75t_L g3760 ( 
.A(n_3603),
.B(n_144),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3616),
.Y(n_3761)
);

OA21x2_ASAP7_75t_L g3762 ( 
.A1(n_3601),
.A2(n_145),
.B(n_146),
.Y(n_3762)
);

INVx3_ASAP7_75t_L g3763 ( 
.A(n_3638),
.Y(n_3763)
);

INVx1_ASAP7_75t_L g3764 ( 
.A(n_3646),
.Y(n_3764)
);

INVx1_ASAP7_75t_L g3765 ( 
.A(n_3648),
.Y(n_3765)
);

BUFx2_ASAP7_75t_L g3766 ( 
.A(n_3603),
.Y(n_3766)
);

OAI22xp33_ASAP7_75t_L g3767 ( 
.A1(n_3654),
.A2(n_145),
.B1(n_146),
.B2(n_147),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3638),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3651),
.Y(n_3769)
);

AND2x2_ASAP7_75t_L g3770 ( 
.A(n_3561),
.B(n_3594),
.Y(n_3770)
);

NAND2x1p5_ASAP7_75t_L g3771 ( 
.A(n_3654),
.B(n_3598),
.Y(n_3771)
);

OAI22xp5_ASAP7_75t_L g3772 ( 
.A1(n_3548),
.A2(n_148),
.B1(n_150),
.B2(n_151),
.Y(n_3772)
);

BUFx10_ASAP7_75t_L g3773 ( 
.A(n_3611),
.Y(n_3773)
);

INVxp67_ASAP7_75t_L g3774 ( 
.A(n_3621),
.Y(n_3774)
);

OAI22xp33_ASAP7_75t_R g3775 ( 
.A1(n_3635),
.A2(n_148),
.B1(n_152),
.B2(n_154),
.Y(n_3775)
);

AOI22xp33_ASAP7_75t_L g3776 ( 
.A1(n_3624),
.A2(n_154),
.B1(n_155),
.B2(n_157),
.Y(n_3776)
);

CKINVDCx11_ASAP7_75t_R g3777 ( 
.A(n_3641),
.Y(n_3777)
);

AOI22xp33_ASAP7_75t_L g3778 ( 
.A1(n_3563),
.A2(n_155),
.B1(n_158),
.B2(n_159),
.Y(n_3778)
);

AOI222xp33_ASAP7_75t_L g3779 ( 
.A1(n_3639),
.A2(n_158),
.B1(n_159),
.B2(n_160),
.C1(n_161),
.C2(n_162),
.Y(n_3779)
);

INVx1_ASAP7_75t_L g3780 ( 
.A(n_3652),
.Y(n_3780)
);

INVx1_ASAP7_75t_L g3781 ( 
.A(n_3659),
.Y(n_3781)
);

INVx2_ASAP7_75t_L g3782 ( 
.A(n_3645),
.Y(n_3782)
);

AOI22xp33_ASAP7_75t_L g3783 ( 
.A1(n_3563),
.A2(n_160),
.B1(n_161),
.B2(n_164),
.Y(n_3783)
);

OAI22xp5_ASAP7_75t_L g3784 ( 
.A1(n_3658),
.A2(n_166),
.B1(n_167),
.B2(n_168),
.Y(n_3784)
);

NAND2x1p5_ASAP7_75t_L g3785 ( 
.A(n_3606),
.B(n_3559),
.Y(n_3785)
);

OAI22xp5_ASAP7_75t_L g3786 ( 
.A1(n_3621),
.A2(n_166),
.B1(n_169),
.B2(n_170),
.Y(n_3786)
);

INVx2_ASAP7_75t_L g3787 ( 
.A(n_3657),
.Y(n_3787)
);

NOR2xp33_ASAP7_75t_L g3788 ( 
.A(n_3636),
.B(n_169),
.Y(n_3788)
);

INVx1_ASAP7_75t_L g3789 ( 
.A(n_3661),
.Y(n_3789)
);

INVx1_ASAP7_75t_L g3790 ( 
.A(n_3575),
.Y(n_3790)
);

HB1xp67_ASAP7_75t_L g3791 ( 
.A(n_3575),
.Y(n_3791)
);

INVx2_ASAP7_75t_L g3792 ( 
.A(n_3641),
.Y(n_3792)
);

INVx1_ASAP7_75t_L g3793 ( 
.A(n_3741),
.Y(n_3793)
);

INVx2_ASAP7_75t_SL g3794 ( 
.A(n_3673),
.Y(n_3794)
);

CKINVDCx14_ASAP7_75t_R g3795 ( 
.A(n_3713),
.Y(n_3795)
);

INVx1_ASAP7_75t_L g3796 ( 
.A(n_3743),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3747),
.Y(n_3797)
);

INVx1_ASAP7_75t_L g3798 ( 
.A(n_3693),
.Y(n_3798)
);

INVx1_ASAP7_75t_L g3799 ( 
.A(n_3695),
.Y(n_3799)
);

AND2x2_ASAP7_75t_L g3800 ( 
.A(n_3683),
.B(n_3568),
.Y(n_3800)
);

INVx1_ASAP7_75t_L g3801 ( 
.A(n_3704),
.Y(n_3801)
);

INVx2_ASAP7_75t_L g3802 ( 
.A(n_3671),
.Y(n_3802)
);

BUFx3_ASAP7_75t_L g3803 ( 
.A(n_3701),
.Y(n_3803)
);

INVx3_ASAP7_75t_L g3804 ( 
.A(n_3673),
.Y(n_3804)
);

OAI22xp5_ASAP7_75t_L g3805 ( 
.A1(n_3719),
.A2(n_3600),
.B1(n_3589),
.B2(n_3558),
.Y(n_3805)
);

OAI21x1_ASAP7_75t_L g3806 ( 
.A1(n_3685),
.A2(n_3546),
.B(n_3571),
.Y(n_3806)
);

INVx1_ASAP7_75t_L g3807 ( 
.A(n_3710),
.Y(n_3807)
);

OAI21x1_ASAP7_75t_L g3808 ( 
.A1(n_3685),
.A2(n_3566),
.B(n_3558),
.Y(n_3808)
);

AO21x2_ASAP7_75t_L g3809 ( 
.A1(n_3767),
.A2(n_3774),
.B(n_3756),
.Y(n_3809)
);

INVx1_ASAP7_75t_L g3810 ( 
.A(n_3714),
.Y(n_3810)
);

BUFx2_ASAP7_75t_L g3811 ( 
.A(n_3699),
.Y(n_3811)
);

INVx1_ASAP7_75t_L g3812 ( 
.A(n_3716),
.Y(n_3812)
);

INVx2_ASAP7_75t_L g3813 ( 
.A(n_3674),
.Y(n_3813)
);

INVx1_ASAP7_75t_L g3814 ( 
.A(n_3718),
.Y(n_3814)
);

INVxp67_ASAP7_75t_L g3815 ( 
.A(n_3753),
.Y(n_3815)
);

OAI21xp5_ASAP7_75t_L g3816 ( 
.A1(n_3772),
.A2(n_3542),
.B(n_3630),
.Y(n_3816)
);

INVx1_ASAP7_75t_L g3817 ( 
.A(n_3732),
.Y(n_3817)
);

INVx1_ASAP7_75t_L g3818 ( 
.A(n_3758),
.Y(n_3818)
);

INVx1_ASAP7_75t_L g3819 ( 
.A(n_3764),
.Y(n_3819)
);

INVx2_ASAP7_75t_L g3820 ( 
.A(n_3688),
.Y(n_3820)
);

INVx2_ASAP7_75t_L g3821 ( 
.A(n_3690),
.Y(n_3821)
);

INVx2_ASAP7_75t_L g3822 ( 
.A(n_3687),
.Y(n_3822)
);

INVx1_ASAP7_75t_L g3823 ( 
.A(n_3765),
.Y(n_3823)
);

INVx8_ASAP7_75t_L g3824 ( 
.A(n_3673),
.Y(n_3824)
);

HB1xp67_ASAP7_75t_L g3825 ( 
.A(n_3739),
.Y(n_3825)
);

CKINVDCx12_ASAP7_75t_R g3826 ( 
.A(n_3759),
.Y(n_3826)
);

INVx2_ASAP7_75t_L g3827 ( 
.A(n_3751),
.Y(n_3827)
);

INVx1_ASAP7_75t_L g3828 ( 
.A(n_3769),
.Y(n_3828)
);

AO21x2_ASAP7_75t_L g3829 ( 
.A1(n_3774),
.A2(n_3653),
.B(n_3620),
.Y(n_3829)
);

OAI22xp5_ASAP7_75t_L g3830 ( 
.A1(n_3719),
.A2(n_3634),
.B1(n_3562),
.B2(n_3549),
.Y(n_3830)
);

INVx1_ASAP7_75t_L g3831 ( 
.A(n_3780),
.Y(n_3831)
);

INVx1_ASAP7_75t_L g3832 ( 
.A(n_3781),
.Y(n_3832)
);

INVx2_ASAP7_75t_L g3833 ( 
.A(n_3751),
.Y(n_3833)
);

INVx1_ASAP7_75t_L g3834 ( 
.A(n_3789),
.Y(n_3834)
);

INVx2_ASAP7_75t_L g3835 ( 
.A(n_3725),
.Y(n_3835)
);

INVx1_ASAP7_75t_L g3836 ( 
.A(n_3730),
.Y(n_3836)
);

OR2x6_ASAP7_75t_L g3837 ( 
.A(n_3680),
.B(n_3665),
.Y(n_3837)
);

INVxp67_ASAP7_75t_L g3838 ( 
.A(n_3753),
.Y(n_3838)
);

INVx1_ASAP7_75t_L g3839 ( 
.A(n_3672),
.Y(n_3839)
);

INVx1_ASAP7_75t_L g3840 ( 
.A(n_3791),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3734),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3734),
.Y(n_3842)
);

INVx3_ASAP7_75t_L g3843 ( 
.A(n_3677),
.Y(n_3843)
);

INVx2_ASAP7_75t_L g3844 ( 
.A(n_3725),
.Y(n_3844)
);

INVx1_ASAP7_75t_L g3845 ( 
.A(n_3790),
.Y(n_3845)
);

INVx1_ASAP7_75t_L g3846 ( 
.A(n_3787),
.Y(n_3846)
);

INVx1_ASAP7_75t_L g3847 ( 
.A(n_3782),
.Y(n_3847)
);

INVx2_ASAP7_75t_L g3848 ( 
.A(n_3762),
.Y(n_3848)
);

OR2x2_ASAP7_75t_L g3849 ( 
.A(n_3707),
.B(n_3549),
.Y(n_3849)
);

INVx2_ASAP7_75t_L g3850 ( 
.A(n_3762),
.Y(n_3850)
);

INVx3_ASAP7_75t_L g3851 ( 
.A(n_3677),
.Y(n_3851)
);

INVx2_ASAP7_75t_L g3852 ( 
.A(n_3729),
.Y(n_3852)
);

INVx2_ASAP7_75t_L g3853 ( 
.A(n_3697),
.Y(n_3853)
);

AND2x2_ASAP7_75t_L g3854 ( 
.A(n_3683),
.B(n_3568),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3785),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3689),
.B(n_3568),
.Y(n_3856)
);

INVx1_ASAP7_75t_L g3857 ( 
.A(n_3744),
.Y(n_3857)
);

INVx2_ASAP7_75t_L g3858 ( 
.A(n_3785),
.Y(n_3858)
);

INVx3_ASAP7_75t_L g3859 ( 
.A(n_3712),
.Y(n_3859)
);

OA21x2_ASAP7_75t_L g3860 ( 
.A1(n_3702),
.A2(n_3644),
.B(n_3640),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3698),
.B(n_3667),
.Y(n_3861)
);

OA21x2_ASAP7_75t_L g3862 ( 
.A1(n_3717),
.A2(n_3581),
.B(n_3609),
.Y(n_3862)
);

INVx1_ASAP7_75t_L g3863 ( 
.A(n_3682),
.Y(n_3863)
);

INVx1_ASAP7_75t_L g3864 ( 
.A(n_3700),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3755),
.Y(n_3865)
);

INVx1_ASAP7_75t_L g3866 ( 
.A(n_3766),
.Y(n_3866)
);

INVx1_ASAP7_75t_L g3867 ( 
.A(n_3792),
.Y(n_3867)
);

HB1xp67_ASAP7_75t_L g3868 ( 
.A(n_3721),
.Y(n_3868)
);

INVx1_ASAP7_75t_L g3869 ( 
.A(n_3679),
.Y(n_3869)
);

INVx2_ASAP7_75t_L g3870 ( 
.A(n_3712),
.Y(n_3870)
);

INVx1_ASAP7_75t_L g3871 ( 
.A(n_3696),
.Y(n_3871)
);

INVx1_ASAP7_75t_L g3872 ( 
.A(n_3705),
.Y(n_3872)
);

AOI22xp33_ASAP7_75t_L g3873 ( 
.A1(n_3772),
.A2(n_3562),
.B1(n_3632),
.B2(n_3583),
.Y(n_3873)
);

AO21x2_ASAP7_75t_L g3874 ( 
.A1(n_3786),
.A2(n_3634),
.B(n_3557),
.Y(n_3874)
);

INVx1_ASAP7_75t_L g3875 ( 
.A(n_3770),
.Y(n_3875)
);

BUFx3_ASAP7_75t_L g3876 ( 
.A(n_3701),
.Y(n_3876)
);

INVx2_ASAP7_75t_L g3877 ( 
.A(n_3686),
.Y(n_3877)
);

INVx2_ASAP7_75t_L g3878 ( 
.A(n_3728),
.Y(n_3878)
);

AOI21x1_ASAP7_75t_L g3879 ( 
.A1(n_3746),
.A2(n_3623),
.B(n_3557),
.Y(n_3879)
);

NAND2xp5_ASAP7_75t_L g3880 ( 
.A(n_3681),
.B(n_3597),
.Y(n_3880)
);

HB1xp67_ASAP7_75t_L g3881 ( 
.A(n_3736),
.Y(n_3881)
);

INVx1_ASAP7_75t_L g3882 ( 
.A(n_3757),
.Y(n_3882)
);

INVx1_ASAP7_75t_L g3883 ( 
.A(n_3757),
.Y(n_3883)
);

CKINVDCx11_ASAP7_75t_R g3884 ( 
.A(n_3703),
.Y(n_3884)
);

HB1xp67_ASAP7_75t_L g3885 ( 
.A(n_3736),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3742),
.Y(n_3886)
);

HB1xp67_ASAP7_75t_L g3887 ( 
.A(n_3736),
.Y(n_3887)
);

INVx1_ASAP7_75t_L g3888 ( 
.A(n_3757),
.Y(n_3888)
);

CKINVDCx5p33_ASAP7_75t_R g3889 ( 
.A(n_3691),
.Y(n_3889)
);

INVx3_ASAP7_75t_L g3890 ( 
.A(n_3689),
.Y(n_3890)
);

HB1xp67_ASAP7_75t_L g3891 ( 
.A(n_3735),
.Y(n_3891)
);

AO21x2_ASAP7_75t_L g3892 ( 
.A1(n_3786),
.A2(n_3660),
.B(n_3649),
.Y(n_3892)
);

AO31x2_ASAP7_75t_L g3893 ( 
.A1(n_3735),
.A2(n_3597),
.A3(n_3580),
.B(n_3559),
.Y(n_3893)
);

INVx2_ASAP7_75t_L g3894 ( 
.A(n_3748),
.Y(n_3894)
);

BUFx8_ASAP7_75t_SL g3895 ( 
.A(n_3759),
.Y(n_3895)
);

AOI222xp33_ASAP7_75t_L g3896 ( 
.A1(n_3775),
.A2(n_3622),
.B1(n_3573),
.B2(n_3590),
.C1(n_3579),
.C2(n_3587),
.Y(n_3896)
);

INVx2_ASAP7_75t_L g3897 ( 
.A(n_3761),
.Y(n_3897)
);

HB1xp67_ASAP7_75t_L g3898 ( 
.A(n_3727),
.Y(n_3898)
);

INVx2_ASAP7_75t_L g3899 ( 
.A(n_3768),
.Y(n_3899)
);

INVx1_ASAP7_75t_L g3900 ( 
.A(n_3709),
.Y(n_3900)
);

INVx1_ASAP7_75t_L g3901 ( 
.A(n_3708),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3675),
.Y(n_3902)
);

INVx1_ASAP7_75t_L g3903 ( 
.A(n_3763),
.Y(n_3903)
);

BUFx6f_ASAP7_75t_L g3904 ( 
.A(n_3777),
.Y(n_3904)
);

BUFx6f_ASAP7_75t_L g3905 ( 
.A(n_3760),
.Y(n_3905)
);

AOI21xp5_ASAP7_75t_L g3906 ( 
.A1(n_3752),
.A2(n_3588),
.B(n_3578),
.Y(n_3906)
);

AOI22xp33_ASAP7_75t_L g3907 ( 
.A1(n_3681),
.A2(n_3564),
.B1(n_3553),
.B2(n_3608),
.Y(n_3907)
);

AOI222xp33_ASAP7_75t_L g3908 ( 
.A1(n_3816),
.A2(n_3750),
.B1(n_3784),
.B2(n_3783),
.C1(n_3778),
.C2(n_3788),
.Y(n_3908)
);

AOI22xp33_ASAP7_75t_L g3909 ( 
.A1(n_3837),
.A2(n_3676),
.B1(n_3720),
.B2(n_3779),
.Y(n_3909)
);

OAI22xp5_ASAP7_75t_L g3910 ( 
.A1(n_3815),
.A2(n_3745),
.B1(n_3691),
.B2(n_3737),
.Y(n_3910)
);

AOI22xp5_ASAP7_75t_L g3911 ( 
.A1(n_3838),
.A2(n_3830),
.B1(n_3809),
.B2(n_3873),
.Y(n_3911)
);

OAI22xp5_ASAP7_75t_L g3912 ( 
.A1(n_3873),
.A2(n_3745),
.B1(n_3737),
.B2(n_3692),
.Y(n_3912)
);

BUFx2_ASAP7_75t_L g3913 ( 
.A(n_3895),
.Y(n_3913)
);

AOI22xp33_ASAP7_75t_L g3914 ( 
.A1(n_3837),
.A2(n_3676),
.B1(n_3720),
.B2(n_3779),
.Y(n_3914)
);

OAI221xp5_ASAP7_75t_L g3915 ( 
.A1(n_3837),
.A2(n_3907),
.B1(n_3906),
.B2(n_3898),
.C(n_3805),
.Y(n_3915)
);

INVx3_ASAP7_75t_L g3916 ( 
.A(n_3904),
.Y(n_3916)
);

AOI21xp5_ASAP7_75t_L g3917 ( 
.A1(n_3837),
.A2(n_3784),
.B(n_3723),
.Y(n_3917)
);

OAI22xp5_ASAP7_75t_L g3918 ( 
.A1(n_3889),
.A2(n_3692),
.B1(n_3684),
.B2(n_3733),
.Y(n_3918)
);

AOI22xp33_ASAP7_75t_L g3919 ( 
.A1(n_3809),
.A2(n_3727),
.B1(n_3723),
.B2(n_3724),
.Y(n_3919)
);

BUFx4f_ASAP7_75t_SL g3920 ( 
.A(n_3904),
.Y(n_3920)
);

AOI22xp33_ASAP7_75t_SL g3921 ( 
.A1(n_3809),
.A2(n_3754),
.B1(n_3760),
.B2(n_3771),
.Y(n_3921)
);

OAI22xp5_ASAP7_75t_L g3922 ( 
.A1(n_3889),
.A2(n_3722),
.B1(n_3706),
.B2(n_3776),
.Y(n_3922)
);

AOI211xp5_ASAP7_75t_L g3923 ( 
.A1(n_3891),
.A2(n_3678),
.B(n_3726),
.C(n_3738),
.Y(n_3923)
);

INVx2_ASAP7_75t_L g3924 ( 
.A(n_3803),
.Y(n_3924)
);

INVx2_ASAP7_75t_SL g3925 ( 
.A(n_3904),
.Y(n_3925)
);

INVx1_ASAP7_75t_L g3926 ( 
.A(n_3793),
.Y(n_3926)
);

OAI22xp5_ASAP7_75t_SL g3927 ( 
.A1(n_3826),
.A2(n_3694),
.B1(n_3771),
.B2(n_3711),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3796),
.Y(n_3928)
);

NAND2xp5_ASAP7_75t_L g3929 ( 
.A(n_3811),
.B(n_3754),
.Y(n_3929)
);

AOI22xp33_ASAP7_75t_L g3930 ( 
.A1(n_3874),
.A2(n_3754),
.B1(n_3773),
.B2(n_3740),
.Y(n_3930)
);

AOI22xp33_ASAP7_75t_L g3931 ( 
.A1(n_3874),
.A2(n_3773),
.B1(n_3715),
.B2(n_3749),
.Y(n_3931)
);

AOI221xp5_ASAP7_75t_L g3932 ( 
.A1(n_3874),
.A2(n_3731),
.B1(n_3763),
.B2(n_173),
.C(n_175),
.Y(n_3932)
);

AOI22xp33_ASAP7_75t_L g3933 ( 
.A1(n_3857),
.A2(n_3860),
.B1(n_3907),
.B2(n_3863),
.Y(n_3933)
);

HB1xp67_ASAP7_75t_L g3934 ( 
.A(n_3825),
.Y(n_3934)
);

AOI22xp33_ASAP7_75t_SL g3935 ( 
.A1(n_3860),
.A2(n_171),
.B1(n_172),
.B2(n_175),
.Y(n_3935)
);

OA21x2_ASAP7_75t_L g3936 ( 
.A1(n_3853),
.A2(n_171),
.B(n_176),
.Y(n_3936)
);

AOI21xp33_ASAP7_75t_L g3937 ( 
.A1(n_3864),
.A2(n_176),
.B(n_177),
.Y(n_3937)
);

AND2x4_ASAP7_75t_L g3938 ( 
.A(n_3794),
.B(n_177),
.Y(n_3938)
);

INVx3_ASAP7_75t_L g3939 ( 
.A(n_3904),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3797),
.Y(n_3940)
);

INVx4_ASAP7_75t_L g3941 ( 
.A(n_3884),
.Y(n_3941)
);

AOI22xp33_ASAP7_75t_L g3942 ( 
.A1(n_3860),
.A2(n_178),
.B1(n_180),
.B2(n_181),
.Y(n_3942)
);

AOI22xp33_ASAP7_75t_L g3943 ( 
.A1(n_3866),
.A2(n_3880),
.B1(n_3901),
.B2(n_3877),
.Y(n_3943)
);

AOI22xp33_ASAP7_75t_SL g3944 ( 
.A1(n_3795),
.A2(n_178),
.B1(n_182),
.B2(n_183),
.Y(n_3944)
);

AOI22xp33_ASAP7_75t_L g3945 ( 
.A1(n_3877),
.A2(n_182),
.B1(n_183),
.B2(n_185),
.Y(n_3945)
);

A2O1A1Ixp33_ASAP7_75t_L g3946 ( 
.A1(n_3795),
.A2(n_3869),
.B(n_3853),
.C(n_3850),
.Y(n_3946)
);

NAND2xp5_ASAP7_75t_L g3947 ( 
.A(n_3865),
.B(n_185),
.Y(n_3947)
);

INVx1_ASAP7_75t_L g3948 ( 
.A(n_3798),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3803),
.Y(n_3949)
);

AOI22xp33_ASAP7_75t_L g3950 ( 
.A1(n_3896),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_3950)
);

INVx1_ASAP7_75t_L g3951 ( 
.A(n_3799),
.Y(n_3951)
);

OAI221xp5_ASAP7_75t_L g3952 ( 
.A1(n_3794),
.A2(n_186),
.B1(n_187),
.B2(n_189),
.C(n_190),
.Y(n_3952)
);

OAI31xp33_ASAP7_75t_L g3953 ( 
.A1(n_3861),
.A2(n_189),
.A3(n_192),
.B(n_195),
.Y(n_3953)
);

OR2x2_ASAP7_75t_L g3954 ( 
.A(n_3841),
.B(n_192),
.Y(n_3954)
);

AOI33xp33_ASAP7_75t_L g3955 ( 
.A1(n_3842),
.A2(n_195),
.A3(n_196),
.B1(n_197),
.B2(n_198),
.B3(n_199),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3801),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3875),
.B(n_196),
.Y(n_3957)
);

OAI22xp33_ASAP7_75t_L g3958 ( 
.A1(n_3879),
.A2(n_198),
.B1(n_201),
.B2(n_203),
.Y(n_3958)
);

OAI221xp5_ASAP7_75t_L g3959 ( 
.A1(n_3881),
.A2(n_203),
.B1(n_204),
.B2(n_207),
.C(n_208),
.Y(n_3959)
);

AOI22xp33_ASAP7_75t_L g3960 ( 
.A1(n_3895),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_3960)
);

AOI22xp33_ASAP7_75t_L g3961 ( 
.A1(n_3892),
.A2(n_213),
.B1(n_214),
.B2(n_215),
.Y(n_3961)
);

INVx3_ASAP7_75t_L g3962 ( 
.A(n_3876),
.Y(n_3962)
);

INVx2_ASAP7_75t_L g3963 ( 
.A(n_3876),
.Y(n_3963)
);

AO21x2_ASAP7_75t_L g3964 ( 
.A1(n_3885),
.A2(n_216),
.B(n_217),
.Y(n_3964)
);

AND2x4_ASAP7_75t_L g3965 ( 
.A(n_3843),
.B(n_3851),
.Y(n_3965)
);

INVx1_ASAP7_75t_L g3966 ( 
.A(n_3807),
.Y(n_3966)
);

OAI221xp5_ASAP7_75t_L g3967 ( 
.A1(n_3887),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.C(n_221),
.Y(n_3967)
);

AND2x2_ASAP7_75t_L g3968 ( 
.A(n_3843),
.B(n_218),
.Y(n_3968)
);

OA21x2_ASAP7_75t_L g3969 ( 
.A1(n_3835),
.A2(n_219),
.B(n_222),
.Y(n_3969)
);

AOI22xp33_ASAP7_75t_L g3970 ( 
.A1(n_3892),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_3970)
);

OAI21xp5_ASAP7_75t_L g3971 ( 
.A1(n_3848),
.A2(n_223),
.B(n_224),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3804),
.Y(n_3972)
);

AOI22xp33_ASAP7_75t_SL g3973 ( 
.A1(n_3868),
.A2(n_225),
.B1(n_227),
.B2(n_228),
.Y(n_3973)
);

NAND2xp5_ASAP7_75t_L g3974 ( 
.A(n_3827),
.B(n_425),
.Y(n_3974)
);

OAI22xp5_ASAP7_75t_L g3975 ( 
.A1(n_3905),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_3975)
);

BUFx2_ASAP7_75t_L g3976 ( 
.A(n_3905),
.Y(n_3976)
);

AOI21xp33_ASAP7_75t_L g3977 ( 
.A1(n_3862),
.A2(n_264),
.B(n_273),
.Y(n_3977)
);

NAND2xp33_ASAP7_75t_L g3978 ( 
.A(n_3905),
.B(n_294),
.Y(n_3978)
);

CKINVDCx14_ASAP7_75t_R g3979 ( 
.A(n_3884),
.Y(n_3979)
);

OAI22xp5_ASAP7_75t_L g3980 ( 
.A1(n_3905),
.A2(n_304),
.B1(n_305),
.B2(n_306),
.Y(n_3980)
);

AND2x2_ASAP7_75t_L g3981 ( 
.A(n_3843),
.B(n_314),
.Y(n_3981)
);

INVx1_ASAP7_75t_L g3982 ( 
.A(n_3810),
.Y(n_3982)
);

INVx2_ASAP7_75t_L g3983 ( 
.A(n_3804),
.Y(n_3983)
);

INVx2_ASAP7_75t_L g3984 ( 
.A(n_3804),
.Y(n_3984)
);

INVx1_ASAP7_75t_L g3985 ( 
.A(n_3812),
.Y(n_3985)
);

AO21x2_ASAP7_75t_L g3986 ( 
.A1(n_3850),
.A2(n_328),
.B(n_330),
.Y(n_3986)
);

BUFx3_ASAP7_75t_L g3987 ( 
.A(n_3851),
.Y(n_3987)
);

AOI222xp33_ASAP7_75t_L g3988 ( 
.A1(n_3839),
.A2(n_3840),
.B1(n_3833),
.B2(n_3827),
.C1(n_3900),
.C2(n_3826),
.Y(n_3988)
);

INVx5_ASAP7_75t_SL g3989 ( 
.A(n_3829),
.Y(n_3989)
);

BUFx2_ASAP7_75t_L g3990 ( 
.A(n_3851),
.Y(n_3990)
);

BUFx8_ASAP7_75t_SL g3991 ( 
.A(n_3882),
.Y(n_3991)
);

BUFx6f_ASAP7_75t_L g3992 ( 
.A(n_3824),
.Y(n_3992)
);

BUFx12f_ASAP7_75t_L g3993 ( 
.A(n_3824),
.Y(n_3993)
);

AND2x2_ASAP7_75t_L g3994 ( 
.A(n_3902),
.B(n_376),
.Y(n_3994)
);

CKINVDCx20_ASAP7_75t_R g3995 ( 
.A(n_3883),
.Y(n_3995)
);

AOI221xp5_ASAP7_75t_L g3996 ( 
.A1(n_3845),
.A2(n_3800),
.B1(n_3856),
.B2(n_3854),
.C(n_3867),
.Y(n_3996)
);

AOI21xp33_ASAP7_75t_L g3997 ( 
.A1(n_3862),
.A2(n_383),
.B(n_384),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_3890),
.Y(n_3998)
);

INVx1_ASAP7_75t_L g3999 ( 
.A(n_3814),
.Y(n_3999)
);

INVx2_ASAP7_75t_L g4000 ( 
.A(n_3890),
.Y(n_4000)
);

INVx1_ASAP7_75t_L g4001 ( 
.A(n_3817),
.Y(n_4001)
);

AOI21x1_ASAP7_75t_L g4002 ( 
.A1(n_3888),
.A2(n_388),
.B(n_389),
.Y(n_4002)
);

AOI22xp33_ASAP7_75t_L g4003 ( 
.A1(n_3800),
.A2(n_3854),
.B1(n_3856),
.B2(n_3847),
.Y(n_4003)
);

INVx4_ASAP7_75t_SL g4004 ( 
.A(n_3893),
.Y(n_4004)
);

BUFx3_ASAP7_75t_L g4005 ( 
.A(n_3890),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3846),
.B(n_421),
.Y(n_4006)
);

AND2x2_ASAP7_75t_L g4007 ( 
.A(n_3878),
.B(n_403),
.Y(n_4007)
);

INVx4_ASAP7_75t_L g4008 ( 
.A(n_3859),
.Y(n_4008)
);

NAND2xp5_ASAP7_75t_L g4009 ( 
.A(n_3911),
.B(n_3878),
.Y(n_4009)
);

INVx1_ASAP7_75t_L g4010 ( 
.A(n_3934),
.Y(n_4010)
);

INVx2_ASAP7_75t_L g4011 ( 
.A(n_4008),
.Y(n_4011)
);

AND2x2_ASAP7_75t_L g4012 ( 
.A(n_3962),
.B(n_3870),
.Y(n_4012)
);

AND2x2_ASAP7_75t_L g4013 ( 
.A(n_3962),
.B(n_3990),
.Y(n_4013)
);

INVx2_ASAP7_75t_L g4014 ( 
.A(n_4008),
.Y(n_4014)
);

AND2x2_ASAP7_75t_L g4015 ( 
.A(n_3965),
.B(n_3870),
.Y(n_4015)
);

NAND2xp5_ASAP7_75t_L g4016 ( 
.A(n_3911),
.B(n_3886),
.Y(n_4016)
);

INVx1_ASAP7_75t_L g4017 ( 
.A(n_3926),
.Y(n_4017)
);

AND2x2_ASAP7_75t_L g4018 ( 
.A(n_3965),
.B(n_3899),
.Y(n_4018)
);

INVx2_ASAP7_75t_L g4019 ( 
.A(n_3998),
.Y(n_4019)
);

OR2x2_ASAP7_75t_L g4020 ( 
.A(n_4003),
.B(n_3849),
.Y(n_4020)
);

AND2x4_ASAP7_75t_SL g4021 ( 
.A(n_3941),
.B(n_3859),
.Y(n_4021)
);

INVx2_ASAP7_75t_L g4022 ( 
.A(n_3998),
.Y(n_4022)
);

INVx1_ASAP7_75t_L g4023 ( 
.A(n_3928),
.Y(n_4023)
);

INVx2_ASAP7_75t_L g4024 ( 
.A(n_3916),
.Y(n_4024)
);

INVx2_ASAP7_75t_SL g4025 ( 
.A(n_3916),
.Y(n_4025)
);

INVx2_ASAP7_75t_L g4026 ( 
.A(n_3939),
.Y(n_4026)
);

INVx1_ASAP7_75t_L g4027 ( 
.A(n_3940),
.Y(n_4027)
);

INVx2_ASAP7_75t_L g4028 ( 
.A(n_3939),
.Y(n_4028)
);

AND2x2_ASAP7_75t_L g4029 ( 
.A(n_3976),
.B(n_3924),
.Y(n_4029)
);

INVxp67_ASAP7_75t_SL g4030 ( 
.A(n_3913),
.Y(n_4030)
);

BUFx2_ASAP7_75t_L g4031 ( 
.A(n_3979),
.Y(n_4031)
);

AND2x2_ASAP7_75t_L g4032 ( 
.A(n_3949),
.B(n_3899),
.Y(n_4032)
);

INVx1_ASAP7_75t_L g4033 ( 
.A(n_3948),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3963),
.B(n_3897),
.Y(n_4034)
);

HB1xp67_ASAP7_75t_L g4035 ( 
.A(n_3969),
.Y(n_4035)
);

INVx2_ASAP7_75t_L g4036 ( 
.A(n_3989),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3951),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3989),
.Y(n_4038)
);

INVx1_ASAP7_75t_L g4039 ( 
.A(n_3956),
.Y(n_4039)
);

HB1xp67_ASAP7_75t_L g4040 ( 
.A(n_3969),
.Y(n_4040)
);

INVx2_ASAP7_75t_L g4041 ( 
.A(n_3989),
.Y(n_4041)
);

AND2x2_ASAP7_75t_L g4042 ( 
.A(n_3987),
.B(n_3897),
.Y(n_4042)
);

OR2x2_ASAP7_75t_L g4043 ( 
.A(n_3972),
.B(n_3849),
.Y(n_4043)
);

BUFx2_ASAP7_75t_L g4044 ( 
.A(n_3941),
.Y(n_4044)
);

INVx1_ASAP7_75t_L g4045 ( 
.A(n_3966),
.Y(n_4045)
);

INVx1_ASAP7_75t_L g4046 ( 
.A(n_3982),
.Y(n_4046)
);

HB1xp67_ASAP7_75t_L g4047 ( 
.A(n_3936),
.Y(n_4047)
);

INVx2_ASAP7_75t_SL g4048 ( 
.A(n_3925),
.Y(n_4048)
);

AND2x4_ASAP7_75t_L g4049 ( 
.A(n_3983),
.B(n_3859),
.Y(n_4049)
);

INVx2_ASAP7_75t_L g4050 ( 
.A(n_4005),
.Y(n_4050)
);

INVx2_ASAP7_75t_L g4051 ( 
.A(n_4004),
.Y(n_4051)
);

HB1xp67_ASAP7_75t_L g4052 ( 
.A(n_3936),
.Y(n_4052)
);

INVx2_ASAP7_75t_L g4053 ( 
.A(n_4004),
.Y(n_4053)
);

AND2x2_ASAP7_75t_L g4054 ( 
.A(n_3921),
.B(n_3894),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_3988),
.B(n_3894),
.Y(n_4055)
);

INVx1_ASAP7_75t_L g4056 ( 
.A(n_3985),
.Y(n_4056)
);

INVx1_ASAP7_75t_L g4057 ( 
.A(n_3999),
.Y(n_4057)
);

INVx2_ASAP7_75t_L g4058 ( 
.A(n_3984),
.Y(n_4058)
);

OAI22xp5_ASAP7_75t_L g4059 ( 
.A1(n_3909),
.A2(n_3844),
.B1(n_3903),
.B2(n_3818),
.Y(n_4059)
);

INVx2_ASAP7_75t_L g4060 ( 
.A(n_3938),
.Y(n_4060)
);

AND2x2_ASAP7_75t_L g4061 ( 
.A(n_3988),
.B(n_3886),
.Y(n_4061)
);

AND2x4_ASAP7_75t_L g4062 ( 
.A(n_4000),
.B(n_3852),
.Y(n_4062)
);

NOR2xp33_ASAP7_75t_L g4063 ( 
.A(n_3920),
.B(n_3872),
.Y(n_4063)
);

BUFx4f_ASAP7_75t_SL g4064 ( 
.A(n_3993),
.Y(n_4064)
);

INVxp67_ASAP7_75t_R g4065 ( 
.A(n_3927),
.Y(n_4065)
);

INVx1_ASAP7_75t_L g4066 ( 
.A(n_4001),
.Y(n_4066)
);

AND2x4_ASAP7_75t_L g4067 ( 
.A(n_3992),
.B(n_3852),
.Y(n_4067)
);

INVx5_ASAP7_75t_L g4068 ( 
.A(n_3992),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_3957),
.Y(n_4069)
);

AND2x4_ASAP7_75t_L g4070 ( 
.A(n_3992),
.B(n_3929),
.Y(n_4070)
);

AND2x2_ASAP7_75t_L g4071 ( 
.A(n_3923),
.B(n_3844),
.Y(n_4071)
);

HB1xp67_ASAP7_75t_L g4072 ( 
.A(n_3938),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_3923),
.B(n_3858),
.Y(n_4073)
);

AND2x4_ASAP7_75t_L g4074 ( 
.A(n_3917),
.B(n_3821),
.Y(n_4074)
);

INVx2_ASAP7_75t_L g4075 ( 
.A(n_3995),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_3954),
.Y(n_4076)
);

INVx1_ASAP7_75t_L g4077 ( 
.A(n_3947),
.Y(n_4077)
);

BUFx6f_ASAP7_75t_L g4078 ( 
.A(n_3964),
.Y(n_4078)
);

OR2x2_ASAP7_75t_L g4079 ( 
.A(n_3914),
.B(n_3836),
.Y(n_4079)
);

INVx1_ASAP7_75t_L g4080 ( 
.A(n_3964),
.Y(n_4080)
);

INVx2_ASAP7_75t_L g4081 ( 
.A(n_3968),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_L g4082 ( 
.A(n_3950),
.B(n_3831),
.Y(n_4082)
);

HB1xp67_ASAP7_75t_L g4083 ( 
.A(n_3991),
.Y(n_4083)
);

AND2x4_ASAP7_75t_SL g4084 ( 
.A(n_3981),
.B(n_3858),
.Y(n_4084)
);

INVx2_ASAP7_75t_L g4085 ( 
.A(n_4007),
.Y(n_4085)
);

INVx3_ASAP7_75t_L g4086 ( 
.A(n_3986),
.Y(n_4086)
);

NOR2x1_ASAP7_75t_SL g4087 ( 
.A(n_3912),
.B(n_3855),
.Y(n_4087)
);

AND2x4_ASAP7_75t_L g4088 ( 
.A(n_3946),
.B(n_3820),
.Y(n_4088)
);

INVx1_ASAP7_75t_L g4089 ( 
.A(n_3974),
.Y(n_4089)
);

OR2x6_ASAP7_75t_L g4090 ( 
.A(n_3927),
.B(n_3806),
.Y(n_4090)
);

INVx2_ASAP7_75t_L g4091 ( 
.A(n_3986),
.Y(n_4091)
);

AND2x4_ASAP7_75t_L g4092 ( 
.A(n_3919),
.B(n_3820),
.Y(n_4092)
);

AND2x2_ASAP7_75t_L g4093 ( 
.A(n_3931),
.B(n_3855),
.Y(n_4093)
);

AND2x2_ASAP7_75t_L g4094 ( 
.A(n_3930),
.B(n_3893),
.Y(n_4094)
);

INVx1_ASAP7_75t_L g4095 ( 
.A(n_4006),
.Y(n_4095)
);

BUFx3_ASAP7_75t_L g4096 ( 
.A(n_3994),
.Y(n_4096)
);

INVx1_ASAP7_75t_L g4097 ( 
.A(n_3996),
.Y(n_4097)
);

NAND2xp5_ASAP7_75t_L g4098 ( 
.A(n_3932),
.B(n_3819),
.Y(n_4098)
);

NAND2x1p5_ASAP7_75t_L g4099 ( 
.A(n_4002),
.B(n_3806),
.Y(n_4099)
);

INVx1_ASAP7_75t_L g4100 ( 
.A(n_3935),
.Y(n_4100)
);

INVx1_ASAP7_75t_L g4101 ( 
.A(n_3955),
.Y(n_4101)
);

AND2x2_ASAP7_75t_L g4102 ( 
.A(n_4030),
.B(n_3943),
.Y(n_4102)
);

AND2x4_ASAP7_75t_L g4103 ( 
.A(n_4021),
.B(n_3821),
.Y(n_4103)
);

INVx3_ASAP7_75t_L g4104 ( 
.A(n_4078),
.Y(n_4104)
);

AND2x2_ASAP7_75t_L g4105 ( 
.A(n_4031),
.B(n_3910),
.Y(n_4105)
);

HB1xp67_ASAP7_75t_L g4106 ( 
.A(n_4072),
.Y(n_4106)
);

HB1xp67_ASAP7_75t_L g4107 ( 
.A(n_4013),
.Y(n_4107)
);

OAI22xp5_ASAP7_75t_L g4108 ( 
.A1(n_4100),
.A2(n_3915),
.B1(n_3933),
.B2(n_3961),
.Y(n_4108)
);

INVx1_ASAP7_75t_L g4109 ( 
.A(n_4078),
.Y(n_4109)
);

NAND2xp5_ASAP7_75t_L g4110 ( 
.A(n_4100),
.B(n_3958),
.Y(n_4110)
);

NAND2xp5_ASAP7_75t_L g4111 ( 
.A(n_4060),
.B(n_3953),
.Y(n_4111)
);

BUFx2_ASAP7_75t_L g4112 ( 
.A(n_4031),
.Y(n_4112)
);

NAND2xp5_ASAP7_75t_L g4113 ( 
.A(n_4060),
.B(n_3953),
.Y(n_4113)
);

AND2x2_ASAP7_75t_L g4114 ( 
.A(n_4013),
.B(n_3893),
.Y(n_4114)
);

AND2x2_ASAP7_75t_L g4115 ( 
.A(n_4083),
.B(n_3893),
.Y(n_4115)
);

INVx1_ASAP7_75t_L g4116 ( 
.A(n_4078),
.Y(n_4116)
);

BUFx2_ASAP7_75t_L g4117 ( 
.A(n_4078),
.Y(n_4117)
);

HB1xp67_ASAP7_75t_L g4118 ( 
.A(n_4048),
.Y(n_4118)
);

INVx2_ASAP7_75t_L g4119 ( 
.A(n_4078),
.Y(n_4119)
);

AND2x2_ASAP7_75t_L g4120 ( 
.A(n_4065),
.B(n_3813),
.Y(n_4120)
);

AND2x2_ASAP7_75t_L g4121 ( 
.A(n_4065),
.B(n_3813),
.Y(n_4121)
);

INVx1_ASAP7_75t_L g4122 ( 
.A(n_4047),
.Y(n_4122)
);

OR2x2_ASAP7_75t_L g4123 ( 
.A(n_4020),
.B(n_4035),
.Y(n_4123)
);

AND2x4_ASAP7_75t_L g4124 ( 
.A(n_4021),
.B(n_3802),
.Y(n_4124)
);

INVx1_ASAP7_75t_L g4125 ( 
.A(n_4052),
.Y(n_4125)
);

INVx2_ASAP7_75t_L g4126 ( 
.A(n_4086),
.Y(n_4126)
);

AND2x4_ASAP7_75t_L g4127 ( 
.A(n_4025),
.B(n_3802),
.Y(n_4127)
);

AND2x2_ASAP7_75t_L g4128 ( 
.A(n_4075),
.B(n_4029),
.Y(n_4128)
);

AND2x2_ASAP7_75t_L g4129 ( 
.A(n_4075),
.B(n_3871),
.Y(n_4129)
);

INVx2_ASAP7_75t_SL g4130 ( 
.A(n_4068),
.Y(n_4130)
);

INVx2_ASAP7_75t_L g4131 ( 
.A(n_4044),
.Y(n_4131)
);

AND2x4_ASAP7_75t_L g4132 ( 
.A(n_4025),
.B(n_3822),
.Y(n_4132)
);

BUFx6f_ASAP7_75t_L g4133 ( 
.A(n_4044),
.Y(n_4133)
);

AND2x2_ASAP7_75t_L g4134 ( 
.A(n_4029),
.B(n_3828),
.Y(n_4134)
);

AND2x2_ASAP7_75t_L g4135 ( 
.A(n_4048),
.B(n_3834),
.Y(n_4135)
);

INVxp67_ASAP7_75t_SL g4136 ( 
.A(n_4087),
.Y(n_4136)
);

INVx1_ASAP7_75t_SL g4137 ( 
.A(n_4064),
.Y(n_4137)
);

BUFx2_ASAP7_75t_L g4138 ( 
.A(n_4040),
.Y(n_4138)
);

INVx1_ASAP7_75t_L g4139 ( 
.A(n_4010),
.Y(n_4139)
);

BUFx2_ASAP7_75t_L g4140 ( 
.A(n_4088),
.Y(n_4140)
);

INVx3_ASAP7_75t_L g4141 ( 
.A(n_4049),
.Y(n_4141)
);

BUFx2_ASAP7_75t_SL g4142 ( 
.A(n_4068),
.Y(n_4142)
);

INVx1_ASAP7_75t_L g4143 ( 
.A(n_4010),
.Y(n_4143)
);

INVx2_ASAP7_75t_L g4144 ( 
.A(n_4049),
.Y(n_4144)
);

OR2x2_ASAP7_75t_L g4145 ( 
.A(n_4020),
.B(n_3832),
.Y(n_4145)
);

AND2x4_ASAP7_75t_L g4146 ( 
.A(n_4068),
.B(n_3822),
.Y(n_4146)
);

OR2x2_ASAP7_75t_L g4147 ( 
.A(n_4080),
.B(n_3823),
.Y(n_4147)
);

INVx1_ASAP7_75t_L g4148 ( 
.A(n_4017),
.Y(n_4148)
);

INVx1_ASAP7_75t_L g4149 ( 
.A(n_4017),
.Y(n_4149)
);

INVx2_ASAP7_75t_L g4150 ( 
.A(n_4086),
.Y(n_4150)
);

INVx1_ASAP7_75t_L g4151 ( 
.A(n_4037),
.Y(n_4151)
);

NAND2xp5_ASAP7_75t_L g4152 ( 
.A(n_4024),
.B(n_3918),
.Y(n_4152)
);

INVx2_ASAP7_75t_L g4153 ( 
.A(n_4086),
.Y(n_4153)
);

INVx2_ASAP7_75t_L g4154 ( 
.A(n_4087),
.Y(n_4154)
);

AND2x2_ASAP7_75t_L g4155 ( 
.A(n_4012),
.B(n_3808),
.Y(n_4155)
);

INVx3_ASAP7_75t_L g4156 ( 
.A(n_4133),
.Y(n_4156)
);

AND2x2_ASAP7_75t_L g4157 ( 
.A(n_4112),
.B(n_4055),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4138),
.Y(n_4158)
);

BUFx3_ASAP7_75t_L g4159 ( 
.A(n_4112),
.Y(n_4159)
);

AND2x2_ASAP7_75t_L g4160 ( 
.A(n_4141),
.B(n_4128),
.Y(n_4160)
);

INVx2_ASAP7_75t_L g4161 ( 
.A(n_4138),
.Y(n_4161)
);

INVx1_ASAP7_75t_L g4162 ( 
.A(n_4117),
.Y(n_4162)
);

INVx2_ASAP7_75t_L g4163 ( 
.A(n_4117),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4106),
.Y(n_4164)
);

INVx2_ASAP7_75t_L g4165 ( 
.A(n_4104),
.Y(n_4165)
);

BUFx2_ASAP7_75t_L g4166 ( 
.A(n_4136),
.Y(n_4166)
);

INVx2_ASAP7_75t_L g4167 ( 
.A(n_4104),
.Y(n_4167)
);

AND2x2_ASAP7_75t_L g4168 ( 
.A(n_4141),
.B(n_4128),
.Y(n_4168)
);

AND2x2_ASAP7_75t_L g4169 ( 
.A(n_4141),
.B(n_4055),
.Y(n_4169)
);

INVx2_ASAP7_75t_L g4170 ( 
.A(n_4104),
.Y(n_4170)
);

AND2x2_ASAP7_75t_L g4171 ( 
.A(n_4141),
.B(n_4061),
.Y(n_4171)
);

AND2x2_ASAP7_75t_L g4172 ( 
.A(n_4154),
.B(n_4061),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4104),
.Y(n_4173)
);

INVx1_ASAP7_75t_L g4174 ( 
.A(n_4133),
.Y(n_4174)
);

AOI33xp33_ASAP7_75t_L g4175 ( 
.A1(n_4102),
.A2(n_4097),
.A3(n_4092),
.B1(n_3944),
.B2(n_4094),
.B3(n_4101),
.Y(n_4175)
);

INVx2_ASAP7_75t_L g4176 ( 
.A(n_4140),
.Y(n_4176)
);

OR2x2_ASAP7_75t_L g4177 ( 
.A(n_4123),
.B(n_4079),
.Y(n_4177)
);

INVx3_ASAP7_75t_L g4178 ( 
.A(n_4133),
.Y(n_4178)
);

AND2x2_ASAP7_75t_L g4179 ( 
.A(n_4154),
.B(n_4107),
.Y(n_4179)
);

INVx2_ASAP7_75t_L g4180 ( 
.A(n_4140),
.Y(n_4180)
);

INVx1_ASAP7_75t_L g4181 ( 
.A(n_4133),
.Y(n_4181)
);

HB1xp67_ASAP7_75t_L g4182 ( 
.A(n_4133),
.Y(n_4182)
);

INVx3_ASAP7_75t_L g4183 ( 
.A(n_4133),
.Y(n_4183)
);

NAND2xp5_ASAP7_75t_L g4184 ( 
.A(n_4131),
.B(n_4122),
.Y(n_4184)
);

HB1xp67_ASAP7_75t_L g4185 ( 
.A(n_4122),
.Y(n_4185)
);

AND2x2_ASAP7_75t_L g4186 ( 
.A(n_4105),
.B(n_4024),
.Y(n_4186)
);

AND2x2_ASAP7_75t_L g4187 ( 
.A(n_4154),
.B(n_4026),
.Y(n_4187)
);

AND2x4_ASAP7_75t_L g4188 ( 
.A(n_4130),
.B(n_4068),
.Y(n_4188)
);

INVxp67_ASAP7_75t_L g4189 ( 
.A(n_4118),
.Y(n_4189)
);

OAI22xp5_ASAP7_75t_L g4190 ( 
.A1(n_4108),
.A2(n_3970),
.B1(n_3942),
.B2(n_4079),
.Y(n_4190)
);

HB1xp67_ASAP7_75t_L g4191 ( 
.A(n_4125),
.Y(n_4191)
);

OAI22xp5_ASAP7_75t_L g4192 ( 
.A1(n_4123),
.A2(n_4098),
.B1(n_4092),
.B2(n_4016),
.Y(n_4192)
);

INVx1_ASAP7_75t_SL g4193 ( 
.A(n_4142),
.Y(n_4193)
);

INVx1_ASAP7_75t_L g4194 ( 
.A(n_4126),
.Y(n_4194)
);

INVx1_ASAP7_75t_L g4195 ( 
.A(n_4126),
.Y(n_4195)
);

INVx1_ASAP7_75t_L g4196 ( 
.A(n_4126),
.Y(n_4196)
);

INVx1_ASAP7_75t_L g4197 ( 
.A(n_4150),
.Y(n_4197)
);

INVx1_ASAP7_75t_L g4198 ( 
.A(n_4150),
.Y(n_4198)
);

AND2x2_ASAP7_75t_L g4199 ( 
.A(n_4105),
.B(n_4026),
.Y(n_4199)
);

AND2x4_ASAP7_75t_L g4200 ( 
.A(n_4130),
.B(n_4068),
.Y(n_4200)
);

INVx4_ASAP7_75t_L g4201 ( 
.A(n_4119),
.Y(n_4201)
);

INVx2_ASAP7_75t_SL g4202 ( 
.A(n_4127),
.Y(n_4202)
);

INVx4_ASAP7_75t_L g4203 ( 
.A(n_4119),
.Y(n_4203)
);

INVx2_ASAP7_75t_L g4204 ( 
.A(n_4125),
.Y(n_4204)
);

INVx2_ASAP7_75t_L g4205 ( 
.A(n_4119),
.Y(n_4205)
);

INVx1_ASAP7_75t_L g4206 ( 
.A(n_4150),
.Y(n_4206)
);

AND2x2_ASAP7_75t_L g4207 ( 
.A(n_4131),
.B(n_4028),
.Y(n_4207)
);

INVx1_ASAP7_75t_L g4208 ( 
.A(n_4182),
.Y(n_4208)
);

AND2x2_ASAP7_75t_L g4209 ( 
.A(n_4186),
.B(n_4137),
.Y(n_4209)
);

OAI21xp5_ASAP7_75t_L g4210 ( 
.A1(n_4192),
.A2(n_4110),
.B(n_4059),
.Y(n_4210)
);

HB1xp67_ASAP7_75t_L g4211 ( 
.A(n_4159),
.Y(n_4211)
);

INVx2_ASAP7_75t_L g4212 ( 
.A(n_4159),
.Y(n_4212)
);

NAND2xp5_ASAP7_75t_L g4213 ( 
.A(n_4186),
.B(n_4102),
.Y(n_4213)
);

OAI21xp33_ASAP7_75t_L g4214 ( 
.A1(n_4175),
.A2(n_4152),
.B(n_4111),
.Y(n_4214)
);

NAND2xp5_ASAP7_75t_L g4215 ( 
.A(n_4199),
.B(n_4120),
.Y(n_4215)
);

NAND2xp5_ASAP7_75t_L g4216 ( 
.A(n_4199),
.B(n_4120),
.Y(n_4216)
);

INVx2_ASAP7_75t_L g4217 ( 
.A(n_4159),
.Y(n_4217)
);

AND2x4_ASAP7_75t_L g4218 ( 
.A(n_4202),
.B(n_4176),
.Y(n_4218)
);

AND2x2_ASAP7_75t_L g4219 ( 
.A(n_4160),
.B(n_4070),
.Y(n_4219)
);

NAND2xp5_ASAP7_75t_L g4220 ( 
.A(n_4157),
.B(n_4121),
.Y(n_4220)
);

AND2x2_ASAP7_75t_L g4221 ( 
.A(n_4160),
.B(n_4121),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4182),
.Y(n_4222)
);

AND2x4_ASAP7_75t_L g4223 ( 
.A(n_4202),
.B(n_4144),
.Y(n_4223)
);

NOR2xp33_ASAP7_75t_L g4224 ( 
.A(n_4166),
.B(n_4113),
.Y(n_4224)
);

INVx2_ASAP7_75t_L g4225 ( 
.A(n_4156),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4176),
.Y(n_4226)
);

NAND2xp67_ASAP7_75t_L g4227 ( 
.A(n_4157),
.B(n_4153),
.Y(n_4227)
);

NAND2xp5_ASAP7_75t_L g4228 ( 
.A(n_4157),
.B(n_4028),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_4156),
.Y(n_4229)
);

AND2x2_ASAP7_75t_L g4230 ( 
.A(n_4160),
.B(n_4070),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4168),
.B(n_4081),
.Y(n_4231)
);

INVx1_ASAP7_75t_L g4232 ( 
.A(n_4176),
.Y(n_4232)
);

INVx2_ASAP7_75t_L g4233 ( 
.A(n_4156),
.Y(n_4233)
);

AND2x4_ASAP7_75t_L g4234 ( 
.A(n_4202),
.B(n_4144),
.Y(n_4234)
);

AND2x4_ASAP7_75t_SL g4235 ( 
.A(n_4168),
.B(n_4103),
.Y(n_4235)
);

INVx2_ASAP7_75t_SL g4236 ( 
.A(n_4156),
.Y(n_4236)
);

OR2x2_ASAP7_75t_L g4237 ( 
.A(n_4177),
.B(n_4009),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4168),
.B(n_4070),
.Y(n_4238)
);

OR2x6_ASAP7_75t_L g4239 ( 
.A(n_4158),
.B(n_4142),
.Y(n_4239)
);

INVx1_ASAP7_75t_L g4240 ( 
.A(n_4180),
.Y(n_4240)
);

INVx1_ASAP7_75t_L g4241 ( 
.A(n_4180),
.Y(n_4241)
);

NAND2xp5_ASAP7_75t_L g4242 ( 
.A(n_4172),
.B(n_4081),
.Y(n_4242)
);

NAND2xp5_ASAP7_75t_L g4243 ( 
.A(n_4172),
.B(n_4169),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4180),
.Y(n_4244)
);

AND2x2_ASAP7_75t_L g4245 ( 
.A(n_4169),
.B(n_4050),
.Y(n_4245)
);

AND2x4_ASAP7_75t_L g4246 ( 
.A(n_4178),
.B(n_4103),
.Y(n_4246)
);

INVx2_ASAP7_75t_L g4247 ( 
.A(n_4218),
.Y(n_4247)
);

AND2x2_ASAP7_75t_L g4248 ( 
.A(n_4209),
.B(n_4219),
.Y(n_4248)
);

NAND3xp33_ASAP7_75t_L g4249 ( 
.A(n_4224),
.B(n_4192),
.C(n_4161),
.Y(n_4249)
);

INVx2_ASAP7_75t_L g4250 ( 
.A(n_4218),
.Y(n_4250)
);

NAND2xp5_ASAP7_75t_SL g4251 ( 
.A(n_4230),
.B(n_4103),
.Y(n_4251)
);

INVx1_ASAP7_75t_L g4252 ( 
.A(n_4211),
.Y(n_4252)
);

AND2x4_ASAP7_75t_SL g4253 ( 
.A(n_4238),
.B(n_4129),
.Y(n_4253)
);

NAND2x1p5_ASAP7_75t_L g4254 ( 
.A(n_4212),
.B(n_4193),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4211),
.Y(n_4255)
);

OR2x2_ASAP7_75t_L g4256 ( 
.A(n_4243),
.B(n_4177),
.Y(n_4256)
);

INVx1_ASAP7_75t_L g4257 ( 
.A(n_4218),
.Y(n_4257)
);

NAND4xp25_ASAP7_75t_L g4258 ( 
.A(n_4214),
.B(n_4164),
.C(n_4190),
.D(n_4166),
.Y(n_4258)
);

NAND2x1p5_ASAP7_75t_L g4259 ( 
.A(n_4212),
.B(n_4193),
.Y(n_4259)
);

HB1xp67_ASAP7_75t_L g4260 ( 
.A(n_4227),
.Y(n_4260)
);

INVxp67_ASAP7_75t_L g4261 ( 
.A(n_4239),
.Y(n_4261)
);

OR2x2_ASAP7_75t_L g4262 ( 
.A(n_4220),
.B(n_4164),
.Y(n_4262)
);

CKINVDCx5p33_ASAP7_75t_R g4263 ( 
.A(n_4239),
.Y(n_4263)
);

AND2x2_ASAP7_75t_L g4264 ( 
.A(n_4245),
.B(n_4169),
.Y(n_4264)
);

AND2x2_ASAP7_75t_L g4265 ( 
.A(n_4221),
.B(n_4171),
.Y(n_4265)
);

BUFx3_ASAP7_75t_L g4266 ( 
.A(n_4235),
.Y(n_4266)
);

OA22x2_ASAP7_75t_L g4267 ( 
.A1(n_4210),
.A2(n_4190),
.B1(n_4172),
.B2(n_4161),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4223),
.Y(n_4268)
);

INVx1_ASAP7_75t_L g4269 ( 
.A(n_4223),
.Y(n_4269)
);

INVx1_ASAP7_75t_L g4270 ( 
.A(n_4223),
.Y(n_4270)
);

NAND3xp33_ASAP7_75t_L g4271 ( 
.A(n_4224),
.B(n_4161),
.C(n_4158),
.Y(n_4271)
);

INVx2_ASAP7_75t_L g4272 ( 
.A(n_4235),
.Y(n_4272)
);

INVx1_ASAP7_75t_L g4273 ( 
.A(n_4268),
.Y(n_4273)
);

AND2x2_ASAP7_75t_L g4274 ( 
.A(n_4248),
.B(n_4221),
.Y(n_4274)
);

INVx1_ASAP7_75t_L g4275 ( 
.A(n_4269),
.Y(n_4275)
);

NAND4xp25_ASAP7_75t_L g4276 ( 
.A(n_4249),
.B(n_4258),
.C(n_4271),
.D(n_4266),
.Y(n_4276)
);

OR2x2_ASAP7_75t_L g4277 ( 
.A(n_4256),
.B(n_4213),
.Y(n_4277)
);

NOR2xp33_ASAP7_75t_L g4278 ( 
.A(n_4254),
.B(n_4259),
.Y(n_4278)
);

AND2x2_ASAP7_75t_L g4279 ( 
.A(n_4264),
.B(n_4129),
.Y(n_4279)
);

OR2x2_ASAP7_75t_L g4280 ( 
.A(n_4254),
.B(n_4228),
.Y(n_4280)
);

AND2x2_ASAP7_75t_L g4281 ( 
.A(n_4265),
.B(n_4171),
.Y(n_4281)
);

INVx1_ASAP7_75t_L g4282 ( 
.A(n_4270),
.Y(n_4282)
);

INVx4_ASAP7_75t_L g4283 ( 
.A(n_4259),
.Y(n_4283)
);

AND2x2_ASAP7_75t_L g4284 ( 
.A(n_4253),
.B(n_4171),
.Y(n_4284)
);

INVx1_ASAP7_75t_L g4285 ( 
.A(n_4257),
.Y(n_4285)
);

AND2x2_ASAP7_75t_L g4286 ( 
.A(n_4272),
.B(n_4179),
.Y(n_4286)
);

NOR2xp33_ASAP7_75t_L g4287 ( 
.A(n_4271),
.B(n_4217),
.Y(n_4287)
);

AND2x2_ASAP7_75t_L g4288 ( 
.A(n_4247),
.B(n_4179),
.Y(n_4288)
);

AND2x4_ASAP7_75t_L g4289 ( 
.A(n_4250),
.B(n_4217),
.Y(n_4289)
);

AND2x2_ASAP7_75t_L g4290 ( 
.A(n_4251),
.B(n_4179),
.Y(n_4290)
);

INVx1_ASAP7_75t_L g4291 ( 
.A(n_4260),
.Y(n_4291)
);

AND2x4_ASAP7_75t_L g4292 ( 
.A(n_4252),
.B(n_4246),
.Y(n_4292)
);

INVx1_ASAP7_75t_L g4293 ( 
.A(n_4292),
.Y(n_4293)
);

INVx2_ASAP7_75t_SL g4294 ( 
.A(n_4292),
.Y(n_4294)
);

INVx1_ASAP7_75t_L g4295 ( 
.A(n_4292),
.Y(n_4295)
);

OAI22xp33_ASAP7_75t_L g4296 ( 
.A1(n_4276),
.A2(n_4090),
.B1(n_4267),
.B2(n_4249),
.Y(n_4296)
);

A2O1A1Ixp33_ASAP7_75t_L g4297 ( 
.A1(n_4287),
.A2(n_4088),
.B(n_4237),
.C(n_4158),
.Y(n_4297)
);

INVx2_ASAP7_75t_SL g4298 ( 
.A(n_4284),
.Y(n_4298)
);

AOI21xp33_ASAP7_75t_L g4299 ( 
.A1(n_4278),
.A2(n_4267),
.B(n_4263),
.Y(n_4299)
);

INVx1_ASAP7_75t_L g4300 ( 
.A(n_4281),
.Y(n_4300)
);

OAI32xp33_ASAP7_75t_L g4301 ( 
.A1(n_4276),
.A2(n_4185),
.A3(n_4191),
.B1(n_4258),
.B2(n_4189),
.Y(n_4301)
);

AOI22xp5_ASAP7_75t_L g4302 ( 
.A1(n_4287),
.A2(n_4189),
.B1(n_4191),
.B2(n_4185),
.Y(n_4302)
);

NAND2xp5_ASAP7_75t_L g4303 ( 
.A(n_4274),
.B(n_4207),
.Y(n_4303)
);

INVx1_ASAP7_75t_L g4304 ( 
.A(n_4288),
.Y(n_4304)
);

INVx2_ASAP7_75t_L g4305 ( 
.A(n_4283),
.Y(n_4305)
);

OAI322xp33_ASAP7_75t_L g4306 ( 
.A1(n_4278),
.A2(n_4261),
.A3(n_4184),
.B1(n_4216),
.B2(n_4215),
.C1(n_4262),
.C2(n_4139),
.Y(n_4306)
);

INVx1_ASAP7_75t_L g4307 ( 
.A(n_4286),
.Y(n_4307)
);

O2A1O1Ixp5_ASAP7_75t_R g4308 ( 
.A1(n_4290),
.A2(n_4242),
.B(n_4231),
.C(n_4184),
.Y(n_4308)
);

INVx1_ASAP7_75t_L g4309 ( 
.A(n_4280),
.Y(n_4309)
);

INVx2_ASAP7_75t_L g4310 ( 
.A(n_4294),
.Y(n_4310)
);

AND2x2_ASAP7_75t_L g4311 ( 
.A(n_4298),
.B(n_4279),
.Y(n_4311)
);

NAND2xp5_ASAP7_75t_L g4312 ( 
.A(n_4293),
.B(n_4178),
.Y(n_4312)
);

AND2x2_ASAP7_75t_L g4313 ( 
.A(n_4300),
.B(n_4289),
.Y(n_4313)
);

AND2x2_ASAP7_75t_L g4314 ( 
.A(n_4307),
.B(n_4289),
.Y(n_4314)
);

OAI33xp33_ASAP7_75t_L g4315 ( 
.A1(n_4296),
.A2(n_4261),
.A3(n_4222),
.B1(n_4208),
.B2(n_4255),
.B3(n_4232),
.Y(n_4315)
);

OR2x2_ASAP7_75t_L g4316 ( 
.A(n_4295),
.B(n_4303),
.Y(n_4316)
);

INVx3_ASAP7_75t_SL g4317 ( 
.A(n_4305),
.Y(n_4317)
);

HB1xp67_ASAP7_75t_L g4318 ( 
.A(n_4302),
.Y(n_4318)
);

AND2x2_ASAP7_75t_L g4319 ( 
.A(n_4304),
.B(n_4283),
.Y(n_4319)
);

AOI21xp5_ASAP7_75t_L g4320 ( 
.A1(n_4297),
.A2(n_4239),
.B(n_4260),
.Y(n_4320)
);

AND2x2_ASAP7_75t_L g4321 ( 
.A(n_4309),
.B(n_4207),
.Y(n_4321)
);

INVx3_ASAP7_75t_SL g4322 ( 
.A(n_4317),
.Y(n_4322)
);

OR2x2_ASAP7_75t_L g4323 ( 
.A(n_4310),
.B(n_4277),
.Y(n_4323)
);

INVx1_ASAP7_75t_SL g4324 ( 
.A(n_4321),
.Y(n_4324)
);

NOR2xp33_ASAP7_75t_L g4325 ( 
.A(n_4315),
.B(n_4306),
.Y(n_4325)
);

OR2x2_ASAP7_75t_L g4326 ( 
.A(n_4316),
.B(n_4273),
.Y(n_4326)
);

NOR2xp33_ASAP7_75t_L g4327 ( 
.A(n_4311),
.B(n_4299),
.Y(n_4327)
);

INVx1_ASAP7_75t_SL g4328 ( 
.A(n_4313),
.Y(n_4328)
);

INVx2_ASAP7_75t_SL g4329 ( 
.A(n_4314),
.Y(n_4329)
);

AOI21xp33_ASAP7_75t_SL g4330 ( 
.A1(n_4322),
.A2(n_4302),
.B(n_4240),
.Y(n_4330)
);

OR2x2_ASAP7_75t_L g4331 ( 
.A(n_4328),
.B(n_4275),
.Y(n_4331)
);

OAI21xp33_ASAP7_75t_L g4332 ( 
.A1(n_4327),
.A2(n_4115),
.B(n_4319),
.Y(n_4332)
);

INVx1_ASAP7_75t_L g4333 ( 
.A(n_4323),
.Y(n_4333)
);

AOI22xp5_ASAP7_75t_L g4334 ( 
.A1(n_4329),
.A2(n_4207),
.B1(n_4050),
.B2(n_4187),
.Y(n_4334)
);

NAND2x1_ASAP7_75t_L g4335 ( 
.A(n_4326),
.B(n_4246),
.Y(n_4335)
);

NAND2xp5_ASAP7_75t_L g4336 ( 
.A(n_4324),
.B(n_4226),
.Y(n_4336)
);

AND2x2_ASAP7_75t_L g4337 ( 
.A(n_4325),
.B(n_4282),
.Y(n_4337)
);

OAI31xp33_ASAP7_75t_L g4338 ( 
.A1(n_4325),
.A2(n_4318),
.A3(n_4241),
.B(n_4244),
.Y(n_4338)
);

INVx2_ASAP7_75t_L g4339 ( 
.A(n_4329),
.Y(n_4339)
);

OR2x2_ASAP7_75t_L g4340 ( 
.A(n_4322),
.B(n_4285),
.Y(n_4340)
);

AND2x2_ASAP7_75t_L g4341 ( 
.A(n_4322),
.B(n_4174),
.Y(n_4341)
);

NAND2xp5_ASAP7_75t_L g4342 ( 
.A(n_4322),
.B(n_4162),
.Y(n_4342)
);

OAI211xp5_ASAP7_75t_L g4343 ( 
.A1(n_4338),
.A2(n_4301),
.B(n_4320),
.C(n_4312),
.Y(n_4343)
);

NAND3xp33_ASAP7_75t_L g4344 ( 
.A(n_4330),
.B(n_4291),
.C(n_4312),
.Y(n_4344)
);

NOR2xp33_ASAP7_75t_L g4345 ( 
.A(n_4334),
.B(n_4308),
.Y(n_4345)
);

INVx1_ASAP7_75t_L g4346 ( 
.A(n_4335),
.Y(n_4346)
);

INVx2_ASAP7_75t_L g4347 ( 
.A(n_4341),
.Y(n_4347)
);

HB1xp67_ASAP7_75t_L g4348 ( 
.A(n_4342),
.Y(n_4348)
);

OAI21xp33_ASAP7_75t_L g4349 ( 
.A1(n_4337),
.A2(n_4187),
.B(n_4115),
.Y(n_4349)
);

OAI211xp5_ASAP7_75t_L g4350 ( 
.A1(n_4332),
.A2(n_4174),
.B(n_4181),
.C(n_4178),
.Y(n_4350)
);

NAND2xp5_ASAP7_75t_L g4351 ( 
.A(n_4333),
.B(n_4162),
.Y(n_4351)
);

NAND2xp5_ASAP7_75t_SL g4352 ( 
.A(n_4336),
.B(n_4246),
.Y(n_4352)
);

AOI32xp33_ASAP7_75t_L g4353 ( 
.A1(n_4339),
.A2(n_4178),
.A3(n_4183),
.B1(n_4181),
.B2(n_4200),
.Y(n_4353)
);

NAND2xp5_ASAP7_75t_L g4354 ( 
.A(n_4340),
.B(n_4234),
.Y(n_4354)
);

INVx1_ASAP7_75t_L g4355 ( 
.A(n_4331),
.Y(n_4355)
);

INVx1_ASAP7_75t_L g4356 ( 
.A(n_4335),
.Y(n_4356)
);

OAI222xp33_ASAP7_75t_L g4357 ( 
.A1(n_4334),
.A2(n_4183),
.B1(n_4236),
.B2(n_4163),
.C1(n_4188),
.C2(n_4200),
.Y(n_4357)
);

NAND2xp5_ASAP7_75t_SL g4358 ( 
.A(n_4334),
.B(n_4188),
.Y(n_4358)
);

AND2x2_ASAP7_75t_L g4359 ( 
.A(n_4341),
.B(n_4234),
.Y(n_4359)
);

INVx2_ASAP7_75t_L g4360 ( 
.A(n_4335),
.Y(n_4360)
);

INVx1_ASAP7_75t_SL g4361 ( 
.A(n_4341),
.Y(n_4361)
);

NAND2xp5_ASAP7_75t_L g4362 ( 
.A(n_4334),
.B(n_4234),
.Y(n_4362)
);

XNOR2x2_ASAP7_75t_L g4363 ( 
.A(n_4342),
.B(n_4163),
.Y(n_4363)
);

INVx1_ASAP7_75t_L g4364 ( 
.A(n_4335),
.Y(n_4364)
);

AND2x4_ASAP7_75t_L g4365 ( 
.A(n_4359),
.B(n_4236),
.Y(n_4365)
);

INVx1_ASAP7_75t_L g4366 ( 
.A(n_4354),
.Y(n_4366)
);

NOR2xp33_ASAP7_75t_L g4367 ( 
.A(n_4349),
.B(n_4357),
.Y(n_4367)
);

INVx2_ASAP7_75t_L g4368 ( 
.A(n_4363),
.Y(n_4368)
);

OR2x2_ASAP7_75t_L g4369 ( 
.A(n_4360),
.B(n_4183),
.Y(n_4369)
);

INVx1_ASAP7_75t_L g4370 ( 
.A(n_4362),
.Y(n_4370)
);

NAND2xp5_ASAP7_75t_SL g4371 ( 
.A(n_4346),
.B(n_4188),
.Y(n_4371)
);

INVx1_ASAP7_75t_L g4372 ( 
.A(n_4356),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4364),
.Y(n_4373)
);

NAND2xp5_ASAP7_75t_L g4374 ( 
.A(n_4353),
.B(n_4183),
.Y(n_4374)
);

INVx1_ASAP7_75t_L g4375 ( 
.A(n_4351),
.Y(n_4375)
);

AND2x2_ASAP7_75t_L g4376 ( 
.A(n_4361),
.B(n_4163),
.Y(n_4376)
);

BUFx2_ASAP7_75t_L g4377 ( 
.A(n_4347),
.Y(n_4377)
);

AND2x2_ASAP7_75t_L g4378 ( 
.A(n_4355),
.B(n_4187),
.Y(n_4378)
);

INVx1_ASAP7_75t_L g4379 ( 
.A(n_4358),
.Y(n_4379)
);

AND2x2_ASAP7_75t_L g4380 ( 
.A(n_4352),
.B(n_4225),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4350),
.B(n_4225),
.Y(n_4381)
);

NAND2xp33_ASAP7_75t_L g4382 ( 
.A(n_4348),
.B(n_4229),
.Y(n_4382)
);

NOR3xp33_ASAP7_75t_SL g4383 ( 
.A(n_4343),
.B(n_4116),
.C(n_4109),
.Y(n_4383)
);

NOR2xp33_ASAP7_75t_L g4384 ( 
.A(n_4344),
.B(n_4229),
.Y(n_4384)
);

AND2x2_ASAP7_75t_L g4385 ( 
.A(n_4345),
.B(n_4233),
.Y(n_4385)
);

NAND2xp5_ASAP7_75t_L g4386 ( 
.A(n_4344),
.B(n_4139),
.Y(n_4386)
);

AND2x2_ASAP7_75t_L g4387 ( 
.A(n_4359),
.B(n_4233),
.Y(n_4387)
);

AND2x2_ASAP7_75t_L g4388 ( 
.A(n_4359),
.B(n_4188),
.Y(n_4388)
);

AOI22xp33_ASAP7_75t_SL g4389 ( 
.A1(n_4359),
.A2(n_4200),
.B1(n_4204),
.B2(n_4109),
.Y(n_4389)
);

NOR2xp33_ASAP7_75t_L g4390 ( 
.A(n_4349),
.B(n_4200),
.Y(n_4390)
);

CKINVDCx16_ASAP7_75t_R g4391 ( 
.A(n_4378),
.Y(n_4391)
);

INVxp67_ASAP7_75t_SL g4392 ( 
.A(n_4371),
.Y(n_4392)
);

INVx2_ASAP7_75t_SL g4393 ( 
.A(n_4365),
.Y(n_4393)
);

OR2x2_ASAP7_75t_L g4394 ( 
.A(n_4365),
.B(n_4388),
.Y(n_4394)
);

NAND2xp5_ASAP7_75t_L g4395 ( 
.A(n_4389),
.B(n_4143),
.Y(n_4395)
);

XNOR2x1_ASAP7_75t_L g4396 ( 
.A(n_4376),
.B(n_4204),
.Y(n_4396)
);

INVx1_ASAP7_75t_L g4397 ( 
.A(n_4387),
.Y(n_4397)
);

INVx1_ASAP7_75t_L g4398 ( 
.A(n_4369),
.Y(n_4398)
);

INVx3_ASAP7_75t_L g4399 ( 
.A(n_4380),
.Y(n_4399)
);

NOR2x1p5_ASAP7_75t_L g4400 ( 
.A(n_4379),
.B(n_4204),
.Y(n_4400)
);

NOR2x1_ASAP7_75t_L g4401 ( 
.A(n_4368),
.B(n_4201),
.Y(n_4401)
);

NAND2xp5_ASAP7_75t_L g4402 ( 
.A(n_4384),
.B(n_4143),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4377),
.Y(n_4403)
);

INVx2_ASAP7_75t_L g4404 ( 
.A(n_4372),
.Y(n_4404)
);

NOR3xp33_ASAP7_75t_L g4405 ( 
.A(n_4373),
.B(n_4203),
.C(n_4201),
.Y(n_4405)
);

NAND2xp5_ASAP7_75t_L g4406 ( 
.A(n_4390),
.B(n_4116),
.Y(n_4406)
);

NAND2xp5_ASAP7_75t_L g4407 ( 
.A(n_4367),
.B(n_4201),
.Y(n_4407)
);

OAI22xp5_ASAP7_75t_L g4408 ( 
.A1(n_4370),
.A2(n_4011),
.B1(n_4014),
.B2(n_4173),
.Y(n_4408)
);

INVx1_ASAP7_75t_L g4409 ( 
.A(n_4381),
.Y(n_4409)
);

INVx2_ASAP7_75t_SL g4410 ( 
.A(n_4374),
.Y(n_4410)
);

INVx1_ASAP7_75t_L g4411 ( 
.A(n_4381),
.Y(n_4411)
);

INVx2_ASAP7_75t_L g4412 ( 
.A(n_4374),
.Y(n_4412)
);

AND2x2_ASAP7_75t_L g4413 ( 
.A(n_4385),
.B(n_4134),
.Y(n_4413)
);

NAND2xp33_ASAP7_75t_SL g4414 ( 
.A(n_4383),
.B(n_4201),
.Y(n_4414)
);

NAND2xp5_ASAP7_75t_L g4415 ( 
.A(n_4413),
.B(n_4382),
.Y(n_4415)
);

AOI211x1_ASAP7_75t_L g4416 ( 
.A1(n_4408),
.A2(n_4386),
.B(n_4366),
.C(n_4173),
.Y(n_4416)
);

INVx1_ASAP7_75t_L g4417 ( 
.A(n_4394),
.Y(n_4417)
);

INVx3_ASAP7_75t_L g4418 ( 
.A(n_4391),
.Y(n_4418)
);

AOI21xp5_ASAP7_75t_L g4419 ( 
.A1(n_4392),
.A2(n_4375),
.B(n_4205),
.Y(n_4419)
);

NOR2x1_ASAP7_75t_L g4420 ( 
.A(n_4400),
.B(n_4203),
.Y(n_4420)
);

INVx1_ASAP7_75t_L g4421 ( 
.A(n_4396),
.Y(n_4421)
);

OAI22xp33_ASAP7_75t_L g4422 ( 
.A1(n_4407),
.A2(n_4393),
.B1(n_4403),
.B2(n_4203),
.Y(n_4422)
);

NAND2xp5_ASAP7_75t_L g4423 ( 
.A(n_4405),
.B(n_4203),
.Y(n_4423)
);

NOR2x1_ASAP7_75t_L g4424 ( 
.A(n_4401),
.B(n_4205),
.Y(n_4424)
);

INVx1_ASAP7_75t_L g4425 ( 
.A(n_4395),
.Y(n_4425)
);

AOI21xp5_ASAP7_75t_L g4426 ( 
.A1(n_4406),
.A2(n_4205),
.B(n_4167),
.Y(n_4426)
);

OA22x2_ASAP7_75t_L g4427 ( 
.A1(n_4397),
.A2(n_4165),
.B1(n_4167),
.B2(n_4170),
.Y(n_4427)
);

OAI21xp33_ASAP7_75t_SL g4428 ( 
.A1(n_4402),
.A2(n_4206),
.B(n_4198),
.Y(n_4428)
);

CKINVDCx5p33_ASAP7_75t_R g4429 ( 
.A(n_4399),
.Y(n_4429)
);

OAI22xp5_ASAP7_75t_L g4430 ( 
.A1(n_4404),
.A2(n_4165),
.B1(n_4167),
.B2(n_4170),
.Y(n_4430)
);

OAI222xp33_ASAP7_75t_L g4431 ( 
.A1(n_4410),
.A2(n_4165),
.B1(n_4170),
.B2(n_4197),
.C1(n_4196),
.C2(n_4195),
.Y(n_4431)
);

INVx1_ASAP7_75t_L g4432 ( 
.A(n_4427),
.Y(n_4432)
);

INVx2_ASAP7_75t_SL g4433 ( 
.A(n_4420),
.Y(n_4433)
);

O2A1O1Ixp33_ASAP7_75t_SL g4434 ( 
.A1(n_4431),
.A2(n_4430),
.B(n_4422),
.C(n_4423),
.Y(n_4434)
);

INVx2_ASAP7_75t_L g4435 ( 
.A(n_4418),
.Y(n_4435)
);

INVx1_ASAP7_75t_SL g4436 ( 
.A(n_4415),
.Y(n_4436)
);

OAI21xp5_ASAP7_75t_L g4437 ( 
.A1(n_4419),
.A2(n_4398),
.B(n_4399),
.Y(n_4437)
);

AOI211xp5_ASAP7_75t_SL g4438 ( 
.A1(n_4417),
.A2(n_4409),
.B(n_4411),
.C(n_4412),
.Y(n_4438)
);

AOI21xp33_ASAP7_75t_L g4439 ( 
.A1(n_4429),
.A2(n_4195),
.B(n_4206),
.Y(n_4439)
);

AOI21xp33_ASAP7_75t_L g4440 ( 
.A1(n_4425),
.A2(n_4198),
.B(n_4197),
.Y(n_4440)
);

OAI21xp5_ASAP7_75t_SL g4441 ( 
.A1(n_4421),
.A2(n_4196),
.B(n_4194),
.Y(n_4441)
);

INVx1_ASAP7_75t_L g4442 ( 
.A(n_4424),
.Y(n_4442)
);

AOI211xp5_ASAP7_75t_L g4443 ( 
.A1(n_4428),
.A2(n_4426),
.B(n_4414),
.C(n_4194),
.Y(n_4443)
);

XOR2x2_ASAP7_75t_L g4444 ( 
.A(n_4416),
.B(n_4063),
.Y(n_4444)
);

INVx1_ASAP7_75t_L g4445 ( 
.A(n_4427),
.Y(n_4445)
);

AOI321xp33_ASAP7_75t_L g4446 ( 
.A1(n_4417),
.A2(n_4153),
.A3(n_4148),
.B1(n_4151),
.B2(n_4149),
.C(n_4036),
.Y(n_4446)
);

AOI221xp5_ASAP7_75t_L g4447 ( 
.A1(n_4439),
.A2(n_4153),
.B1(n_4151),
.B2(n_4149),
.C(n_4148),
.Y(n_4447)
);

AOI22xp5_ASAP7_75t_L g4448 ( 
.A1(n_4435),
.A2(n_4051),
.B1(n_4053),
.B2(n_4014),
.Y(n_4448)
);

AOI22xp5_ASAP7_75t_L g4449 ( 
.A1(n_4436),
.A2(n_4051),
.B1(n_4053),
.B2(n_4011),
.Y(n_4449)
);

AOI21xp33_ASAP7_75t_L g4450 ( 
.A1(n_4433),
.A2(n_4437),
.B(n_4442),
.Y(n_4450)
);

OAI21x1_ASAP7_75t_SL g4451 ( 
.A1(n_4441),
.A2(n_4038),
.B(n_4036),
.Y(n_4451)
);

AOI22xp5_ASAP7_75t_L g4452 ( 
.A1(n_4444),
.A2(n_4041),
.B1(n_4038),
.B2(n_4103),
.Y(n_4452)
);

NOR3xp33_ASAP7_75t_L g4453 ( 
.A(n_4434),
.B(n_4077),
.C(n_4041),
.Y(n_4453)
);

INVx1_ASAP7_75t_SL g4454 ( 
.A(n_4440),
.Y(n_4454)
);

AOI33xp33_ASAP7_75t_L g4455 ( 
.A1(n_4432),
.A2(n_4146),
.A3(n_4124),
.B1(n_4114),
.B2(n_4088),
.B3(n_4073),
.Y(n_4455)
);

AOI221xp5_ASAP7_75t_L g4456 ( 
.A1(n_4445),
.A2(n_4146),
.B1(n_4124),
.B2(n_4114),
.C(n_4067),
.Y(n_4456)
);

OAI211xp5_ASAP7_75t_L g4457 ( 
.A1(n_4443),
.A2(n_4145),
.B(n_4147),
.C(n_4073),
.Y(n_4457)
);

NOR3xp33_ASAP7_75t_L g4458 ( 
.A(n_4438),
.B(n_4145),
.C(n_4094),
.Y(n_4458)
);

AOI22xp5_ASAP7_75t_L g4459 ( 
.A1(n_4446),
.A2(n_4124),
.B1(n_4146),
.B2(n_4067),
.Y(n_4459)
);

AOI221xp5_ASAP7_75t_L g4460 ( 
.A1(n_4439),
.A2(n_4146),
.B1(n_4124),
.B2(n_4067),
.C(n_4039),
.Y(n_4460)
);

AOI22xp33_ASAP7_75t_SL g4461 ( 
.A1(n_4435),
.A2(n_4071),
.B1(n_4054),
.B2(n_4092),
.Y(n_4461)
);

NAND2x1_ASAP7_75t_L g4462 ( 
.A(n_4442),
.B(n_4127),
.Y(n_4462)
);

OAI222xp33_ASAP7_75t_L g4463 ( 
.A1(n_4436),
.A2(n_4090),
.B1(n_4147),
.B2(n_4058),
.C1(n_4019),
.C2(n_4022),
.Y(n_4463)
);

INVx1_ASAP7_75t_L g4464 ( 
.A(n_4446),
.Y(n_4464)
);

INVx1_ASAP7_75t_L g4465 ( 
.A(n_4462),
.Y(n_4465)
);

NOR2xp67_ASAP7_75t_L g4466 ( 
.A(n_4459),
.B(n_4076),
.Y(n_4466)
);

NOR2x1_ASAP7_75t_L g4467 ( 
.A(n_4464),
.B(n_4090),
.Y(n_4467)
);

NAND4xp75_ASAP7_75t_L g4468 ( 
.A(n_4450),
.B(n_4071),
.C(n_4054),
.D(n_4135),
.Y(n_4468)
);

INVx1_ASAP7_75t_SL g4469 ( 
.A(n_4454),
.Y(n_4469)
);

OAI22x1_ASAP7_75t_L g4470 ( 
.A1(n_4449),
.A2(n_4058),
.B1(n_4074),
.B2(n_4127),
.Y(n_4470)
);

AOI21x1_ASAP7_75t_L g4471 ( 
.A1(n_4451),
.A2(n_4127),
.B(n_4132),
.Y(n_4471)
);

NAND3xp33_ASAP7_75t_L g4472 ( 
.A(n_4453),
.B(n_4039),
.C(n_4037),
.Y(n_4472)
);

AND4x1_ASAP7_75t_L g4473 ( 
.A(n_4458),
.B(n_3960),
.C(n_4134),
.D(n_4135),
.Y(n_4473)
);

INVx1_ASAP7_75t_L g4474 ( 
.A(n_4448),
.Y(n_4474)
);

AOI22xp5_ASAP7_75t_L g4475 ( 
.A1(n_4452),
.A2(n_4132),
.B1(n_4019),
.B2(n_4022),
.Y(n_4475)
);

INVx1_ASAP7_75t_L g4476 ( 
.A(n_4457),
.Y(n_4476)
);

NOR4xp25_ASAP7_75t_L g4477 ( 
.A(n_4447),
.B(n_4046),
.C(n_4045),
.D(n_4033),
.Y(n_4477)
);

NOR2x1_ASAP7_75t_L g4478 ( 
.A(n_4463),
.B(n_4090),
.Y(n_4478)
);

NAND2xp5_ASAP7_75t_L g4479 ( 
.A(n_4461),
.B(n_4069),
.Y(n_4479)
);

AND2x4_ASAP7_75t_L g4480 ( 
.A(n_4460),
.B(n_4132),
.Y(n_4480)
);

INVxp67_ASAP7_75t_L g4481 ( 
.A(n_4456),
.Y(n_4481)
);

OAI21xp5_ASAP7_75t_L g4482 ( 
.A1(n_4466),
.A2(n_4455),
.B(n_4093),
.Y(n_4482)
);

AOI21xp33_ASAP7_75t_L g4483 ( 
.A1(n_4465),
.A2(n_4027),
.B(n_4056),
.Y(n_4483)
);

AOI221xp5_ASAP7_75t_L g4484 ( 
.A1(n_4480),
.A2(n_4132),
.B1(n_4023),
.B2(n_4066),
.C(n_4057),
.Y(n_4484)
);

NAND4xp25_ASAP7_75t_SL g4485 ( 
.A(n_4467),
.B(n_4093),
.C(n_4091),
.D(n_4155),
.Y(n_4485)
);

NOR3x1_ASAP7_75t_SL g4486 ( 
.A(n_4481),
.B(n_4074),
.C(n_4091),
.Y(n_4486)
);

NOR3xp33_ASAP7_75t_L g4487 ( 
.A(n_4476),
.B(n_4474),
.C(n_4469),
.Y(n_4487)
);

NAND2xp5_ASAP7_75t_L g4488 ( 
.A(n_4468),
.B(n_4480),
.Y(n_4488)
);

AOI211xp5_ASAP7_75t_L g4489 ( 
.A1(n_4479),
.A2(n_4155),
.B(n_4074),
.C(n_3959),
.Y(n_4489)
);

NAND2xp5_ASAP7_75t_SL g4490 ( 
.A(n_4478),
.B(n_4049),
.Y(n_4490)
);

NOR5xp2_ASAP7_75t_L g4491 ( 
.A(n_4472),
.B(n_4089),
.C(n_4095),
.D(n_3967),
.E(n_3952),
.Y(n_4491)
);

NAND2xp5_ASAP7_75t_L g4492 ( 
.A(n_4477),
.B(n_4034),
.Y(n_4492)
);

INVxp67_ASAP7_75t_L g4493 ( 
.A(n_4488),
.Y(n_4493)
);

NOR2x1_ASAP7_75t_L g4494 ( 
.A(n_4490),
.B(n_4471),
.Y(n_4494)
);

AOI31xp33_ASAP7_75t_L g4495 ( 
.A1(n_4482),
.A2(n_4475),
.A3(n_4473),
.B(n_4470),
.Y(n_4495)
);

AND2x2_ASAP7_75t_L g4496 ( 
.A(n_4487),
.B(n_4492),
.Y(n_4496)
);

INVx2_ASAP7_75t_SL g4497 ( 
.A(n_4486),
.Y(n_4497)
);

AND2x4_ASAP7_75t_L g4498 ( 
.A(n_4483),
.B(n_4018),
.Y(n_4498)
);

NOR4xp25_ASAP7_75t_SL g4499 ( 
.A(n_4494),
.B(n_4484),
.C(n_4485),
.D(n_4491),
.Y(n_4499)
);

NOR4xp25_ASAP7_75t_L g4500 ( 
.A(n_4497),
.B(n_4495),
.C(n_4493),
.D(n_4496),
.Y(n_4500)
);

NOR3xp33_ASAP7_75t_L g4501 ( 
.A(n_4498),
.B(n_4489),
.C(n_4082),
.Y(n_4501)
);

AOI22xp5_ASAP7_75t_L g4502 ( 
.A1(n_4501),
.A2(n_4500),
.B1(n_4499),
.B2(n_4012),
.Y(n_4502)
);

AOI22xp33_ASAP7_75t_L g4503 ( 
.A1(n_4501),
.A2(n_4062),
.B1(n_4015),
.B2(n_4032),
.Y(n_4503)
);

INVx1_ASAP7_75t_L g4504 ( 
.A(n_4502),
.Y(n_4504)
);

AOI22xp5_ASAP7_75t_L g4505 ( 
.A1(n_4504),
.A2(n_4503),
.B1(n_4062),
.B2(n_4015),
.Y(n_4505)
);

NOR2x1_ASAP7_75t_L g4506 ( 
.A(n_4505),
.B(n_4096),
.Y(n_4506)
);

NOR3xp33_ASAP7_75t_L g4507 ( 
.A(n_4506),
.B(n_3937),
.C(n_3971),
.Y(n_4507)
);

INVx1_ASAP7_75t_L g4508 ( 
.A(n_4507),
.Y(n_4508)
);

NAND4xp25_ASAP7_75t_L g4509 ( 
.A(n_4508),
.B(n_3973),
.C(n_3945),
.D(n_3908),
.Y(n_4509)
);

AOI21xp33_ASAP7_75t_SL g4510 ( 
.A1(n_4509),
.A2(n_4099),
.B(n_410),
.Y(n_4510)
);

NAND2xp5_ASAP7_75t_SL g4511 ( 
.A(n_4510),
.B(n_4062),
.Y(n_4511)
);

NAND3xp33_ASAP7_75t_L g4512 ( 
.A(n_4511),
.B(n_3908),
.C(n_3978),
.Y(n_4512)
);

OAI22xp5_ASAP7_75t_L g4513 ( 
.A1(n_4512),
.A2(n_4043),
.B1(n_4085),
.B2(n_4018),
.Y(n_4513)
);

NAND2xp5_ASAP7_75t_L g4514 ( 
.A(n_4512),
.B(n_4034),
.Y(n_4514)
);

INVxp67_ASAP7_75t_L g4515 ( 
.A(n_4514),
.Y(n_4515)
);

INVx1_ASAP7_75t_L g4516 ( 
.A(n_4513),
.Y(n_4516)
);

OA21x2_ASAP7_75t_L g4517 ( 
.A1(n_4516),
.A2(n_4042),
.B(n_4032),
.Y(n_4517)
);

OA21x2_ASAP7_75t_L g4518 ( 
.A1(n_4515),
.A2(n_4042),
.B(n_4085),
.Y(n_4518)
);

AOI221xp5_ASAP7_75t_L g4519 ( 
.A1(n_4517),
.A2(n_3922),
.B1(n_4099),
.B2(n_4096),
.C(n_3997),
.Y(n_4519)
);

AOI22xp5_ASAP7_75t_L g4520 ( 
.A1(n_4519),
.A2(n_4518),
.B1(n_4099),
.B2(n_4084),
.Y(n_4520)
);

AOI211xp5_ASAP7_75t_L g4521 ( 
.A1(n_4520),
.A2(n_3977),
.B(n_3975),
.C(n_3980),
.Y(n_4521)
);


endmodule