module fake_jpeg_3136_n_307 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_307);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_307;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_208;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx5_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_9),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx6_ASAP7_75t_SL g39 ( 
.A(n_9),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_2),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_15),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g133 ( 
.A(n_44),
.Y(n_133)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_46),
.Y(n_90)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g130 ( 
.A(n_47),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_35),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_48),
.B(n_55),
.Y(n_98)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g102 ( 
.A(n_51),
.Y(n_102)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_28),
.Y(n_53)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_53),
.Y(n_87)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_21),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_35),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_30),
.A2(n_15),
.B1(n_4),
.B2(n_5),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_57),
.A2(n_41),
.B1(n_38),
.B2(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_17),
.B(n_10),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_58),
.B(n_64),
.Y(n_105)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_59),
.Y(n_107)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_40),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_62),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_19),
.B(n_10),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_40),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_65),
.B(n_68),
.Y(n_115)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_66),
.Y(n_113)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_67),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_21),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_71),
.B(n_78),
.Y(n_92)
);

BUFx12f_ASAP7_75t_SL g72 ( 
.A(n_19),
.Y(n_72)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_29),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_26),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_73),
.B(n_76),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_26),
.B(n_31),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_74),
.B(n_75),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_33),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_33),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_17),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_79),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_16),
.Y(n_79)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_21),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_80),
.A2(n_83),
.B1(n_43),
.B2(n_23),
.Y(n_91)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_43),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_16),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_23),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_43),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_84),
.Y(n_104)
);

OAI21xp33_ASAP7_75t_L g85 ( 
.A1(n_72),
.A2(n_42),
.B(n_37),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_85),
.A2(n_13),
.B(n_123),
.Y(n_156)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_86),
.B(n_84),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_88),
.B(n_94),
.C(n_96),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g155 ( 
.A1(n_91),
.A2(n_47),
.B1(n_12),
.B2(n_13),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_81),
.A2(n_42),
.B1(n_37),
.B2(n_34),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_95),
.A2(n_118),
.B1(n_121),
.B2(n_124),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_53),
.B(n_20),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_29),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_97),
.B(n_116),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_48),
.A2(n_20),
.B1(n_34),
.B2(n_24),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g150 ( 
.A1(n_99),
.A2(n_111),
.B1(n_127),
.B2(n_133),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_110),
.A2(n_122),
.B1(n_126),
.B2(n_54),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_55),
.A2(n_24),
.B1(n_38),
.B2(n_36),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_78),
.B(n_25),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g118 ( 
.A1(n_79),
.A2(n_82),
.B1(n_62),
.B2(n_61),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_65),
.A2(n_25),
.B1(n_22),
.B2(n_41),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_46),
.A2(n_10),
.B1(n_6),
.B2(n_7),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_77),
.B(n_1),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_123),
.B(n_131),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_73),
.A2(n_76),
.B1(n_63),
.B2(n_50),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_56),
.A2(n_1),
.B(n_6),
.Y(n_125)
);

O2A1O1Ixp33_ASAP7_75t_SL g138 ( 
.A1(n_125),
.A2(n_67),
.B(n_51),
.C(n_83),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_52),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_49),
.A2(n_7),
.B1(n_8),
.B2(n_11),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_70),
.B(n_8),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_60),
.B(n_12),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_12),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_117),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_134),
.B(n_147),
.Y(n_192)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_135),
.B(n_136),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_71),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_137),
.A2(n_150),
.B1(n_173),
.B2(n_133),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_138),
.A2(n_156),
.B(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_120),
.B(n_83),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_142),
.B(n_151),
.Y(n_177)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_89),
.Y(n_143)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_143),
.Y(n_194)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_144),
.Y(n_175)
);

BUFx12_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_145),
.Y(n_180)
);

HB1xp67_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_146),
.Y(n_183)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_148),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_87),
.B(n_69),
.C(n_71),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_103),
.C(n_102),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_128),
.B(n_45),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_90),
.Y(n_152)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_152),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_97),
.A2(n_80),
.B1(n_66),
.B2(n_44),
.Y(n_154)
);

OR2x2_ASAP7_75t_L g191 ( 
.A(n_154),
.B(n_155),
.Y(n_191)
);

OAI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_116),
.A2(n_96),
.B1(n_125),
.B2(n_88),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_157),
.A2(n_139),
.B1(n_141),
.B2(n_153),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_98),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_160),
.Y(n_179)
);

OR2x4_ASAP7_75t_L g159 ( 
.A(n_85),
.B(n_131),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_159),
.A2(n_172),
.B(n_155),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_105),
.B(n_107),
.Y(n_160)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_161),
.Y(n_206)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_130),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_162),
.B(n_166),
.Y(n_182)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_106),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_126),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_122),
.A2(n_92),
.B1(n_104),
.B2(n_113),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_100),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_112),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_169),
.Y(n_199)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_95),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_168),
.B(n_170),
.Y(n_181)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_109),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_92),
.B(n_109),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_92),
.B(n_113),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_101),
.Y(n_172)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_103),
.A2(n_133),
.B1(n_101),
.B2(n_100),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_114),
.Y(n_174)
);

NOR3xp33_ASAP7_75t_SL g189 ( 
.A(n_174),
.B(n_130),
.C(n_108),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_186),
.A2(n_187),
.B1(n_193),
.B2(n_195),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_164),
.A2(n_119),
.B1(n_114),
.B2(n_108),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_188),
.B(n_190),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g213 ( 
.A(n_189),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_141),
.B(n_93),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_137),
.A2(n_119),
.B1(n_90),
.B2(n_93),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_139),
.A2(n_165),
.B1(n_168),
.B2(n_159),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_136),
.A2(n_138),
.B(n_135),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_196),
.A2(n_203),
.B(n_145),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_155),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_135),
.A2(n_136),
.B1(n_154),
.B2(n_147),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_200),
.A2(n_201),
.B1(n_152),
.B2(n_162),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_171),
.A2(n_140),
.B1(n_170),
.B2(n_163),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_149),
.B(n_156),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g211 ( 
.A(n_202),
.B(n_155),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_161),
.B(n_167),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_143),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_207),
.B(n_216),
.Y(n_234)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_204),
.Y(n_208)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_208),
.Y(n_237)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_199),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_211),
.B(n_197),
.C(n_198),
.Y(n_243)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_206),
.Y(n_212)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_212),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_183),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_148),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_217),
.Y(n_235)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_206),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_218),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g245 ( 
.A(n_219),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_196),
.A2(n_145),
.B1(n_176),
.B2(n_181),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_220),
.A2(n_226),
.B1(n_227),
.B2(n_228),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_221),
.Y(n_246)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_222),
.B(n_225),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_203),
.A2(n_181),
.B(n_195),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_230),
.B(n_178),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_182),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_224),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_179),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_191),
.A2(n_184),
.B1(n_201),
.B2(n_178),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_192),
.B(n_175),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_205),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_229),
.A2(n_218),
.B1(n_212),
.B2(n_227),
.Y(n_249)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_191),
.B1(n_184),
.B2(n_178),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_226),
.B1(n_211),
.B2(n_220),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_SL g260 ( 
.A1(n_233),
.A2(n_236),
.B(n_238),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_221),
.A2(n_200),
.B(n_202),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_223),
.A2(n_188),
.B(n_177),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_210),
.B(n_190),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_240),
.B(n_243),
.C(n_216),
.Y(n_254)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_249),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_250),
.A2(n_238),
.B1(n_232),
.B2(n_243),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_247),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_251),
.B(n_253),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_240),
.B(n_210),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_252),
.B(n_254),
.C(n_261),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_248),
.B(n_175),
.Y(n_253)
);

AND2x2_ASAP7_75t_L g255 ( 
.A(n_248),
.B(n_224),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g269 ( 
.A(n_255),
.B(n_262),
.Y(n_269)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_247),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_256),
.B(n_258),
.Y(n_274)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_249),
.Y(n_258)
);

CKINVDCx16_ASAP7_75t_R g259 ( 
.A(n_233),
.Y(n_259)
);

BUFx2_ASAP7_75t_L g276 ( 
.A(n_259),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_240),
.B(n_208),
.C(n_209),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_239),
.Y(n_262)
);

AOI322xp5_ASAP7_75t_L g263 ( 
.A1(n_235),
.A2(n_207),
.A3(n_177),
.B1(n_198),
.B2(n_213),
.C1(n_193),
.C2(n_187),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_263),
.A2(n_231),
.B(n_244),
.Y(n_273)
);

OAI22xp33_ASAP7_75t_L g264 ( 
.A1(n_245),
.A2(n_189),
.B1(n_185),
.B2(n_222),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_264),
.A2(n_231),
.B1(n_244),
.B2(n_241),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_237),
.Y(n_265)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_265),
.A2(n_234),
.B(n_237),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_266),
.A2(n_272),
.B1(n_273),
.B2(n_274),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_250),
.A2(n_246),
.B(n_236),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_265),
.B(n_262),
.Y(n_282)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_241),
.C(n_180),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_275),
.B(n_261),
.C(n_255),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_273),
.A2(n_258),
.B1(n_257),
.B2(n_260),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_277),
.A2(n_279),
.B1(n_285),
.B2(n_276),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_254),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_278),
.B(n_280),
.Y(n_287)
);

OAI22x1_ASAP7_75t_SL g279 ( 
.A1(n_272),
.A2(n_257),
.B1(n_255),
.B2(n_264),
.Y(n_279)
);

MAJx2_ASAP7_75t_L g290 ( 
.A(n_282),
.B(n_276),
.C(n_275),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_283),
.A2(n_281),
.B1(n_269),
.B2(n_279),
.Y(n_286)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_284),
.Y(n_292)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_269),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_289),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g288 ( 
.A1(n_282),
.A2(n_267),
.B(n_269),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_288),
.A2(n_229),
.B(n_185),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_290),
.B(n_291),
.C(n_242),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_242),
.B1(n_268),
.B2(n_180),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_287),
.B(n_278),
.C(n_280),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_293),
.B(n_294),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g299 ( 
.A(n_295),
.B(n_297),
.Y(n_299)
);

INVx11_ASAP7_75t_L g297 ( 
.A(n_286),
.Y(n_297)
);

OAI21x1_ASAP7_75t_SL g298 ( 
.A1(n_296),
.A2(n_292),
.B(n_290),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_298),
.B(n_301),
.Y(n_302)
);

AOI211xp5_ASAP7_75t_L g301 ( 
.A1(n_297),
.A2(n_291),
.B(n_183),
.C(n_230),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_L g305 ( 
.A1(n_303),
.A2(n_293),
.B(n_301),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_302),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_304),
.B(n_305),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_306),
.B(n_302),
.Y(n_307)
);


endmodule