module fake_ibex_1833_n_22 (n_3, n_1, n_5, n_4, n_2, n_0, n_6, n_22);

input n_3;
input n_1;
input n_5;
input n_4;
input n_2;
input n_0;
input n_6;

output n_22;



endmodule