module fake_jpeg_12116_n_496 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_496);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_496;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_490;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_16),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx14_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_SL g32 ( 
.A(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_1),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_3),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_13),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_49),
.Y(n_118)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_18),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_51),
.Y(n_133)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

INVx2_ASAP7_75t_SL g108 ( 
.A(n_53),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_20),
.B(n_16),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_54),
.B(n_63),
.Y(n_129)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_48),
.Y(n_55)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_55),
.Y(n_140)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g116 ( 
.A(n_56),
.Y(n_116)
);

BUFx5_ASAP7_75t_L g57 ( 
.A(n_31),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g142 ( 
.A(n_57),
.Y(n_142)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_58),
.Y(n_107)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_59),
.Y(n_104)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_60),
.Y(n_120)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_61),
.Y(n_109)
);

BUFx16f_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVxp67_ASAP7_75t_SL g148 ( 
.A(n_62),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_20),
.B(n_16),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g141 ( 
.A(n_64),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_18),
.Y(n_65)
);

INVx6_ASAP7_75t_L g153 ( 
.A(n_65),
.Y(n_153)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_66),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_67),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx8_ASAP7_75t_L g135 ( 
.A(n_68),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_69),
.Y(n_106)
);

INVx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g124 ( 
.A(n_70),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_71),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_72),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_32),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_80),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_30),
.Y(n_74)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_74),
.Y(n_139)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_75),
.Y(n_125)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_36),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_40),
.Y(n_77)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_77),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_78),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_79),
.Y(n_146)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_27),
.B(n_15),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_28),
.Y(n_81)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_81),
.Y(n_122)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_82),
.Y(n_136)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_40),
.Y(n_83)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_30),
.Y(n_84)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_93),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_42),
.Y(n_86)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_32),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_87),
.B(n_89),
.Y(n_111)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_88),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_24),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_24),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_39),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_39),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_92),
.B(n_94),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_42),
.Y(n_93)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_42),
.Y(n_94)
);

BUFx4f_ASAP7_75t_SL g95 ( 
.A(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_95),
.B(n_96),
.Y(n_130)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_23),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_36),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_97),
.B(n_44),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_80),
.A2(n_41),
.B1(n_46),
.B2(n_42),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g175 ( 
.A1(n_98),
.A2(n_69),
.B1(n_68),
.B2(n_65),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_96),
.A2(n_23),
.B1(n_27),
.B2(n_46),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_99),
.A2(n_149),
.B1(n_74),
.B2(n_29),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_50),
.B(n_47),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_102),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_55),
.B(n_47),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_95),
.B(n_43),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_103),
.B(n_137),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_51),
.A2(n_41),
.B1(n_46),
.B2(n_22),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_105),
.A2(n_117),
.B1(n_152),
.B2(n_29),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_58),
.A2(n_41),
.B1(n_46),
.B2(n_27),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_64),
.B(n_38),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_126),
.B(n_128),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g127 ( 
.A(n_88),
.B(n_41),
.C(n_38),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_56),
.C(n_78),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_45),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_83),
.B(n_45),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_134),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_94),
.B(n_26),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g143 ( 
.A(n_95),
.B(n_44),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_19),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_53),
.A2(n_29),
.B1(n_43),
.B2(n_37),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_49),
.A2(n_37),
.B1(n_19),
.B2(n_26),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_62),
.B(n_25),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_155),
.B(n_84),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_156),
.B(n_184),
.Y(n_236)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_131),
.Y(n_158)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_158),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_170),
.Y(n_229)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_161),
.Y(n_223)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_101),
.Y(n_163)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_163),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_118),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_165),
.A2(n_212),
.B1(n_151),
.B2(n_124),
.Y(n_217)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_109),
.Y(n_166)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_166),
.Y(n_225)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_167),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_78),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_179),
.C(n_204),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_169),
.Y(n_227)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_98),
.A2(n_70),
.B1(n_21),
.B2(n_25),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_171),
.Y(n_230)
);

AO22x2_ASAP7_75t_L g172 ( 
.A1(n_107),
.A2(n_93),
.B1(n_86),
.B2(n_85),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_172),
.B(n_200),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_129),
.B(n_21),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_173),
.B(n_178),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_102),
.A2(n_79),
.B1(n_72),
.B2(n_71),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_174),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g216 ( 
.A1(n_175),
.A2(n_182),
.B1(n_191),
.B2(n_105),
.Y(n_216)
);

FAx1_ASAP7_75t_SL g176 ( 
.A(n_126),
.B(n_14),
.CI(n_13),
.CON(n_176),
.SN(n_176)
);

A2O1A1Ixp33_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_187),
.B(n_189),
.C(n_167),
.Y(n_214)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_119),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_130),
.B(n_12),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_180),
.Y(n_244)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_124),
.Y(n_181)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_181),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_114),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_182)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

BUFx2_ASAP7_75t_L g248 ( 
.A(n_183),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_115),
.B(n_1),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_146),
.Y(n_185)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_185),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_111),
.B(n_2),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_186),
.B(n_196),
.Y(n_251)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_128),
.B(n_2),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_189),
.B(n_197),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_118),
.Y(n_190)
);

INVx4_ASAP7_75t_SL g222 ( 
.A(n_190),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_114),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_121),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_192),
.Y(n_226)
);

INVx13_ASAP7_75t_L g193 ( 
.A(n_148),
.Y(n_193)
);

BUFx24_ASAP7_75t_L g242 ( 
.A(n_193),
.Y(n_242)
);

INVx2_ASAP7_75t_SL g194 ( 
.A(n_150),
.Y(n_194)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_195),
.Y(n_258)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_153),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_154),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_104),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_198),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_110),
.B(n_3),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_199),
.B(n_203),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g200 ( 
.A(n_113),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_138),
.Y(n_201)
);

OR2x2_ASAP7_75t_L g256 ( 
.A(n_201),
.B(n_202),
.Y(n_256)
);

OR2x2_ASAP7_75t_SL g202 ( 
.A(n_104),
.B(n_4),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_120),
.B(n_125),
.Y(n_204)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_139),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_205),
.B(n_208),
.Y(n_241)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_122),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_206),
.B(n_9),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_127),
.B(n_4),
.C(n_5),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_207),
.B(n_6),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_120),
.B(n_5),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_136),
.B(n_6),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_209),
.B(n_211),
.Y(n_252)
);

BUFx24_ASAP7_75t_L g210 ( 
.A(n_108),
.Y(n_210)
);

O2A1O1Ixp33_ASAP7_75t_L g253 ( 
.A1(n_210),
.A2(n_116),
.B(n_141),
.C(n_140),
.Y(n_253)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_117),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_212)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_214),
.A2(n_193),
.B(n_172),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_216),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_217),
.A2(n_220),
.B1(n_245),
.B2(n_210),
.Y(n_262)
);

MAJx2_ASAP7_75t_L g218 ( 
.A(n_157),
.B(n_138),
.C(n_108),
.Y(n_218)
);

A2O1A1O1Ixp25_ASAP7_75t_L g279 ( 
.A1(n_218),
.A2(n_260),
.B(n_213),
.C(n_219),
.D(n_241),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_195),
.A2(n_107),
.B1(n_153),
.B2(n_133),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_159),
.A2(n_133),
.B1(n_124),
.B2(n_135),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_221),
.A2(n_228),
.B1(n_237),
.B2(n_243),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_159),
.A2(n_135),
.B1(n_144),
.B2(n_106),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g237 ( 
.A1(n_187),
.A2(n_144),
.B1(n_123),
.B2(n_106),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_157),
.A2(n_123),
.B1(n_108),
.B2(n_116),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_156),
.A2(n_116),
.B1(n_141),
.B2(n_140),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_247),
.B(n_211),
.Y(n_288)
);

AO21x1_ASAP7_75t_SL g306 ( 
.A1(n_253),
.A2(n_215),
.B(n_225),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_207),
.A2(n_147),
.B1(n_142),
.B2(n_9),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_254),
.A2(n_255),
.B1(n_181),
.B2(n_190),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_168),
.A2(n_147),
.B1(n_142),
.B2(n_9),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_179),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_259),
.A2(n_210),
.B(n_179),
.Y(n_266)
);

MAJx2_ASAP7_75t_L g260 ( 
.A(n_202),
.B(n_7),
.C(n_8),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_261),
.B(n_208),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_L g313 ( 
.A1(n_262),
.A2(n_303),
.B1(n_304),
.B2(n_306),
.Y(n_313)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_223),
.Y(n_263)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_263),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_226),
.B(n_162),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g341 ( 
.A(n_264),
.B(n_272),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_265),
.B(n_274),
.Y(n_326)
);

INVxp67_ASAP7_75t_L g334 ( 
.A(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_223),
.Y(n_267)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_267),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_242),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_268),
.B(n_276),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g270 ( 
.A1(n_227),
.A2(n_176),
.B(n_205),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_229),
.B(n_176),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_SL g273 ( 
.A1(n_250),
.A2(n_172),
.B1(n_161),
.B2(n_194),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_273),
.A2(n_293),
.B1(n_228),
.B2(n_237),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_231),
.B(n_197),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_257),
.Y(n_275)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_275),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_242),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_241),
.B(n_204),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_277),
.B(n_280),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_256),
.A2(n_204),
.B(n_194),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_278),
.B(n_291),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g328 ( 
.A(n_279),
.B(n_288),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_242),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_257),
.Y(n_281)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_281),
.Y(n_312)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_261),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_282),
.B(n_284),
.Y(n_319)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_235),
.Y(n_283)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_283),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_233),
.Y(n_284)
);

BUFx2_ASAP7_75t_L g285 ( 
.A(n_246),
.Y(n_285)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_285),
.Y(n_345)
);

OAI32xp33_ASAP7_75t_L g286 ( 
.A1(n_214),
.A2(n_198),
.A3(n_177),
.B1(n_158),
.B2(n_180),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_290),
.Y(n_329)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_231),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_287),
.A2(n_259),
.B1(n_248),
.B2(n_249),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_289),
.A2(n_294),
.B1(n_302),
.B2(n_217),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_188),
.Y(n_290)
);

A2O1A1O1Ixp25_ASAP7_75t_L g292 ( 
.A1(n_213),
.A2(n_256),
.B(n_258),
.C(n_234),
.D(n_218),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_300),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_250),
.A2(n_172),
.B1(n_196),
.B2(n_185),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_239),
.A2(n_183),
.B1(n_164),
.B2(n_12),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_235),
.Y(n_295)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_295),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_251),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_296),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g297 ( 
.A(n_246),
.Y(n_297)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_297),
.Y(n_344)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_238),
.Y(n_298)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_298),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_SL g299 ( 
.A1(n_260),
.A2(n_11),
.B(n_12),
.Y(n_299)
);

AOI22x1_ASAP7_75t_L g321 ( 
.A1(n_299),
.A2(n_255),
.B1(n_254),
.B2(n_236),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_236),
.A2(n_230),
.B(n_227),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_238),
.Y(n_301)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_301),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_240),
.B(n_234),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_232),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_236),
.A2(n_230),
.B(n_239),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_305),
.B(n_300),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_316),
.A2(n_325),
.B1(n_342),
.B2(n_262),
.Y(n_355)
);

CKINVDCx20_ASAP7_75t_R g318 ( 
.A(n_284),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_318),
.B(n_332),
.Y(n_351)
);

OA22x2_ASAP7_75t_L g374 ( 
.A1(n_320),
.A2(n_295),
.B1(n_301),
.B2(n_283),
.Y(n_374)
);

CKINVDCx16_ASAP7_75t_R g346 ( 
.A(n_321),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_288),
.B(n_258),
.C(n_247),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_322),
.B(n_327),
.C(n_333),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_324),
.B(n_299),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_L g325 ( 
.A1(n_269),
.A2(n_252),
.B1(n_220),
.B2(n_245),
.Y(n_325)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_252),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_268),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_292),
.B(n_251),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_269),
.A2(n_221),
.B1(n_251),
.B2(n_253),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_336),
.A2(n_289),
.B1(n_294),
.B2(n_275),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_SL g373 ( 
.A(n_337),
.B(n_285),
.Y(n_373)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_280),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_338),
.B(n_339),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_290),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_263),
.Y(n_340)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_340),
.B(n_281),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g342 ( 
.A1(n_271),
.A2(n_224),
.B1(n_248),
.B2(n_249),
.Y(n_342)
);

A2O1A1O1Ixp25_ASAP7_75t_L g347 ( 
.A1(n_328),
.A2(n_305),
.B(n_278),
.C(n_277),
.D(n_286),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g405 ( 
.A(n_347),
.B(n_372),
.Y(n_405)
);

INVx5_ASAP7_75t_L g348 ( 
.A(n_344),
.Y(n_348)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_348),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_314),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_349),
.B(n_353),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_328),
.B(n_327),
.C(n_315),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_352),
.B(n_375),
.C(n_378),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_310),
.A2(n_270),
.B(n_306),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_308),
.Y(n_354)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_354),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_355),
.A2(n_364),
.B1(n_366),
.B2(n_373),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_334),
.A2(n_309),
.B(n_311),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_SL g403 ( 
.A(n_356),
.B(n_349),
.Y(n_403)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_310),
.A2(n_276),
.B(n_296),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_358),
.Y(n_395)
);

AOI21xp5_ASAP7_75t_L g358 ( 
.A1(n_329),
.A2(n_266),
.B(n_271),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_308),
.Y(n_359)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_359),
.Y(n_379)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_312),
.Y(n_360)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_360),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_319),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_361),
.B(n_365),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_320),
.A2(n_329),
.B1(n_313),
.B2(n_336),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g401 ( 
.A1(n_363),
.A2(n_367),
.B1(n_345),
.B2(n_344),
.Y(n_401)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_307),
.A2(n_293),
.B1(n_273),
.B2(n_334),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_319),
.Y(n_365)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_311),
.A2(n_282),
.B1(n_272),
.B2(n_267),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_312),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_368),
.B(n_377),
.Y(n_381)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_369),
.Y(n_383)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_317),
.Y(n_370)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_370),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_304),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_SL g404 ( 
.A(n_371),
.B(n_222),
.Y(n_404)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_374),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_315),
.B(n_298),
.C(n_303),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_317),
.Y(n_376)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_376),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_324),
.A2(n_285),
.B(n_297),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_322),
.B(n_297),
.C(n_224),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_350),
.B(n_333),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_380),
.B(n_386),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_350),
.B(n_321),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_352),
.B(n_321),
.Y(n_388)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_388),
.B(n_358),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_375),
.B(n_330),
.C(n_331),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_389),
.B(n_399),
.C(n_377),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_351),
.B(n_326),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_390),
.B(n_402),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_346),
.A2(n_337),
.B1(n_323),
.B2(n_335),
.Y(n_393)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_393),
.A2(n_367),
.B1(n_363),
.B2(n_373),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_355),
.A2(n_323),
.B1(n_335),
.B2(n_343),
.Y(n_396)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_396),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g399 ( 
.A(n_378),
.B(n_343),
.C(n_345),
.Y(n_399)
);

HB1xp67_ASAP7_75t_L g414 ( 
.A(n_401),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_362),
.B(n_222),
.Y(n_402)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_403),
.A2(n_347),
.B(n_360),
.Y(n_428)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_404),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_361),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_406),
.B(n_365),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

XNOR2xp5_ASAP7_75t_L g411 ( 
.A(n_385),
.B(n_356),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_L g441 ( 
.A(n_411),
.B(n_413),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_385),
.B(n_357),
.Y(n_413)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_415),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_416),
.B(n_419),
.Y(n_437)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_417),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_426),
.C(n_405),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_353),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_398),
.Y(n_420)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_420),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_383),
.B(n_368),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_421),
.B(n_422),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_389),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_379),
.Y(n_423)
);

BUFx2_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g424 ( 
.A(n_388),
.B(n_372),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g444 ( 
.A(n_424),
.B(n_425),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_386),
.B(n_366),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_399),
.B(n_364),
.C(n_374),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_397),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_427),
.B(n_348),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_428),
.A2(n_395),
.B(n_384),
.Y(n_430)
);

INVx11_ASAP7_75t_L g429 ( 
.A(n_381),
.Y(n_429)
);

INVx13_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

XOR2x2_ASAP7_75t_L g450 ( 
.A(n_430),
.B(n_432),
.Y(n_450)
);

HAxp5_ASAP7_75t_SL g432 ( 
.A(n_429),
.B(n_395),
.CON(n_432),
.SN(n_432)
);

AOI22xp5_ASAP7_75t_SL g434 ( 
.A1(n_426),
.A2(n_391),
.B1(n_384),
.B2(n_392),
.Y(n_434)
);

OAI21xp33_ASAP7_75t_L g454 ( 
.A1(n_434),
.A2(n_439),
.B(n_425),
.Y(n_454)
);

AOI21xp33_ASAP7_75t_L g435 ( 
.A1(n_410),
.A2(n_409),
.B(n_428),
.Y(n_435)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_435),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_411),
.B(n_400),
.Y(n_436)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_436),
.B(n_442),
.Y(n_456)
);

AOI22xp5_ASAP7_75t_SL g439 ( 
.A1(n_414),
.A2(n_392),
.B1(n_393),
.B2(n_405),
.Y(n_439)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_407),
.B(n_401),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_443),
.B(n_415),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_418),
.C(n_412),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g449 ( 
.A(n_444),
.B(n_419),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g463 ( 
.A(n_449),
.B(n_454),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_451),
.B(n_430),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g452 ( 
.A(n_431),
.Y(n_452)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_452),
.Y(n_465)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_413),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g467 ( 
.A(n_453),
.B(n_459),
.Y(n_467)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_437),
.B(n_412),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_458),
.C(n_439),
.Y(n_468)
);

OAI21x1_ASAP7_75t_L g457 ( 
.A1(n_433),
.A2(n_374),
.B(n_424),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_457),
.B(n_445),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_437),
.B(n_444),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_441),
.B(n_416),
.C(n_374),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_461),
.B(n_462),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_L g462 ( 
.A1(n_447),
.A2(n_379),
.B(n_387),
.Y(n_462)
);

NOR2xp33_ASAP7_75t_L g464 ( 
.A(n_456),
.B(n_431),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_464),
.B(n_466),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g477 ( 
.A(n_468),
.B(n_469),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_452),
.B(n_438),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_438),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_471),
.B(n_472),
.C(n_473),
.Y(n_475)
);

OAI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_461),
.A2(n_434),
.B1(n_446),
.B2(n_445),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_450),
.B(n_446),
.Y(n_473)
);

A2O1A1Ixp33_ASAP7_75t_L g476 ( 
.A1(n_474),
.A2(n_450),
.B(n_432),
.C(n_440),
.Y(n_476)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_476),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_467),
.B(n_458),
.C(n_455),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_478),
.B(n_479),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_470),
.B(n_449),
.C(n_440),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_468),
.B(n_448),
.C(n_454),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_481),
.A2(n_482),
.B(n_477),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_472),
.B(n_448),
.C(n_382),
.Y(n_482)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_484),
.Y(n_489)
);

NOR2xp67_ASAP7_75t_L g486 ( 
.A(n_475),
.B(n_465),
.Y(n_486)
);

AOI21x1_ASAP7_75t_L g488 ( 
.A1(n_486),
.A2(n_487),
.B(n_463),
.Y(n_488)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_480),
.A2(n_474),
.B(n_463),
.Y(n_487)
);

A2O1A1O1Ixp25_ASAP7_75t_L g491 ( 
.A1(n_488),
.A2(n_485),
.B(n_394),
.C(n_370),
.D(n_376),
.Y(n_491)
);

OAI22xp5_ASAP7_75t_L g490 ( 
.A1(n_483),
.A2(n_448),
.B1(n_382),
.B2(n_387),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_490),
.B(n_394),
.C(n_354),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_491),
.B(n_492),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g494 ( 
.A(n_493),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_494),
.B(n_489),
.Y(n_495)
);

HAxp5_ASAP7_75t_SL g496 ( 
.A(n_495),
.B(n_359),
.CON(n_496),
.SN(n_496)
);


endmodule