module fake_netlist_6_1978_n_72 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_6, n_15, n_3, n_14, n_0, n_4, n_13, n_11, n_17, n_12, n_20, n_7, n_2, n_5, n_19, n_72);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_6;
input n_15;
input n_3;
input n_14;
input n_0;
input n_4;
input n_13;
input n_11;
input n_17;
input n_12;
input n_20;
input n_7;
input n_2;
input n_5;
input n_19;

output n_72;

wire n_41;
wire n_52;
wire n_45;
wire n_46;
wire n_34;
wire n_42;
wire n_70;
wire n_24;
wire n_71;
wire n_37;
wire n_33;
wire n_54;
wire n_67;
wire n_27;
wire n_38;
wire n_61;
wire n_39;
wire n_63;
wire n_60;
wire n_59;
wire n_32;
wire n_66;
wire n_36;
wire n_22;
wire n_26;
wire n_68;
wire n_55;
wire n_35;
wire n_28;
wire n_23;
wire n_58;
wire n_69;
wire n_50;
wire n_64;
wire n_30;
wire n_49;
wire n_43;
wire n_47;
wire n_48;
wire n_29;
wire n_62;
wire n_31;
wire n_65;
wire n_40;
wire n_57;
wire n_25;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_12),
.A2(n_15),
.B1(n_16),
.B2(n_19),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_7),
.B(n_5),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22x1_ASAP7_75t_SL g25 ( 
.A1(n_20),
.A2(n_0),
.B1(n_17),
.B2(n_21),
.Y(n_25)
);

OAI21x1_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_5),
.B(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_18),
.B(n_3),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

AND2x4_ASAP7_75t_L g35 ( 
.A(n_6),
.B(n_2),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_33),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_29),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_30),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

OAI21x1_ASAP7_75t_L g44 ( 
.A1(n_38),
.A2(n_26),
.B(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_33),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_33),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_43),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_39),
.Y(n_48)
);

OAI21x1_ASAP7_75t_L g49 ( 
.A1(n_44),
.A2(n_26),
.B(n_42),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_47),
.B(n_41),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_48),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_41),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g56 ( 
.A(n_54),
.B(n_39),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_52),
.Y(n_57)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_54),
.B(n_40),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_57),
.B(n_53),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_58),
.B(n_53),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_58),
.B(n_50),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_61),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_59),
.A2(n_55),
.B(n_56),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_56),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_51),
.Y(n_65)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_31),
.C(n_34),
.Y(n_66)
);

NOR3xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_22),
.C(n_24),
.Y(n_67)
);

AND2x4_ASAP7_75t_L g68 ( 
.A(n_67),
.B(n_66),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_67),
.A2(n_65),
.B1(n_25),
.B2(n_35),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_68),
.A2(n_25),
.B1(n_49),
.B2(n_55),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_69),
.Y(n_71)
);

OR2x6_ASAP7_75t_L g72 ( 
.A(n_71),
.B(n_55),
.Y(n_72)
);


endmodule