module fake_jpeg_22599_n_75 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_75);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_75;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_73;
wire n_19;
wire n_20;
wire n_18;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_71;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_65;
wire n_63;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_72;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_9;
wire n_36;
wire n_74;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_29;
wire n_43;
wire n_50;
wire n_37;
wire n_12;
wire n_32;
wire n_70;
wire n_15;
wire n_66;

INVx2_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_5),
.Y(n_10)
);

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_4),
.B(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_10),
.B(n_13),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_20),
.B(n_22),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_9),
.Y(n_27)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_24),
.A2(n_25),
.B1(n_19),
.B2(n_12),
.Y(n_28)
);

INVx11_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_13),
.B(n_0),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_26),
.B(n_12),
.C(n_17),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g45 ( 
.A(n_27),
.B(n_14),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

XNOR2xp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_20),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_26),
.B(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_31),
.A2(n_23),
.B(n_26),
.Y(n_35)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_35),
.A2(n_44),
.B(n_32),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_31),
.A2(n_22),
.B1(n_25),
.B2(n_24),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_36),
.B(n_43),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_42),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_23),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_34),
.A2(n_25),
.B1(n_21),
.B2(n_22),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g53 ( 
.A1(n_45),
.A2(n_14),
.B(n_15),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_30),
.C(n_32),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_51),
.C(n_39),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_48),
.A2(n_18),
.B1(n_11),
.B2(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_17),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_11),
.Y(n_57)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_53),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_30),
.C(n_21),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_47),
.A2(n_40),
.B1(n_44),
.B2(n_19),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_54),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g55 ( 
.A(n_46),
.B(n_40),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_55),
.B(n_59),
.C(n_52),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_57),
.Y(n_63)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_51),
.Y(n_60)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_60),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_61),
.B(n_65),
.C(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_0),
.Y(n_66)
);

OAI21xp5_ASAP7_75t_L g65 ( 
.A1(n_59),
.A2(n_0),
.B(n_1),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_66),
.B(n_68),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_67),
.B(n_61),
.C(n_62),
.Y(n_69)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

OAI21xp33_ASAP7_75t_L g71 ( 
.A1(n_69),
.A2(n_58),
.B(n_65),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_72),
.B(n_3),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_70),
.A2(n_54),
.B1(n_64),
.B2(n_2),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_3),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g75 ( 
.A(n_74),
.B(n_3),
.Y(n_75)
);


endmodule