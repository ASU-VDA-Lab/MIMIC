module real_aes_6523_n_100 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_100);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_100;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_726;
wire n_369;
wire n_343;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_119;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_552;
wire n_402;
wire n_617;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_148;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_349;
wire n_336;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g551 ( .A1(n_0), .A2(n_158), .B(n_552), .C(n_555), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_1), .B(n_496), .Y(n_556) );
INVx1_ASAP7_75t_L g106 ( .A(n_2), .Y(n_106) );
INVx1_ASAP7_75t_L g192 ( .A(n_3), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g530 ( .A(n_4), .B(n_150), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g489 ( .A1(n_5), .A2(n_465), .B(n_490), .Y(n_489) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_6), .A2(n_135), .B(n_481), .Y(n_480) );
AOI22xp33_ASAP7_75t_L g221 ( .A1(n_7), .A2(n_36), .B1(n_144), .B2(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_8), .B(n_135), .Y(n_161) );
AND2x6_ASAP7_75t_L g159 ( .A(n_9), .B(n_160), .Y(n_159) );
A2O1A1Ixp33_ASAP7_75t_L g454 ( .A1(n_10), .A2(n_159), .B(n_455), .C(n_457), .Y(n_454) );
INVx1_ASAP7_75t_L g104 ( .A(n_11), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_11), .B(n_37), .Y(n_121) );
INVx1_ASAP7_75t_L g140 ( .A(n_12), .Y(n_140) );
INVx1_ASAP7_75t_L g185 ( .A(n_13), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_14), .B(n_148), .Y(n_228) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_15), .B(n_150), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_16), .B(n_136), .Y(n_197) );
AO32x2_ASAP7_75t_L g219 ( .A1(n_17), .A2(n_135), .A3(n_165), .B1(n_176), .B2(n_220), .Y(n_219) );
NAND2xp5_ASAP7_75t_SL g232 ( .A(n_18), .B(n_144), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_19), .B(n_136), .Y(n_194) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_20), .A2(n_53), .B1(n_144), .B2(n_222), .Y(n_223) );
AOI22xp33_ASAP7_75t_SL g244 ( .A1(n_21), .A2(n_80), .B1(n_144), .B2(n_148), .Y(n_244) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_22), .B(n_144), .Y(n_214) );
A2O1A1Ixp33_ASAP7_75t_L g515 ( .A1(n_23), .A2(n_176), .B(n_455), .C(n_516), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g100 ( .A1(n_24), .A2(n_101), .B1(n_102), .B2(n_110), .Y(n_100) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_25), .A2(n_176), .B(n_455), .C(n_484), .Y(n_483) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_26), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_27), .B(n_178), .Y(n_177) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_28), .Y(n_122) );
AOI21xp5_ASAP7_75t_L g548 ( .A1(n_29), .A2(n_465), .B(n_549), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_30), .B(n_178), .Y(n_216) );
INVx2_ASAP7_75t_L g146 ( .A(n_31), .Y(n_146) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_32), .A2(n_467), .B(n_475), .C(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g168 ( .A(n_33), .B(n_144), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_34), .B(n_178), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_35), .B(n_230), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g103 ( .A(n_37), .B(n_104), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_38), .B(n_514), .Y(n_513) );
CKINVDCx20_ASAP7_75t_R g461 ( .A(n_39), .Y(n_461) );
AOI222xp33_ASAP7_75t_SL g123 ( .A1(n_40), .A2(n_78), .B1(n_124), .B2(n_730), .C1(n_731), .C2(n_735), .Y(n_123) );
CKINVDCx16_ASAP7_75t_R g730 ( .A(n_40), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_41), .B(n_150), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_42), .B(n_465), .Y(n_482) );
OAI22xp5_ASAP7_75t_SL g745 ( .A1(n_43), .A2(n_77), .B1(n_438), .B2(n_746), .Y(n_745) );
CKINVDCx20_ASAP7_75t_R g746 ( .A(n_43), .Y(n_746) );
A2O1A1Ixp33_ASAP7_75t_L g466 ( .A1(n_44), .A2(n_467), .B(n_469), .C(n_475), .Y(n_466) );
NAND2xp5_ASAP7_75t_SL g143 ( .A(n_45), .B(n_144), .Y(n_143) );
INVx1_ASAP7_75t_L g553 ( .A(n_46), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_47), .A2(n_89), .B1(n_222), .B2(n_243), .Y(n_242) );
INVx1_ASAP7_75t_L g470 ( .A(n_48), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g154 ( .A(n_49), .B(n_144), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_50), .B(n_144), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_51), .B(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_52), .B(n_156), .Y(n_155) );
AOI22xp33_ASAP7_75t_SL g201 ( .A1(n_54), .A2(n_58), .B1(n_144), .B2(n_148), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g521 ( .A(n_55), .Y(n_521) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_56), .B(n_144), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g227 ( .A(n_57), .B(n_144), .Y(n_227) );
INVx1_ASAP7_75t_L g160 ( .A(n_59), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_60), .B(n_465), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_61), .B(n_496), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_62), .A2(n_156), .B(n_188), .C(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_63), .B(n_144), .Y(n_193) );
INVx1_ASAP7_75t_L g139 ( .A(n_64), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_65), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_66), .B(n_150), .Y(n_506) );
AO32x2_ASAP7_75t_L g240 ( .A1(n_67), .A2(n_135), .A3(n_176), .B1(n_241), .B2(n_245), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_68), .B(n_151), .Y(n_458) );
INVx1_ASAP7_75t_L g171 ( .A(n_69), .Y(n_171) );
INVx1_ASAP7_75t_L g211 ( .A(n_70), .Y(n_211) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_71), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_72), .B(n_472), .Y(n_517) );
A2O1A1Ixp33_ASAP7_75t_L g527 ( .A1(n_73), .A2(n_455), .B(n_475), .C(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_74), .B(n_148), .Y(n_212) );
CKINVDCx16_ASAP7_75t_R g491 ( .A(n_75), .Y(n_491) );
INVx1_ASAP7_75t_L g109 ( .A(n_76), .Y(n_109) );
OAI22xp5_ASAP7_75t_SL g126 ( .A1(n_77), .A2(n_127), .B1(n_437), .B2(n_438), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_77), .Y(n_438) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_79), .B(n_471), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_81), .B(n_222), .Y(n_233) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_82), .Y(n_508) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_83), .B(n_148), .Y(n_215) );
INVx2_ASAP7_75t_L g137 ( .A(n_84), .Y(n_137) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_85), .Y(n_534) );
NAND2xp5_ASAP7_75t_SL g459 ( .A(n_86), .B(n_175), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_87), .B(n_148), .Y(n_147) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_88), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g118 ( .A(n_88), .B(n_119), .Y(n_118) );
OR2x2_ASAP7_75t_L g441 ( .A(n_88), .B(n_120), .Y(n_441) );
INVx2_ASAP7_75t_L g729 ( .A(n_88), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g200 ( .A1(n_90), .A2(n_99), .B1(n_148), .B2(n_149), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_91), .B(n_465), .Y(n_502) );
INVx1_ASAP7_75t_L g505 ( .A(n_92), .Y(n_505) );
INVxp67_ASAP7_75t_L g494 ( .A(n_93), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_94), .B(n_148), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_95), .B(n_109), .Y(n_108) );
INVx1_ASAP7_75t_L g451 ( .A(n_96), .Y(n_451) );
INVx1_ASAP7_75t_L g529 ( .A(n_97), .Y(n_529) );
AND2x2_ASAP7_75t_L g477 ( .A(n_98), .B(n_178), .Y(n_477) );
INVx1_ASAP7_75t_L g101 ( .A(n_102), .Y(n_101) );
OR2x4_ASAP7_75t_L g102 ( .A(n_103), .B(n_105), .Y(n_102) );
AND2x2_ASAP7_75t_L g120 ( .A(n_106), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_123), .B1(n_738), .B2(n_739), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_116), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_SL g738 ( .A(n_114), .Y(n_738) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g739 ( .A1(n_116), .A2(n_740), .B(n_747), .Y(n_739) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_122), .Y(n_116) );
HB1xp67_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_SL g748 ( .A(n_118), .Y(n_748) );
NOR2x2_ASAP7_75t_L g737 ( .A(n_119), .B(n_729), .Y(n_737) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g728 ( .A(n_120), .B(n_729), .Y(n_728) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_439), .B1(n_442), .B2(n_726), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_SL g731 ( .A1(n_126), .A2(n_732), .B1(n_733), .B2(n_734), .Y(n_731) );
INVx2_ASAP7_75t_L g437 ( .A(n_127), .Y(n_437) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_127), .A2(n_437), .B1(n_744), .B2(n_745), .Y(n_743) );
NAND2x1p5_ASAP7_75t_L g127 ( .A(n_128), .B(n_361), .Y(n_127) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_319), .Y(n_128) );
NOR4xp25_ASAP7_75t_L g129 ( .A(n_130), .B(n_259), .C(n_295), .D(n_309), .Y(n_129) );
OAI221xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_203), .B1(n_235), .B2(n_246), .C(n_250), .Y(n_130) );
NAND2xp5_ASAP7_75t_SL g393 ( .A(n_131), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g131 ( .A(n_132), .B(n_179), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
AND2x2_ASAP7_75t_L g133 ( .A(n_134), .B(n_162), .Y(n_133) );
AND2x2_ASAP7_75t_L g256 ( .A(n_134), .B(n_163), .Y(n_256) );
INVx3_ASAP7_75t_L g264 ( .A(n_134), .Y(n_264) );
AND2x2_ASAP7_75t_L g318 ( .A(n_134), .B(n_182), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_134), .B(n_181), .Y(n_354) );
AND2x2_ASAP7_75t_L g412 ( .A(n_134), .B(n_274), .Y(n_412) );
OA21x2_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_141), .B(n_161), .Y(n_134) );
INVx4_ASAP7_75t_L g202 ( .A(n_135), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_135), .A2(n_482), .B(n_483), .Y(n_481) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_135), .Y(n_488) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g165 ( .A(n_136), .Y(n_165) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_137), .B(n_138), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
OAI21xp5_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_153), .B(n_159), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g142 ( .A1(n_143), .A2(n_147), .B(n_150), .Y(n_142) );
INVx3_ASAP7_75t_L g210 ( .A(n_144), .Y(n_210) );
HB1xp67_ASAP7_75t_L g531 ( .A(n_144), .Y(n_531) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g222 ( .A(n_145), .Y(n_222) );
BUFx3_ASAP7_75t_L g243 ( .A(n_145), .Y(n_243) );
AND2x6_ASAP7_75t_L g455 ( .A(n_145), .B(n_456), .Y(n_455) );
INVx2_ASAP7_75t_L g145 ( .A(n_146), .Y(n_145) );
INVx1_ASAP7_75t_L g149 ( .A(n_146), .Y(n_149) );
INVx1_ASAP7_75t_L g157 ( .A(n_146), .Y(n_157) );
INVx2_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx3_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g158 ( .A(n_150), .Y(n_158) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_150), .A2(n_168), .B(n_169), .Y(n_167) );
O2A1O1Ixp5_ASAP7_75t_SL g209 ( .A1(n_150), .A2(n_210), .B(n_211), .C(n_212), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_150), .B(n_494), .Y(n_493) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI22xp5_ASAP7_75t_SL g241 ( .A1(n_151), .A2(n_175), .B1(n_242), .B2(n_244), .Y(n_241) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_152), .Y(n_175) );
BUFx6f_ASAP7_75t_L g190 ( .A(n_152), .Y(n_190) );
INVx1_ASAP7_75t_L g230 ( .A(n_152), .Y(n_230) );
AND2x2_ASAP7_75t_L g453 ( .A(n_152), .B(n_157), .Y(n_453) );
INVx1_ASAP7_75t_L g456 ( .A(n_152), .Y(n_456) );
AOI21xp5_ASAP7_75t_L g153 ( .A1(n_154), .A2(n_155), .B(n_158), .Y(n_153) );
INVx2_ASAP7_75t_L g172 ( .A(n_156), .Y(n_172) );
INVx1_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
O2A1O1Ixp33_ASAP7_75t_L g191 ( .A1(n_158), .A2(n_172), .B(n_192), .C(n_193), .Y(n_191) );
OAI22xp5_ASAP7_75t_L g199 ( .A1(n_158), .A2(n_175), .B1(n_200), .B2(n_201), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g220 ( .A1(n_158), .A2(n_175), .B1(n_221), .B2(n_223), .Y(n_220) );
BUFx3_ASAP7_75t_L g176 ( .A(n_159), .Y(n_176) );
OAI21xp5_ASAP7_75t_L g183 ( .A1(n_159), .A2(n_184), .B(n_191), .Y(n_183) );
OAI21xp5_ASAP7_75t_L g208 ( .A1(n_159), .A2(n_209), .B(n_213), .Y(n_208) );
OAI21xp5_ASAP7_75t_L g225 ( .A1(n_159), .A2(n_226), .B(n_231), .Y(n_225) );
NAND2x1p5_ASAP7_75t_L g452 ( .A(n_159), .B(n_453), .Y(n_452) );
AND2x4_ASAP7_75t_L g465 ( .A(n_159), .B(n_453), .Y(n_465) );
INVx4_ASAP7_75t_SL g476 ( .A(n_159), .Y(n_476) );
AND2x2_ASAP7_75t_L g247 ( .A(n_162), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g261 ( .A(n_162), .B(n_182), .Y(n_261) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_163), .B(n_182), .Y(n_276) );
AND2x2_ASAP7_75t_L g288 ( .A(n_163), .B(n_264), .Y(n_288) );
OR2x2_ASAP7_75t_L g290 ( .A(n_163), .B(n_248), .Y(n_290) );
AND2x2_ASAP7_75t_L g325 ( .A(n_163), .B(n_248), .Y(n_325) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_163), .Y(n_370) );
INVx1_ASAP7_75t_L g378 ( .A(n_163), .Y(n_378) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_166), .B(n_177), .Y(n_163) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_164), .A2(n_183), .B(n_194), .Y(n_182) );
INVx2_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_165), .B(n_461), .Y(n_460) );
OAI21xp5_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_170), .B(n_176), .Y(n_166) );
O2A1O1Ixp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_172), .B(n_173), .C(n_174), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_172), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g231 ( .A1(n_174), .A2(n_232), .B(n_233), .Y(n_231) );
INVx2_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
INVx4_ASAP7_75t_L g554 ( .A(n_175), .Y(n_554) );
NAND3xp33_ASAP7_75t_L g198 ( .A(n_176), .B(n_199), .C(n_202), .Y(n_198) );
OA21x2_ASAP7_75t_L g207 ( .A1(n_178), .A2(n_208), .B(n_216), .Y(n_207) );
OA21x2_ASAP7_75t_L g224 ( .A1(n_178), .A2(n_225), .B(n_234), .Y(n_224) );
INVx2_ASAP7_75t_L g245 ( .A(n_178), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_178), .A2(n_464), .B(n_466), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_178), .A2(n_502), .B(n_503), .Y(n_501) );
INVx1_ASAP7_75t_L g522 ( .A(n_178), .Y(n_522) );
OAI221xp5_ASAP7_75t_L g295 ( .A1(n_179), .A2(n_296), .B1(n_300), .B2(n_304), .C(n_305), .Y(n_295) );
INVx1_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
AND2x2_ASAP7_75t_L g255 ( .A(n_180), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_195), .Y(n_180) );
INVx2_ASAP7_75t_L g254 ( .A(n_181), .Y(n_254) );
AND2x2_ASAP7_75t_L g307 ( .A(n_181), .B(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g326 ( .A(n_181), .B(n_264), .Y(n_326) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AND2x2_ASAP7_75t_L g389 ( .A(n_182), .B(n_264), .Y(n_389) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_185), .A2(n_186), .B(n_187), .C(n_188), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g457 ( .A1(n_186), .A2(n_458), .B(n_459), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_186), .A2(n_485), .B(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g528 ( .A1(n_188), .A2(n_529), .B(n_530), .C(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_189), .A2(n_214), .B(n_215), .Y(n_213) );
INVx4_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
INVx2_ASAP7_75t_L g472 ( .A(n_190), .Y(n_472) );
AND2x2_ASAP7_75t_L g311 ( .A(n_195), .B(n_256), .Y(n_311) );
OAI322xp33_ASAP7_75t_L g379 ( .A1(n_195), .A2(n_335), .A3(n_380), .B1(n_382), .B2(n_385), .C1(n_387), .C2(n_391), .Y(n_379) );
INVx3_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
NOR2x1_ASAP7_75t_L g262 ( .A(n_196), .B(n_263), .Y(n_262) );
INVx2_ASAP7_75t_L g275 ( .A(n_196), .Y(n_275) );
AND2x2_ASAP7_75t_L g384 ( .A(n_196), .B(n_264), .Y(n_384) );
AND2x2_ASAP7_75t_L g416 ( .A(n_196), .B(n_288), .Y(n_416) );
OR2x2_ASAP7_75t_L g419 ( .A(n_196), .B(n_420), .Y(n_419) );
AND2x4_ASAP7_75t_L g196 ( .A(n_197), .B(n_198), .Y(n_196) );
INVx1_ASAP7_75t_L g249 ( .A(n_197), .Y(n_249) );
AO21x1_ASAP7_75t_L g248 ( .A1(n_199), .A2(n_202), .B(n_249), .Y(n_248) );
AO21x2_ASAP7_75t_L g449 ( .A1(n_202), .A2(n_450), .B(n_460), .Y(n_449) );
INVx3_ASAP7_75t_L g496 ( .A(n_202), .Y(n_496) );
NOR2xp33_ASAP7_75t_L g507 ( .A(n_202), .B(n_508), .Y(n_507) );
AO21x2_ASAP7_75t_L g525 ( .A1(n_202), .A2(n_526), .B(n_533), .Y(n_525) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_202), .B(n_534), .Y(n_533) );
INVx1_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_217), .Y(n_204) );
INVx1_ASAP7_75t_L g432 ( .A(n_205), .Y(n_432) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g237 ( .A(n_206), .B(n_224), .Y(n_237) );
INVx2_ASAP7_75t_L g272 ( .A(n_206), .Y(n_272) );
INVx2_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
INVx2_ASAP7_75t_L g294 ( .A(n_207), .Y(n_294) );
HB1xp67_ASAP7_75t_L g302 ( .A(n_207), .Y(n_302) );
OR2x2_ASAP7_75t_L g426 ( .A(n_207), .B(n_427), .Y(n_426) );
AND2x2_ASAP7_75t_L g251 ( .A(n_217), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g291 ( .A(n_217), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g343 ( .A(n_217), .B(n_344), .Y(n_343) );
AND2x2_ASAP7_75t_L g217 ( .A(n_218), .B(n_224), .Y(n_217) );
AND2x2_ASAP7_75t_L g238 ( .A(n_218), .B(n_239), .Y(n_238) );
NOR2xp67_ASAP7_75t_L g298 ( .A(n_218), .B(n_299), .Y(n_298) );
AND2x2_ASAP7_75t_L g352 ( .A(n_218), .B(n_240), .Y(n_352) );
OR2x2_ASAP7_75t_L g360 ( .A(n_218), .B(n_294), .Y(n_360) );
INVx2_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
BUFx2_ASAP7_75t_L g269 ( .A(n_219), .Y(n_269) );
AND2x2_ASAP7_75t_L g279 ( .A(n_219), .B(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g303 ( .A(n_219), .B(n_224), .Y(n_303) );
AND2x2_ASAP7_75t_L g367 ( .A(n_219), .B(n_240), .Y(n_367) );
NOR2xp33_ASAP7_75t_L g257 ( .A(n_224), .B(n_258), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_224), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g280 ( .A(n_224), .Y(n_280) );
INVx1_ASAP7_75t_L g285 ( .A(n_224), .Y(n_285) );
AND2x2_ASAP7_75t_L g297 ( .A(n_224), .B(n_298), .Y(n_297) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_224), .Y(n_375) );
INVx1_ASAP7_75t_L g427 ( .A(n_224), .Y(n_427) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_228), .B(n_229), .Y(n_226) );
INVx1_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g235 ( .A(n_236), .B(n_238), .Y(n_235) );
AND2x2_ASAP7_75t_L g404 ( .A(n_236), .B(n_313), .Y(n_404) );
INVx2_ASAP7_75t_SL g236 ( .A(n_237), .Y(n_236) );
AND2x2_ASAP7_75t_L g331 ( .A(n_238), .B(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g430 ( .A(n_238), .B(n_365), .Y(n_430) );
INVx1_ASAP7_75t_L g252 ( .A(n_239), .Y(n_252) );
AND2x2_ASAP7_75t_L g278 ( .A(n_239), .B(n_272), .Y(n_278) );
BUFx2_ASAP7_75t_L g337 ( .A(n_239), .Y(n_337) );
INVx1_ASAP7_75t_L g239 ( .A(n_240), .Y(n_239) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_240), .Y(n_258) );
INVx1_ASAP7_75t_L g268 ( .A(n_240), .Y(n_268) );
HB1xp67_ASAP7_75t_L g474 ( .A(n_243), .Y(n_474) );
INVx2_ASAP7_75t_L g555 ( .A(n_243), .Y(n_555) );
INVx1_ASAP7_75t_L g519 ( .A(n_245), .Y(n_519) );
NOR2xp67_ASAP7_75t_L g406 ( .A(n_246), .B(n_253), .Y(n_406) );
INVx2_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AOI32xp33_ASAP7_75t_L g250 ( .A1(n_247), .A2(n_251), .A3(n_253), .B1(n_255), .B2(n_257), .Y(n_250) );
AND2x2_ASAP7_75t_L g390 ( .A(n_247), .B(n_263), .Y(n_390) );
AND2x2_ASAP7_75t_L g428 ( .A(n_247), .B(n_326), .Y(n_428) );
INVx1_ASAP7_75t_L g308 ( .A(n_248), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_252), .B(n_314), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_253), .B(n_288), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_253), .B(n_256), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g407 ( .A(n_253), .B(n_325), .Y(n_407) );
OR2x2_ASAP7_75t_L g421 ( .A(n_253), .B(n_290), .Y(n_421) );
INVx3_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g348 ( .A(n_254), .B(n_256), .Y(n_348) );
OR2x2_ASAP7_75t_L g357 ( .A(n_254), .B(n_344), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_256), .B(n_307), .Y(n_329) );
INVx2_ASAP7_75t_L g344 ( .A(n_258), .Y(n_344) );
OR2x2_ASAP7_75t_L g359 ( .A(n_258), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g374 ( .A(n_258), .B(n_375), .Y(n_374) );
A2O1A1Ixp33_ASAP7_75t_L g431 ( .A1(n_258), .A2(n_351), .B(n_432), .C(n_433), .Y(n_431) );
OAI321xp33_ASAP7_75t_L g259 ( .A1(n_260), .A2(n_265), .A3(n_270), .B1(n_273), .B2(n_277), .C(n_281), .Y(n_259) );
INVx1_ASAP7_75t_L g372 ( .A(n_260), .Y(n_372) );
NAND2x1p5_ASAP7_75t_L g260 ( .A(n_261), .B(n_262), .Y(n_260) );
AND2x2_ASAP7_75t_L g383 ( .A(n_261), .B(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g335 ( .A(n_263), .Y(n_335) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_264), .B(n_378), .Y(n_395) );
OAI221xp5_ASAP7_75t_L g402 ( .A1(n_265), .A2(n_403), .B1(n_405), .B2(n_407), .C(n_408), .Y(n_402) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
AND2x2_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g340 ( .A(n_267), .B(n_314), .Y(n_340) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_268), .B(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g313 ( .A(n_269), .Y(n_313) );
A2O1A1Ixp33_ASAP7_75t_L g355 ( .A1(n_270), .A2(n_311), .B(n_356), .C(n_358), .Y(n_355) );
INVx1_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
AND2x2_ASAP7_75t_L g322 ( .A(n_272), .B(n_279), .Y(n_322) );
BUFx2_ASAP7_75t_L g332 ( .A(n_272), .Y(n_332) );
INVx1_ASAP7_75t_L g347 ( .A(n_272), .Y(n_347) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
NOR2xp33_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
OR2x2_ASAP7_75t_L g353 ( .A(n_275), .B(n_354), .Y(n_353) );
INVx1_ASAP7_75t_L g436 ( .A(n_275), .Y(n_436) );
INVx1_ASAP7_75t_L g429 ( .A(n_276), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_278), .B(n_279), .Y(n_277) );
AND2x2_ASAP7_75t_L g282 ( .A(n_278), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g386 ( .A(n_278), .B(n_303), .Y(n_386) );
INVx1_ASAP7_75t_L g315 ( .A(n_279), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_286), .B1(n_289), .B2(n_291), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_283), .B(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g351 ( .A(n_284), .B(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g284 ( .A(n_285), .Y(n_284) );
AND2x2_ASAP7_75t_SL g314 ( .A(n_285), .B(n_294), .Y(n_314) );
INVx1_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g306 ( .A(n_288), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g316 ( .A(n_290), .B(n_317), .Y(n_316) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
OAI221xp5_ASAP7_75t_L g410 ( .A1(n_293), .A2(n_411), .B1(n_413), .B2(n_414), .C(n_415), .Y(n_410) );
INVx1_ASAP7_75t_L g299 ( .A(n_294), .Y(n_299) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_294), .Y(n_365) );
INVx1_ASAP7_75t_SL g296 ( .A(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_297), .B(n_416), .Y(n_415) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_298), .A2(n_303), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_301), .B(n_311), .Y(n_408) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
INVx1_ASAP7_75t_L g377 ( .A(n_302), .Y(n_377) );
AND2x2_ASAP7_75t_L g336 ( .A(n_303), .B(n_337), .Y(n_336) );
INVx2_ASAP7_75t_L g425 ( .A(n_303), .Y(n_425) );
INVx1_ASAP7_75t_L g341 ( .A(n_306), .Y(n_341) );
INVx1_ASAP7_75t_L g396 ( .A(n_307), .Y(n_396) );
OAI22xp5_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_312), .B1(n_315), .B2(n_316), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_313), .B(n_347), .Y(n_346) );
INVx2_ASAP7_75t_L g381 ( .A(n_314), .Y(n_381) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_314), .B(n_352), .Y(n_418) );
OR2x2_ASAP7_75t_L g391 ( .A(n_315), .B(n_344), .Y(n_391) );
INVx1_ASAP7_75t_L g330 ( .A(n_316), .Y(n_330) );
INVx1_ASAP7_75t_SL g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_318), .B(n_369), .Y(n_368) );
NOR3xp33_ASAP7_75t_L g319 ( .A(n_320), .B(n_338), .C(n_349), .Y(n_319) );
OAI211xp5_ASAP7_75t_L g320 ( .A1(n_321), .A2(n_323), .B(n_327), .C(n_333), .Y(n_320) );
INVxp67_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
AOI221xp5_ASAP7_75t_L g392 ( .A1(n_322), .A2(n_393), .B1(n_397), .B2(n_400), .C(n_402), .Y(n_392) );
INVx1_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
AND2x2_ASAP7_75t_L g334 ( .A(n_325), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g388 ( .A(n_325), .B(n_389), .Y(n_388) );
OAI211xp5_ASAP7_75t_L g373 ( .A1(n_326), .A2(n_374), .B(n_376), .C(n_378), .Y(n_373) );
INVx2_ASAP7_75t_L g420 ( .A(n_326), .Y(n_420) );
OAI21xp5_ASAP7_75t_SL g327 ( .A1(n_328), .A2(n_330), .B(n_331), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g399 ( .A(n_332), .B(n_352), .Y(n_399) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_334), .B(n_336), .Y(n_333) );
OAI21xp5_ASAP7_75t_SL g338 ( .A1(n_339), .A2(n_341), .B(n_342), .Y(n_338) );
INVxp67_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
OAI21xp5_ASAP7_75t_SL g342 ( .A1(n_343), .A2(n_345), .B(n_348), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_343), .B(n_372), .Y(n_371) );
INVxp67_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_348), .B(n_435), .Y(n_434) );
OAI21xp33_ASAP7_75t_L g349 ( .A1(n_350), .A2(n_353), .B(n_355), .Y(n_349) );
INVx1_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g376 ( .A(n_352), .B(n_377), .Y(n_376) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
AND4x1_ASAP7_75t_L g361 ( .A(n_362), .B(n_392), .C(n_409), .D(n_431), .Y(n_361) );
NOR2xp33_ASAP7_75t_L g362 ( .A(n_363), .B(n_379), .Y(n_362) );
OAI211xp5_ASAP7_75t_SL g363 ( .A1(n_364), .A2(n_368), .B(n_371), .C(n_373), .Y(n_363) );
OR2x2_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
INVx1_ASAP7_75t_SL g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_367), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_378), .B(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_388), .B(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g413 ( .A(n_388), .Y(n_413) );
INVx2_ASAP7_75t_SL g401 ( .A(n_389), .Y(n_401) );
OR2x2_ASAP7_75t_L g394 ( .A(n_395), .B(n_396), .Y(n_394) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g414 ( .A(n_399), .Y(n_414) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NOR2xp33_ASAP7_75t_SL g409 ( .A(n_410), .B(n_417), .Y(n_409) );
INVx1_ASAP7_75t_SL g411 ( .A(n_412), .Y(n_411) );
OAI221xp5_ASAP7_75t_SL g417 ( .A1(n_418), .A2(n_419), .B1(n_421), .B2(n_422), .C(n_423), .Y(n_417) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_424), .A2(n_428), .B1(n_429), .B2(n_430), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g424 ( .A(n_425), .B(n_426), .Y(n_424) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx2_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g732 ( .A(n_440), .Y(n_732) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g733 ( .A(n_442), .Y(n_733) );
OR3x1_ASAP7_75t_L g442 ( .A(n_443), .B(n_624), .C(n_689), .Y(n_442) );
NAND4xp25_ASAP7_75t_SL g443 ( .A(n_444), .B(n_565), .C(n_591), .D(n_614), .Y(n_443) );
AOI221xp5_ASAP7_75t_L g444 ( .A1(n_445), .A2(n_497), .B1(n_535), .B2(n_542), .C(n_557), .Y(n_444) );
CKINVDCx14_ASAP7_75t_R g445 ( .A(n_446), .Y(n_445) );
OAI22xp5_ASAP7_75t_L g712 ( .A1(n_446), .A2(n_558), .B1(n_582), .B2(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g446 ( .A(n_447), .B(n_478), .Y(n_446) );
INVx1_ASAP7_75t_SL g618 ( .A(n_447), .Y(n_618) );
OR2x2_ASAP7_75t_L g447 ( .A(n_448), .B(n_462), .Y(n_447) );
OR2x2_ASAP7_75t_L g540 ( .A(n_448), .B(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g560 ( .A(n_448), .B(n_479), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_448), .B(n_487), .Y(n_573) );
AND2x2_ASAP7_75t_L g590 ( .A(n_448), .B(n_462), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g612 ( .A(n_448), .B(n_538), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_448), .B(n_589), .Y(n_701) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_448), .B(n_478), .Y(n_711) );
AOI211xp5_ASAP7_75t_SL g722 ( .A1(n_448), .A2(n_628), .B(n_723), .C(n_724), .Y(n_722) );
INVx5_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g594 ( .A(n_449), .B(n_479), .Y(n_594) );
AND2x2_ASAP7_75t_L g597 ( .A(n_449), .B(n_480), .Y(n_597) );
OR2x2_ASAP7_75t_L g642 ( .A(n_449), .B(n_479), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_449), .B(n_487), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_451), .A2(n_452), .B(n_454), .Y(n_450) );
INVx5_ASAP7_75t_L g468 ( .A(n_455), .Y(n_468) );
INVx5_ASAP7_75t_SL g541 ( .A(n_462), .Y(n_541) );
AND2x2_ASAP7_75t_L g559 ( .A(n_462), .B(n_560), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_462), .B(n_642), .Y(n_641) );
AND2x2_ASAP7_75t_L g645 ( .A(n_462), .B(n_646), .Y(n_645) );
AND2x2_ASAP7_75t_L g677 ( .A(n_462), .B(n_487), .Y(n_677) );
OR2x2_ASAP7_75t_L g683 ( .A(n_462), .B(n_573), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_462), .B(n_633), .Y(n_692) );
OR2x6_ASAP7_75t_L g462 ( .A(n_463), .B(n_477), .Y(n_462) );
BUFx2_ASAP7_75t_L g514 ( .A(n_465), .Y(n_514) );
INVx2_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
O2A1O1Ixp33_ASAP7_75t_L g490 ( .A1(n_468), .A2(n_476), .B(n_491), .C(n_492), .Y(n_490) );
O2A1O1Ixp33_ASAP7_75t_SL g549 ( .A1(n_468), .A2(n_476), .B(n_550), .C(n_551), .Y(n_549) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_473), .C(n_474), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_471), .A2(n_474), .B(n_505), .C(n_506), .Y(n_504) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g478 ( .A(n_479), .B(n_487), .Y(n_478) );
AND2x2_ASAP7_75t_L g574 ( .A(n_479), .B(n_541), .Y(n_574) );
INVx1_ASAP7_75t_SL g587 ( .A(n_479), .Y(n_587) );
OR2x2_ASAP7_75t_L g622 ( .A(n_479), .B(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g628 ( .A(n_479), .B(n_487), .Y(n_628) );
AND2x2_ASAP7_75t_L g686 ( .A(n_479), .B(n_538), .Y(n_686) );
INVx2_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_480), .B(n_541), .Y(n_613) );
INVx3_ASAP7_75t_L g538 ( .A(n_487), .Y(n_538) );
OR2x2_ASAP7_75t_L g579 ( .A(n_487), .B(n_541), .Y(n_579) );
AND2x2_ASAP7_75t_L g589 ( .A(n_487), .B(n_587), .Y(n_589) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_487), .Y(n_637) );
AND2x2_ASAP7_75t_L g646 ( .A(n_487), .B(n_560), .Y(n_646) );
OA21x2_ASAP7_75t_L g487 ( .A1(n_488), .A2(n_489), .B(n_495), .Y(n_487) );
OA21x2_ASAP7_75t_L g547 ( .A1(n_496), .A2(n_548), .B(n_556), .Y(n_547) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_497), .A2(n_663), .B1(n_665), .B2(n_667), .C(n_670), .Y(n_662) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_509), .Y(n_498) );
AND2x2_ASAP7_75t_L g636 ( .A(n_499), .B(n_617), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_499), .B(n_695), .Y(n_699) );
OR2x2_ASAP7_75t_L g720 ( .A(n_499), .B(n_721), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_499), .B(n_725), .Y(n_724) );
BUFx2_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx5_ASAP7_75t_L g567 ( .A(n_500), .Y(n_567) );
AND2x2_ASAP7_75t_L g644 ( .A(n_500), .B(n_511), .Y(n_644) );
AND2x2_ASAP7_75t_L g705 ( .A(n_500), .B(n_584), .Y(n_705) );
AND2x2_ASAP7_75t_L g718 ( .A(n_500), .B(n_538), .Y(n_718) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_507), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_510), .B(n_523), .Y(n_509) );
AND2x4_ASAP7_75t_L g545 ( .A(n_510), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g563 ( .A(n_510), .B(n_564), .Y(n_563) );
INVx2_ASAP7_75t_L g570 ( .A(n_510), .Y(n_570) );
AND2x2_ASAP7_75t_L g639 ( .A(n_510), .B(n_617), .Y(n_639) );
AND2x2_ASAP7_75t_L g649 ( .A(n_510), .B(n_567), .Y(n_649) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_510), .Y(n_657) );
AND2x2_ASAP7_75t_L g669 ( .A(n_510), .B(n_547), .Y(n_669) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_510), .B(n_601), .Y(n_673) );
AND2x2_ASAP7_75t_L g710 ( .A(n_510), .B(n_705), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_510), .B(n_584), .Y(n_721) );
OR2x2_ASAP7_75t_L g723 ( .A(n_510), .B(n_659), .Y(n_723) );
INVx5_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g609 ( .A(n_511), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g619 ( .A(n_511), .B(n_564), .Y(n_619) );
AND2x2_ASAP7_75t_L g631 ( .A(n_511), .B(n_547), .Y(n_631) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_511), .Y(n_661) );
AND2x4_ASAP7_75t_L g695 ( .A(n_511), .B(n_546), .Y(n_695) );
OR2x6_ASAP7_75t_L g511 ( .A(n_512), .B(n_520), .Y(n_511) );
AOI21xp5_ASAP7_75t_SL g512 ( .A1(n_513), .A2(n_515), .B(n_519), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_522), .Y(n_520) );
BUFx2_ASAP7_75t_L g544 ( .A(n_523), .Y(n_544) );
HB1xp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g584 ( .A(n_524), .Y(n_584) );
AND2x2_ASAP7_75t_L g617 ( .A(n_524), .B(n_547), .Y(n_617) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
AND2x2_ASAP7_75t_L g564 ( .A(n_525), .B(n_547), .Y(n_564) );
BUFx2_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_527), .B(n_532), .Y(n_526) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_539), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_537), .B(n_618), .Y(n_697) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_538), .B(n_560), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_538), .B(n_541), .Y(n_599) );
AND2x2_ASAP7_75t_L g654 ( .A(n_538), .B(n_590), .Y(n_654) );
AOI221xp5_ASAP7_75t_SL g591 ( .A1(n_539), .A2(n_592), .B1(n_600), .B2(n_602), .C(n_606), .Y(n_591) );
INVx2_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
OR2x2_ASAP7_75t_L g586 ( .A(n_540), .B(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g627 ( .A(n_540), .B(n_628), .Y(n_627) );
OAI321xp33_ASAP7_75t_L g634 ( .A1(n_540), .A2(n_593), .A3(n_635), .B1(n_637), .B2(n_638), .C(n_640), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_541), .B(n_686), .Y(n_685) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_544), .B(n_545), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_544), .B(n_695), .Y(n_713) );
AND2x2_ASAP7_75t_L g600 ( .A(n_545), .B(n_601), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_545), .B(n_604), .Y(n_603) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_546), .Y(n_576) );
AND2x2_ASAP7_75t_L g583 ( .A(n_546), .B(n_584), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_546), .B(n_658), .Y(n_688) );
INVx1_ASAP7_75t_L g725 ( .A(n_546), .Y(n_725) );
INVx2_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_562), .Y(n_557) );
INVx1_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
A2O1A1Ixp33_ASAP7_75t_L g717 ( .A1(n_559), .A2(n_669), .B(n_718), .C(n_719), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_560), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_560), .B(n_598), .Y(n_664) );
INVx1_ASAP7_75t_SL g562 ( .A(n_563), .Y(n_562) );
INVx1_ASAP7_75t_L g607 ( .A(n_564), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_564), .B(n_567), .Y(n_621) );
NOR2xp33_ASAP7_75t_L g630 ( .A(n_564), .B(n_631), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_564), .B(n_649), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_566), .A2(n_568), .B1(n_580), .B2(n_585), .Y(n_565) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
OR2x2_ASAP7_75t_L g581 ( .A(n_567), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g604 ( .A(n_567), .B(n_605), .Y(n_604) );
AND2x2_ASAP7_75t_L g616 ( .A(n_567), .B(n_617), .Y(n_616) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_567), .B(n_610), .Y(n_652) );
OR2x2_ASAP7_75t_L g659 ( .A(n_567), .B(n_584), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_567), .B(n_669), .Y(n_668) );
AND2x2_ASAP7_75t_L g709 ( .A(n_567), .B(n_695), .Y(n_709) );
OAI22xp33_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_571), .B1(n_575), .B2(n_577), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
AND2x2_ASAP7_75t_L g615 ( .A(n_570), .B(n_616), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_572), .B(n_574), .Y(n_571) );
INVx1_ASAP7_75t_SL g572 ( .A(n_573), .Y(n_572) );
OAI22xp33_ASAP7_75t_L g655 ( .A1(n_573), .A2(n_588), .B1(n_656), .B2(n_660), .Y(n_655) );
INVx1_ASAP7_75t_L g703 ( .A(n_574), .Y(n_703) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g614 ( .A1(n_578), .A2(n_615), .B1(n_618), .B2(n_619), .C(n_620), .Y(n_614) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OR2x2_ASAP7_75t_L g593 ( .A(n_579), .B(n_594), .Y(n_593) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
INVx1_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_583), .B(n_649), .Y(n_681) );
HB1xp67_ASAP7_75t_L g601 ( .A(n_584), .Y(n_601) );
INVx1_ASAP7_75t_L g605 ( .A(n_584), .Y(n_605) );
NAND2xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_588), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
INVx1_ASAP7_75t_L g623 ( .A(n_590), .Y(n_623) );
AND2x2_ASAP7_75t_L g632 ( .A(n_590), .B(n_633), .Y(n_632) );
NAND2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
INVx2_ASAP7_75t_SL g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AND2x2_ASAP7_75t_L g676 ( .A(n_597), .B(n_677), .Y(n_676) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
AOI221xp5_ASAP7_75t_L g625 ( .A1(n_600), .A2(n_626), .B1(n_629), .B2(n_632), .C(n_634), .Y(n_625) );
INVx1_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_604), .B(n_661), .Y(n_660) );
AOI21xp33_ASAP7_75t_SL g606 ( .A1(n_607), .A2(n_608), .B(n_611), .Y(n_606) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
CKINVDCx16_ASAP7_75t_R g708 ( .A(n_611), .Y(n_708) );
OR2x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_613), .Y(n_611) );
OR2x2_ASAP7_75t_L g650 ( .A(n_613), .B(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g671 ( .A(n_616), .Y(n_671) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_616), .B(n_676), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_619), .B(n_641), .Y(n_640) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
NAND4xp25_ASAP7_75t_L g624 ( .A(n_625), .B(n_643), .C(n_662), .D(n_675), .Y(n_624) );
INVx1_ASAP7_75t_SL g626 ( .A(n_627), .Y(n_626) );
INVx1_ASAP7_75t_SL g633 ( .A(n_628), .Y(n_633) );
INVxp67_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
OR2x2_ASAP7_75t_L g666 ( .A(n_637), .B(n_642), .Y(n_666) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AOI211xp5_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_647), .C(n_655), .Y(n_643) );
AOI211xp5_ASAP7_75t_L g714 ( .A1(n_645), .A2(n_687), .B(n_715), .C(n_722), .Y(n_714) );
INVx1_ASAP7_75t_SL g674 ( .A(n_646), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_648), .A2(n_650), .B1(n_652), .B2(n_653), .Y(n_647) );
INVx1_ASAP7_75t_L g678 ( .A(n_652), .Y(n_678) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_657), .B(n_658), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_658), .B(n_695), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_658), .B(n_669), .Y(n_702) );
INVx2_ASAP7_75t_SL g658 ( .A(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
INVx1_ASAP7_75t_L g679 ( .A(n_669), .Y(n_679) );
AOI21xp33_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_672), .B(n_674), .Y(n_670) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
AOI322xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_678), .A3(n_679), .B1(n_680), .B2(n_682), .C1(n_684), .C2(n_687), .Y(n_675) );
INVxp67_ASAP7_75t_L g680 ( .A(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NAND3xp33_ASAP7_75t_SL g689 ( .A(n_690), .B(n_707), .C(n_714), .Y(n_689) );
AOI221xp5_ASAP7_75t_L g690 ( .A1(n_691), .A2(n_693), .B1(n_696), .B2(n_698), .C(n_700), .Y(n_690) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g706 ( .A(n_695), .Y(n_706) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVxp67_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
OAI22xp33_ASAP7_75t_L g700 ( .A1(n_701), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_706), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_708), .A2(n_709), .B1(n_710), .B2(n_711), .C(n_712), .Y(n_707) );
NAND2xp33_ASAP7_75t_L g715 ( .A(n_716), .B(n_717), .Y(n_715) );
INVxp67_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx2_ASAP7_75t_L g734 ( .A(n_727), .Y(n_734) );
INVx1_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx3_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVxp67_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
HB1xp67_ASAP7_75t_L g741 ( .A(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_SL g747 ( .A(n_748), .Y(n_747) );
endmodule