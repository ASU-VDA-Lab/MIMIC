module fake_jpeg_25605_n_341 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_18;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_9),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

BUFx8_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_16),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_36),
.B(n_37),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_33),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_38),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_33),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_45),
.Y(n_58)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_41),
.Y(n_51)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_14),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_17),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_46),
.B(n_47),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_20),
.Y(n_47)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_53),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_42),
.A2(n_26),
.B1(n_19),
.B2(n_17),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_54),
.A2(n_42),
.B1(n_41),
.B2(n_38),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_55),
.Y(n_75)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_56),
.Y(n_79)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_65),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_40),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_66),
.B(n_68),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_36),
.B(n_46),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_67),
.B(n_21),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_40),
.Y(n_68)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_69),
.Y(n_125)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_77),
.Y(n_111)
);

BUFx10_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx5_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_37),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_76),
.B(n_82),
.Y(n_124)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_78),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_48),
.B(n_58),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_63),
.Y(n_83)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_83),
.Y(n_135)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_53),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_84),
.B(n_88),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_57),
.A2(n_26),
.B1(n_36),
.B2(n_37),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_85),
.A2(n_87),
.B1(n_92),
.B2(n_93),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_86),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_57),
.A2(n_26),
.B1(n_38),
.B2(n_41),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_60),
.B(n_47),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_47),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

OA22x2_ASAP7_75t_SL g90 ( 
.A1(n_61),
.A2(n_41),
.B1(n_38),
.B2(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_90),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_46),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_91),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_57),
.A2(n_21),
.B1(n_24),
.B2(n_30),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_63),
.B(n_45),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g94 ( 
.A(n_49),
.Y(n_94)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_94),
.Y(n_120)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_59),
.B(n_45),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_95),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_65),
.Y(n_96)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

INVx5_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx3_ASAP7_75t_L g128 ( 
.A(n_97),
.Y(n_128)
);

CKINVDCx12_ASAP7_75t_R g98 ( 
.A(n_49),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_98),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_55),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_55),
.Y(n_100)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_100),
.Y(n_121)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_64),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_59),
.Y(n_103)
);

AND2x2_ASAP7_75t_SL g105 ( 
.A(n_64),
.B(n_43),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_43),
.C(n_44),
.Y(n_115)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_106),
.B(n_108),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_48),
.A2(n_42),
.B1(n_41),
.B2(n_21),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_107),
.A2(n_102),
.B1(n_90),
.B2(n_83),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_20),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_62),
.B(n_22),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_29),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_130),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_115),
.B(n_133),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_43),
.C(n_44),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_117),
.B(n_86),
.C(n_81),
.Y(n_147)
);

XOR2xp5_ASAP7_75t_L g123 ( 
.A(n_67),
.B(n_22),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_132),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_43),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_138),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g132 ( 
.A(n_92),
.B(n_24),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_105),
.B(n_44),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_105),
.B(n_19),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_140),
.B(n_28),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_124),
.B(n_74),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_141),
.B(n_161),
.Y(n_183)
);

OA22x2_ASAP7_75t_SL g142 ( 
.A1(n_113),
.A2(n_90),
.B1(n_87),
.B2(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_142),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_133),
.A2(n_0),
.B(n_1),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_140),
.B(n_110),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_113),
.A2(n_70),
.B1(n_104),
.B2(n_71),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_144),
.A2(n_158),
.B1(n_163),
.B2(n_136),
.Y(n_174)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_146),
.B(n_149),
.Y(n_172)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_138),
.Y(n_178)
);

INVx13_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_134),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_151),
.B(n_159),
.Y(n_182)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_111),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_152),
.B(n_157),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g153 ( 
.A1(n_116),
.A2(n_70),
.B1(n_104),
.B2(n_97),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_153),
.A2(n_164),
.B1(n_23),
.B2(n_28),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_116),
.A2(n_101),
.B1(n_73),
.B2(n_75),
.Y(n_154)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_154),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_139),
.A2(n_75),
.B1(n_80),
.B2(n_73),
.Y(n_158)
);

INVx13_ASAP7_75t_L g159 ( 
.A(n_135),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_160),
.B(n_166),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_112),
.B(n_94),
.Y(n_161)
);

OAI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_137),
.A2(n_80),
.B1(n_84),
.B2(n_100),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_162),
.A2(n_134),
.B1(n_128),
.B2(n_114),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g163 ( 
.A1(n_139),
.A2(n_72),
.B1(n_106),
.B2(n_19),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_137),
.A2(n_30),
.B1(n_24),
.B2(n_32),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_112),
.B(n_94),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_165),
.B(n_25),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_115),
.Y(n_166)
);

AND2x6_ASAP7_75t_L g167 ( 
.A(n_123),
.B(n_14),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_167),
.B(n_11),
.Y(n_201)
);

BUFx24_ASAP7_75t_L g168 ( 
.A(n_125),
.Y(n_168)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_168),
.Y(n_181)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_122),
.Y(n_169)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_171),
.B(n_189),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_174),
.A2(n_175),
.B1(n_184),
.B2(n_190),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_155),
.A2(n_117),
.B1(n_131),
.B2(n_132),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_176),
.A2(n_177),
.B(n_180),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_SL g177 ( 
.A(n_156),
.B(n_118),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_178),
.B(n_188),
.C(n_195),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_143),
.A2(n_114),
.B1(n_128),
.B2(n_125),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_179),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_155),
.A2(n_129),
.B(n_119),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_155),
.A2(n_129),
.B1(n_119),
.B2(n_121),
.Y(n_184)
);

OAI22x1_ASAP7_75t_L g186 ( 
.A1(n_163),
.A2(n_72),
.B1(n_34),
.B2(n_130),
.Y(n_186)
);

OA21x2_ASAP7_75t_L g230 ( 
.A1(n_186),
.A2(n_199),
.B(n_34),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_156),
.B(n_127),
.C(n_121),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_144),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_79),
.B1(n_30),
.B2(n_127),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_158),
.A2(n_32),
.B1(n_29),
.B2(n_28),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_191),
.A2(n_194),
.B1(n_202),
.B2(n_169),
.Y(n_211)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_193),
.B(n_164),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_142),
.A2(n_145),
.B1(n_160),
.B2(n_163),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_147),
.B(n_22),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_200),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_148),
.B(n_35),
.C(n_27),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_151),
.C(n_150),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_163),
.A2(n_165),
.B(n_161),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_141),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_200),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_142),
.A2(n_23),
.B1(n_18),
.B2(n_27),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_192),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_203),
.B(n_216),
.Y(n_238)
);

CKINVDCx12_ASAP7_75t_R g204 ( 
.A(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_204),
.B(n_208),
.Y(n_254)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_182),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_209),
.B(n_213),
.Y(n_234)
);

OAI32xp33_ASAP7_75t_L g210 ( 
.A1(n_173),
.A2(n_142),
.A3(n_167),
.B1(n_152),
.B2(n_148),
.Y(n_210)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_210),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_211),
.A2(n_222),
.B1(n_227),
.B2(n_185),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_212),
.B(n_230),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_199),
.B(n_169),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_172),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_214),
.B(n_221),
.Y(n_249)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_183),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_218),
.B(n_232),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g219 ( 
.A(n_180),
.B(n_146),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

INVx5_ASAP7_75t_L g220 ( 
.A(n_186),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_183),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_173),
.A2(n_194),
.B1(n_174),
.B2(n_184),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_187),
.B(n_159),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_223),
.B(n_224),
.Y(n_250)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_170),
.Y(n_224)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_190),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_229),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_175),
.A2(n_159),
.B1(n_149),
.B2(n_151),
.Y(n_227)
);

INVx13_ASAP7_75t_L g228 ( 
.A(n_192),
.Y(n_228)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_228),
.Y(n_245)
);

OAI31xp33_ASAP7_75t_L g229 ( 
.A1(n_202),
.A2(n_31),
.A3(n_149),
.B(n_34),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_197),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_197),
.B(n_198),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_178),
.C(n_195),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_241),
.C(n_209),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_235),
.A2(n_237),
.B1(n_243),
.B2(n_252),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_185),
.B1(n_176),
.B2(n_188),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_206),
.B(n_196),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_248),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_212),
.B(n_181),
.C(n_191),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_205),
.A2(n_181),
.B1(n_168),
.B2(n_23),
.Y(n_243)
);

OAI32xp33_ASAP7_75t_L g247 ( 
.A1(n_226),
.A2(n_18),
.A3(n_35),
.B1(n_27),
.B2(n_168),
.Y(n_247)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_247),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_225),
.B(n_210),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_205),
.A2(n_168),
.B1(n_35),
.B2(n_18),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_213),
.A2(n_0),
.B(n_1),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_253),
.A2(n_230),
.B(n_208),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_25),
.C(n_18),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_255),
.B(n_31),
.Y(n_275)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_258),
.B(n_266),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_260),
.A2(n_265),
.B1(n_269),
.B2(n_271),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_256),
.A2(n_219),
.B(n_230),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_261),
.A2(n_276),
.B(n_253),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_246),
.A2(n_256),
.B1(n_239),
.B2(n_220),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_207),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_236),
.A2(n_215),
.B1(n_217),
.B2(n_207),
.Y(n_264)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_264),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_235),
.A2(n_211),
.B1(n_227),
.B2(n_215),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_250),
.B(n_223),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_242),
.B(n_214),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_267),
.B(n_270),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_251),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_244),
.A2(n_208),
.B1(n_229),
.B2(n_203),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g271 ( 
.A(n_234),
.B(n_251),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_244),
.A2(n_228),
.B1(n_35),
.B2(n_25),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_272),
.B(n_274),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_233),
.B(n_31),
.C(n_13),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_273),
.B(n_255),
.C(n_241),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_237),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_275),
.B(n_31),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_249),
.B(n_2),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_278),
.B(n_275),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_257),
.A2(n_254),
.B1(n_248),
.B2(n_252),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_279),
.A2(n_272),
.B1(n_276),
.B2(n_5),
.Y(n_307)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_281),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_240),
.C(n_234),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_283),
.B(n_289),
.C(n_31),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_285),
.B(n_286),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_SL g286 ( 
.A(n_259),
.B(n_243),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_259),
.B(n_245),
.C(n_247),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_13),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_294),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_293),
.B(n_295),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_260),
.B(n_13),
.Y(n_294)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_273),
.B(n_12),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_257),
.B1(n_277),
.B2(n_265),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_296),
.A2(n_304),
.B1(n_308),
.B2(n_294),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_280),
.A2(n_271),
.B1(n_277),
.B2(n_269),
.Y(n_298)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_298),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_291),
.B(n_258),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_299),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_300),
.B(n_307),
.Y(n_319)
);

INVx2_ASAP7_75t_R g303 ( 
.A(n_286),
.Y(n_303)
);

OAI21xp33_ASAP7_75t_L g313 ( 
.A1(n_303),
.A2(n_292),
.B(n_283),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_288),
.A2(n_274),
.B1(n_266),
.B2(n_263),
.Y(n_304)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_282),
.A2(n_284),
.B(n_285),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_306),
.B(n_309),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_279),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_302),
.A2(n_290),
.B1(n_289),
.B2(n_278),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_311),
.B(n_317),
.C(n_305),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_312),
.Y(n_327)
);

INVxp33_ASAP7_75t_L g325 ( 
.A(n_313),
.Y(n_325)
);

BUFx24_ASAP7_75t_SL g316 ( 
.A(n_297),
.Y(n_316)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_316),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_296),
.A2(n_295),
.B1(n_12),
.B2(n_7),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_309),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g321 ( 
.A1(n_318),
.A2(n_303),
.B1(n_308),
.B2(n_301),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_321),
.A2(n_322),
.B1(n_5),
.B2(n_6),
.Y(n_332)
);

OAI21x1_ASAP7_75t_SL g322 ( 
.A1(n_313),
.A2(n_298),
.B(n_301),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_297),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_326),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_315),
.C(n_318),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_310),
.B(n_305),
.Y(n_326)
);

OAI31xp67_ASAP7_75t_L g328 ( 
.A1(n_327),
.A2(n_314),
.A3(n_312),
.B(n_304),
.Y(n_328)
);

NOR2x1_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_332),
.Y(n_334)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_329),
.B(n_330),
.Y(n_333)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_12),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_333),
.B(n_330),
.Y(n_335)
);

NOR2x1_ASAP7_75t_SL g336 ( 
.A(n_335),
.B(n_334),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_331),
.B(n_327),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_337),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_338),
.B(n_328),
.C(n_320),
.Y(n_339)
);

AOI321xp33_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_325),
.A3(n_7),
.B1(n_8),
.B2(n_10),
.C(n_6),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_6),
.B(n_8),
.Y(n_341)
);


endmodule