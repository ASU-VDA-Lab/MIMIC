module real_jpeg_22688_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx13_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_1),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_1),
.A2(n_25),
.B1(n_27),
.B2(n_169),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_1),
.A2(n_43),
.B1(n_44),
.B2(n_169),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_1),
.A2(n_48),
.B1(n_49),
.B2(n_169),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_137),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_3),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_3),
.A2(n_25),
.B1(n_27),
.B2(n_137),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_137),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_3),
.A2(n_43),
.B1(n_44),
.B2(n_137),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_4),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_24),
.Y(n_195)
);

AOI21xp33_ASAP7_75t_L g217 ( 
.A1(n_4),
.A2(n_12),
.B(n_49),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_4),
.A2(n_43),
.B1(n_44),
.B2(n_167),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_4),
.A2(n_81),
.B1(n_83),
.B2(n_226),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_4),
.B(n_199),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_4),
.B(n_27),
.Y(n_250)
);

AOI21xp33_ASAP7_75t_L g254 ( 
.A1(n_4),
.A2(n_27),
.B(n_250),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_5),
.B(n_48),
.Y(n_82)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_5),
.Y(n_83)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_5),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_6),
.A2(n_43),
.B1(n_44),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_6),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_6),
.A2(n_48),
.B1(n_49),
.B2(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_6),
.A2(n_25),
.B1(n_27),
.B2(n_53),
.Y(n_105)
);

BUFx8_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_8),
.A2(n_25),
.B1(n_27),
.B2(n_163),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_8),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_163),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_163),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_8),
.A2(n_43),
.B1(n_44),
.B2(n_163),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_9),
.A2(n_25),
.B1(n_27),
.B2(n_65),
.Y(n_64)
);

CKINVDCx14_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_9),
.A2(n_43),
.B1(n_44),
.B2(n_65),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_65),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_9),
.A2(n_48),
.B1(n_49),
.B2(n_65),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g28 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_11),
.A2(n_25),
.B1(n_27),
.B2(n_32),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_11),
.A2(n_32),
.B1(n_43),
.B2(n_44),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_11),
.A2(n_32),
.B1(n_48),
.B2(n_49),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g42 ( 
.A1(n_12),
.A2(n_43),
.B(n_46),
.C(n_47),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_12),
.B(n_43),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_12),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_13),
.A2(n_25),
.B1(n_26),
.B2(n_27),
.Y(n_24)
);

INVx13_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

OAI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_14),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_35),
.Y(n_67)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_14),
.A2(n_35),
.B1(n_43),
.B2(n_44),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_14),
.A2(n_35),
.B1(n_48),
.B2(n_49),
.Y(n_128)
);

INVx11_ASAP7_75t_SL g45 ( 
.A(n_15),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_114),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_112),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_95),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_19),
.B(n_95),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_68),
.C(n_77),
.Y(n_19)
);

FAx1_ASAP7_75t_SL g141 ( 
.A(n_20),
.B(n_68),
.CI(n_77),
.CON(n_141),
.SN(n_141)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_38),
.B2(n_39),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_21),
.A2(n_22),
.B1(n_97),
.B2(n_110),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_22),
.B(n_40),
.C(n_55),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_28),
.B(n_33),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_23),
.A2(n_28),
.B1(n_91),
.B2(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_23),
.A2(n_91),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_23),
.A2(n_91),
.B1(n_136),
.B2(n_180),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

O2A1O1Ixp33_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_26),
.B(n_30),
.C(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_24),
.B(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_24),
.B(n_93),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_24),
.A2(n_36),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_25),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_25),
.A2(n_37),
.B1(n_166),
.B2(n_173),
.Y(n_172)
);

AOI32xp33_ASAP7_75t_L g249 ( 
.A1(n_25),
.A2(n_43),
.A3(n_62),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_26),
.B(n_30),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_26),
.B(n_27),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_27),
.A2(n_58),
.B(n_60),
.C(n_61),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_27),
.B(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

HAxp5_ASAP7_75t_SL g166 ( 
.A(n_30),
.B(n_167),
.CON(n_166),
.SN(n_166)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_36),
.Y(n_33)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g39 ( 
.A1(n_40),
.A2(n_41),
.B1(n_54),
.B2(n_55),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_40),
.A2(n_41),
.B1(n_102),
.B2(n_108),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

AOI21xp5_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_47),
.B(n_51),
.Y(n_41)
);

INVxp67_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_87),
.B(n_88),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_42),
.A2(n_47),
.B1(n_87),
.B2(n_133),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_42),
.A2(n_51),
.B(n_88),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_42),
.A2(n_47),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_42),
.A2(n_47),
.B1(n_221),
.B2(n_241),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_42),
.A2(n_47),
.B1(n_241),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_42),
.A2(n_72),
.B(n_257),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_43),
.A2(n_44),
.B1(n_58),
.B2(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_44),
.A2(n_50),
.B(n_167),
.C(n_217),
.Y(n_216)
);

NAND2xp33_ASAP7_75t_SL g251 ( 
.A(n_44),
.B(n_58),
.Y(n_251)
);

INVx11_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_47),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_47),
.A2(n_74),
.B(n_133),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_47),
.B(n_167),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_48),
.B(n_230),
.Y(n_229)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_52),
.B(n_73),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_63),
.B(n_66),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_56),
.B(n_107),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_56),
.A2(n_104),
.B(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_56),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_56),
.A2(n_66),
.B(n_296),
.Y(n_295)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_57),
.A2(n_61),
.B1(n_64),
.B2(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_57),
.A2(n_61),
.B1(n_162),
.B2(n_164),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_57),
.A2(n_61),
.B1(n_198),
.B2(n_254),
.Y(n_253)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_61),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_61),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_61),
.A2(n_70),
.B(n_106),
.Y(n_140)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_61),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_64),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_67),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g121 ( 
.A1(n_68),
.A2(n_69),
.B(n_71),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_74),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_73),
.B(n_75),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_89),
.B(n_90),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_78),
.A2(n_79),
.B1(n_118),
.B2(n_119),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_86),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_80),
.A2(n_89),
.B1(n_90),
.B2(n_120),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g309 ( 
.A1(n_80),
.A2(n_86),
.B1(n_89),
.B2(n_310),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_83),
.B(n_84),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_81),
.A2(n_152),
.B(n_153),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_81),
.A2(n_83),
.B1(n_152),
.B2(n_175),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_81),
.A2(n_131),
.B1(n_210),
.B2(n_226),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_81),
.A2(n_129),
.B(n_213),
.Y(n_242)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_82),
.B(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_82),
.A2(n_209),
.B1(n_211),
.B2(n_212),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_82),
.A2(n_85),
.B(n_154),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_83),
.B(n_128),
.Y(n_154)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_83),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_83),
.B(n_167),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_85),
.B(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g310 ( 
.A(n_86),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_90),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_91),
.A2(n_92),
.B(n_94),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_91),
.A2(n_136),
.B(n_138),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_111),
.Y(n_95)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_109),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_98),
.Y(n_109)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_102),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_106),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_105),
.Y(n_296)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g114 ( 
.A1(n_115),
.A2(n_142),
.B(n_319),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_141),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_116),
.B(n_141),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.C(n_122),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_117),
.B(n_121),
.Y(n_317)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_122),
.A2(n_123),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_123),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_134),
.C(n_139),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_124),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_132),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g286 ( 
.A(n_125),
.B(n_132),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

OAI21x1_ASAP7_75t_SL g193 ( 
.A1(n_126),
.A2(n_175),
.B(n_194),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_130),
.Y(n_194)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_134),
.A2(n_135),
.B1(n_139),
.B2(n_140),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_140),
.Y(n_139)
);

BUFx24_ASAP7_75t_SL g321 ( 
.A(n_141),
.Y(n_321)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_313),
.B(n_318),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_301),
.B(n_312),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_201),
.B(n_280),
.C(n_300),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_185),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_146),
.B(n_185),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_147),
.A2(n_148),
.B1(n_170),
.B2(n_184),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_149),
.B(n_157),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_149),
.B(n_157),
.C(n_184),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_150),
.A2(n_151),
.B1(n_155),
.B2(n_156),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_150),
.B(n_156),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_155),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_160),
.C(n_165),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_158),
.A2(n_159),
.B1(n_160),
.B2(n_161),
.Y(n_187)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_162),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_164),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_165),
.B(n_187),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_168),
.Y(n_179)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_170),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_176),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_171),
.B(n_177),
.C(n_182),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_174),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_181),
.B2(n_182),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g181 ( 
.A(n_182),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_188),
.C(n_190),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_186),
.B(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_188),
.A2(n_189),
.B1(n_190),
.B2(n_191),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_191),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_195),
.C(n_196),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_192),
.A2(n_193),
.B1(n_195),
.B2(n_268),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_195),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g266 ( 
.A(n_196),
.B(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_279),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_274),
.B(n_278),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_262),
.B(n_273),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_244),
.B(n_261),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_233),
.B(n_243),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_222),
.B(n_232),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_214),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_208),
.B(n_214),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_215),
.A2(n_216),
.B1(n_218),
.B2(n_219),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_216),
.B(n_218),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_227),
.B(n_231),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_225),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_224),
.B(n_225),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_234),
.B(n_235),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_246),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_252),
.B1(n_259),
.B2(n_260),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_247),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_252),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g252 ( 
.A1(n_253),
.A2(n_255),
.B1(n_256),
.B2(n_258),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_253),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_255),
.B(n_258),
.C(n_259),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_263),
.B(n_264),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_269),
.B2(n_270),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_265),
.B(n_271),
.C(n_272),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_266),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_270),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_275),
.B(n_276),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_281),
.B(n_282),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_298),
.B2(n_299),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g284 ( 
.A1(n_285),
.A2(n_286),
.B1(n_287),
.B2(n_288),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_285),
.B(n_288),
.C(n_299),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_286),
.Y(n_285)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_291),
.B2(n_297),
.Y(n_288)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_289),
.Y(n_297)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_292),
.A2(n_293),
.B1(n_294),
.B2(n_295),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_292),
.B(n_295),
.C(n_297),
.Y(n_311)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_303),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_302),
.B(n_303),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_311),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_305),
.A2(n_306),
.B1(n_308),
.B2(n_309),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_305),
.B(n_309),
.C(n_311),
.Y(n_314)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

CKINVDCx14_ASAP7_75t_R g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g318 ( 
.A(n_314),
.B(n_315),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);


endmodule