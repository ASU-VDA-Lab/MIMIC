module real_aes_336_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_287;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_754;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_713;
wire n_735;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_300;
wire n_252;
wire n_741;
wire n_314;
wire n_283;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_183;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_762;
wire n_210;
wire n_212;
wire n_325;
wire n_575;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_639;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g251 ( .A(n_0), .B(n_158), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g116 ( .A(n_1), .B(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_2), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_3), .B(n_147), .Y(n_522) );
NAND2xp5_ASAP7_75t_L g486 ( .A(n_4), .B(n_156), .Y(n_486) );
INVx1_ASAP7_75t_L g146 ( .A(n_5), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_6), .B(n_147), .Y(n_204) );
NAND2xp33_ASAP7_75t_SL g197 ( .A(n_7), .B(n_153), .Y(n_197) );
INVx1_ASAP7_75t_L g177 ( .A(n_8), .Y(n_177) );
CKINVDCx16_ASAP7_75t_R g117 ( .A(n_9), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g748 ( .A(n_10), .Y(n_748) );
AND2x2_ASAP7_75t_L g202 ( .A(n_11), .B(n_137), .Y(n_202) );
AND2x2_ASAP7_75t_L g479 ( .A(n_12), .B(n_194), .Y(n_479) );
AND2x2_ASAP7_75t_L g488 ( .A(n_13), .B(n_169), .Y(n_488) );
INVx2_ASAP7_75t_L g138 ( .A(n_14), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_15), .B(n_156), .Y(n_541) );
CKINVDCx16_ASAP7_75t_R g109 ( .A(n_16), .Y(n_109) );
AOI221x1_ASAP7_75t_L g191 ( .A1(n_17), .A2(n_141), .B1(n_192), .B2(n_194), .C(n_196), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g164 ( .A(n_18), .B(n_147), .Y(n_164) );
NAND2xp5_ASAP7_75t_SL g526 ( .A(n_19), .B(n_147), .Y(n_526) );
INVx1_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_21), .A2(n_90), .B1(n_147), .B2(n_179), .Y(n_467) );
AOI221xp5_ASAP7_75t_SL g140 ( .A1(n_22), .A2(n_37), .B1(n_141), .B2(n_147), .C(n_154), .Y(n_140) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_23), .A2(n_141), .B(n_206), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_24), .B(n_158), .Y(n_207) );
OR2x2_ASAP7_75t_L g139 ( .A(n_25), .B(n_89), .Y(n_139) );
OA21x2_ASAP7_75t_L g170 ( .A1(n_25), .A2(n_89), .B(n_138), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_26), .B(n_156), .Y(n_168) );
INVxp67_ASAP7_75t_L g190 ( .A(n_27), .Y(n_190) );
AND2x2_ASAP7_75t_L g240 ( .A(n_28), .B(n_136), .Y(n_240) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_29), .A2(n_141), .B(n_250), .Y(n_249) );
AO21x2_ASAP7_75t_L g536 ( .A1(n_30), .A2(n_194), .B(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_31), .B(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_32), .A2(n_141), .B(n_484), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_33), .B(n_156), .Y(n_521) );
AND2x2_ASAP7_75t_L g142 ( .A(n_34), .B(n_143), .Y(n_142) );
AND2x2_ASAP7_75t_L g153 ( .A(n_34), .B(n_146), .Y(n_153) );
INVx1_ASAP7_75t_L g186 ( .A(n_34), .Y(n_186) );
OR2x6_ASAP7_75t_L g111 ( .A(n_35), .B(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g765 ( .A(n_36), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_38), .B(n_147), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g224 ( .A1(n_39), .A2(n_82), .B1(n_141), .B2(n_184), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_40), .B(n_156), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_41), .B(n_147), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_42), .B(n_158), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_43), .A2(n_141), .B(n_475), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_44), .A2(n_72), .B1(n_740), .B2(n_741), .Y(n_739) );
CKINVDCx20_ASAP7_75t_R g740 ( .A(n_44), .Y(n_740) );
AND2x2_ASAP7_75t_L g254 ( .A(n_45), .B(n_136), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_46), .B(n_158), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_47), .B(n_136), .Y(n_160) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_48), .B(n_147), .Y(n_538) );
INVx1_ASAP7_75t_L g145 ( .A(n_49), .Y(n_145) );
INVx1_ASAP7_75t_L g150 ( .A(n_49), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_50), .B(n_156), .Y(n_477) );
AND2x2_ASAP7_75t_L g507 ( .A(n_51), .B(n_136), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_52), .B(n_147), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g476 ( .A(n_53), .B(n_158), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_54), .B(n_158), .Y(n_520) );
AND2x2_ASAP7_75t_L g218 ( .A(n_55), .B(n_136), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g478 ( .A(n_56), .B(n_147), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_57), .B(n_156), .Y(n_252) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_58), .B(n_147), .Y(n_509) );
AOI21xp5_ASAP7_75t_L g518 ( .A1(n_59), .A2(n_141), .B(n_519), .Y(n_518) );
AND2x2_ASAP7_75t_SL g171 ( .A(n_60), .B(n_137), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_61), .B(n_158), .Y(n_215) );
AND2x2_ASAP7_75t_L g532 ( .A(n_62), .B(n_137), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g235 ( .A1(n_63), .A2(n_141), .B(n_236), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_64), .B(n_156), .Y(n_208) );
AND2x2_ASAP7_75t_SL g225 ( .A(n_65), .B(n_169), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_66), .B(n_158), .Y(n_513) );
OAI22xp5_ASAP7_75t_SL g754 ( .A1(n_67), .A2(n_70), .B1(n_755), .B2(n_756), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_67), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_68), .B(n_158), .Y(n_542) );
AOI22xp5_ASAP7_75t_L g468 ( .A1(n_69), .A2(n_92), .B1(n_141), .B2(n_184), .Y(n_468) );
INVx1_ASAP7_75t_L g756 ( .A(n_70), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_71), .B(n_156), .Y(n_529) );
INVx1_ASAP7_75t_L g741 ( .A(n_72), .Y(n_741) );
INVx1_ASAP7_75t_L g143 ( .A(n_73), .Y(n_143) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_74), .B(n_158), .Y(n_485) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_75), .A2(n_141), .B(n_511), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_76), .A2(n_141), .B(n_497), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_77), .A2(n_141), .B(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g523 ( .A(n_78), .B(n_137), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_79), .B(n_136), .Y(n_465) );
NAND2xp5_ASAP7_75t_SL g216 ( .A(n_80), .B(n_147), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g223 ( .A1(n_81), .A2(n_84), .B1(n_147), .B2(n_179), .Y(n_223) );
INVx1_ASAP7_75t_L g114 ( .A(n_83), .Y(n_114) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_85), .B(n_158), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_86), .B(n_158), .Y(n_157) );
AND2x2_ASAP7_75t_L g500 ( .A(n_87), .B(n_169), .Y(n_500) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_88), .A2(n_141), .B(n_213), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_91), .B(n_156), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g527 ( .A1(n_93), .A2(n_141), .B(n_528), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_94), .B(n_156), .Y(n_498) );
INVxp67_ASAP7_75t_L g193 ( .A(n_95), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_96), .B(n_147), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g237 ( .A(n_97), .B(n_156), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g165 ( .A1(n_98), .A2(n_141), .B(n_166), .Y(n_165) );
BUFx2_ASAP7_75t_L g531 ( .A(n_99), .Y(n_531) );
BUFx2_ASAP7_75t_L g122 ( .A(n_100), .Y(n_122) );
BUFx2_ASAP7_75t_SL g752 ( .A(n_100), .Y(n_752) );
AOI21xp5_ASAP7_75t_L g101 ( .A1(n_102), .A2(n_118), .B(n_764), .Y(n_101) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx20_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx1_ASAP7_75t_SL g767 ( .A(n_104), .Y(n_767) );
INVx2_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
NAND2xp5_ASAP7_75t_SL g105 ( .A(n_106), .B(n_115), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_107), .Y(n_106) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
BUFx3_ASAP7_75t_L g126 ( .A(n_108), .Y(n_126) );
BUFx2_ASAP7_75t_L g763 ( .A(n_108), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_109), .B(n_110), .Y(n_108) );
AND2x6_ASAP7_75t_SL g450 ( .A(n_109), .B(n_111), .Y(n_450) );
OR2x6_ASAP7_75t_SL g453 ( .A(n_109), .B(n_110), .Y(n_453) );
OR2x2_ASAP7_75t_L g747 ( .A(n_109), .B(n_111), .Y(n_747) );
CKINVDCx5p33_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
NAND2xp5_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
INVx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OA21x2_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_127), .B(n_749), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_120), .B(n_123), .Y(n_119) );
HB1xp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
HB1xp67_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
OAI21xp5_ASAP7_75t_L g760 ( .A1(n_123), .A2(n_754), .B(n_759), .Y(n_760) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_123), .B(n_762), .Y(n_761) );
BUFx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI222xp33_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_738), .B1(n_739), .B2(n_742), .C1(n_745), .C2(n_748), .Y(n_127) );
OA22x2_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_447), .B1(n_451), .B2(n_454), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
OAI22xp5_ASAP7_75t_SL g743 ( .A1(n_130), .A2(n_451), .B1(n_455), .B2(n_744), .Y(n_743) );
INVx4_ASAP7_75t_L g759 ( .A(n_130), .Y(n_759) );
OR2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_360), .Y(n_130) );
NAND3xp33_ASAP7_75t_SL g131 ( .A(n_132), .B(n_270), .C(n_310), .Y(n_131) );
O2A1O1Ixp33_ASAP7_75t_L g132 ( .A1(n_133), .A2(n_172), .B(n_199), .C(n_226), .Y(n_132) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_133), .B(n_275), .Y(n_309) );
NOR2x1p5_ASAP7_75t_L g133 ( .A(n_134), .B(n_161), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g245 ( .A(n_135), .Y(n_245) );
INVx2_ASAP7_75t_L g261 ( .A(n_135), .Y(n_261) );
OR2x2_ASAP7_75t_L g273 ( .A(n_135), .B(n_162), .Y(n_273) );
AND2x2_ASAP7_75t_L g287 ( .A(n_135), .B(n_246), .Y(n_287) );
INVx1_ASAP7_75t_L g315 ( .A(n_135), .Y(n_315) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_135), .Y(n_376) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_135), .B(n_162), .Y(n_421) );
OA21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_160), .Y(n_135) );
CKINVDCx5p33_ASAP7_75t_R g217 ( .A(n_136), .Y(n_217) );
AO21x2_ASAP7_75t_L g466 ( .A1(n_136), .A2(n_467), .B(n_468), .Y(n_466) );
AOI21xp5_ASAP7_75t_L g494 ( .A1(n_136), .A2(n_495), .B(n_496), .Y(n_494) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
AND2x2_ASAP7_75t_SL g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x4_ASAP7_75t_L g178 ( .A(n_138), .B(n_139), .Y(n_178) );
AND2x6_ASAP7_75t_L g141 ( .A(n_142), .B(n_144), .Y(n_141) );
BUFx3_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
AND2x6_ASAP7_75t_L g158 ( .A(n_143), .B(n_149), .Y(n_158) );
INVx2_ASAP7_75t_L g188 ( .A(n_143), .Y(n_188) );
AND2x4_ASAP7_75t_L g184 ( .A(n_144), .B(n_185), .Y(n_184) );
AND2x2_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
AND2x4_ASAP7_75t_L g156 ( .A(n_145), .B(n_151), .Y(n_156) );
INVx2_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
HB1xp67_ASAP7_75t_L g182 ( .A(n_146), .Y(n_182) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
INVx1_ASAP7_75t_L g198 ( .A(n_148), .Y(n_198) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g159 ( .A(n_153), .Y(n_159) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_157), .B(n_159), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_158), .B(n_531), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g166 ( .A1(n_159), .A2(n_167), .B(n_168), .Y(n_166) );
AOI21xp5_ASAP7_75t_L g206 ( .A1(n_159), .A2(n_207), .B(n_208), .Y(n_206) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_159), .A2(n_214), .B(n_215), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g236 ( .A1(n_159), .A2(n_237), .B(n_238), .Y(n_236) );
AOI21xp5_ASAP7_75t_L g250 ( .A1(n_159), .A2(n_251), .B(n_252), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_159), .A2(n_476), .B(n_477), .Y(n_475) );
AOI21xp5_ASAP7_75t_L g484 ( .A1(n_159), .A2(n_485), .B(n_486), .Y(n_484) );
AOI21xp5_ASAP7_75t_L g497 ( .A1(n_159), .A2(n_498), .B(n_499), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_159), .A2(n_512), .B(n_513), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_159), .A2(n_520), .B(n_521), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g528 ( .A1(n_159), .A2(n_529), .B(n_530), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g540 ( .A1(n_159), .A2(n_541), .B(n_542), .Y(n_540) );
OR2x2_ASAP7_75t_L g242 ( .A(n_161), .B(n_243), .Y(n_242) );
HB1xp67_ASAP7_75t_L g377 ( .A(n_161), .Y(n_377) );
AND2x2_ASAP7_75t_L g382 ( .A(n_161), .B(n_244), .Y(n_382) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
AND2x4_ASAP7_75t_L g172 ( .A(n_162), .B(n_173), .Y(n_172) );
OR2x2_ASAP7_75t_L g241 ( .A(n_162), .B(n_174), .Y(n_241) );
OR2x2_ASAP7_75t_L g260 ( .A(n_162), .B(n_261), .Y(n_260) );
INVx2_ASAP7_75t_L g289 ( .A(n_162), .Y(n_289) );
AND2x4_ASAP7_75t_SL g328 ( .A(n_162), .B(n_174), .Y(n_328) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_162), .Y(n_332) );
OR2x2_ASAP7_75t_L g349 ( .A(n_162), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g359 ( .A(n_162), .B(n_266), .Y(n_359) );
INVx1_ASAP7_75t_L g388 ( .A(n_162), .Y(n_388) );
OR2x6_ASAP7_75t_L g162 ( .A(n_163), .B(n_171), .Y(n_162) );
AOI21xp5_ASAP7_75t_L g163 ( .A1(n_164), .A2(n_165), .B(n_169), .Y(n_163) );
INVx2_ASAP7_75t_SL g221 ( .A(n_169), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_169), .A2(n_526), .B(n_527), .Y(n_525) );
BUFx4f_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx3_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_172), .B(n_317), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g263 ( .A(n_173), .B(n_246), .Y(n_263) );
AND2x2_ASAP7_75t_L g275 ( .A(n_173), .B(n_276), .Y(n_275) );
OR2x2_ASAP7_75t_L g293 ( .A(n_173), .B(n_260), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_173), .B(n_314), .Y(n_313) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
AND2x4_ASAP7_75t_L g266 ( .A(n_174), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g288 ( .A(n_174), .B(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g323 ( .A(n_174), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g347 ( .A(n_174), .B(n_246), .Y(n_347) );
AND2x4_ASAP7_75t_L g174 ( .A(n_175), .B(n_191), .Y(n_174) );
AOI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_179), .B1(n_184), .B2(n_189), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_178), .B(n_190), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g192 ( .A(n_178), .B(n_193), .Y(n_192) );
NOR3xp33_ASAP7_75t_L g196 ( .A(n_178), .B(n_197), .C(n_198), .Y(n_196) );
AOI21xp5_ASAP7_75t_L g203 ( .A1(n_178), .A2(n_204), .B(n_205), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_178), .A2(n_509), .B(n_510), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_178), .A2(n_538), .B(n_539), .Y(n_537) );
AND2x4_ASAP7_75t_L g179 ( .A(n_180), .B(n_183), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
NOR2x1p5_ASAP7_75t_L g185 ( .A(n_186), .B(n_187), .Y(n_185) );
INVx3_ASAP7_75t_L g187 ( .A(n_188), .Y(n_187) );
INVx3_ASAP7_75t_L g516 ( .A(n_194), .Y(n_516) );
INVx4_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
AOI21x1_ASAP7_75t_L g247 ( .A1(n_195), .A2(n_248), .B(n_254), .Y(n_247) );
AO21x2_ASAP7_75t_L g472 ( .A1(n_195), .A2(n_473), .B(n_479), .Y(n_472) );
AND2x2_ASAP7_75t_L g199 ( .A(n_200), .B(n_209), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_200), .B(n_279), .Y(n_278) );
AND2x4_ASAP7_75t_L g296 ( .A(n_200), .B(n_297), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_200), .B(n_210), .Y(n_301) );
NAND3xp33_ASAP7_75t_L g316 ( .A(n_200), .B(n_317), .C(n_318), .Y(n_316) );
AND2x2_ASAP7_75t_L g364 ( .A(n_200), .B(n_269), .Y(n_364) );
INVx5_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g231 ( .A(n_201), .B(n_232), .Y(n_231) );
AND2x4_ASAP7_75t_SL g268 ( .A(n_201), .B(n_269), .Y(n_268) );
INVx2_ASAP7_75t_L g284 ( .A(n_201), .Y(n_284) );
OR2x2_ASAP7_75t_L g307 ( .A(n_201), .B(n_297), .Y(n_307) );
HB1xp67_ASAP7_75t_L g324 ( .A(n_201), .Y(n_324) );
AND2x2_ASAP7_75t_SL g342 ( .A(n_201), .B(n_230), .Y(n_342) );
AND2x4_ASAP7_75t_L g357 ( .A(n_201), .B(n_233), .Y(n_357) );
AND2x2_ASAP7_75t_L g371 ( .A(n_201), .B(n_210), .Y(n_371) );
OR2x2_ASAP7_75t_L g392 ( .A(n_201), .B(n_219), .Y(n_392) );
OR2x6_ASAP7_75t_L g201 ( .A(n_202), .B(n_203), .Y(n_201) );
AND2x2_ASAP7_75t_L g446 ( .A(n_209), .B(n_324), .Y(n_446) );
AND2x2_ASAP7_75t_L g209 ( .A(n_210), .B(n_219), .Y(n_209) );
AND2x4_ASAP7_75t_L g269 ( .A(n_210), .B(n_232), .Y(n_269) );
INVx2_ASAP7_75t_L g280 ( .A(n_210), .Y(n_280) );
AND2x2_ASAP7_75t_L g285 ( .A(n_210), .B(n_230), .Y(n_285) );
HB1xp67_ASAP7_75t_L g318 ( .A(n_210), .Y(n_318) );
OR2x2_ASAP7_75t_L g341 ( .A(n_210), .B(n_233), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_210), .B(n_233), .Y(n_344) );
INVx1_ASAP7_75t_L g353 ( .A(n_210), .Y(n_353) );
AO21x2_ASAP7_75t_L g210 ( .A1(n_211), .A2(n_217), .B(n_218), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_212), .B(n_216), .Y(n_211) );
AO21x2_ASAP7_75t_L g233 ( .A1(n_217), .A2(n_234), .B(n_240), .Y(n_233) );
AO21x2_ASAP7_75t_L g297 ( .A1(n_217), .A2(n_234), .B(n_240), .Y(n_297) );
AOI21x1_ASAP7_75t_L g481 ( .A1(n_217), .A2(n_482), .B(n_488), .Y(n_481) );
AND2x2_ASAP7_75t_L g256 ( .A(n_219), .B(n_233), .Y(n_256) );
BUFx2_ASAP7_75t_L g305 ( .A(n_219), .Y(n_305) );
AND2x2_ASAP7_75t_L g400 ( .A(n_219), .B(n_280), .Y(n_400) );
INVx2_ASAP7_75t_L g219 ( .A(n_220), .Y(n_219) );
BUFx6f_ASAP7_75t_L g230 ( .A(n_220), .Y(n_230) );
AOI21x1_ASAP7_75t_L g220 ( .A1(n_221), .A2(n_222), .B(n_225), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_223), .B(n_224), .Y(n_222) );
OAI221xp5_ASAP7_75t_L g226 ( .A1(n_227), .A2(n_241), .B1(n_242), .B2(n_255), .C(n_257), .Y(n_226) );
INVx1_ASAP7_75t_SL g227 ( .A(n_228), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_231), .Y(n_228) );
NOR2x1_ASAP7_75t_L g302 ( .A(n_229), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_229), .B(n_296), .Y(n_336) );
OR2x2_ASAP7_75t_L g348 ( .A(n_229), .B(n_344), .Y(n_348) );
OR2x2_ASAP7_75t_L g351 ( .A(n_229), .B(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_L g440 ( .A(n_229), .B(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g229 ( .A(n_230), .Y(n_229) );
AND2x4_ASAP7_75t_L g279 ( .A(n_230), .B(n_280), .Y(n_279) );
OA33x2_ASAP7_75t_L g312 ( .A1(n_230), .A2(n_273), .A3(n_313), .B1(n_316), .B2(n_319), .B3(n_322), .Y(n_312) );
OR2x2_ASAP7_75t_L g343 ( .A(n_230), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g367 ( .A(n_230), .B(n_368), .Y(n_367) );
OR2x2_ASAP7_75t_L g375 ( .A(n_230), .B(n_376), .Y(n_375) );
AND2x2_ASAP7_75t_L g395 ( .A(n_230), .B(n_269), .Y(n_395) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_230), .B(n_284), .Y(n_433) );
INVx2_ASAP7_75t_L g303 ( .A(n_231), .Y(n_303) );
AOI322xp5_ASAP7_75t_L g373 ( .A1(n_231), .A2(n_286), .A3(n_374), .B1(n_377), .B2(n_378), .C1(n_380), .C2(n_382), .Y(n_373) );
INVx2_ASAP7_75t_L g232 ( .A(n_233), .Y(n_232) );
HB1xp67_ASAP7_75t_L g402 ( .A(n_233), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_239), .Y(n_234) );
OR2x2_ASAP7_75t_L g355 ( .A(n_241), .B(n_334), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_241), .B(n_408), .Y(n_407) );
INVx1_ASAP7_75t_SL g428 ( .A(n_241), .Y(n_428) );
INVx1_ASAP7_75t_SL g294 ( .A(n_242), .Y(n_294) );
INVx1_ASAP7_75t_L g243 ( .A(n_244), .Y(n_243) );
AND2x2_ASAP7_75t_L g327 ( .A(n_244), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_246), .Y(n_244) );
INVx2_ASAP7_75t_L g267 ( .A(n_246), .Y(n_267) );
INVx1_ASAP7_75t_L g276 ( .A(n_246), .Y(n_276) );
INVx1_ASAP7_75t_L g317 ( .A(n_246), .Y(n_317) );
OR2x2_ASAP7_75t_L g334 ( .A(n_246), .B(n_261), .Y(n_334) );
HB1xp67_ASAP7_75t_L g409 ( .A(n_246), .Y(n_409) );
INVx3_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_253), .Y(n_248) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_SL g378 ( .A(n_256), .B(n_379), .Y(n_378) );
OAI21xp5_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_264), .B(n_268), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g331 ( .A1(n_258), .A2(n_332), .B(n_333), .C(n_335), .Y(n_331) );
AND2x4_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g396 ( .A(n_260), .B(n_397), .Y(n_396) );
HB1xp67_ASAP7_75t_L g265 ( .A(n_261), .Y(n_265) );
INVx1_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g420 ( .A(n_263), .B(n_421), .Y(n_420) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
AND2x2_ASAP7_75t_SL g389 ( .A(n_266), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g397 ( .A(n_266), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_266), .B(n_388), .Y(n_405) );
INVx3_ASAP7_75t_SL g330 ( .A(n_269), .Y(n_330) );
AOI221xp5_ASAP7_75t_L g270 ( .A1(n_271), .A2(n_277), .B1(n_281), .B2(n_286), .C(n_290), .Y(n_270) );
INVx1_ASAP7_75t_SL g271 ( .A(n_272), .Y(n_271) );
OR2x2_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
HB1xp67_ASAP7_75t_L g321 ( .A(n_276), .Y(n_321) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_279), .A2(n_306), .B(n_378), .Y(n_384) );
AND2x2_ASAP7_75t_L g410 ( .A(n_279), .B(n_357), .Y(n_410) );
HB1xp67_ASAP7_75t_L g298 ( .A(n_280), .Y(n_298) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_283), .B(n_285), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_284), .B(n_400), .Y(n_399) );
OR2x2_ASAP7_75t_L g419 ( .A(n_284), .B(n_341), .Y(n_419) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
INVx2_ASAP7_75t_L g368 ( .A(n_287), .Y(n_368) );
OAI21xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_295), .B(n_299), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx1_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_296), .B(n_298), .Y(n_295) );
INVx2_ASAP7_75t_L g441 ( .A(n_296), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_297), .B(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_L g370 ( .A(n_297), .B(n_371), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_298), .B(n_320), .Y(n_319) );
OAI31xp33_ASAP7_75t_SL g299 ( .A1(n_300), .A2(n_302), .A3(n_304), .B(n_308), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_303), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
OR2x2_ASAP7_75t_L g381 ( .A(n_305), .B(n_307), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_305), .B(n_357), .Y(n_436) );
INVx1_ASAP7_75t_SL g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR5xp2_ASAP7_75t_L g310 ( .A(n_311), .B(n_325), .C(n_337), .D(n_346), .E(n_354), .Y(n_310) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_315), .B(n_317), .Y(n_350) );
INVx1_ASAP7_75t_L g390 ( .A(n_315), .Y(n_390) );
INVxp67_ASAP7_75t_SL g427 ( .A(n_315), .Y(n_427) );
INVx1_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
NAND2xp33_ASAP7_75t_SL g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OAI321xp33_ASAP7_75t_L g362 ( .A1(n_323), .A2(n_363), .A3(n_365), .B1(n_369), .B2(n_372), .C(n_373), .Y(n_362) );
INVx1_ASAP7_75t_L g416 ( .A(n_324), .Y(n_416) );
OAI21xp33_ASAP7_75t_L g325 ( .A1(n_326), .A2(n_329), .B(n_331), .Y(n_325) );
INVx1_ASAP7_75t_SL g326 ( .A(n_327), .Y(n_326) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_327), .A2(n_400), .B1(n_407), .B2(n_410), .Y(n_406) );
AND2x2_ASAP7_75t_L g435 ( .A(n_328), .B(n_409), .Y(n_435) );
INVx1_ASAP7_75t_L g345 ( .A(n_333), .Y(n_345) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_338), .A2(n_343), .B(n_345), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g339 ( .A(n_340), .B(n_342), .Y(n_339) );
INVx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
OAI22xp5_ASAP7_75t_L g354 ( .A1(n_344), .A2(n_355), .B1(n_356), .B2(n_358), .Y(n_354) );
INVx1_ASAP7_75t_L g417 ( .A(n_344), .Y(n_417) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_348), .B1(n_349), .B2(n_351), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_353), .B(n_357), .Y(n_356) );
OAI221xp5_ASAP7_75t_L g431 ( .A1(n_355), .A2(n_432), .B1(n_434), .B2(n_436), .C(n_437), .Y(n_431) );
INVx1_ASAP7_75t_L g438 ( .A(n_355), .Y(n_438) );
OAI221xp5_ASAP7_75t_L g412 ( .A1(n_356), .A2(n_413), .B1(n_420), .B2(n_422), .C(n_423), .Y(n_412) );
OAI21xp5_ASAP7_75t_L g383 ( .A1(n_358), .A2(n_384), .B(n_385), .Y(n_383) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_361), .B(n_411), .Y(n_360) );
NOR3xp33_ASAP7_75t_L g361 ( .A(n_362), .B(n_383), .C(n_401), .Y(n_361) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
HB1xp67_ASAP7_75t_L g430 ( .A(n_364), .Y(n_430) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx1_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g429 ( .A(n_372), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_374), .B(n_404), .Y(n_403) );
INVx1_ASAP7_75t_SL g374 ( .A(n_375), .Y(n_374) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g422 ( .A(n_382), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_391), .B(n_393), .Y(n_385) );
INVxp67_ASAP7_75t_L g443 ( .A(n_386), .Y(n_443) );
AND2x2_ASAP7_75t_L g386 ( .A(n_387), .B(n_389), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx2_ASAP7_75t_SL g398 ( .A(n_389), .Y(n_398) );
INVx1_ASAP7_75t_SL g391 ( .A(n_392), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g393 ( .A1(n_394), .A2(n_396), .B1(n_398), .B2(n_399), .Y(n_393) );
INVx2_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI21xp33_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_403), .B(n_406), .Y(n_401) );
INVx1_ASAP7_75t_SL g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g444 ( .A(n_407), .Y(n_444) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR3xp33_ASAP7_75t_L g411 ( .A(n_412), .B(n_431), .C(n_442), .Y(n_411) );
NOR2xp33_ASAP7_75t_L g413 ( .A(n_414), .B(n_418), .Y(n_413) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
NAND2xp5_ASAP7_75t_SL g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g418 ( .A(n_419), .Y(n_418) );
OAI21xp5_ASAP7_75t_SL g423 ( .A1(n_424), .A2(n_429), .B(n_430), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_428), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
OAI21xp5_ASAP7_75t_L g437 ( .A1(n_435), .A2(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
AOI21xp33_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_445), .Y(n_442) );
INVx1_ASAP7_75t_SL g445 ( .A(n_446), .Y(n_445) );
CKINVDCx6p67_ASAP7_75t_R g447 ( .A(n_448), .Y(n_447) );
INVx4_ASAP7_75t_SL g744 ( .A(n_448), .Y(n_744) );
INVx3_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
CKINVDCx5p33_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
CKINVDCx11_ASAP7_75t_R g452 ( .A(n_453), .Y(n_452) );
INVx4_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OR2x6_ASAP7_75t_L g455 ( .A(n_456), .B(n_675), .Y(n_455) );
NAND3xp33_ASAP7_75t_L g456 ( .A(n_457), .B(n_591), .C(n_628), .Y(n_456) );
NOR3xp33_ASAP7_75t_L g457 ( .A(n_458), .B(n_559), .C(n_574), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_504), .B1(n_533), .B2(n_545), .C(n_546), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_461), .B(n_489), .Y(n_460) );
OAI22xp33_ASAP7_75t_SL g619 ( .A1(n_461), .A2(n_583), .B1(n_620), .B2(n_623), .Y(n_619) );
OR2x2_ASAP7_75t_L g461 ( .A(n_462), .B(n_469), .Y(n_461) );
OAI21xp33_ASAP7_75t_SL g629 ( .A1(n_462), .A2(n_630), .B(n_636), .Y(n_629) );
OR2x2_ASAP7_75t_L g658 ( .A(n_462), .B(n_491), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_462), .B(n_578), .Y(n_659) );
INVx2_ASAP7_75t_L g690 ( .A(n_462), .Y(n_690) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_463), .B(n_550), .Y(n_671) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
OR2x2_ASAP7_75t_L g545 ( .A(n_464), .B(n_472), .Y(n_545) );
BUFx3_ASAP7_75t_L g571 ( .A(n_464), .Y(n_571) );
AND2x2_ASAP7_75t_L g707 ( .A(n_464), .B(n_708), .Y(n_707) );
AND2x2_ASAP7_75t_L g730 ( .A(n_464), .B(n_492), .Y(n_730) );
AND2x4_ASAP7_75t_L g464 ( .A(n_465), .B(n_466), .Y(n_464) );
AND2x4_ASAP7_75t_L g503 ( .A(n_465), .B(n_466), .Y(n_503) );
INVx1_ASAP7_75t_SL g469 ( .A(n_470), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_470), .B(n_492), .Y(n_650) );
INVx1_ASAP7_75t_L g687 ( .A(n_470), .Y(n_687) );
AND2x2_ASAP7_75t_L g470 ( .A(n_471), .B(n_480), .Y(n_470) );
AND2x2_ASAP7_75t_L g502 ( .A(n_471), .B(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g708 ( .A(n_471), .Y(n_708) );
INVx2_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g551 ( .A(n_472), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_472), .B(n_480), .Y(n_552) );
AND2x2_ASAP7_75t_L g573 ( .A(n_472), .B(n_493), .Y(n_573) );
AND2x2_ASAP7_75t_L g655 ( .A(n_472), .B(n_481), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_474), .B(n_478), .Y(n_473) );
AND2x4_ASAP7_75t_SL g548 ( .A(n_480), .B(n_493), .Y(n_548) );
INVx1_ASAP7_75t_L g579 ( .A(n_480), .Y(n_579) );
INVx2_ASAP7_75t_L g587 ( .A(n_480), .Y(n_587) );
HB1xp67_ASAP7_75t_L g611 ( .A(n_480), .Y(n_611) );
INVx3_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_481), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_490), .B(n_502), .Y(n_489) );
AND2x2_ASAP7_75t_L g726 ( .A(n_490), .B(n_589), .Y(n_726) );
INVx1_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_492), .B(n_501), .Y(n_491) );
NAND2x1p5_ASAP7_75t_L g585 ( .A(n_492), .B(n_586), .Y(n_585) );
AND2x2_ASAP7_75t_L g637 ( .A(n_492), .B(n_552), .Y(n_637) );
AND2x2_ASAP7_75t_L g654 ( .A(n_492), .B(n_655), .Y(n_654) );
INVx4_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g578 ( .A(n_493), .B(n_579), .Y(n_578) );
INVx1_ASAP7_75t_L g594 ( .A(n_493), .Y(n_594) );
AND2x2_ASAP7_75t_L g638 ( .A(n_493), .B(n_639), .Y(n_638) );
OR2x2_ASAP7_75t_L g645 ( .A(n_493), .B(n_646), .Y(n_645) );
NOR2x1_ASAP7_75t_L g660 ( .A(n_493), .B(n_551), .Y(n_660) );
BUFx2_ASAP7_75t_L g670 ( .A(n_493), .Y(n_670) );
AND2x2_ASAP7_75t_L g695 ( .A(n_493), .B(n_655), .Y(n_695) );
AND2x2_ASAP7_75t_L g716 ( .A(n_493), .B(n_717), .Y(n_716) );
OR2x6_ASAP7_75t_L g493 ( .A(n_494), .B(n_500), .Y(n_493) );
INVx1_ASAP7_75t_L g647 ( .A(n_501), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_502), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g677 ( .A(n_502), .B(n_548), .Y(n_677) );
INVx3_ASAP7_75t_L g584 ( .A(n_503), .Y(n_584) );
AND2x2_ASAP7_75t_L g717 ( .A(n_503), .B(n_639), .Y(n_717) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
AOI22xp5_ASAP7_75t_L g546 ( .A1(n_505), .A2(n_547), .B1(n_552), .B2(n_553), .Y(n_546) );
AND2x2_ASAP7_75t_L g505 ( .A(n_506), .B(n_514), .Y(n_505) );
INVx4_ASAP7_75t_L g544 ( .A(n_506), .Y(n_544) );
INVx2_ASAP7_75t_L g581 ( .A(n_506), .Y(n_581) );
NAND2x1_ASAP7_75t_L g607 ( .A(n_506), .B(n_524), .Y(n_607) );
OR2x2_ASAP7_75t_L g622 ( .A(n_506), .B(n_557), .Y(n_622) );
OR2x2_ASAP7_75t_SL g649 ( .A(n_506), .B(n_621), .Y(n_649) );
AND2x2_ASAP7_75t_L g662 ( .A(n_506), .B(n_536), .Y(n_662) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_506), .Y(n_683) );
OR2x6_ASAP7_75t_L g506 ( .A(n_507), .B(n_508), .Y(n_506) );
INVx2_ASAP7_75t_L g562 ( .A(n_514), .Y(n_562) );
AND2x2_ASAP7_75t_L g694 ( .A(n_514), .B(n_668), .Y(n_694) );
NOR2x1_ASAP7_75t_SL g514 ( .A(n_515), .B(n_524), .Y(n_514) );
AND2x2_ASAP7_75t_L g535 ( .A(n_515), .B(n_536), .Y(n_535) );
AND2x2_ASAP7_75t_L g711 ( .A(n_515), .B(n_634), .Y(n_711) );
AO21x1_ASAP7_75t_SL g515 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_515) );
AO21x2_ASAP7_75t_L g558 ( .A1(n_516), .A2(n_517), .B(n_523), .Y(n_558) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_518), .B(n_522), .Y(n_517) );
OR2x2_ASAP7_75t_L g543 ( .A(n_524), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g554 ( .A(n_524), .B(n_544), .Y(n_554) );
AND2x2_ASAP7_75t_L g600 ( .A(n_524), .B(n_557), .Y(n_600) );
OR2x2_ASAP7_75t_L g621 ( .A(n_524), .B(n_536), .Y(n_621) );
INVx2_ASAP7_75t_SL g627 ( .A(n_524), .Y(n_627) );
AND2x2_ASAP7_75t_L g633 ( .A(n_524), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g643 ( .A(n_524), .B(n_626), .Y(n_643) );
BUFx2_ASAP7_75t_L g665 ( .A(n_524), .Y(n_665) );
OR2x6_ASAP7_75t_L g524 ( .A(n_525), .B(n_532), .Y(n_524) );
INVx2_ASAP7_75t_L g712 ( .A(n_533), .Y(n_712) );
OR2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_543), .Y(n_533) );
OR2x2_ASAP7_75t_L g737 ( .A(n_534), .B(n_581), .Y(n_737) );
INVx2_ASAP7_75t_SL g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_535), .B(n_544), .Y(n_603) );
AND2x2_ASAP7_75t_L g674 ( .A(n_535), .B(n_554), .Y(n_674) );
INVx1_ASAP7_75t_L g556 ( .A(n_536), .Y(n_556) );
HB1xp67_ASAP7_75t_L g565 ( .A(n_536), .Y(n_565) );
INVx1_ASAP7_75t_L g598 ( .A(n_536), .Y(n_598) );
INVx2_ASAP7_75t_L g634 ( .A(n_536), .Y(n_634) );
NOR2xp67_ASAP7_75t_L g564 ( .A(n_544), .B(n_565), .Y(n_564) );
BUFx2_ASAP7_75t_L g624 ( .A(n_544), .Y(n_624) );
INVx2_ASAP7_75t_SL g700 ( .A(n_545), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g601 ( .A1(n_547), .A2(n_602), .B1(n_604), .B2(n_608), .Y(n_601) );
AND2x2_ASAP7_75t_SL g547 ( .A(n_548), .B(n_549), .Y(n_547) );
AND2x2_ASAP7_75t_L g728 ( .A(n_548), .B(n_584), .Y(n_728) );
INVx1_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_550), .B(n_594), .Y(n_673) );
INVx1_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
AND2x2_ASAP7_75t_L g639 ( .A(n_551), .B(n_587), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_552), .B(n_689), .Y(n_688) );
INVx1_ASAP7_75t_L g582 ( .A(n_553), .Y(n_582) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_553), .A2(n_697), .B1(n_701), .B2(n_703), .C(n_705), .Y(n_696) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g566 ( .A(n_554), .B(n_567), .Y(n_566) );
INVxp67_ASAP7_75t_SL g590 ( .A(n_554), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_554), .B(n_597), .Y(n_652) );
INVx1_ASAP7_75t_SL g648 ( .A(n_555), .Y(n_648) );
AOI221xp5_ASAP7_75t_SL g676 ( .A1(n_555), .A2(n_566), .B1(n_677), .B2(n_678), .C(n_681), .Y(n_676) );
AOI322xp5_ASAP7_75t_L g709 ( .A1(n_555), .A2(n_627), .A3(n_654), .B1(n_710), .B2(n_712), .C1(n_713), .C2(n_716), .Y(n_709) );
AND2x2_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
BUFx2_ASAP7_75t_L g576 ( .A(n_556), .Y(n_576) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_557), .Y(n_568) );
INVx2_ASAP7_75t_L g626 ( .A(n_557), .Y(n_626) );
AND2x2_ASAP7_75t_L g667 ( .A(n_557), .B(n_668), .Y(n_667) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OA21x2_ASAP7_75t_SL g559 ( .A1(n_560), .A2(n_566), .B(n_569), .Y(n_559) );
AOI211xp5_ASAP7_75t_L g729 ( .A1(n_560), .A2(n_730), .B(n_731), .C(n_735), .Y(n_729) );
INVx1_ASAP7_75t_SL g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OR2x2_ASAP7_75t_L g618 ( .A(n_562), .B(n_580), .Y(n_618) );
OR2x2_ASAP7_75t_L g702 ( .A(n_562), .B(n_597), .Y(n_702) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g642 ( .A(n_564), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g720 ( .A(n_567), .Y(n_720) );
INVx1_ASAP7_75t_L g567 ( .A(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g606 ( .A(n_568), .Y(n_606) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
OR2x2_ASAP7_75t_L g575 ( .A(n_571), .B(n_576), .Y(n_575) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g610 ( .A(n_573), .B(n_611), .Y(n_610) );
OAI322xp33_ASAP7_75t_L g574 ( .A1(n_575), .A2(n_577), .A3(n_580), .B1(n_582), .B2(n_583), .C1(n_588), .C2(n_590), .Y(n_574) );
INVx1_ASAP7_75t_L g616 ( .A(n_575), .Y(n_616) );
OR2x2_ASAP7_75t_L g588 ( .A(n_577), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_577), .B(n_715), .Y(n_714) );
INVx2_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
AND2x2_ASAP7_75t_L g599 ( .A(n_581), .B(n_600), .Y(n_599) );
OAI32xp33_ASAP7_75t_L g644 ( .A1(n_581), .A2(n_645), .A3(n_648), .B1(n_649), .B2(n_650), .Y(n_644) );
OR2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_585), .Y(n_583) );
INVx2_ASAP7_75t_L g589 ( .A(n_584), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_584), .B(n_647), .Y(n_646) );
NOR2x1_ASAP7_75t_L g686 ( .A(n_584), .B(n_687), .Y(n_686) );
AND2x2_ASAP7_75t_L g710 ( .A(n_584), .B(n_711), .Y(n_710) );
INVx1_ASAP7_75t_L g631 ( .A(n_585), .Y(n_631) );
INVx1_ASAP7_75t_SL g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_589), .B(n_655), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_592), .B(n_612), .Y(n_591) );
OAI21xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_595), .B(n_601), .Y(n_592) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x4_ASAP7_75t_SL g596 ( .A(n_597), .B(n_599), .Y(n_596) );
INVx3_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g661 ( .A(n_600), .B(n_662), .Y(n_661) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g724 ( .A1(n_603), .A2(n_623), .B1(n_725), .B2(n_727), .Y(n_724) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
A2O1A1Ixp33_ASAP7_75t_L g651 ( .A1(n_605), .A2(n_652), .B(n_653), .C(n_656), .Y(n_651) );
OR2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_607), .Y(n_605) );
INVx3_ASAP7_75t_L g733 ( .A(n_607), .Y(n_733) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g614 ( .A(n_611), .Y(n_614) );
AO21x1_ASAP7_75t_L g612 ( .A1(n_613), .A2(n_615), .B(n_619), .Y(n_612) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
INVx2_ASAP7_75t_L g679 ( .A(n_614), .Y(n_679) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g705 ( .A(n_620), .B(n_706), .Y(n_705) );
OR2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_622), .Y(n_620) );
INVx1_ASAP7_75t_L g635 ( .A(n_622), .Y(n_635) );
OR2x2_ASAP7_75t_L g623 ( .A(n_624), .B(n_625), .Y(n_623) );
INVx1_ASAP7_75t_L g692 ( .A(n_625), .Y(n_692) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
NOR3xp33_ASAP7_75t_L g628 ( .A(n_629), .B(n_651), .C(n_663), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_632), .Y(n_630) );
OAI21xp5_ASAP7_75t_SL g693 ( .A1(n_632), .A2(n_694), .B(n_695), .Y(n_693) );
AND2x4_ASAP7_75t_L g632 ( .A(n_633), .B(n_635), .Y(n_632) );
INVx1_ASAP7_75t_L g668 ( .A(n_634), .Y(n_668) );
O2A1O1Ixp5_ASAP7_75t_SL g636 ( .A1(n_637), .A2(n_638), .B(n_640), .C(n_644), .Y(n_636) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx2_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
HB1xp67_ASAP7_75t_L g736 ( .A(n_646), .Y(n_736) );
INVx2_ASAP7_75t_L g721 ( .A(n_649), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g735 ( .A1(n_650), .A2(n_736), .B(n_737), .Y(n_735) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g715 ( .A(n_655), .Y(n_715) );
OAI31xp33_ASAP7_75t_L g656 ( .A1(n_657), .A2(n_659), .A3(n_660), .B(n_661), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g734 ( .A(n_662), .Y(n_734) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_669), .B(n_672), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_665), .B(n_666), .Y(n_664) );
BUFx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g684 ( .A(n_667), .Y(n_684) );
AOI21xp33_ASAP7_75t_SL g731 ( .A1(n_669), .A2(n_732), .B(n_734), .Y(n_731) );
OR2x2_ASAP7_75t_L g669 ( .A(n_670), .B(n_671), .Y(n_669) );
INVx2_ASAP7_75t_L g699 ( .A(n_670), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_670), .B(n_690), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_670), .B(n_707), .Y(n_706) );
INVx2_ASAP7_75t_L g680 ( .A(n_671), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_673), .B(n_674), .Y(n_672) );
NAND5xp2_ASAP7_75t_L g675 ( .A(n_676), .B(n_696), .C(n_709), .D(n_718), .E(n_729), .Y(n_675) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_680), .Y(n_678) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_682), .A2(n_685), .B1(n_688), .B2(n_691), .C(n_693), .Y(n_681) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_684), .Y(n_682) );
INVx1_ASAP7_75t_L g685 ( .A(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_SL g689 ( .A(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
INVxp67_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_722), .B(n_724), .Y(n_718) );
AND2x4_ASAP7_75t_L g719 ( .A(n_720), .B(n_721), .Y(n_719) );
INVx1_ASAP7_75t_SL g722 ( .A(n_723), .Y(n_722) );
INVx1_ASAP7_75t_SL g725 ( .A(n_726), .Y(n_725) );
INVxp67_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
INVx1_ASAP7_75t_L g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx3_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_753), .Y(n_749) );
HB1xp67_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
CKINVDCx5p33_ASAP7_75t_R g751 ( .A(n_752), .Y(n_751) );
A2O1A1Ixp33_ASAP7_75t_L g753 ( .A1(n_754), .A2(n_757), .B(n_760), .C(n_761), .Y(n_753) );
INVxp67_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g762 ( .A(n_763), .Y(n_762) );
NOR2xp33_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .Y(n_764) );
INVx1_ASAP7_75t_SL g766 ( .A(n_767), .Y(n_766) );
endmodule