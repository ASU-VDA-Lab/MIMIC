module real_aes_5995_n_8 (n_4, n_0, n_3, n_5, n_2, n_7, n_6, n_1, n_8);
input n_4;
input n_0;
input n_3;
input n_5;
input n_2;
input n_7;
input n_6;
input n_1;
output n_8;
wire n_17;
wire n_28;
wire n_22;
wire n_13;
wire n_24;
wire n_34;
wire n_12;
wire n_19;
wire n_25;
wire n_32;
wire n_30;
wire n_14;
wire n_11;
wire n_16;
wire n_35;
wire n_15;
wire n_27;
wire n_9;
wire n_23;
wire n_29;
wire n_20;
wire n_18;
wire n_26;
wire n_21;
wire n_31;
wire n_10;
wire n_33;
HB1xp67_ASAP7_75t_L g11 ( .A(n_0), .Y(n_11) );
NOR2xp33_ASAP7_75t_L g20 ( .A(n_0), .B(n_5), .Y(n_20) );
AND2x4_ASAP7_75t_L g14 ( .A(n_1), .B(n_3), .Y(n_14) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_1), .Y(n_22) );
AND2x4_ASAP7_75t_L g34 ( .A(n_1), .B(n_35), .Y(n_34) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_2), .B(n_25), .Y(n_24) );
INVx1_ASAP7_75t_L g35 ( .A(n_3), .Y(n_35) );
BUFx6f_ASAP7_75t_L g28 ( .A(n_4), .Y(n_28) );
AOI21xp5_ASAP7_75t_L g8 ( .A1(n_5), .A2(n_9), .B(n_17), .Y(n_8) );
INVx2_ASAP7_75t_L g16 ( .A(n_6), .Y(n_16) );
AND2x4_ASAP7_75t_L g15 ( .A(n_7), .B(n_16), .Y(n_15) );
INVx1_ASAP7_75t_SL g31 ( .A(n_7), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g9 ( .A(n_10), .B(n_12), .Y(n_9) );
CKINVDCx5p33_ASAP7_75t_R g10 ( .A(n_11), .Y(n_10) );
BUFx2_ASAP7_75t_L g12 ( .A(n_13), .Y(n_12) );
AND2x4_ASAP7_75t_L g13 ( .A(n_14), .B(n_15), .Y(n_13) );
HB1xp67_ASAP7_75t_L g33 ( .A(n_16), .Y(n_33) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_18), .Y(n_17) );
OAI21xp33_ASAP7_75t_L g18 ( .A1(n_19), .A2(n_21), .B(n_23), .Y(n_18) );
HB1xp67_ASAP7_75t_L g19 ( .A(n_20), .Y(n_19) );
AOI211xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_24), .B(n_29), .C(n_34), .Y(n_23) );
INVx1_ASAP7_75t_L g21 ( .A(n_22), .Y(n_21) );
AOI21xp5_ASAP7_75t_L g30 ( .A1(n_22), .A2(n_31), .B(n_32), .Y(n_30) );
INVx2_ASAP7_75t_SL g25 ( .A(n_26), .Y(n_25) );
BUFx2_ASAP7_75t_L g26 ( .A(n_27), .Y(n_26) );
HB1xp67_ASAP7_75t_L g27 ( .A(n_28), .Y(n_27) );
INVxp67_ASAP7_75t_SL g29 ( .A(n_30), .Y(n_29) );
INVx1_ASAP7_75t_L g32 ( .A(n_33), .Y(n_32) );
endmodule