module fake_netlist_6_435_n_1933 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1933);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1933;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1691;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_658;
wire n_616;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1875;
wire n_1865;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_268;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1135;
wire n_1179;
wire n_1169;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1321;
wire n_1241;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1741;
wire n_1325;
wire n_1002;
wire n_1746;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_535;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1890;
wire n_1632;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_151),
.Y(n_185)
);

BUFx4f_ASAP7_75t_SL g186 ( 
.A(n_155),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_78),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_117),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_90),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_115),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_136),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_40),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_135),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_48),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_92),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_1),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_12),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_132),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_55),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_121),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_111),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_112),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_89),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_181),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_104),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_93),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_50),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_69),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_152),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_38),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_40),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_41),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_47),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_87),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_156),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_119),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_154),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_37),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_56),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_74),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_41),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_85),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_39),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_164),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_143),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_38),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_12),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_43),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_9),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_65),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_53),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_52),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_55),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g235 ( 
.A(n_4),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_37),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_32),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_149),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_75),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_113),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_57),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_83),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_120),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_163),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_47),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_67),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_61),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_9),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_165),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_105),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_146),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_126),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_56),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_184),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_179),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_25),
.Y(n_257)
);

INVx1_ASAP7_75t_SL g258 ( 
.A(n_0),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_53),
.Y(n_259)
);

INVx1_ASAP7_75t_SL g260 ( 
.A(n_180),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_158),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_36),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_11),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_18),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_161),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_32),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_110),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_60),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_49),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_23),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_58),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_2),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_86),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_42),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_60),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_20),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_114),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_63),
.Y(n_279)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_98),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_177),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_28),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_21),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_80),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_43),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_175),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_68),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_31),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_19),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_162),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_1),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_107),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_103),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_169),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_17),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_160),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_59),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_128),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_138),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_18),
.Y(n_300)
);

INVx3_ASAP7_75t_L g301 ( 
.A(n_30),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_150),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_54),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_3),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_52),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g306 ( 
.A(n_178),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_33),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_153),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_39),
.Y(n_309)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_174),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_33),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_6),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_157),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_44),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_4),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_145),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_109),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_182),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_72),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_26),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_25),
.Y(n_321)
);

CKINVDCx11_ASAP7_75t_R g322 ( 
.A(n_2),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g323 ( 
.A(n_10),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_168),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_124),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_123),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_102),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_166),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_140),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_13),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_141),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_116),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_159),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_48),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_58),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_91),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_100),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_95),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_65),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_42),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_70),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_101),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_27),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_46),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_8),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_46),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_20),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_15),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_127),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_71),
.Y(n_350)
);

BUFx3_ASAP7_75t_L g351 ( 
.A(n_76),
.Y(n_351)
);

BUFx6f_ASAP7_75t_L g352 ( 
.A(n_97),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_59),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_7),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g355 ( 
.A(n_129),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_106),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_24),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_17),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_67),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_3),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_144),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_57),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_130),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_79),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g365 ( 
.A(n_31),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_24),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_7),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_125),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_301),
.Y(n_369)
);

BUFx2_ASAP7_75t_L g370 ( 
.A(n_227),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_322),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_301),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_301),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_301),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_187),
.Y(n_375)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_196),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_231),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_231),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_351),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_208),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_282),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_188),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_189),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_282),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_196),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_214),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_249),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_323),
.B(n_0),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_190),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_193),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_195),
.Y(n_391)
);

INVxp67_ASAP7_75t_SL g392 ( 
.A(n_351),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_198),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_269),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_200),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_210),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_351),
.Y(n_397)
);

INVxp67_ASAP7_75t_L g398 ( 
.A(n_210),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_220),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_202),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_220),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g402 ( 
.A(n_281),
.Y(n_402)
);

OR2x2_ASAP7_75t_L g403 ( 
.A(n_222),
.B(n_5),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_287),
.Y(n_404)
);

INVxp67_ASAP7_75t_SL g405 ( 
.A(n_215),
.Y(n_405)
);

INVxp67_ASAP7_75t_L g406 ( 
.A(n_222),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_298),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_203),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_280),
.B(n_5),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_230),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g411 ( 
.A(n_326),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_280),
.B(n_6),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_185),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_230),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_349),
.Y(n_416)
);

INVxp67_ASAP7_75t_L g417 ( 
.A(n_237),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_364),
.B(n_8),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_237),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_264),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_191),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_227),
.Y(n_422)
);

HB1xp67_ASAP7_75t_L g423 ( 
.A(n_269),
.Y(n_423)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_318),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_205),
.Y(n_425)
);

CKINVDCx14_ASAP7_75t_R g426 ( 
.A(n_241),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_264),
.Y(n_427)
);

CKINVDCx20_ASAP7_75t_R g428 ( 
.A(n_318),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_206),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_270),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_216),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_270),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_186),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_194),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_291),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_291),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_295),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_295),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_221),
.Y(n_439)
);

INVxp33_ASAP7_75t_SL g440 ( 
.A(n_197),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_223),
.Y(n_441)
);

BUFx10_ASAP7_75t_L g442 ( 
.A(n_364),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_225),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_297),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_226),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_238),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_239),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_297),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_R g449 ( 
.A(n_242),
.B(n_176),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g450 ( 
.A(n_241),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_315),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_243),
.Y(n_452)
);

INVxp33_ASAP7_75t_L g453 ( 
.A(n_315),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_321),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_321),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_335),
.Y(n_456)
);

NOR2xp33_ASAP7_75t_L g457 ( 
.A(n_191),
.B(n_10),
.Y(n_457)
);

CKINVDCx5p33_ASAP7_75t_R g458 ( 
.A(n_244),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_335),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_252),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_413),
.Y(n_461)
);

BUFx2_ASAP7_75t_L g462 ( 
.A(n_424),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_413),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

INVx3_ASAP7_75t_L g465 ( 
.A(n_421),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_369),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_369),
.Y(n_467)
);

BUFx2_ASAP7_75t_L g468 ( 
.A(n_428),
.Y(n_468)
);

OA21x2_ASAP7_75t_L g469 ( 
.A1(n_372),
.A2(n_348),
.B(n_340),
.Y(n_469)
);

BUFx6f_ASAP7_75t_L g470 ( 
.A(n_421),
.Y(n_470)
);

HB1xp67_ASAP7_75t_L g471 ( 
.A(n_394),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_372),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_385),
.Y(n_473)
);

BUFx12f_ASAP7_75t_L g474 ( 
.A(n_371),
.Y(n_474)
);

AND2x2_ASAP7_75t_SL g475 ( 
.A(n_409),
.B(n_185),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_385),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_379),
.B(n_253),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_396),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_373),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_379),
.B(n_368),
.Y(n_480)
);

BUFx8_ASAP7_75t_L g481 ( 
.A(n_370),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_373),
.Y(n_482)
);

INVxp67_ASAP7_75t_L g483 ( 
.A(n_423),
.Y(n_483)
);

BUFx6f_ASAP7_75t_L g484 ( 
.A(n_374),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_374),
.Y(n_485)
);

AND2x4_ASAP7_75t_L g486 ( 
.A(n_379),
.B(n_251),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_377),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_377),
.Y(n_488)
);

BUFx6f_ASAP7_75t_L g489 ( 
.A(n_378),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_381),
.Y(n_491)
);

BUFx6f_ASAP7_75t_L g492 ( 
.A(n_381),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_384),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_384),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_392),
.B(n_255),
.Y(n_495)
);

HB1xp67_ASAP7_75t_L g496 ( 
.A(n_370),
.Y(n_496)
);

AND2x2_ASAP7_75t_L g497 ( 
.A(n_397),
.B(n_422),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_396),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_SL g499 ( 
.A1(n_450),
.A2(n_272),
.B1(n_365),
.B2(n_212),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_399),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_399),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_412),
.B(n_261),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g503 ( 
.A(n_418),
.B(n_265),
.Y(n_503)
);

AND2x2_ASAP7_75t_L g504 ( 
.A(n_401),
.B(n_201),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_401),
.B(n_201),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_410),
.Y(n_506)
);

BUFx6f_ASAP7_75t_L g507 ( 
.A(n_410),
.Y(n_507)
);

HB1xp67_ASAP7_75t_L g508 ( 
.A(n_434),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_415),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_415),
.Y(n_510)
);

NOR2xp33_ASAP7_75t_SL g511 ( 
.A(n_450),
.B(n_241),
.Y(n_511)
);

AND2x4_ASAP7_75t_L g512 ( 
.A(n_419),
.B(n_251),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_419),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_420),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_420),
.Y(n_515)
);

INVxp67_ASAP7_75t_L g516 ( 
.A(n_405),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g517 ( 
.A(n_457),
.B(n_278),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_430),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_430),
.Y(n_519)
);

INVx2_ASAP7_75t_L g520 ( 
.A(n_435),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_435),
.B(n_436),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_436),
.B(n_284),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_437),
.Y(n_523)
);

BUFx6f_ASAP7_75t_L g524 ( 
.A(n_437),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_438),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_438),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_444),
.B(n_290),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_444),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_448),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_448),
.Y(n_530)
);

HB1xp67_ASAP7_75t_L g531 ( 
.A(n_388),
.Y(n_531)
);

AND2x4_ASAP7_75t_L g532 ( 
.A(n_454),
.B(n_267),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_454),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_426),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_455),
.Y(n_535)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_455),
.B(n_292),
.Y(n_536)
);

INVx2_ASAP7_75t_L g537 ( 
.A(n_456),
.Y(n_537)
);

AND2x6_ASAP7_75t_L g538 ( 
.A(n_456),
.B(n_185),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_459),
.B(n_204),
.Y(n_539)
);

NAND2xp33_ASAP7_75t_L g540 ( 
.A(n_517),
.B(n_531),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_463),
.Y(n_541)
);

BUFx10_ASAP7_75t_L g542 ( 
.A(n_475),
.Y(n_542)
);

NOR2xp33_ASAP7_75t_SL g543 ( 
.A(n_511),
.B(n_433),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_486),
.Y(n_544)
);

INVx2_ASAP7_75t_L g545 ( 
.A(n_463),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_516),
.B(n_440),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_SL g547 ( 
.A(n_511),
.B(n_445),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_497),
.B(n_459),
.Y(n_548)
);

AND2x4_ASAP7_75t_L g549 ( 
.A(n_504),
.B(n_204),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_463),
.Y(n_550)
);

AOI22xp5_ASAP7_75t_L g551 ( 
.A1(n_531),
.A2(n_447),
.B1(n_382),
.B2(n_383),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_475),
.A2(n_403),
.B1(n_340),
.B2(n_367),
.Y(n_552)
);

INVx3_ASAP7_75t_L g553 ( 
.A(n_484),
.Y(n_553)
);

BUFx10_ASAP7_75t_L g554 ( 
.A(n_475),
.Y(n_554)
);

INVx3_ASAP7_75t_L g555 ( 
.A(n_484),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_463),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_461),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_534),
.B(n_375),
.Y(n_558)
);

BUFx6f_ASAP7_75t_SL g559 ( 
.A(n_475),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

INVx1_ASAP7_75t_SL g561 ( 
.A(n_462),
.Y(n_561)
);

BUFx6f_ASAP7_75t_L g562 ( 
.A(n_507),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_496),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_461),
.Y(n_564)
);

AOI22xp33_ASAP7_75t_L g565 ( 
.A1(n_517),
.A2(n_403),
.B1(n_348),
.B2(n_367),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_496),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_484),
.Y(n_567)
);

NAND3xp33_ASAP7_75t_SL g568 ( 
.A(n_502),
.B(n_229),
.C(n_192),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_461),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_497),
.A2(n_267),
.B1(n_361),
.B2(n_453),
.Y(n_570)
);

NOR2x1p5_ASAP7_75t_L g571 ( 
.A(n_474),
.B(n_199),
.Y(n_571)
);

INVx3_ASAP7_75t_L g572 ( 
.A(n_484),
.Y(n_572)
);

INVx2_ASAP7_75t_SL g573 ( 
.A(n_497),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_486),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_486),
.Y(n_575)
);

INVx4_ASAP7_75t_L g576 ( 
.A(n_470),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_464),
.Y(n_577)
);

BUFx2_ASAP7_75t_L g578 ( 
.A(n_481),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_464),
.Y(n_579)
);

AND2x6_ASAP7_75t_L g580 ( 
.A(n_486),
.B(n_185),
.Y(n_580)
);

NOR2x1p5_ASAP7_75t_L g581 ( 
.A(n_474),
.B(n_207),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_464),
.Y(n_582)
);

AOI22xp5_ASAP7_75t_L g583 ( 
.A1(n_516),
.A2(n_460),
.B1(n_458),
.B2(n_452),
.Y(n_583)
);

OAI22xp33_ASAP7_75t_L g584 ( 
.A1(n_502),
.A2(n_258),
.B1(n_303),
.B2(n_362),
.Y(n_584)
);

INVx3_ASAP7_75t_L g585 ( 
.A(n_484),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_495),
.B(n_389),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_464),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_464),
.Y(n_589)
);

INVx2_ASAP7_75t_SL g590 ( 
.A(n_508),
.Y(n_590)
);

INVx3_ASAP7_75t_L g591 ( 
.A(n_484),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_469),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_495),
.B(n_390),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_L g594 ( 
.A(n_477),
.B(n_391),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_469),
.Y(n_595)
);

INVx4_ASAP7_75t_L g596 ( 
.A(n_470),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_462),
.Y(n_597)
);

BUFx10_ASAP7_75t_L g598 ( 
.A(n_508),
.Y(n_598)
);

AOI22xp33_ASAP7_75t_L g599 ( 
.A1(n_503),
.A2(n_361),
.B1(n_209),
.B2(n_217),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_477),
.B(n_393),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_SL g601 ( 
.A(n_534),
.B(n_395),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_484),
.Y(n_602)
);

OR2x6_ASAP7_75t_L g603 ( 
.A(n_474),
.B(n_209),
.Y(n_603)
);

BUFx3_ASAP7_75t_L g604 ( 
.A(n_469),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_480),
.B(n_400),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_466),
.Y(n_606)
);

HAxp5_ASAP7_75t_SL g607 ( 
.A(n_499),
.B(n_217),
.CON(n_607),
.SN(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_480),
.B(n_408),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_469),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_466),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_466),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_503),
.B(n_425),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_469),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_466),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_469),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_472),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_472),
.Y(n_617)
);

AND3x2_ASAP7_75t_L g618 ( 
.A(n_534),
.B(n_235),
.C(n_218),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_498),
.Y(n_619)
);

NOR2xp33_ASAP7_75t_L g620 ( 
.A(n_522),
.B(n_429),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_498),
.Y(n_621)
);

OAI22xp5_ASAP7_75t_L g622 ( 
.A1(n_483),
.A2(n_431),
.B1(n_446),
.B2(n_443),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_472),
.Y(n_623)
);

BUFx3_ASAP7_75t_L g624 ( 
.A(n_467),
.Y(n_624)
);

AND2x2_ASAP7_75t_L g625 ( 
.A(n_504),
.B(n_442),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_512),
.A2(n_328),
.B1(n_218),
.B2(n_240),
.Y(n_626)
);

INVx2_ASAP7_75t_L g627 ( 
.A(n_472),
.Y(n_627)
);

AND2x2_ASAP7_75t_L g628 ( 
.A(n_504),
.B(n_442),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_SL g629 ( 
.A(n_481),
.B(n_439),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_481),
.B(n_441),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_485),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_522),
.B(n_442),
.Y(n_632)
);

BUFx10_ASAP7_75t_L g633 ( 
.A(n_471),
.Y(n_633)
);

INVx1_ASAP7_75t_SL g634 ( 
.A(n_462),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_485),
.Y(n_635)
);

AOI22xp5_ASAP7_75t_L g636 ( 
.A1(n_483),
.A2(n_266),
.B1(n_320),
.B2(n_236),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_481),
.B(n_442),
.Y(n_637)
);

AND2x6_ASAP7_75t_L g638 ( 
.A(n_505),
.B(n_185),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_498),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_485),
.Y(n_640)
);

INVx4_ASAP7_75t_L g641 ( 
.A(n_470),
.Y(n_641)
);

AND2x2_ASAP7_75t_L g642 ( 
.A(n_505),
.B(n_376),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_481),
.B(n_449),
.Y(n_643)
);

INVx1_ASAP7_75t_SL g644 ( 
.A(n_468),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_SL g645 ( 
.A(n_481),
.B(n_250),
.Y(n_645)
);

AND2x6_ASAP7_75t_L g646 ( 
.A(n_505),
.B(n_185),
.Y(n_646)
);

AND2x4_ASAP7_75t_L g647 ( 
.A(n_539),
.B(n_240),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_L g648 ( 
.A(n_527),
.B(n_260),
.Y(n_648)
);

BUFx10_ASAP7_75t_L g649 ( 
.A(n_471),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_527),
.B(n_306),
.Y(n_650)
);

AND2x2_ASAP7_75t_L g651 ( 
.A(n_539),
.B(n_500),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_500),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_536),
.B(n_355),
.Y(n_653)
);

INVx4_ASAP7_75t_L g654 ( 
.A(n_470),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_485),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_L g656 ( 
.A(n_536),
.B(n_380),
.Y(n_656)
);

INVx3_ASAP7_75t_L g657 ( 
.A(n_484),
.Y(n_657)
);

INVx1_ASAP7_75t_SL g658 ( 
.A(n_468),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_500),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_530),
.B(n_386),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_512),
.B(n_250),
.Y(n_661)
);

AND2x2_ASAP7_75t_L g662 ( 
.A(n_539),
.B(n_398),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_482),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_482),
.Y(n_664)
);

NOR2xp33_ASAP7_75t_L g665 ( 
.A(n_530),
.B(n_387),
.Y(n_665)
);

AND2x4_ASAP7_75t_L g666 ( 
.A(n_512),
.B(n_256),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_482),
.Y(n_667)
);

BUFx3_ASAP7_75t_L g668 ( 
.A(n_467),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_530),
.B(n_402),
.Y(n_669)
);

INVx3_ASAP7_75t_L g670 ( 
.A(n_470),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_482),
.B(n_293),
.Y(n_671)
);

BUFx10_ASAP7_75t_L g672 ( 
.A(n_512),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_482),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_474),
.Y(n_674)
);

BUFx3_ASAP7_75t_L g675 ( 
.A(n_467),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_507),
.Y(n_676)
);

NOR2xp33_ASAP7_75t_L g677 ( 
.A(n_530),
.B(n_404),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_507),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_514),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_514),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_468),
.Y(n_681)
);

AND2x4_ASAP7_75t_SL g682 ( 
.A(n_512),
.B(n_250),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_514),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_515),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_507),
.Y(n_685)
);

INVx3_ASAP7_75t_L g686 ( 
.A(n_470),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_515),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_507),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_507),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_507),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_521),
.B(n_406),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_507),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_563),
.B(n_499),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_541),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_620),
.B(n_530),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_573),
.B(n_211),
.Y(n_696)
);

INVx2_ASAP7_75t_L g697 ( 
.A(n_541),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_544),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_560),
.Y(n_699)
);

HB1xp67_ASAP7_75t_L g700 ( 
.A(n_563),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_573),
.B(n_509),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_566),
.B(n_417),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_560),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_612),
.B(n_509),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_574),
.Y(n_705)
);

AND2x4_ASAP7_75t_L g706 ( 
.A(n_651),
.B(n_473),
.Y(n_706)
);

INVxp67_ASAP7_75t_L g707 ( 
.A(n_546),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_574),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_651),
.B(n_473),
.Y(n_709)
);

INVx2_ASAP7_75t_L g710 ( 
.A(n_604),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_625),
.B(n_509),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_SL g712 ( 
.A(n_542),
.B(n_310),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_625),
.B(n_509),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_628),
.B(n_509),
.Y(n_714)
);

BUFx8_ASAP7_75t_L g715 ( 
.A(n_590),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_575),
.Y(n_716)
);

NOR2xp33_ASAP7_75t_L g717 ( 
.A(n_648),
.B(n_213),
.Y(n_717)
);

AO22x2_ASAP7_75t_L g718 ( 
.A1(n_607),
.A2(n_350),
.B1(n_313),
.B2(n_316),
.Y(n_718)
);

AND2x2_ASAP7_75t_L g719 ( 
.A(n_628),
.B(n_407),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_604),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_542),
.B(n_310),
.Y(n_721)
);

NOR2xp33_ASAP7_75t_L g722 ( 
.A(n_650),
.B(n_653),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_542),
.B(n_310),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_L g724 ( 
.A(n_586),
.B(n_509),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_587),
.Y(n_725)
);

INVx8_ASAP7_75t_L g726 ( 
.A(n_603),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_593),
.B(n_509),
.Y(n_727)
);

AND2x2_ASAP7_75t_L g728 ( 
.A(n_590),
.B(n_566),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_594),
.B(n_509),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_587),
.Y(n_730)
);

NAND2x1p5_ASAP7_75t_L g731 ( 
.A(n_604),
.B(n_256),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_542),
.B(n_554),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_600),
.B(n_524),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_605),
.B(n_524),
.Y(n_734)
);

OR2x2_ASAP7_75t_L g735 ( 
.A(n_691),
.B(n_427),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_541),
.Y(n_736)
);

AOI22xp33_ASAP7_75t_L g737 ( 
.A1(n_552),
.A2(n_512),
.B1(n_532),
.B2(n_479),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_624),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_608),
.B(n_524),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_554),
.B(n_310),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_624),
.Y(n_741)
);

AND2x2_ASAP7_75t_L g742 ( 
.A(n_642),
.B(n_411),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_615),
.A2(n_532),
.B1(n_479),
.B2(n_299),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_668),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_559),
.A2(n_416),
.B1(n_414),
.B2(n_329),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_545),
.Y(n_746)
);

NAND2xp5_ASAP7_75t_L g747 ( 
.A(n_668),
.B(n_675),
.Y(n_747)
);

AOI221xp5_ASAP7_75t_L g748 ( 
.A1(n_584),
.A2(n_432),
.B1(n_451),
.B2(n_343),
.C(n_358),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_668),
.B(n_524),
.Y(n_749)
);

OR2x2_ASAP7_75t_SL g750 ( 
.A(n_568),
.B(n_273),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_675),
.Y(n_751)
);

INVx2_ASAP7_75t_SL g752 ( 
.A(n_633),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_675),
.B(n_524),
.Y(n_753)
);

BUFx6f_ASAP7_75t_L g754 ( 
.A(n_615),
.Y(n_754)
);

NOR2xp33_ASAP7_75t_SL g755 ( 
.A(n_547),
.B(n_250),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_619),
.Y(n_756)
);

AND2x4_ASAP7_75t_L g757 ( 
.A(n_549),
.B(n_476),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_548),
.B(n_524),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_540),
.B(n_219),
.Y(n_759)
);

NAND2xp5_ASAP7_75t_L g760 ( 
.A(n_548),
.B(n_524),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_691),
.B(n_224),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_636),
.A2(n_314),
.B1(n_312),
.B2(n_311),
.Y(n_762)
);

NOR2xp33_ASAP7_75t_R g763 ( 
.A(n_674),
.B(n_296),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_545),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_554),
.B(n_615),
.Y(n_765)
);

NAND2xp33_ASAP7_75t_L g766 ( 
.A(n_632),
.B(n_302),
.Y(n_766)
);

NOR2x1p5_ASAP7_75t_SL g767 ( 
.A(n_592),
.B(n_479),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_619),
.B(n_524),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_633),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_642),
.B(n_521),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_559),
.A2(n_656),
.B1(n_665),
.B2(n_660),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_622),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_621),
.B(n_532),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_621),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_671),
.A2(n_465),
.B(n_470),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_583),
.B(n_228),
.Y(n_776)
);

NOR2xp33_ASAP7_75t_SL g777 ( 
.A(n_578),
.B(n_241),
.Y(n_777)
);

BUFx12f_ASAP7_75t_SL g778 ( 
.A(n_603),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_554),
.B(n_310),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_592),
.A2(n_465),
.B(n_470),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_639),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_639),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_652),
.B(n_532),
.Y(n_783)
);

OR2x2_ASAP7_75t_SL g784 ( 
.A(n_607),
.B(n_273),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_652),
.B(n_532),
.Y(n_785)
);

INVx1_ASAP7_75t_SL g786 ( 
.A(n_561),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_672),
.B(n_595),
.Y(n_787)
);

OAI22xp5_ASAP7_75t_L g788 ( 
.A1(n_559),
.A2(n_286),
.B1(n_328),
.B2(n_327),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_659),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_669),
.B(n_232),
.Y(n_790)
);

NAND3xp33_ASAP7_75t_L g791 ( 
.A(n_565),
.B(n_234),
.C(n_233),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_659),
.B(n_679),
.Y(n_792)
);

NAND3xp33_ASAP7_75t_L g793 ( 
.A(n_570),
.B(n_246),
.C(n_245),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_SL g794 ( 
.A(n_672),
.B(n_310),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_679),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_680),
.B(n_532),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_680),
.B(n_510),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_683),
.Y(n_798)
);

AOI22xp5_ASAP7_75t_L g799 ( 
.A1(n_559),
.A2(n_341),
.B1(n_338),
.B2(n_337),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_SL g800 ( 
.A(n_672),
.B(n_352),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_684),
.B(n_510),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_684),
.B(n_687),
.Y(n_802)
);

AOI22xp5_ASAP7_75t_L g803 ( 
.A1(n_677),
.A2(n_317),
.B1(n_319),
.B2(n_324),
.Y(n_803)
);

BUFx3_ASAP7_75t_L g804 ( 
.A(n_666),
.Y(n_804)
);

NOR2xp33_ASAP7_75t_L g805 ( 
.A(n_551),
.B(n_247),
.Y(n_805)
);

OR2x2_ASAP7_75t_L g806 ( 
.A(n_597),
.B(n_634),
.Y(n_806)
);

XOR2xp5_ASAP7_75t_L g807 ( 
.A(n_636),
.B(n_325),
.Y(n_807)
);

INVx2_ASAP7_75t_SL g808 ( 
.A(n_633),
.Y(n_808)
);

OR2x2_ASAP7_75t_L g809 ( 
.A(n_644),
.B(n_476),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_687),
.B(n_510),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_663),
.Y(n_811)
);

AOI22xp33_ASAP7_75t_L g812 ( 
.A1(n_595),
.A2(n_286),
.B1(n_294),
.B2(n_363),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_SL g813 ( 
.A(n_672),
.B(n_352),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_662),
.B(n_248),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_609),
.B(n_613),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_663),
.Y(n_816)
);

INVx2_ASAP7_75t_L g817 ( 
.A(n_609),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_613),
.B(n_352),
.Y(n_818)
);

A2O1A1Ixp33_ASAP7_75t_L g819 ( 
.A1(n_662),
.A2(n_515),
.B(n_518),
.C(n_535),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_558),
.B(n_254),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_SL g821 ( 
.A(n_549),
.B(n_647),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_549),
.B(n_510),
.Y(n_822)
);

INVx2_ASAP7_75t_SL g823 ( 
.A(n_633),
.Y(n_823)
);

AND2x2_ASAP7_75t_L g824 ( 
.A(n_598),
.B(n_478),
.Y(n_824)
);

BUFx3_ASAP7_75t_L g825 ( 
.A(n_666),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_SL g826 ( 
.A(n_578),
.B(n_331),
.Y(n_826)
);

AOI22xp5_ASAP7_75t_L g827 ( 
.A1(n_549),
.A2(n_336),
.B1(n_333),
.B2(n_294),
.Y(n_827)
);

INVxp67_ASAP7_75t_L g828 ( 
.A(n_543),
.Y(n_828)
);

AOI21xp5_ASAP7_75t_L g829 ( 
.A1(n_647),
.A2(n_465),
.B(n_537),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_647),
.B(n_513),
.Y(n_830)
);

NOR2xp33_ASAP7_75t_L g831 ( 
.A(n_601),
.B(n_257),
.Y(n_831)
);

O2A1O1Ixp33_ASAP7_75t_L g832 ( 
.A1(n_661),
.A2(n_478),
.B(n_501),
.C(n_506),
.Y(n_832)
);

INVx2_ASAP7_75t_L g833 ( 
.A(n_545),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_550),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_663),
.Y(n_835)
);

INVx2_ASAP7_75t_L g836 ( 
.A(n_550),
.Y(n_836)
);

NAND3xp33_ASAP7_75t_L g837 ( 
.A(n_599),
.B(n_276),
.C(n_288),
.Y(n_837)
);

O2A1O1Ixp33_ASAP7_75t_L g838 ( 
.A1(n_647),
.A2(n_501),
.B(n_506),
.C(n_519),
.Y(n_838)
);

INVx2_ASAP7_75t_L g839 ( 
.A(n_550),
.Y(n_839)
);

AOI22xp5_ASAP7_75t_L g840 ( 
.A1(n_645),
.A2(n_299),
.B1(n_363),
.B2(n_350),
.Y(n_840)
);

NOR2xp33_ASAP7_75t_L g841 ( 
.A(n_682),
.B(n_259),
.Y(n_841)
);

INVx1_ASAP7_75t_L g842 ( 
.A(n_664),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_682),
.B(n_513),
.Y(n_843)
);

NAND3xp33_ASAP7_75t_L g844 ( 
.A(n_626),
.B(n_271),
.C(n_274),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_556),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_664),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_664),
.Y(n_847)
);

O2A1O1Ixp5_ASAP7_75t_L g848 ( 
.A1(n_666),
.A2(n_308),
.B(n_329),
.C(n_356),
.Y(n_848)
);

OAI22xp5_ASAP7_75t_L g849 ( 
.A1(n_682),
.A2(n_308),
.B1(n_332),
.B2(n_327),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_666),
.B(n_513),
.Y(n_850)
);

NAND2xp5_ASAP7_75t_L g851 ( 
.A(n_667),
.B(n_513),
.Y(n_851)
);

NAND2xp5_ASAP7_75t_L g852 ( 
.A(n_667),
.B(n_520),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_667),
.B(n_520),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_673),
.Y(n_854)
);

AND2x4_ASAP7_75t_L g855 ( 
.A(n_603),
.B(n_519),
.Y(n_855)
);

NAND2xp33_ASAP7_75t_L g856 ( 
.A(n_638),
.B(n_352),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_673),
.B(n_352),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_673),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_557),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_629),
.B(n_262),
.Y(n_860)
);

HB1xp67_ASAP7_75t_L g861 ( 
.A(n_700),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_722),
.B(n_770),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_722),
.B(n_717),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_717),
.B(n_630),
.Y(n_864)
);

AO21x1_ASAP7_75t_L g865 ( 
.A1(n_712),
.A2(n_637),
.B(n_643),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_771),
.A2(n_603),
.B1(n_646),
.B2(n_638),
.Y(n_866)
);

AO21x1_ASAP7_75t_L g867 ( 
.A1(n_712),
.A2(n_316),
.B(n_313),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_711),
.A2(n_678),
.B(n_676),
.Y(n_868)
);

OAI21xp33_ASAP7_75t_L g869 ( 
.A1(n_761),
.A2(n_814),
.B(n_805),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_728),
.B(n_598),
.Y(n_870)
);

O2A1O1Ixp33_ASAP7_75t_L g871 ( 
.A1(n_819),
.A2(n_332),
.B(n_356),
.C(n_569),
.Y(n_871)
);

AOI21xp5_ASAP7_75t_L g872 ( 
.A1(n_713),
.A2(n_678),
.B(n_676),
.Y(n_872)
);

CKINVDCx5p33_ASAP7_75t_R g873 ( 
.A(n_763),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_781),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_754),
.B(n_638),
.Y(n_875)
);

AOI21xp5_ASAP7_75t_L g876 ( 
.A1(n_714),
.A2(n_678),
.B(n_676),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_781),
.Y(n_877)
);

OAI22xp5_ASAP7_75t_L g878 ( 
.A1(n_743),
.A2(n_603),
.B1(n_681),
.B2(n_658),
.Y(n_878)
);

INVx11_ASAP7_75t_L g879 ( 
.A(n_715),
.Y(n_879)
);

NOR3xp33_ASAP7_75t_L g880 ( 
.A(n_805),
.B(n_525),
.C(n_523),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_821),
.A2(n_765),
.B(n_760),
.Y(n_881)
);

OAI21x1_ASAP7_75t_L g882 ( 
.A1(n_780),
.A2(n_686),
.B(n_670),
.Y(n_882)
);

OAI21xp5_ASAP7_75t_L g883 ( 
.A1(n_818),
.A2(n_688),
.B(n_685),
.Y(n_883)
);

OAI21x1_ASAP7_75t_L g884 ( 
.A1(n_749),
.A2(n_686),
.B(n_670),
.Y(n_884)
);

AND2x4_ASAP7_75t_L g885 ( 
.A(n_706),
.B(n_709),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_707),
.B(n_553),
.Y(n_886)
);

OAI21xp5_ASAP7_75t_L g887 ( 
.A1(n_818),
.A2(n_688),
.B(n_685),
.Y(n_887)
);

OAI21xp5_ASAP7_75t_L g888 ( 
.A1(n_721),
.A2(n_740),
.B(n_723),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_821),
.A2(n_688),
.B(n_685),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_843),
.A2(n_596),
.B(n_576),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_700),
.B(n_598),
.Y(n_891)
);

O2A1O1Ixp33_ASAP7_75t_L g892 ( 
.A1(n_819),
.A2(n_557),
.B(n_564),
.C(n_569),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_790),
.B(n_553),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_790),
.B(n_553),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_706),
.B(n_553),
.Y(n_895)
);

AOI22xp33_ASAP7_75t_L g896 ( 
.A1(n_757),
.A2(n_646),
.B1(n_638),
.B2(n_580),
.Y(n_896)
);

AND2x4_ASAP7_75t_L g897 ( 
.A(n_709),
.B(n_571),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_782),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_695),
.B(n_757),
.Y(n_899)
);

INVx1_ASAP7_75t_SL g900 ( 
.A(n_786),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_806),
.B(n_598),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_828),
.B(n_649),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_696),
.B(n_555),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_696),
.B(n_555),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_754),
.B(n_649),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_L g906 ( 
.A(n_735),
.B(n_649),
.Y(n_906)
);

NAND2x1p5_ASAP7_75t_L g907 ( 
.A(n_754),
.B(n_555),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_743),
.B(n_555),
.Y(n_908)
);

OAI22xp5_ASAP7_75t_L g909 ( 
.A1(n_812),
.A2(n_690),
.B1(n_689),
.B2(n_692),
.Y(n_909)
);

AOI21xp5_ASAP7_75t_L g910 ( 
.A1(n_765),
.A2(n_690),
.B(n_689),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_710),
.B(n_567),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_758),
.A2(n_690),
.B(n_689),
.Y(n_912)
);

AOI21xp5_ASAP7_75t_L g913 ( 
.A1(n_729),
.A2(n_692),
.B(n_596),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_733),
.A2(n_692),
.B(n_596),
.Y(n_914)
);

AOI21xp5_ASAP7_75t_L g915 ( 
.A1(n_734),
.A2(n_596),
.B(n_576),
.Y(n_915)
);

INVx2_ASAP7_75t_SL g916 ( 
.A(n_809),
.Y(n_916)
);

HB1xp67_ASAP7_75t_L g917 ( 
.A(n_742),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_754),
.B(n_649),
.Y(n_918)
);

INVx5_ASAP7_75t_L g919 ( 
.A(n_815),
.Y(n_919)
);

OAI21xp5_ASAP7_75t_L g920 ( 
.A1(n_721),
.A2(n_610),
.B(n_606),
.Y(n_920)
);

O2A1O1Ixp33_ASAP7_75t_L g921 ( 
.A1(n_788),
.A2(n_564),
.B(n_569),
.C(n_557),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_804),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_710),
.B(n_567),
.Y(n_923)
);

HB1xp67_ASAP7_75t_L g924 ( 
.A(n_824),
.Y(n_924)
);

AND2x4_ASAP7_75t_L g925 ( 
.A(n_804),
.B(n_571),
.Y(n_925)
);

AOI21x1_ASAP7_75t_L g926 ( 
.A1(n_794),
.A2(n_610),
.B(n_606),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_698),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_825),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_699),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_739),
.A2(n_641),
.B(n_576),
.Y(n_930)
);

NOR2xp33_ASAP7_75t_L g931 ( 
.A(n_776),
.B(n_618),
.Y(n_931)
);

NOR2x1_ASAP7_75t_R g932 ( 
.A(n_772),
.B(n_752),
.Y(n_932)
);

O2A1O1Ixp33_ASAP7_75t_L g933 ( 
.A1(n_723),
.A2(n_564),
.B(n_525),
.C(n_523),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_720),
.B(n_567),
.Y(n_934)
);

NOR2xp33_ASAP7_75t_L g935 ( 
.A(n_776),
.B(n_263),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_720),
.B(n_812),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_755),
.B(n_562),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_740),
.A2(n_528),
.B(n_518),
.C(n_535),
.Y(n_938)
);

INVxp67_ASAP7_75t_L g939 ( 
.A(n_702),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_704),
.A2(n_641),
.B(n_576),
.Y(n_940)
);

AOI21xp33_ASAP7_75t_L g941 ( 
.A1(n_759),
.A2(n_275),
.B(n_268),
.Y(n_941)
);

BUFx6f_ASAP7_75t_L g942 ( 
.A(n_825),
.Y(n_942)
);

AOI21xp5_ASAP7_75t_L g943 ( 
.A1(n_724),
.A2(n_641),
.B(n_654),
.Y(n_943)
);

NAND2x1p5_ASAP7_75t_L g944 ( 
.A(n_732),
.B(n_567),
.Y(n_944)
);

AND2x2_ASAP7_75t_L g945 ( 
.A(n_761),
.B(n_581),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_703),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_817),
.B(n_572),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_855),
.B(n_562),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_817),
.B(n_572),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_756),
.B(n_572),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_855),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_774),
.B(n_789),
.Y(n_952)
);

OAI21xp5_ASAP7_75t_L g953 ( 
.A1(n_779),
.A2(n_627),
.B(n_606),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_727),
.A2(n_641),
.B(n_654),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_822),
.A2(n_654),
.B(n_562),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_830),
.A2(n_654),
.B(n_562),
.Y(n_956)
);

INVx2_ASAP7_75t_L g957 ( 
.A(n_705),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_747),
.A2(n_562),
.B(n_686),
.Y(n_958)
);

AOI21xp5_ASAP7_75t_L g959 ( 
.A1(n_701),
.A2(n_562),
.B(n_686),
.Y(n_959)
);

OR2x6_ASAP7_75t_L g960 ( 
.A(n_726),
.B(n_581),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_719),
.B(n_528),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_795),
.B(n_572),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_798),
.B(n_585),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_850),
.A2(n_670),
.B(n_657),
.Y(n_964)
);

AOI21x1_ASAP7_75t_L g965 ( 
.A1(n_794),
.A2(n_813),
.B(n_800),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_787),
.A2(n_670),
.B(n_657),
.Y(n_966)
);

AND2x2_ASAP7_75t_L g967 ( 
.A(n_814),
.B(n_518),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_693),
.B(n_820),
.Y(n_968)
);

AOI21xp5_ASAP7_75t_L g969 ( 
.A1(n_787),
.A2(n_657),
.B(n_585),
.Y(n_969)
);

O2A1O1Ixp33_ASAP7_75t_L g970 ( 
.A1(n_779),
.A2(n_535),
.B(n_655),
.C(n_611),
.Y(n_970)
);

A2O1A1Ixp33_ASAP7_75t_L g971 ( 
.A1(n_759),
.A2(n_657),
.B(n_591),
.C(n_602),
.Y(n_971)
);

NAND2x1p5_ASAP7_75t_L g972 ( 
.A(n_732),
.B(n_585),
.Y(n_972)
);

AOI21xp5_ASAP7_75t_L g973 ( 
.A1(n_773),
.A2(n_655),
.B(n_610),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_860),
.B(n_841),
.Y(n_974)
);

AOI21xp5_ASAP7_75t_L g975 ( 
.A1(n_783),
.A2(n_655),
.B(n_611),
.Y(n_975)
);

AOI21xp5_ASAP7_75t_L g976 ( 
.A1(n_785),
.A2(n_623),
.B(n_640),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_708),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_716),
.Y(n_978)
);

INVx1_ASAP7_75t_L g979 ( 
.A(n_725),
.Y(n_979)
);

OAI22xp5_ASAP7_75t_L g980 ( 
.A1(n_731),
.A2(n_591),
.B1(n_602),
.B2(n_585),
.Y(n_980)
);

BUFx4f_ASAP7_75t_L g981 ( 
.A(n_726),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_730),
.B(n_591),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_726),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_738),
.B(n_591),
.Y(n_984)
);

AOI22xp5_ASAP7_75t_L g985 ( 
.A1(n_860),
.A2(n_646),
.B1(n_638),
.B2(n_580),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_841),
.B(n_602),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_741),
.B(n_602),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_796),
.A2(n_753),
.B(n_800),
.Y(n_988)
);

AO21x1_ASAP7_75t_L g989 ( 
.A1(n_731),
.A2(n_617),
.B(n_640),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_715),
.Y(n_990)
);

A2O1A1Ixp33_ASAP7_75t_L g991 ( 
.A1(n_838),
.A2(n_831),
.B(n_820),
.C(n_767),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_815),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_744),
.B(n_751),
.Y(n_993)
);

AND2x2_ASAP7_75t_L g994 ( 
.A(n_769),
.B(n_808),
.Y(n_994)
);

HB1xp67_ASAP7_75t_L g995 ( 
.A(n_745),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_815),
.B(n_611),
.Y(n_996)
);

AOI21xp5_ASAP7_75t_L g997 ( 
.A1(n_813),
.A2(n_623),
.B(n_640),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_737),
.A2(n_617),
.B(n_614),
.Y(n_998)
);

INVx3_ASAP7_75t_L g999 ( 
.A(n_815),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_737),
.A2(n_617),
.B(n_614),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_792),
.A2(n_616),
.B(n_614),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_L g1002 ( 
.A(n_815),
.B(n_616),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_802),
.A2(n_616),
.B1(n_635),
.B2(n_631),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_859),
.B(n_623),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_858),
.B(n_627),
.Y(n_1005)
);

INVx2_ASAP7_75t_L g1006 ( 
.A(n_811),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_816),
.Y(n_1007)
);

O2A1O1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_849),
.A2(n_627),
.B(n_631),
.C(n_635),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_840),
.A2(n_768),
.B(n_797),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_835),
.Y(n_1010)
);

A2O1A1Ixp33_ASAP7_75t_L g1011 ( 
.A1(n_831),
.A2(n_635),
.B(n_631),
.C(n_577),
.Y(n_1011)
);

OAI22xp5_ASAP7_75t_L g1012 ( 
.A1(n_799),
.A2(n_577),
.B1(n_589),
.B2(n_588),
.Y(n_1012)
);

AOI21xp5_ASAP7_75t_L g1013 ( 
.A1(n_801),
.A2(n_589),
.B(n_588),
.Y(n_1013)
);

INVxp67_ASAP7_75t_L g1014 ( 
.A(n_793),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_777),
.B(n_352),
.Y(n_1015)
);

INVxp67_ASAP7_75t_L g1016 ( 
.A(n_791),
.Y(n_1016)
);

BUFx6f_ASAP7_75t_L g1017 ( 
.A(n_823),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_718),
.A2(n_646),
.B1(n_638),
.B2(n_580),
.Y(n_1018)
);

AOI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_810),
.A2(n_589),
.B(n_588),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_842),
.B(n_646),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_L g1021 ( 
.A(n_846),
.B(n_646),
.Y(n_1021)
);

AND2x2_ASAP7_75t_L g1022 ( 
.A(n_748),
.B(n_488),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_847),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_854),
.Y(n_1024)
);

OAI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_829),
.A2(n_556),
.B(n_582),
.Y(n_1025)
);

INVx2_ASAP7_75t_L g1026 ( 
.A(n_694),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_851),
.A2(n_577),
.B(n_582),
.Y(n_1027)
);

O2A1O1Ixp33_ASAP7_75t_L g1028 ( 
.A1(n_832),
.A2(n_529),
.B(n_520),
.C(n_533),
.Y(n_1028)
);

INVx2_ASAP7_75t_L g1029 ( 
.A(n_697),
.Y(n_1029)
);

INVx2_ASAP7_75t_L g1030 ( 
.A(n_736),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_803),
.B(n_638),
.Y(n_1031)
);

AO21x1_ASAP7_75t_L g1032 ( 
.A1(n_857),
.A2(n_582),
.B(n_579),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_746),
.B(n_646),
.Y(n_1033)
);

NOR2xp33_ASAP7_75t_L g1034 ( 
.A(n_807),
.B(n_277),
.Y(n_1034)
);

INVx4_ASAP7_75t_L g1035 ( 
.A(n_764),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_833),
.B(n_638),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_834),
.B(n_646),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_836),
.B(n_556),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_852),
.A2(n_579),
.B(n_465),
.Y(n_1039)
);

NOR2xp33_ASAP7_75t_L g1040 ( 
.A(n_750),
.B(n_279),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_839),
.Y(n_1041)
);

AOI21xp5_ASAP7_75t_L g1042 ( 
.A1(n_853),
.A2(n_579),
.B(n_465),
.Y(n_1042)
);

NOR3xp33_ASAP7_75t_L g1043 ( 
.A(n_762),
.B(n_353),
.C(n_285),
.Y(n_1043)
);

AOI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_775),
.A2(n_845),
.B(n_857),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_856),
.A2(n_529),
.B(n_520),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_827),
.B(n_526),
.Y(n_1046)
);

AOI21xp5_ASAP7_75t_L g1047 ( 
.A1(n_848),
.A2(n_537),
.B(n_533),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_766),
.B(n_526),
.Y(n_1048)
);

NAND3xp33_ASAP7_75t_L g1049 ( 
.A(n_869),
.B(n_837),
.C(n_826),
.Y(n_1049)
);

AND2x2_ASAP7_75t_L g1050 ( 
.A(n_968),
.B(n_718),
.Y(n_1050)
);

CKINVDCx5p33_ASAP7_75t_R g1051 ( 
.A(n_873),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_877),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_863),
.B(n_784),
.Y(n_1053)
);

A2O1A1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_935),
.A2(n_844),
.B(n_718),
.C(n_778),
.Y(n_1054)
);

OAI22xp5_ASAP7_75t_L g1055 ( 
.A1(n_862),
.A2(n_357),
.B1(n_289),
.B2(n_300),
.Y(n_1055)
);

AOI22xp33_ASAP7_75t_SL g1056 ( 
.A1(n_1034),
.A2(n_763),
.B1(n_354),
.B2(n_347),
.Y(n_1056)
);

NAND2xp5_ASAP7_75t_L g1057 ( 
.A(n_967),
.B(n_526),
.Y(n_1057)
);

AO21x2_ASAP7_75t_L g1058 ( 
.A1(n_888),
.A2(n_493),
.B(n_488),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_899),
.A2(n_526),
.B(n_537),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_864),
.B(n_529),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_939),
.B(n_283),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_900),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_885),
.B(n_488),
.Y(n_1063)
);

NOR3xp33_ASAP7_75t_SL g1064 ( 
.A(n_931),
.B(n_304),
.C(n_305),
.Y(n_1064)
);

INVx2_ASAP7_75t_SL g1065 ( 
.A(n_916),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_1022),
.B(n_529),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_974),
.A2(n_580),
.B1(n_493),
.B2(n_537),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_915),
.A2(n_533),
.B(n_487),
.Y(n_1068)
);

BUFx6f_ASAP7_75t_L g1069 ( 
.A(n_983),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_924),
.B(n_906),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_983),
.Y(n_1071)
);

INVx5_ASAP7_75t_L g1072 ( 
.A(n_983),
.Y(n_1072)
);

INVx2_ASAP7_75t_L g1073 ( 
.A(n_874),
.Y(n_1073)
);

A2O1A1Ixp33_ASAP7_75t_L g1074 ( 
.A1(n_881),
.A2(n_493),
.B(n_307),
.C(n_359),
.Y(n_1074)
);

O2A1O1Ixp5_ASAP7_75t_L g1075 ( 
.A1(n_865),
.A2(n_533),
.B(n_494),
.C(n_491),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_898),
.Y(n_1076)
);

NOR2xp33_ASAP7_75t_L g1077 ( 
.A(n_995),
.B(n_309),
.Y(n_1077)
);

NOR2xp33_ASAP7_75t_L g1078 ( 
.A(n_917),
.B(n_330),
.Y(n_1078)
);

AOI21xp5_ASAP7_75t_L g1079 ( 
.A1(n_915),
.A2(n_494),
.B(n_491),
.Y(n_1079)
);

INVx6_ASAP7_75t_L g1080 ( 
.A(n_1017),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_941),
.B(n_366),
.C(n_339),
.Y(n_1081)
);

BUFx6f_ASAP7_75t_L g1082 ( 
.A(n_951),
.Y(n_1082)
);

OAI22xp5_ASAP7_75t_SL g1083 ( 
.A1(n_901),
.A2(n_334),
.B1(n_344),
.B2(n_345),
.Y(n_1083)
);

INVx4_ASAP7_75t_L g1084 ( 
.A(n_922),
.Y(n_1084)
);

NOR2xp33_ASAP7_75t_R g1085 ( 
.A(n_981),
.B(n_346),
.Y(n_1085)
);

OAI21xp33_ASAP7_75t_SL g1086 ( 
.A1(n_936),
.A2(n_487),
.B(n_491),
.Y(n_1086)
);

NOR2xp33_ASAP7_75t_L g1087 ( 
.A(n_902),
.B(n_360),
.Y(n_1087)
);

BUFx6f_ASAP7_75t_L g1088 ( 
.A(n_951),
.Y(n_1088)
);

AO32x1_ASAP7_75t_L g1089 ( 
.A1(n_1012),
.A2(n_494),
.A3(n_491),
.B1(n_487),
.B2(n_580),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_881),
.A2(n_991),
.B(n_1016),
.C(n_1014),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1017),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_952),
.B(n_929),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_861),
.B(n_11),
.Y(n_1093)
);

BUFx3_ASAP7_75t_L g1094 ( 
.A(n_1017),
.Y(n_1094)
);

AOI21xp5_ASAP7_75t_L g1095 ( 
.A1(n_930),
.A2(n_494),
.B(n_487),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_SL g1096 ( 
.A1(n_1040),
.A2(n_580),
.B(n_538),
.C(n_77),
.Y(n_1096)
);

NOR3xp33_ASAP7_75t_L g1097 ( 
.A(n_945),
.B(n_13),
.C(n_14),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_977),
.B(n_580),
.Y(n_1098)
);

AOI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_930),
.A2(n_489),
.B(n_492),
.Y(n_1099)
);

AOI21xp5_ASAP7_75t_L g1100 ( 
.A1(n_940),
.A2(n_489),
.B(n_492),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_919),
.A2(n_489),
.B1(n_490),
.B2(n_492),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_979),
.B(n_927),
.Y(n_1102)
);

AND2x6_ASAP7_75t_L g1103 ( 
.A(n_999),
.B(n_489),
.Y(n_1103)
);

OAI22xp5_ASAP7_75t_L g1104 ( 
.A1(n_919),
.A2(n_908),
.B1(n_957),
.B2(n_946),
.Y(n_1104)
);

BUFx2_ASAP7_75t_L g1105 ( 
.A(n_891),
.Y(n_1105)
);

BUFx2_ASAP7_75t_L g1106 ( 
.A(n_885),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_940),
.A2(n_489),
.B(n_492),
.Y(n_1107)
);

BUFx2_ASAP7_75t_L g1108 ( 
.A(n_925),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_1006),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_919),
.A2(n_489),
.B1(n_490),
.B2(n_492),
.Y(n_1110)
);

OR2x2_ASAP7_75t_L g1111 ( 
.A(n_961),
.B(n_489),
.Y(n_1111)
);

BUFx6f_ASAP7_75t_L g1112 ( 
.A(n_951),
.Y(n_1112)
);

NOR2xp33_ASAP7_75t_R g1113 ( 
.A(n_981),
.B(n_73),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_L g1114 ( 
.A(n_978),
.B(n_492),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_L g1115 ( 
.A(n_878),
.B(n_14),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_954),
.A2(n_489),
.B(n_492),
.Y(n_1116)
);

INVx2_ASAP7_75t_L g1117 ( 
.A(n_1007),
.Y(n_1117)
);

AOI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_880),
.A2(n_897),
.B1(n_925),
.B2(n_870),
.Y(n_1118)
);

NOR3xp33_ASAP7_75t_SL g1119 ( 
.A(n_1015),
.B(n_15),
.C(n_16),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_993),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_SL g1121 ( 
.A(n_922),
.B(n_490),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_SL g1122 ( 
.A(n_922),
.B(n_490),
.Y(n_1122)
);

BUFx6f_ASAP7_75t_SL g1123 ( 
.A(n_990),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_960),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_988),
.A2(n_490),
.B(n_19),
.C(n_21),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_886),
.B(n_490),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_919),
.A2(n_490),
.B1(n_22),
.B2(n_23),
.Y(n_1127)
);

BUFx2_ASAP7_75t_L g1128 ( 
.A(n_897),
.Y(n_1128)
);

AO32x2_ASAP7_75t_L g1129 ( 
.A1(n_909),
.A2(n_16),
.A3(n_22),
.B1(n_26),
.B2(n_27),
.Y(n_1129)
);

A2O1A1Ixp33_ASAP7_75t_L g1130 ( 
.A1(n_988),
.A2(n_28),
.B(n_29),
.C(n_30),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_992),
.A2(n_29),
.B1(n_34),
.B2(n_35),
.Y(n_1131)
);

AND2x2_ASAP7_75t_L g1132 ( 
.A(n_994),
.B(n_34),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_893),
.B(n_538),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1010),
.Y(n_1134)
);

A2O1A1Ixp33_ASAP7_75t_SL g1135 ( 
.A1(n_871),
.A2(n_538),
.B(n_96),
.C(n_99),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_894),
.B(n_538),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_954),
.A2(n_94),
.B(n_173),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_903),
.B(n_538),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_928),
.B(n_88),
.Y(n_1139)
);

BUFx2_ASAP7_75t_L g1140 ( 
.A(n_928),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_SL g1141 ( 
.A(n_928),
.B(n_108),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_942),
.B(n_36),
.Y(n_1142)
);

AOI33xp33_ASAP7_75t_L g1143 ( 
.A1(n_938),
.A2(n_1018),
.A3(n_933),
.B1(n_1023),
.B2(n_892),
.B3(n_1029),
.Y(n_1143)
);

AND2x4_ASAP7_75t_L g1144 ( 
.A(n_942),
.B(n_960),
.Y(n_1144)
);

BUFx8_ASAP7_75t_SL g1145 ( 
.A(n_960),
.Y(n_1145)
);

AND2x4_ASAP7_75t_L g1146 ( 
.A(n_942),
.B(n_118),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_943),
.A2(n_84),
.B(n_172),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_890),
.A2(n_82),
.B(n_171),
.Y(n_1148)
);

NAND2xp5_ASAP7_75t_L g1149 ( 
.A(n_904),
.B(n_538),
.Y(n_1149)
);

BUFx3_ASAP7_75t_L g1150 ( 
.A(n_992),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1026),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1043),
.B(n_44),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1030),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1046),
.A2(n_45),
.B(n_49),
.C(n_50),
.Y(n_1154)
);

OAI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_998),
.A2(n_538),
.B(n_131),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_992),
.B(n_122),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_1024),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_1041),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_895),
.Y(n_1159)
);

NOR3xp33_ASAP7_75t_SL g1160 ( 
.A(n_905),
.B(n_45),
.C(n_51),
.Y(n_1160)
);

INVx2_ASAP7_75t_SL g1161 ( 
.A(n_879),
.Y(n_1161)
);

BUFx3_ASAP7_75t_L g1162 ( 
.A(n_1024),
.Y(n_1162)
);

OAI22xp5_ASAP7_75t_L g1163 ( 
.A1(n_866),
.A2(n_51),
.B1(n_54),
.B2(n_61),
.Y(n_1163)
);

OAI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_999),
.A2(n_62),
.B1(n_63),
.B2(n_64),
.Y(n_1164)
);

AND2x2_ASAP7_75t_L g1165 ( 
.A(n_918),
.B(n_948),
.Y(n_1165)
);

INVx4_ASAP7_75t_L g1166 ( 
.A(n_907),
.Y(n_1166)
);

AOI221xp5_ASAP7_75t_L g1167 ( 
.A1(n_937),
.A2(n_62),
.B1(n_64),
.B2(n_66),
.C(n_81),
.Y(n_1167)
);

O2A1O1Ixp33_ASAP7_75t_L g1168 ( 
.A1(n_986),
.A2(n_66),
.B(n_538),
.C(n_134),
.Y(n_1168)
);

BUFx6f_ASAP7_75t_L g1169 ( 
.A(n_907),
.Y(n_1169)
);

INVx2_ASAP7_75t_SL g1170 ( 
.A(n_1035),
.Y(n_1170)
);

NAND3xp33_ASAP7_75t_L g1171 ( 
.A(n_1011),
.B(n_133),
.C(n_139),
.Y(n_1171)
);

BUFx3_ASAP7_75t_L g1172 ( 
.A(n_944),
.Y(n_1172)
);

NOR3xp33_ASAP7_75t_SL g1173 ( 
.A(n_971),
.B(n_932),
.C(n_889),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1005),
.Y(n_1174)
);

INVx2_ASAP7_75t_L g1175 ( 
.A(n_1004),
.Y(n_1175)
);

A2O1A1Ixp33_ASAP7_75t_L g1176 ( 
.A1(n_889),
.A2(n_142),
.B(n_147),
.C(n_148),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_911),
.B(n_167),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_996),
.B(n_170),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_SL g1179 ( 
.A(n_1031),
.B(n_1002),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_955),
.A2(n_956),
.B(n_875),
.Y(n_1180)
);

BUFx8_ASAP7_75t_L g1181 ( 
.A(n_867),
.Y(n_1181)
);

BUFx3_ASAP7_75t_L g1182 ( 
.A(n_944),
.Y(n_1182)
);

AND2x6_ASAP7_75t_L g1183 ( 
.A(n_985),
.B(n_934),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_913),
.A2(n_914),
.B(n_923),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_947),
.B(n_949),
.Y(n_1185)
);

OAI22xp5_ASAP7_75t_SL g1186 ( 
.A1(n_972),
.A2(n_896),
.B1(n_963),
.B2(n_962),
.Y(n_1186)
);

O2A1O1Ixp33_ASAP7_75t_L g1187 ( 
.A1(n_950),
.A2(n_921),
.B(n_982),
.C(n_1008),
.Y(n_1187)
);

INVx5_ASAP7_75t_L g1188 ( 
.A(n_989),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_1038),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1000),
.B(n_912),
.Y(n_1190)
);

A2O1A1Ixp33_ASAP7_75t_L g1191 ( 
.A1(n_964),
.A2(n_910),
.B(n_912),
.C(n_876),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_913),
.A2(n_914),
.B(n_958),
.Y(n_1192)
);

NAND3xp33_ASAP7_75t_SL g1193 ( 
.A(n_1009),
.B(n_972),
.C(n_1048),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_959),
.A2(n_1044),
.B(n_980),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_984),
.Y(n_1195)
);

BUFx6f_ASAP7_75t_L g1196 ( 
.A(n_987),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1028),
.Y(n_1197)
);

O2A1O1Ixp33_ASAP7_75t_L g1198 ( 
.A1(n_970),
.A2(n_1003),
.B(n_953),
.C(n_920),
.Y(n_1198)
);

AOI21xp5_ASAP7_75t_L g1199 ( 
.A1(n_1044),
.A2(n_868),
.B(n_872),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_926),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_882),
.Y(n_1201)
);

NAND2xp5_ASAP7_75t_L g1202 ( 
.A(n_1001),
.B(n_868),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_SL g1203 ( 
.A(n_965),
.B(n_1020),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_SL g1204 ( 
.A(n_1021),
.B(n_1033),
.Y(n_1204)
);

NAND2xp5_ASAP7_75t_L g1205 ( 
.A(n_872),
.B(n_876),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1052),
.Y(n_1206)
);

OAI21x1_ASAP7_75t_SL g1207 ( 
.A1(n_1137),
.A2(n_1032),
.B(n_910),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_SL g1208 ( 
.A(n_1062),
.B(n_1037),
.Y(n_1208)
);

AOI21xp5_ASAP7_75t_L g1209 ( 
.A1(n_1180),
.A2(n_1025),
.B(n_1001),
.Y(n_1209)
);

HB1xp67_ASAP7_75t_L g1210 ( 
.A(n_1105),
.Y(n_1210)
);

HB1xp67_ASAP7_75t_L g1211 ( 
.A(n_1065),
.Y(n_1211)
);

AOI21xp5_ASAP7_75t_L g1212 ( 
.A1(n_1190),
.A2(n_973),
.B(n_976),
.Y(n_1212)
);

AO31x2_ASAP7_75t_L g1213 ( 
.A1(n_1191),
.A2(n_1047),
.A3(n_976),
.B(n_975),
.Y(n_1213)
);

INVx5_ASAP7_75t_L g1214 ( 
.A(n_1069),
.Y(n_1214)
);

NAND2x1p5_ASAP7_75t_L g1215 ( 
.A(n_1072),
.B(n_884),
.Y(n_1215)
);

A2O1A1Ixp33_ASAP7_75t_L g1216 ( 
.A1(n_1053),
.A2(n_969),
.B(n_966),
.C(n_1013),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1090),
.A2(n_1202),
.B(n_1192),
.Y(n_1217)
);

BUFx3_ASAP7_75t_L g1218 ( 
.A(n_1091),
.Y(n_1218)
);

AOI21xp5_ASAP7_75t_L g1219 ( 
.A1(n_1202),
.A2(n_1205),
.B(n_1184),
.Y(n_1219)
);

AND2x4_ASAP7_75t_L g1220 ( 
.A(n_1144),
.B(n_883),
.Y(n_1220)
);

OAI21xp33_ASAP7_75t_L g1221 ( 
.A1(n_1077),
.A2(n_1036),
.B(n_887),
.Y(n_1221)
);

OAI21xp33_ASAP7_75t_SL g1222 ( 
.A1(n_1155),
.A2(n_973),
.B(n_975),
.Y(n_1222)
);

AOI221xp5_ASAP7_75t_SL g1223 ( 
.A1(n_1115),
.A2(n_997),
.B1(n_1013),
.B2(n_1019),
.C(n_1039),
.Y(n_1223)
);

AND2x4_ASAP7_75t_L g1224 ( 
.A(n_1144),
.B(n_1019),
.Y(n_1224)
);

AOI221x1_ASAP7_75t_L g1225 ( 
.A1(n_1163),
.A2(n_1047),
.B1(n_997),
.B2(n_1045),
.C(n_1042),
.Y(n_1225)
);

NOR3xp33_ASAP7_75t_L g1226 ( 
.A(n_1081),
.B(n_1027),
.C(n_1045),
.Y(n_1226)
);

AOI21xp5_ASAP7_75t_L g1227 ( 
.A1(n_1194),
.A2(n_1057),
.B(n_1199),
.Y(n_1227)
);

BUFx2_ASAP7_75t_R g1228 ( 
.A(n_1145),
.Y(n_1228)
);

OAI22xp5_ASAP7_75t_L g1229 ( 
.A1(n_1092),
.A2(n_1120),
.B1(n_1054),
.B2(n_1049),
.Y(n_1229)
);

BUFx10_ASAP7_75t_L g1230 ( 
.A(n_1051),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1161),
.B(n_1124),
.Y(n_1231)
);

NOR2xp33_ASAP7_75t_L g1232 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1232)
);

AO31x2_ASAP7_75t_L g1233 ( 
.A1(n_1104),
.A2(n_1074),
.A3(n_1201),
.B(n_1125),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1069),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1092),
.A2(n_1050),
.B1(n_1102),
.B2(n_1170),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1068),
.A2(n_1095),
.B(n_1079),
.Y(n_1236)
);

AO21x1_ASAP7_75t_L g1237 ( 
.A1(n_1104),
.A2(n_1155),
.B(n_1163),
.Y(n_1237)
);

AOI21xp5_ASAP7_75t_L g1238 ( 
.A1(n_1193),
.A2(n_1060),
.B(n_1198),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1174),
.B(n_1175),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1179),
.A2(n_1178),
.B(n_1195),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1060),
.A2(n_1185),
.B(n_1187),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_L g1242 ( 
.A(n_1159),
.B(n_1189),
.Y(n_1242)
);

AO21x1_ASAP7_75t_L g1243 ( 
.A1(n_1127),
.A2(n_1197),
.B(n_1148),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1106),
.Y(n_1244)
);

AOI21xp5_ASAP7_75t_SL g1245 ( 
.A1(n_1176),
.A2(n_1146),
.B(n_1066),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1073),
.Y(n_1246)
);

HB1xp67_ASAP7_75t_L g1247 ( 
.A(n_1140),
.Y(n_1247)
);

AOI21xp5_ASAP7_75t_L g1248 ( 
.A1(n_1203),
.A2(n_1177),
.B(n_1186),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1099),
.A2(n_1100),
.A3(n_1116),
.B(n_1107),
.Y(n_1249)
);

AND2x6_ASAP7_75t_L g1250 ( 
.A(n_1146),
.B(n_1157),
.Y(n_1250)
);

NAND3xp33_ASAP7_75t_L g1251 ( 
.A(n_1081),
.B(n_1056),
.C(n_1097),
.Y(n_1251)
);

BUFx6f_ASAP7_75t_L g1252 ( 
.A(n_1069),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1126),
.A2(n_1204),
.B(n_1133),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1063),
.B(n_1132),
.Y(n_1254)
);

NOR2xp67_ASAP7_75t_SL g1255 ( 
.A(n_1072),
.B(n_1157),
.Y(n_1255)
);

NAND3xp33_ASAP7_75t_L g1256 ( 
.A(n_1064),
.B(n_1078),
.C(n_1061),
.Y(n_1256)
);

OAI21x1_ASAP7_75t_SL g1257 ( 
.A1(n_1147),
.A2(n_1168),
.B(n_1131),
.Y(n_1257)
);

OAI21x1_ASAP7_75t_L g1258 ( 
.A1(n_1200),
.A2(n_1075),
.B(n_1059),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1169),
.Y(n_1259)
);

A2O1A1Ixp33_ASAP7_75t_L g1260 ( 
.A1(n_1173),
.A2(n_1171),
.B(n_1118),
.C(n_1167),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1063),
.B(n_1109),
.Y(n_1261)
);

OAI21xp33_ASAP7_75t_SL g1262 ( 
.A1(n_1143),
.A2(n_1076),
.B(n_1127),
.Y(n_1262)
);

OAI21x1_ASAP7_75t_L g1263 ( 
.A1(n_1114),
.A2(n_1138),
.B(n_1149),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1117),
.B(n_1134),
.Y(n_1264)
);

OR2x4_ASAP7_75t_L g1265 ( 
.A(n_1093),
.B(n_1082),
.Y(n_1265)
);

AO21x1_ASAP7_75t_L g1266 ( 
.A1(n_1131),
.A2(n_1164),
.B(n_1156),
.Y(n_1266)
);

O2A1O1Ixp33_ASAP7_75t_L g1267 ( 
.A1(n_1154),
.A2(n_1130),
.B(n_1055),
.C(n_1152),
.Y(n_1267)
);

OAI21x1_ASAP7_75t_L g1268 ( 
.A1(n_1136),
.A2(n_1110),
.B(n_1101),
.Y(n_1268)
);

AO32x2_ASAP7_75t_L g1269 ( 
.A1(n_1164),
.A2(n_1055),
.A3(n_1129),
.B1(n_1083),
.B2(n_1166),
.Y(n_1269)
);

AO31x2_ASAP7_75t_L g1270 ( 
.A1(n_1101),
.A2(n_1110),
.A3(n_1089),
.B(n_1098),
.Y(n_1270)
);

AND2x2_ASAP7_75t_L g1271 ( 
.A(n_1108),
.B(n_1128),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1162),
.A2(n_1172),
.B1(n_1182),
.B2(n_1157),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1072),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1142),
.B(n_1158),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1151),
.B(n_1153),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1058),
.Y(n_1276)
);

OAI21x1_ASAP7_75t_L g1277 ( 
.A1(n_1121),
.A2(n_1122),
.B(n_1171),
.Y(n_1277)
);

NOR2xp67_ASAP7_75t_SL g1278 ( 
.A(n_1071),
.B(n_1094),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1165),
.B(n_1196),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_SL g1280 ( 
.A(n_1082),
.B(n_1112),
.Y(n_1280)
);

NAND2x1p5_ASAP7_75t_L g1281 ( 
.A(n_1071),
.B(n_1084),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1058),
.Y(n_1282)
);

NAND3xp33_ASAP7_75t_L g1283 ( 
.A(n_1160),
.B(n_1119),
.C(n_1181),
.Y(n_1283)
);

AOI21xp5_ASAP7_75t_L g1284 ( 
.A1(n_1089),
.A2(n_1188),
.B(n_1086),
.Y(n_1284)
);

AOI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1089),
.A2(n_1188),
.B(n_1196),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1196),
.B(n_1084),
.Y(n_1286)
);

OAI21xp5_ASAP7_75t_SL g1287 ( 
.A1(n_1139),
.A2(n_1141),
.B(n_1067),
.Y(n_1287)
);

OA21x2_ASAP7_75t_L g1288 ( 
.A1(n_1111),
.A2(n_1188),
.B(n_1183),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_SL g1289 ( 
.A1(n_1080),
.A2(n_1150),
.B1(n_1088),
.B2(n_1082),
.Y(n_1289)
);

AO31x2_ASAP7_75t_L g1290 ( 
.A1(n_1166),
.A2(n_1129),
.A3(n_1183),
.B(n_1135),
.Y(n_1290)
);

OAI21x1_ASAP7_75t_L g1291 ( 
.A1(n_1183),
.A2(n_1103),
.B(n_1096),
.Y(n_1291)
);

INVx4_ASAP7_75t_L g1292 ( 
.A(n_1088),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1129),
.Y(n_1293)
);

AND2x4_ASAP7_75t_L g1294 ( 
.A(n_1088),
.B(n_1112),
.Y(n_1294)
);

AO31x2_ASAP7_75t_L g1295 ( 
.A1(n_1183),
.A2(n_1181),
.A3(n_1103),
.B(n_1113),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_1103),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1112),
.B(n_1085),
.Y(n_1297)
);

BUFx3_ASAP7_75t_L g1298 ( 
.A(n_1080),
.Y(n_1298)
);

AOI221x1_ASAP7_75t_L g1299 ( 
.A1(n_1103),
.A2(n_869),
.B1(n_1163),
.B2(n_935),
.C(n_718),
.Y(n_1299)
);

NOR2xp33_ASAP7_75t_SL g1300 ( 
.A(n_1123),
.B(n_786),
.Y(n_1300)
);

OAI22xp33_ASAP7_75t_L g1301 ( 
.A1(n_1123),
.A2(n_547),
.B1(n_755),
.B2(n_863),
.Y(n_1301)
);

OAI22x1_ASAP7_75t_L g1302 ( 
.A1(n_1115),
.A2(n_968),
.B1(n_1053),
.B2(n_935),
.Y(n_1302)
);

OAI21x1_ASAP7_75t_L g1303 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1053),
.B(n_735),
.Y(n_1304)
);

O2A1O1Ixp5_ASAP7_75t_L g1305 ( 
.A1(n_1087),
.A2(n_935),
.B(n_863),
.C(n_864),
.Y(n_1305)
);

AO31x2_ASAP7_75t_L g1306 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1306)
);

OAI21x1_ASAP7_75t_L g1307 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1053),
.B(n_742),
.Y(n_1308)
);

OAI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1092),
.A2(n_863),
.B1(n_869),
.B2(n_968),
.Y(n_1309)
);

BUFx3_ASAP7_75t_L g1310 ( 
.A(n_1062),
.Y(n_1310)
);

INVx1_ASAP7_75t_L g1311 ( 
.A(n_1052),
.Y(n_1311)
);

OAI21x1_ASAP7_75t_L g1312 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1312)
);

AO31x2_ASAP7_75t_L g1313 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1075),
.A2(n_1199),
.B(n_1192),
.Y(n_1314)
);

OR2x6_ASAP7_75t_L g1315 ( 
.A(n_1161),
.B(n_726),
.Y(n_1315)
);

AOI21xp5_ASAP7_75t_L g1316 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1316)
);

O2A1O1Ixp33_ASAP7_75t_L g1317 ( 
.A1(n_1054),
.A2(n_869),
.B(n_935),
.C(n_863),
.Y(n_1317)
);

AOI21xp5_ASAP7_75t_L g1318 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1318)
);

AOI21xp5_ASAP7_75t_L g1319 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1319)
);

AO31x2_ASAP7_75t_L g1320 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1320)
);

A2O1A1Ixp33_ASAP7_75t_L g1321 ( 
.A1(n_1053),
.A2(n_869),
.B(n_863),
.C(n_935),
.Y(n_1321)
);

INVx1_ASAP7_75t_L g1322 ( 
.A(n_1052),
.Y(n_1322)
);

BUFx3_ASAP7_75t_L g1323 ( 
.A(n_1062),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1053),
.B(n_862),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1053),
.B(n_742),
.Y(n_1325)
);

O2A1O1Ixp33_ASAP7_75t_SL g1326 ( 
.A1(n_1054),
.A2(n_864),
.B(n_863),
.C(n_974),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1053),
.B(n_862),
.Y(n_1327)
);

OAI22xp5_ASAP7_75t_L g1328 ( 
.A1(n_1092),
.A2(n_863),
.B1(n_869),
.B2(n_968),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1090),
.A2(n_863),
.B(n_869),
.Y(n_1330)
);

AOI21x1_ASAP7_75t_L g1331 ( 
.A1(n_1190),
.A2(n_1202),
.B(n_1179),
.Y(n_1331)
);

AO21x2_ASAP7_75t_L g1332 ( 
.A1(n_1193),
.A2(n_1199),
.B(n_1192),
.Y(n_1332)
);

AOI21xp5_ASAP7_75t_L g1333 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1333)
);

AOI21xp5_ASAP7_75t_L g1334 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1053),
.A2(n_869),
.B1(n_968),
.B2(n_935),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1062),
.Y(n_1336)
);

AO31x2_ASAP7_75t_L g1337 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1087),
.B(n_935),
.C(n_869),
.Y(n_1339)
);

INVx2_ASAP7_75t_SL g1340 ( 
.A(n_1080),
.Y(n_1340)
);

AOI21xp33_ASAP7_75t_L g1341 ( 
.A1(n_1053),
.A2(n_935),
.B(n_869),
.Y(n_1341)
);

NOR2xp67_ASAP7_75t_L g1342 ( 
.A(n_1049),
.B(n_573),
.Y(n_1342)
);

NOR2xp67_ASAP7_75t_SL g1343 ( 
.A(n_1072),
.B(n_578),
.Y(n_1343)
);

AOI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1344)
);

AO31x2_ASAP7_75t_L g1345 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1345)
);

NOR2xp33_ASAP7_75t_L g1346 ( 
.A(n_1053),
.B(n_707),
.Y(n_1346)
);

AOI22x1_ASAP7_75t_L g1347 ( 
.A1(n_1197),
.A2(n_967),
.B1(n_945),
.B2(n_1180),
.Y(n_1347)
);

OAI21x1_ASAP7_75t_L g1348 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1053),
.B(n_707),
.Y(n_1349)
);

AOI221xp5_ASAP7_75t_SL g1350 ( 
.A1(n_1115),
.A2(n_869),
.B1(n_935),
.B2(n_784),
.C(n_968),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1052),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1052),
.Y(n_1352)
);

AOI21xp5_ASAP7_75t_L g1353 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1354)
);

OAI21x1_ASAP7_75t_L g1355 ( 
.A1(n_1068),
.A2(n_884),
.B(n_1079),
.Y(n_1355)
);

INVx5_ASAP7_75t_L g1356 ( 
.A(n_1069),
.Y(n_1356)
);

OR2x2_ASAP7_75t_L g1357 ( 
.A(n_1053),
.B(n_735),
.Y(n_1357)
);

AND2x6_ASAP7_75t_L g1358 ( 
.A(n_1146),
.B(n_992),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1052),
.Y(n_1359)
);

AOI21xp5_ASAP7_75t_L g1360 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1361)
);

AO31x2_ASAP7_75t_L g1362 ( 
.A1(n_1191),
.A2(n_1104),
.A3(n_1090),
.B(n_1199),
.Y(n_1362)
);

O2A1O1Ixp33_ASAP7_75t_SL g1363 ( 
.A1(n_1054),
.A2(n_864),
.B(n_863),
.C(n_974),
.Y(n_1363)
);

AOI21xp5_ASAP7_75t_L g1364 ( 
.A1(n_1180),
.A2(n_863),
.B(n_1190),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1206),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_L g1366 ( 
.A(n_1324),
.B(n_1327),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1335),
.A2(n_1328),
.B1(n_1309),
.B2(n_1232),
.Y(n_1367)
);

CKINVDCx20_ASAP7_75t_R g1368 ( 
.A(n_1310),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1302),
.A2(n_1341),
.B1(n_1339),
.B2(n_1335),
.Y(n_1369)
);

CKINVDCx11_ASAP7_75t_R g1370 ( 
.A(n_1230),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1346),
.B(n_1349),
.Y(n_1371)
);

AOI22xp33_ASAP7_75t_L g1372 ( 
.A1(n_1251),
.A2(n_1330),
.B1(n_1237),
.B2(n_1266),
.Y(n_1372)
);

BUFx3_ASAP7_75t_L g1373 ( 
.A(n_1298),
.Y(n_1373)
);

AOI22xp33_ASAP7_75t_L g1374 ( 
.A1(n_1256),
.A2(n_1308),
.B1(n_1325),
.B2(n_1283),
.Y(n_1374)
);

BUFx6f_ASAP7_75t_SL g1375 ( 
.A(n_1230),
.Y(n_1375)
);

OAI22xp5_ASAP7_75t_L g1376 ( 
.A1(n_1321),
.A2(n_1304),
.B1(n_1357),
.B2(n_1260),
.Y(n_1376)
);

CKINVDCx6p67_ASAP7_75t_R g1377 ( 
.A(n_1323),
.Y(n_1377)
);

AOI22xp33_ASAP7_75t_SL g1378 ( 
.A1(n_1300),
.A2(n_1229),
.B1(n_1257),
.B2(n_1347),
.Y(n_1378)
);

CKINVDCx8_ASAP7_75t_R g1379 ( 
.A(n_1214),
.Y(n_1379)
);

INVx6_ASAP7_75t_L g1380 ( 
.A(n_1214),
.Y(n_1380)
);

CKINVDCx20_ASAP7_75t_R g1381 ( 
.A(n_1336),
.Y(n_1381)
);

CKINVDCx20_ASAP7_75t_R g1382 ( 
.A(n_1265),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1206),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1275),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1301),
.A2(n_1243),
.B1(n_1274),
.B2(n_1235),
.Y(n_1385)
);

NAND2x1p5_ASAP7_75t_L g1386 ( 
.A(n_1255),
.B(n_1356),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1342),
.A2(n_1242),
.B1(n_1224),
.B2(n_1240),
.Y(n_1387)
);

OAI22xp5_ASAP7_75t_L g1388 ( 
.A1(n_1254),
.A2(n_1317),
.B1(n_1239),
.B2(n_1279),
.Y(n_1388)
);

CKINVDCx14_ASAP7_75t_R g1389 ( 
.A(n_1271),
.Y(n_1389)
);

AOI22xp33_ASAP7_75t_L g1390 ( 
.A1(n_1342),
.A2(n_1224),
.B1(n_1350),
.B2(n_1238),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1262),
.A2(n_1217),
.B1(n_1226),
.B2(n_1210),
.Y(n_1391)
);

INVx6_ASAP7_75t_L g1392 ( 
.A(n_1356),
.Y(n_1392)
);

BUFx3_ASAP7_75t_L g1393 ( 
.A(n_1218),
.Y(n_1393)
);

BUFx4f_ASAP7_75t_SL g1394 ( 
.A(n_1234),
.Y(n_1394)
);

OAI22xp5_ASAP7_75t_L g1395 ( 
.A1(n_1245),
.A2(n_1244),
.B1(n_1261),
.B2(n_1220),
.Y(n_1395)
);

INVx1_ASAP7_75t_SL g1396 ( 
.A(n_1211),
.Y(n_1396)
);

OAI22xp33_ASAP7_75t_SL g1397 ( 
.A1(n_1208),
.A2(n_1352),
.B1(n_1322),
.B2(n_1351),
.Y(n_1397)
);

NAND2x1p5_ASAP7_75t_L g1398 ( 
.A(n_1273),
.B(n_1278),
.Y(n_1398)
);

BUFx3_ASAP7_75t_L g1399 ( 
.A(n_1294),
.Y(n_1399)
);

AOI22xp33_ASAP7_75t_SL g1400 ( 
.A1(n_1250),
.A2(n_1358),
.B1(n_1262),
.B2(n_1297),
.Y(n_1400)
);

AOI22xp33_ASAP7_75t_SL g1401 ( 
.A1(n_1250),
.A2(n_1358),
.B1(n_1220),
.B2(n_1299),
.Y(n_1401)
);

INVx1_ASAP7_75t_SL g1402 ( 
.A(n_1247),
.Y(n_1402)
);

OAI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1311),
.A2(n_1322),
.B1(n_1359),
.B2(n_1352),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1234),
.Y(n_1404)
);

INVx1_ASAP7_75t_SL g1405 ( 
.A(n_1340),
.Y(n_1405)
);

BUFx3_ASAP7_75t_L g1406 ( 
.A(n_1231),
.Y(n_1406)
);

INVx1_ASAP7_75t_SL g1407 ( 
.A(n_1228),
.Y(n_1407)
);

AOI22xp33_ASAP7_75t_L g1408 ( 
.A1(n_1221),
.A2(n_1311),
.B1(n_1359),
.B2(n_1351),
.Y(n_1408)
);

OAI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1267),
.A2(n_1287),
.B1(n_1315),
.B2(n_1286),
.Y(n_1409)
);

OAI21xp5_ASAP7_75t_L g1410 ( 
.A1(n_1305),
.A2(n_1248),
.B(n_1241),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1264),
.B(n_1250),
.Y(n_1411)
);

CKINVDCx5p33_ASAP7_75t_R g1412 ( 
.A(n_1231),
.Y(n_1412)
);

AO22x1_ASAP7_75t_L g1413 ( 
.A1(n_1250),
.A2(n_1358),
.B1(n_1273),
.B2(n_1272),
.Y(n_1413)
);

BUFx12f_ASAP7_75t_L g1414 ( 
.A(n_1252),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1358),
.B(n_1326),
.Y(n_1415)
);

BUFx6f_ASAP7_75t_L g1416 ( 
.A(n_1252),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1246),
.A2(n_1364),
.B1(n_1318),
.B2(n_1316),
.Y(n_1417)
);

OAI22xp33_ASAP7_75t_L g1418 ( 
.A1(n_1293),
.A2(n_1315),
.B1(n_1319),
.B2(n_1333),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1280),
.Y(n_1419)
);

INVx6_ASAP7_75t_L g1420 ( 
.A(n_1252),
.Y(n_1420)
);

AOI22xp33_ASAP7_75t_SL g1421 ( 
.A1(n_1293),
.A2(n_1289),
.B1(n_1222),
.B2(n_1288),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1259),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1334),
.A2(n_1353),
.B1(n_1344),
.B2(n_1338),
.Y(n_1423)
);

AOI22xp33_ASAP7_75t_SL g1424 ( 
.A1(n_1222),
.A2(n_1288),
.B1(n_1269),
.B2(n_1291),
.Y(n_1424)
);

AOI22xp33_ASAP7_75t_L g1425 ( 
.A1(n_1360),
.A2(n_1332),
.B1(n_1276),
.B2(n_1282),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1363),
.B(n_1331),
.Y(n_1426)
);

OAI21xp5_ASAP7_75t_SL g1427 ( 
.A1(n_1216),
.A2(n_1209),
.B(n_1219),
.Y(n_1427)
);

BUFx3_ASAP7_75t_L g1428 ( 
.A(n_1281),
.Y(n_1428)
);

INVx3_ASAP7_75t_L g1429 ( 
.A(n_1292),
.Y(n_1429)
);

AOI22xp33_ASAP7_75t_L g1430 ( 
.A1(n_1332),
.A2(n_1253),
.B1(n_1212),
.B2(n_1343),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1269),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1269),
.Y(n_1432)
);

CKINVDCx14_ASAP7_75t_R g1433 ( 
.A(n_1292),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_1296),
.Y(n_1434)
);

AOI22xp33_ASAP7_75t_SL g1435 ( 
.A1(n_1207),
.A2(n_1277),
.B1(n_1296),
.B2(n_1285),
.Y(n_1435)
);

AOI22xp5_ASAP7_75t_SL g1436 ( 
.A1(n_1295),
.A2(n_1284),
.B1(n_1215),
.B2(n_1314),
.Y(n_1436)
);

BUFx2_ASAP7_75t_L g1437 ( 
.A(n_1295),
.Y(n_1437)
);

AOI22xp33_ASAP7_75t_L g1438 ( 
.A1(n_1227),
.A2(n_1314),
.B1(n_1263),
.B2(n_1258),
.Y(n_1438)
);

CKINVDCx8_ASAP7_75t_R g1439 ( 
.A(n_1295),
.Y(n_1439)
);

BUFx6f_ASAP7_75t_L g1440 ( 
.A(n_1268),
.Y(n_1440)
);

AOI22xp33_ASAP7_75t_L g1441 ( 
.A1(n_1236),
.A2(n_1312),
.B1(n_1303),
.B2(n_1355),
.Y(n_1441)
);

OAI22xp33_ASAP7_75t_SL g1442 ( 
.A1(n_1290),
.A2(n_1313),
.B1(n_1361),
.B2(n_1345),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1306),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_SL g1444 ( 
.A1(n_1290),
.A2(n_1313),
.B1(n_1361),
.B2(n_1345),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1307),
.A2(n_1354),
.B1(n_1348),
.B2(n_1329),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1306),
.Y(n_1446)
);

INVx8_ASAP7_75t_L g1447 ( 
.A(n_1223),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1290),
.B(n_1313),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1306),
.Y(n_1449)
);

AOI22xp33_ASAP7_75t_SL g1450 ( 
.A1(n_1320),
.A2(n_1362),
.B1(n_1337),
.B2(n_1361),
.Y(n_1450)
);

AOI22xp33_ASAP7_75t_L g1451 ( 
.A1(n_1320),
.A2(n_1362),
.B1(n_1345),
.B2(n_1337),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1225),
.Y(n_1452)
);

CKINVDCx11_ASAP7_75t_R g1453 ( 
.A(n_1233),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1233),
.A2(n_1213),
.B1(n_1249),
.B2(n_1270),
.Y(n_1454)
);

AOI21xp5_ASAP7_75t_L g1455 ( 
.A1(n_1249),
.A2(n_1213),
.B(n_1270),
.Y(n_1455)
);

CKINVDCx11_ASAP7_75t_R g1456 ( 
.A(n_1213),
.Y(n_1456)
);

CKINVDCx20_ASAP7_75t_R g1457 ( 
.A(n_1249),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_L g1458 ( 
.A1(n_1270),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1458)
);

CKINVDCx6p67_ASAP7_75t_R g1459 ( 
.A(n_1310),
.Y(n_1459)
);

INVxp67_ASAP7_75t_L g1460 ( 
.A(n_1210),
.Y(n_1460)
);

AND2x2_ASAP7_75t_L g1461 ( 
.A(n_1308),
.B(n_1325),
.Y(n_1461)
);

AOI22xp33_ASAP7_75t_L g1462 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1462)
);

BUFx6f_ASAP7_75t_L g1463 ( 
.A(n_1214),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_1230),
.Y(n_1464)
);

AOI22xp33_ASAP7_75t_L g1465 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1465)
);

BUFx6f_ASAP7_75t_L g1466 ( 
.A(n_1214),
.Y(n_1466)
);

BUFx10_ASAP7_75t_L g1467 ( 
.A(n_1265),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_L g1468 ( 
.A(n_1324),
.B(n_1327),
.Y(n_1468)
);

CKINVDCx11_ASAP7_75t_R g1469 ( 
.A(n_1230),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1230),
.Y(n_1470)
);

CKINVDCx6p67_ASAP7_75t_R g1471 ( 
.A(n_1310),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_1336),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1206),
.Y(n_1474)
);

AOI22xp33_ASAP7_75t_L g1475 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1477)
);

INVx4_ASAP7_75t_L g1478 ( 
.A(n_1214),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1335),
.B(n_1339),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1302),
.A2(n_935),
.B1(n_1053),
.B2(n_968),
.Y(n_1480)
);

AOI22xp33_ASAP7_75t_L g1481 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1481)
);

BUFx3_ASAP7_75t_L g1482 ( 
.A(n_1218),
.Y(n_1482)
);

INVx1_ASAP7_75t_SL g1483 ( 
.A(n_1336),
.Y(n_1483)
);

CKINVDCx11_ASAP7_75t_R g1484 ( 
.A(n_1230),
.Y(n_1484)
);

NAND2xp5_ASAP7_75t_L g1485 ( 
.A(n_1324),
.B(n_1327),
.Y(n_1485)
);

CKINVDCx11_ASAP7_75t_R g1486 ( 
.A(n_1230),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_SL g1487 ( 
.A1(n_1339),
.A2(n_547),
.B1(n_935),
.B2(n_755),
.Y(n_1487)
);

AND2x4_ASAP7_75t_L g1488 ( 
.A(n_1294),
.B(n_1144),
.Y(n_1488)
);

AOI22xp33_ASAP7_75t_SL g1489 ( 
.A1(n_1339),
.A2(n_547),
.B1(n_935),
.B2(n_755),
.Y(n_1489)
);

AOI22xp33_ASAP7_75t_L g1490 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1490)
);

INVx6_ASAP7_75t_L g1491 ( 
.A(n_1214),
.Y(n_1491)
);

INVx4_ASAP7_75t_L g1492 ( 
.A(n_1214),
.Y(n_1492)
);

AOI22xp33_ASAP7_75t_SL g1493 ( 
.A1(n_1339),
.A2(n_547),
.B1(n_935),
.B2(n_755),
.Y(n_1493)
);

CKINVDCx20_ASAP7_75t_R g1494 ( 
.A(n_1310),
.Y(n_1494)
);

BUFx10_ASAP7_75t_L g1495 ( 
.A(n_1265),
.Y(n_1495)
);

AOI22xp33_ASAP7_75t_L g1496 ( 
.A1(n_1302),
.A2(n_869),
.B1(n_968),
.B2(n_1053),
.Y(n_1496)
);

AO21x2_ASAP7_75t_L g1497 ( 
.A1(n_1410),
.A2(n_1418),
.B(n_1427),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1443),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1446),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1449),
.Y(n_1500)
);

AOI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1479),
.A2(n_1426),
.B(n_1455),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1487),
.A2(n_1493),
.B1(n_1489),
.B2(n_1479),
.Y(n_1502)
);

AND2x2_ASAP7_75t_L g1503 ( 
.A(n_1431),
.B(n_1432),
.Y(n_1503)
);

AND2x4_ASAP7_75t_SL g1504 ( 
.A(n_1387),
.B(n_1440),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1369),
.A2(n_1376),
.B1(n_1374),
.B2(n_1367),
.Y(n_1505)
);

NAND2xp33_ASAP7_75t_L g1506 ( 
.A(n_1371),
.B(n_1464),
.Y(n_1506)
);

OAI21x1_ASAP7_75t_L g1507 ( 
.A1(n_1445),
.A2(n_1441),
.B(n_1423),
.Y(n_1507)
);

BUFx2_ASAP7_75t_L g1508 ( 
.A(n_1437),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1403),
.Y(n_1509)
);

CKINVDCx20_ASAP7_75t_R g1510 ( 
.A(n_1368),
.Y(n_1510)
);

BUFx3_ASAP7_75t_L g1511 ( 
.A(n_1434),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1403),
.Y(n_1512)
);

HB1xp67_ASAP7_75t_L g1513 ( 
.A(n_1460),
.Y(n_1513)
);

AO21x1_ASAP7_75t_SL g1514 ( 
.A1(n_1372),
.A2(n_1415),
.B(n_1385),
.Y(n_1514)
);

INVx1_ASAP7_75t_L g1515 ( 
.A(n_1365),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1418),
.A2(n_1454),
.B(n_1448),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1440),
.Y(n_1517)
);

CKINVDCx5p33_ASAP7_75t_R g1518 ( 
.A(n_1370),
.Y(n_1518)
);

INVx3_ASAP7_75t_L g1519 ( 
.A(n_1439),
.Y(n_1519)
);

INVx2_ASAP7_75t_L g1520 ( 
.A(n_1447),
.Y(n_1520)
);

OA21x2_ASAP7_75t_L g1521 ( 
.A1(n_1425),
.A2(n_1438),
.B(n_1417),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1447),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1383),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1447),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1474),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1452),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1444),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1456),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1457),
.Y(n_1529)
);

INVx2_ASAP7_75t_L g1530 ( 
.A(n_1453),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1366),
.B(n_1468),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1442),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1458),
.B(n_1372),
.Y(n_1533)
);

OAI21x1_ASAP7_75t_L g1534 ( 
.A1(n_1425),
.A2(n_1430),
.B(n_1451),
.Y(n_1534)
);

AND2x2_ASAP7_75t_L g1535 ( 
.A(n_1458),
.B(n_1421),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1450),
.Y(n_1536)
);

BUFx2_ASAP7_75t_L g1537 ( 
.A(n_1384),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1424),
.B(n_1451),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1408),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1485),
.B(n_1385),
.Y(n_1540)
);

OAI21xp5_ASAP7_75t_L g1541 ( 
.A1(n_1369),
.A2(n_1496),
.B(n_1477),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1408),
.Y(n_1542)
);

INVx1_ASAP7_75t_L g1543 ( 
.A(n_1436),
.Y(n_1543)
);

OAI21x1_ASAP7_75t_L g1544 ( 
.A1(n_1430),
.A2(n_1391),
.B(n_1390),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1397),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1435),
.Y(n_1546)
);

INVx1_ASAP7_75t_SL g1547 ( 
.A(n_1402),
.Y(n_1547)
);

BUFx2_ASAP7_75t_L g1548 ( 
.A(n_1395),
.Y(n_1548)
);

BUFx2_ASAP7_75t_L g1549 ( 
.A(n_1409),
.Y(n_1549)
);

BUFx6f_ASAP7_75t_L g1550 ( 
.A(n_1463),
.Y(n_1550)
);

AOI31xp33_ASAP7_75t_L g1551 ( 
.A1(n_1480),
.A2(n_1378),
.A3(n_1490),
.B(n_1462),
.Y(n_1551)
);

AND2x4_ASAP7_75t_L g1552 ( 
.A(n_1390),
.B(n_1391),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1462),
.A2(n_1496),
.B(n_1465),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1461),
.B(n_1387),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1388),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1419),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1396),
.Y(n_1557)
);

BUFx6f_ASAP7_75t_L g1558 ( 
.A(n_1463),
.Y(n_1558)
);

OAI21x1_ASAP7_75t_L g1559 ( 
.A1(n_1411),
.A2(n_1476),
.B(n_1490),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1401),
.B(n_1476),
.Y(n_1560)
);

CKINVDCx5p33_ASAP7_75t_R g1561 ( 
.A(n_1469),
.Y(n_1561)
);

NOR2x1_ASAP7_75t_L g1562 ( 
.A(n_1478),
.B(n_1492),
.Y(n_1562)
);

BUFx2_ASAP7_75t_L g1563 ( 
.A(n_1399),
.Y(n_1563)
);

OAI21x1_ASAP7_75t_L g1564 ( 
.A1(n_1465),
.A2(n_1473),
.B(n_1477),
.Y(n_1564)
);

BUFx3_ASAP7_75t_L g1565 ( 
.A(n_1406),
.Y(n_1565)
);

OAI21x1_ASAP7_75t_L g1566 ( 
.A1(n_1473),
.A2(n_1481),
.B(n_1475),
.Y(n_1566)
);

OR2x2_ASAP7_75t_L g1567 ( 
.A(n_1374),
.B(n_1475),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1413),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1398),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1400),
.Y(n_1570)
);

INVx2_ASAP7_75t_SL g1571 ( 
.A(n_1380),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1481),
.B(n_1399),
.Y(n_1572)
);

AO21x2_ASAP7_75t_L g1573 ( 
.A1(n_1488),
.A2(n_1386),
.B(n_1422),
.Y(n_1573)
);

BUFx3_ASAP7_75t_L g1574 ( 
.A(n_1470),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1472),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1488),
.B(n_1389),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1483),
.Y(n_1577)
);

NAND3xp33_ASAP7_75t_L g1578 ( 
.A(n_1389),
.B(n_1484),
.C(n_1486),
.Y(n_1578)
);

NAND2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1428),
.B(n_1466),
.Y(n_1579)
);

OA21x2_ASAP7_75t_L g1580 ( 
.A1(n_1412),
.A2(n_1405),
.B(n_1491),
.Y(n_1580)
);

OAI21x1_ASAP7_75t_L g1581 ( 
.A1(n_1429),
.A2(n_1375),
.B(n_1392),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1529),
.B(n_1495),
.Y(n_1582)
);

AND2x4_ASAP7_75t_L g1583 ( 
.A(n_1581),
.B(n_1482),
.Y(n_1583)
);

NOR2xp33_ASAP7_75t_L g1584 ( 
.A(n_1531),
.B(n_1381),
.Y(n_1584)
);

AOI221x1_ASAP7_75t_SL g1585 ( 
.A1(n_1531),
.A2(n_1495),
.B1(n_1467),
.B2(n_1382),
.C(n_1375),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1505),
.A2(n_1379),
.B1(n_1377),
.B2(n_1459),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1529),
.B(n_1467),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1545),
.Y(n_1588)
);

OR2x6_ASAP7_75t_L g1589 ( 
.A(n_1544),
.B(n_1580),
.Y(n_1589)
);

AND2x2_ASAP7_75t_L g1590 ( 
.A(n_1528),
.B(n_1416),
.Y(n_1590)
);

NOR2xp33_ASAP7_75t_L g1591 ( 
.A(n_1551),
.B(n_1433),
.Y(n_1591)
);

O2A1O1Ixp33_ASAP7_75t_L g1592 ( 
.A1(n_1551),
.A2(n_1433),
.B(n_1482),
.C(n_1407),
.Y(n_1592)
);

OA21x2_ASAP7_75t_L g1593 ( 
.A1(n_1534),
.A2(n_1491),
.B(n_1420),
.Y(n_1593)
);

AOI21xp5_ASAP7_75t_L g1594 ( 
.A1(n_1497),
.A2(n_1521),
.B(n_1544),
.Y(n_1594)
);

OR2x2_ASAP7_75t_L g1595 ( 
.A(n_1528),
.B(n_1471),
.Y(n_1595)
);

OA21x2_ASAP7_75t_L g1596 ( 
.A1(n_1534),
.A2(n_1491),
.B(n_1420),
.Y(n_1596)
);

AND2x4_ASAP7_75t_SL g1597 ( 
.A(n_1510),
.B(n_1494),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_SL g1598 ( 
.A1(n_1552),
.A2(n_1393),
.B(n_1404),
.Y(n_1598)
);

O2A1O1Ixp33_ASAP7_75t_SL g1599 ( 
.A1(n_1541),
.A2(n_1394),
.B(n_1414),
.C(n_1420),
.Y(n_1599)
);

BUFx2_ASAP7_75t_SL g1600 ( 
.A(n_1511),
.Y(n_1600)
);

AOI21xp5_ASAP7_75t_L g1601 ( 
.A1(n_1497),
.A2(n_1404),
.B(n_1416),
.Y(n_1601)
);

NOR2xp33_ASAP7_75t_L g1602 ( 
.A(n_1506),
.B(n_1373),
.Y(n_1602)
);

INVxp67_ASAP7_75t_L g1603 ( 
.A(n_1545),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1554),
.B(n_1394),
.Y(n_1604)
);

OR2x2_ASAP7_75t_L g1605 ( 
.A(n_1537),
.B(n_1525),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1530),
.B(n_1572),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1530),
.B(n_1572),
.Y(n_1607)
);

NOR2xp33_ASAP7_75t_L g1608 ( 
.A(n_1540),
.B(n_1549),
.Y(n_1608)
);

AOI21xp33_ASAP7_75t_L g1609 ( 
.A1(n_1541),
.A2(n_1553),
.B(n_1555),
.Y(n_1609)
);

OAI21x1_ASAP7_75t_SL g1610 ( 
.A1(n_1553),
.A2(n_1540),
.B(n_1524),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1511),
.B(n_1577),
.Y(n_1611)
);

OAI22xp5_ASAP7_75t_L g1612 ( 
.A1(n_1502),
.A2(n_1567),
.B1(n_1552),
.B2(n_1570),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1515),
.Y(n_1613)
);

AO32x1_ASAP7_75t_L g1614 ( 
.A1(n_1560),
.A2(n_1535),
.A3(n_1524),
.B1(n_1546),
.B2(n_1527),
.Y(n_1614)
);

AND2x4_ASAP7_75t_L g1615 ( 
.A(n_1581),
.B(n_1569),
.Y(n_1615)
);

HB1xp67_ASAP7_75t_L g1616 ( 
.A(n_1508),
.Y(n_1616)
);

OAI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1564),
.A2(n_1566),
.B(n_1544),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1515),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1581),
.B(n_1569),
.Y(n_1619)
);

NOR2x1_ASAP7_75t_SL g1620 ( 
.A(n_1573),
.B(n_1497),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1523),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1526),
.B(n_1576),
.Y(n_1622)
);

NAND2xp5_ASAP7_75t_L g1623 ( 
.A(n_1539),
.B(n_1542),
.Y(n_1623)
);

OAI21xp5_ASAP7_75t_L g1624 ( 
.A1(n_1564),
.A2(n_1566),
.B(n_1549),
.Y(n_1624)
);

NOR2x1_ASAP7_75t_SL g1625 ( 
.A(n_1573),
.B(n_1497),
.Y(n_1625)
);

AO32x2_ASAP7_75t_L g1626 ( 
.A1(n_1571),
.A2(n_1532),
.A3(n_1503),
.B1(n_1508),
.B2(n_1536),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1539),
.B(n_1542),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1548),
.B(n_1563),
.Y(n_1628)
);

OAI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1564),
.A2(n_1566),
.B(n_1559),
.Y(n_1629)
);

OAI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1559),
.A2(n_1552),
.B(n_1567),
.Y(n_1630)
);

OAI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1559),
.A2(n_1552),
.B(n_1533),
.Y(n_1631)
);

INVx8_ASAP7_75t_L g1632 ( 
.A(n_1550),
.Y(n_1632)
);

AOI211xp5_ASAP7_75t_L g1633 ( 
.A1(n_1543),
.A2(n_1548),
.B(n_1533),
.C(n_1570),
.Y(n_1633)
);

NOR2xp33_ASAP7_75t_L g1634 ( 
.A(n_1511),
.B(n_1577),
.Y(n_1634)
);

OA21x2_ASAP7_75t_L g1635 ( 
.A1(n_1507),
.A2(n_1543),
.B(n_1501),
.Y(n_1635)
);

AOI22xp5_ASAP7_75t_L g1636 ( 
.A1(n_1520),
.A2(n_1522),
.B1(n_1568),
.B2(n_1519),
.Y(n_1636)
);

NAND2xp5_ASAP7_75t_L g1637 ( 
.A(n_1509),
.B(n_1512),
.Y(n_1637)
);

O2A1O1Ixp33_ASAP7_75t_L g1638 ( 
.A1(n_1513),
.A2(n_1575),
.B(n_1557),
.C(n_1547),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1521),
.A2(n_1516),
.B(n_1504),
.Y(n_1639)
);

NOR2x1_ASAP7_75t_SL g1640 ( 
.A(n_1573),
.B(n_1514),
.Y(n_1640)
);

NOR2x1_ASAP7_75t_R g1641 ( 
.A(n_1518),
.B(n_1561),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1509),
.B(n_1512),
.Y(n_1642)
);

NOR2xp33_ASAP7_75t_L g1643 ( 
.A(n_1547),
.B(n_1578),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1617),
.B(n_1516),
.Y(n_1644)
);

HB1xp67_ASAP7_75t_L g1645 ( 
.A(n_1588),
.Y(n_1645)
);

AOI22xp33_ASAP7_75t_L g1646 ( 
.A1(n_1609),
.A2(n_1514),
.B1(n_1536),
.B2(n_1538),
.Y(n_1646)
);

OR2x2_ASAP7_75t_L g1647 ( 
.A(n_1589),
.B(n_1516),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1617),
.B(n_1516),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1629),
.B(n_1521),
.Y(n_1649)
);

INVx1_ASAP7_75t_L g1650 ( 
.A(n_1613),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1589),
.B(n_1603),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1618),
.Y(n_1652)
);

BUFx3_ASAP7_75t_L g1653 ( 
.A(n_1615),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1609),
.A2(n_1538),
.B1(n_1568),
.B2(n_1578),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1619),
.Y(n_1655)
);

BUFx2_ASAP7_75t_L g1656 ( 
.A(n_1626),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1621),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1616),
.Y(n_1658)
);

AOI22xp33_ASAP7_75t_SL g1659 ( 
.A1(n_1612),
.A2(n_1519),
.B1(n_1504),
.B2(n_1580),
.Y(n_1659)
);

BUFx3_ASAP7_75t_L g1660 ( 
.A(n_1593),
.Y(n_1660)
);

INVx3_ASAP7_75t_L g1661 ( 
.A(n_1593),
.Y(n_1661)
);

INVxp67_ASAP7_75t_L g1662 ( 
.A(n_1606),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_L g1663 ( 
.A(n_1638),
.B(n_1580),
.Y(n_1663)
);

AND2x2_ASAP7_75t_L g1664 ( 
.A(n_1631),
.B(n_1503),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1626),
.Y(n_1665)
);

AND2x2_ASAP7_75t_L g1666 ( 
.A(n_1631),
.B(n_1500),
.Y(n_1666)
);

AND2x4_ASAP7_75t_L g1667 ( 
.A(n_1640),
.B(n_1517),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1605),
.Y(n_1668)
);

AND2x2_ASAP7_75t_L g1669 ( 
.A(n_1626),
.B(n_1498),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1612),
.A2(n_1520),
.B1(n_1522),
.B2(n_1519),
.Y(n_1670)
);

INVxp67_ASAP7_75t_SL g1671 ( 
.A(n_1620),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1626),
.B(n_1498),
.Y(n_1672)
);

NAND2xp5_ASAP7_75t_L g1673 ( 
.A(n_1623),
.B(n_1627),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1596),
.B(n_1499),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1596),
.Y(n_1675)
);

AOI221xp5_ASAP7_75t_L g1676 ( 
.A1(n_1654),
.A2(n_1608),
.B1(n_1592),
.B2(n_1586),
.C(n_1633),
.Y(n_1676)
);

INVx1_ASAP7_75t_L g1677 ( 
.A(n_1650),
.Y(n_1677)
);

INVx2_ASAP7_75t_L g1678 ( 
.A(n_1674),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1650),
.Y(n_1679)
);

HB1xp67_ASAP7_75t_L g1680 ( 
.A(n_1658),
.Y(n_1680)
);

OAI31xp33_ASAP7_75t_L g1681 ( 
.A1(n_1654),
.A2(n_1586),
.A3(n_1592),
.B(n_1591),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1650),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_SL g1683 ( 
.A1(n_1644),
.A2(n_1591),
.B1(n_1624),
.B2(n_1630),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1664),
.B(n_1607),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1652),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1653),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1673),
.B(n_1630),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1673),
.B(n_1624),
.Y(n_1688)
);

AND2x2_ASAP7_75t_L g1689 ( 
.A(n_1664),
.B(n_1625),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1652),
.Y(n_1690)
);

INVx4_ASAP7_75t_L g1691 ( 
.A(n_1667),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1645),
.B(n_1668),
.Y(n_1692)
);

AOI22xp5_ASAP7_75t_L g1693 ( 
.A1(n_1646),
.A2(n_1643),
.B1(n_1584),
.B2(n_1634),
.Y(n_1693)
);

AOI221xp5_ASAP7_75t_L g1694 ( 
.A1(n_1646),
.A2(n_1638),
.B1(n_1585),
.B2(n_1594),
.C(n_1610),
.Y(n_1694)
);

AND2x2_ASAP7_75t_L g1695 ( 
.A(n_1664),
.B(n_1639),
.Y(n_1695)
);

NAND4xp25_ASAP7_75t_SL g1696 ( 
.A(n_1663),
.B(n_1598),
.C(n_1639),
.D(n_1636),
.Y(n_1696)
);

OAI221xp5_ASAP7_75t_SL g1697 ( 
.A1(n_1670),
.A2(n_1594),
.B1(n_1595),
.B2(n_1611),
.C(n_1614),
.Y(n_1697)
);

AOI211xp5_ASAP7_75t_L g1698 ( 
.A1(n_1644),
.A2(n_1599),
.B(n_1602),
.C(n_1582),
.Y(n_1698)
);

HB1xp67_ASAP7_75t_L g1699 ( 
.A(n_1645),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1651),
.B(n_1635),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1675),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1662),
.B(n_1628),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1657),
.Y(n_1703)
);

INVx2_ASAP7_75t_L g1704 ( 
.A(n_1675),
.Y(n_1704)
);

AOI221xp5_ASAP7_75t_L g1705 ( 
.A1(n_1644),
.A2(n_1642),
.B1(n_1637),
.B2(n_1587),
.C(n_1556),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1666),
.B(n_1642),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1657),
.Y(n_1707)
);

AND2x4_ASAP7_75t_SL g1708 ( 
.A(n_1667),
.B(n_1583),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1655),
.B(n_1622),
.Y(n_1709)
);

NAND2x1_ASAP7_75t_SL g1710 ( 
.A(n_1695),
.B(n_1663),
.Y(n_1710)
);

NAND2xp33_ASAP7_75t_R g1711 ( 
.A(n_1686),
.B(n_1580),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1695),
.B(n_1656),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1677),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1688),
.B(n_1669),
.Y(n_1714)
);

INVxp33_ASAP7_75t_L g1715 ( 
.A(n_1693),
.Y(n_1715)
);

NAND3xp33_ASAP7_75t_SL g1716 ( 
.A(n_1681),
.B(n_1659),
.C(n_1670),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1680),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1689),
.B(n_1656),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1689),
.B(n_1691),
.Y(n_1719)
);

AND2x4_ASAP7_75t_L g1720 ( 
.A(n_1691),
.B(n_1660),
.Y(n_1720)
);

INVx3_ASAP7_75t_SL g1721 ( 
.A(n_1708),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1701),
.Y(n_1722)
);

AND2x4_ASAP7_75t_L g1723 ( 
.A(n_1691),
.B(n_1660),
.Y(n_1723)
);

OR2x2_ASAP7_75t_L g1724 ( 
.A(n_1678),
.B(n_1656),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1677),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1691),
.B(n_1665),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1679),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1679),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1678),
.B(n_1665),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1682),
.Y(n_1730)
);

INVx2_ASAP7_75t_L g1731 ( 
.A(n_1701),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1688),
.B(n_1669),
.Y(n_1732)
);

BUFx2_ASAP7_75t_L g1733 ( 
.A(n_1699),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1678),
.B(n_1665),
.Y(n_1734)
);

AND2x4_ASAP7_75t_L g1735 ( 
.A(n_1708),
.B(n_1660),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1682),
.Y(n_1736)
);

NAND2xp5_ASAP7_75t_L g1737 ( 
.A(n_1687),
.B(n_1669),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1687),
.B(n_1672),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1685),
.Y(n_1739)
);

INVx1_ASAP7_75t_L g1740 ( 
.A(n_1690),
.Y(n_1740)
);

INVx4_ASAP7_75t_L g1741 ( 
.A(n_1686),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1690),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1708),
.B(n_1660),
.Y(n_1743)
);

INVx2_ASAP7_75t_L g1744 ( 
.A(n_1701),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1704),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1704),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1721),
.B(n_1684),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1715),
.B(n_1694),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1733),
.B(n_1694),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1713),
.Y(n_1750)
);

AND2x4_ASAP7_75t_SL g1751 ( 
.A(n_1735),
.B(n_1583),
.Y(n_1751)
);

INVxp33_ASAP7_75t_L g1752 ( 
.A(n_1716),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1721),
.B(n_1684),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1713),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1716),
.B(n_1641),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1725),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1725),
.Y(n_1757)
);

NOR2xp67_ASAP7_75t_L g1758 ( 
.A(n_1741),
.B(n_1696),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1727),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1733),
.B(n_1705),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1727),
.Y(n_1761)
);

AND2x2_ASAP7_75t_L g1762 ( 
.A(n_1721),
.B(n_1735),
.Y(n_1762)
);

NAND2xp5_ASAP7_75t_L g1763 ( 
.A(n_1710),
.B(n_1705),
.Y(n_1763)
);

AND3x1_ASAP7_75t_L g1764 ( 
.A(n_1726),
.B(n_1698),
.C(n_1681),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1717),
.Y(n_1765)
);

AND2x2_ASAP7_75t_L g1766 ( 
.A(n_1735),
.B(n_1743),
.Y(n_1766)
);

INVxp67_ASAP7_75t_L g1767 ( 
.A(n_1717),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1735),
.B(n_1686),
.Y(n_1768)
);

NAND2xp67_ASAP7_75t_L g1769 ( 
.A(n_1719),
.B(n_1597),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1728),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1710),
.B(n_1706),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1728),
.Y(n_1772)
);

NAND2xp33_ASAP7_75t_L g1773 ( 
.A(n_1712),
.B(n_1676),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1724),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1735),
.B(n_1686),
.Y(n_1775)
);

OR2x6_ASAP7_75t_L g1776 ( 
.A(n_1741),
.B(n_1600),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1743),
.B(n_1683),
.Y(n_1777)
);

OAI21xp33_ASAP7_75t_L g1778 ( 
.A1(n_1737),
.A2(n_1683),
.B(n_1696),
.Y(n_1778)
);

INVx1_ASAP7_75t_L g1779 ( 
.A(n_1730),
.Y(n_1779)
);

INVx2_ASAP7_75t_SL g1780 ( 
.A(n_1743),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1730),
.Y(n_1781)
);

OR2x6_ASAP7_75t_L g1782 ( 
.A(n_1741),
.B(n_1601),
.Y(n_1782)
);

O2A1O1Ixp5_ASAP7_75t_SL g1783 ( 
.A1(n_1736),
.A2(n_1661),
.B(n_1707),
.C(n_1703),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1743),
.Y(n_1784)
);

NAND2xp5_ASAP7_75t_L g1785 ( 
.A(n_1737),
.B(n_1706),
.Y(n_1785)
);

INVx1_ASAP7_75t_L g1786 ( 
.A(n_1736),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1739),
.Y(n_1787)
);

AND2x2_ASAP7_75t_L g1788 ( 
.A(n_1743),
.B(n_1709),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1724),
.Y(n_1789)
);

NAND2xp5_ASAP7_75t_L g1790 ( 
.A(n_1748),
.B(n_1693),
.Y(n_1790)
);

AND3x2_ASAP7_75t_L g1791 ( 
.A(n_1755),
.B(n_1698),
.C(n_1676),
.Y(n_1791)
);

NAND2x1p5_ASAP7_75t_L g1792 ( 
.A(n_1764),
.B(n_1580),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1752),
.B(n_1712),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1749),
.B(n_1712),
.Y(n_1794)
);

INVx2_ASAP7_75t_L g1795 ( 
.A(n_1774),
.Y(n_1795)
);

INVx1_ASAP7_75t_L g1796 ( 
.A(n_1770),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1762),
.B(n_1719),
.Y(n_1797)
);

INVxp67_ASAP7_75t_SL g1798 ( 
.A(n_1758),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1765),
.B(n_1738),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_L g1800 ( 
.A(n_1773),
.B(n_1738),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1762),
.B(n_1719),
.Y(n_1801)
);

OR2x2_ASAP7_75t_L g1802 ( 
.A(n_1767),
.B(n_1714),
.Y(n_1802)
);

AND2x4_ASAP7_75t_L g1803 ( 
.A(n_1766),
.B(n_1726),
.Y(n_1803)
);

NAND2xp5_ASAP7_75t_L g1804 ( 
.A(n_1773),
.B(n_1714),
.Y(n_1804)
);

INVx1_ASAP7_75t_SL g1805 ( 
.A(n_1777),
.Y(n_1805)
);

OAI32xp33_ASAP7_75t_L g1806 ( 
.A1(n_1763),
.A2(n_1711),
.A3(n_1647),
.B1(n_1732),
.B2(n_1724),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1778),
.B(n_1732),
.Y(n_1807)
);

INVxp33_ASAP7_75t_L g1808 ( 
.A(n_1777),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1750),
.Y(n_1809)
);

AND2x2_ASAP7_75t_L g1810 ( 
.A(n_1747),
.B(n_1753),
.Y(n_1810)
);

AOI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1760),
.A2(n_1697),
.B(n_1648),
.C(n_1647),
.Y(n_1811)
);

NAND2x1_ASAP7_75t_L g1812 ( 
.A(n_1776),
.B(n_1741),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1747),
.B(n_1718),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1771),
.B(n_1702),
.Y(n_1814)
);

AND2x2_ASAP7_75t_L g1815 ( 
.A(n_1753),
.B(n_1766),
.Y(n_1815)
);

OAI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1783),
.A2(n_1697),
.B(n_1648),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1774),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1750),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1756),
.Y(n_1819)
);

INVx1_ASAP7_75t_SL g1820 ( 
.A(n_1751),
.Y(n_1820)
);

AND2x4_ASAP7_75t_L g1821 ( 
.A(n_1780),
.B(n_1726),
.Y(n_1821)
);

INVxp67_ASAP7_75t_L g1822 ( 
.A(n_1780),
.Y(n_1822)
);

INVx2_ASAP7_75t_SL g1823 ( 
.A(n_1784),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1788),
.B(n_1718),
.Y(n_1824)
);

OR2x2_ASAP7_75t_L g1825 ( 
.A(n_1789),
.B(n_1692),
.Y(n_1825)
);

INVx2_ASAP7_75t_L g1826 ( 
.A(n_1803),
.Y(n_1826)
);

AOI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1791),
.A2(n_1648),
.B1(n_1784),
.B2(n_1788),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1809),
.Y(n_1828)
);

INVxp67_ASAP7_75t_L g1829 ( 
.A(n_1798),
.Y(n_1829)
);

NAND2x1p5_ASAP7_75t_L g1830 ( 
.A(n_1812),
.B(n_1741),
.Y(n_1830)
);

AO21x1_ASAP7_75t_L g1831 ( 
.A1(n_1792),
.A2(n_1757),
.B(n_1756),
.Y(n_1831)
);

AOI22xp5_ASAP7_75t_L g1832 ( 
.A1(n_1811),
.A2(n_1776),
.B1(n_1751),
.B2(n_1775),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1823),
.B(n_1768),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1809),
.Y(n_1834)
);

OAI221xp5_ASAP7_75t_L g1835 ( 
.A1(n_1816),
.A2(n_1776),
.B1(n_1782),
.B2(n_1789),
.C(n_1659),
.Y(n_1835)
);

AND2x2_ASAP7_75t_L g1836 ( 
.A(n_1815),
.B(n_1768),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1805),
.B(n_1790),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1807),
.B(n_1754),
.Y(n_1838)
);

OAI32xp33_ASAP7_75t_L g1839 ( 
.A1(n_1792),
.A2(n_1804),
.A3(n_1800),
.B1(n_1793),
.B2(n_1808),
.Y(n_1839)
);

NOR2xp33_ASAP7_75t_L g1840 ( 
.A(n_1794),
.B(n_1769),
.Y(n_1840)
);

INVx2_ASAP7_75t_SL g1841 ( 
.A(n_1823),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1796),
.B(n_1786),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1818),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1803),
.Y(n_1844)
);

NAND3xp33_ASAP7_75t_L g1845 ( 
.A(n_1822),
.B(n_1783),
.C(n_1776),
.Y(n_1845)
);

AOI31xp33_ASAP7_75t_L g1846 ( 
.A1(n_1792),
.A2(n_1775),
.A3(n_1604),
.B(n_1579),
.Y(n_1846)
);

AOI21xp5_ASAP7_75t_L g1847 ( 
.A1(n_1806),
.A2(n_1782),
.B(n_1785),
.Y(n_1847)
);

OAI22x1_ASAP7_75t_L g1848 ( 
.A1(n_1820),
.A2(n_1720),
.B1(n_1723),
.B2(n_1787),
.Y(n_1848)
);

INVx1_ASAP7_75t_L g1849 ( 
.A(n_1818),
.Y(n_1849)
);

AOI21xp5_ASAP7_75t_L g1850 ( 
.A1(n_1806),
.A2(n_1782),
.B(n_1759),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1814),
.B(n_1769),
.Y(n_1851)
);

INVx1_ASAP7_75t_SL g1852 ( 
.A(n_1796),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1829),
.B(n_1837),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1828),
.Y(n_1854)
);

INVxp67_ASAP7_75t_L g1855 ( 
.A(n_1841),
.Y(n_1855)
);

AND2x2_ASAP7_75t_L g1856 ( 
.A(n_1836),
.B(n_1815),
.Y(n_1856)
);

NAND2x1p5_ASAP7_75t_L g1857 ( 
.A(n_1852),
.B(n_1812),
.Y(n_1857)
);

AND2x2_ASAP7_75t_L g1858 ( 
.A(n_1826),
.B(n_1810),
.Y(n_1858)
);

NAND2xp5_ASAP7_75t_L g1859 ( 
.A(n_1852),
.B(n_1810),
.Y(n_1859)
);

BUFx2_ASAP7_75t_L g1860 ( 
.A(n_1844),
.Y(n_1860)
);

NAND3xp33_ASAP7_75t_L g1861 ( 
.A(n_1835),
.B(n_1827),
.C(n_1845),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1833),
.Y(n_1862)
);

AOI22xp5_ASAP7_75t_L g1863 ( 
.A1(n_1831),
.A2(n_1801),
.B1(n_1797),
.B2(n_1803),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1834),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1832),
.A2(n_1803),
.B1(n_1824),
.B2(n_1813),
.Y(n_1865)
);

NAND2xp5_ASAP7_75t_L g1866 ( 
.A(n_1838),
.B(n_1813),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1839),
.A2(n_1799),
.B(n_1802),
.C(n_1801),
.Y(n_1867)
);

NOR4xp25_ASAP7_75t_SL g1868 ( 
.A(n_1843),
.B(n_1819),
.C(n_1757),
.D(n_1761),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1849),
.Y(n_1869)
);

AOI31xp33_ASAP7_75t_L g1870 ( 
.A1(n_1830),
.A2(n_1797),
.A3(n_1802),
.B(n_1799),
.Y(n_1870)
);

INVx1_ASAP7_75t_SL g1871 ( 
.A(n_1833),
.Y(n_1871)
);

INVxp67_ASAP7_75t_L g1872 ( 
.A(n_1840),
.Y(n_1872)
);

OAI21xp33_ASAP7_75t_L g1873 ( 
.A1(n_1851),
.A2(n_1824),
.B(n_1817),
.Y(n_1873)
);

A2O1A1Ixp33_ASAP7_75t_L g1874 ( 
.A1(n_1861),
.A2(n_1847),
.B(n_1850),
.C(n_1838),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1862),
.B(n_1842),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1870),
.A2(n_1846),
.B(n_1830),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1860),
.Y(n_1877)
);

AOI222xp33_ASAP7_75t_L g1878 ( 
.A1(n_1853),
.A2(n_1848),
.B1(n_1842),
.B2(n_1819),
.C1(n_1821),
.C2(n_1817),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1859),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1856),
.B(n_1821),
.Y(n_1880)
);

OAI21xp5_ASAP7_75t_L g1881 ( 
.A1(n_1863),
.A2(n_1846),
.B(n_1795),
.Y(n_1881)
);

O2A1O1Ixp33_ASAP7_75t_L g1882 ( 
.A1(n_1855),
.A2(n_1795),
.B(n_1782),
.C(n_1825),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1858),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1854),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1869),
.Y(n_1885)
);

INVx2_ASAP7_75t_L g1886 ( 
.A(n_1857),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1877),
.Y(n_1887)
);

NOR3xp33_ASAP7_75t_L g1888 ( 
.A(n_1874),
.B(n_1872),
.C(n_1855),
.Y(n_1888)
);

OAI21xp33_ASAP7_75t_L g1889 ( 
.A1(n_1874),
.A2(n_1873),
.B(n_1871),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1883),
.B(n_1866),
.Y(n_1890)
);

NAND2xp5_ASAP7_75t_SL g1891 ( 
.A(n_1876),
.B(n_1857),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1875),
.Y(n_1892)
);

INVxp67_ASAP7_75t_L g1893 ( 
.A(n_1886),
.Y(n_1893)
);

INVx1_ASAP7_75t_L g1894 ( 
.A(n_1886),
.Y(n_1894)
);

NAND4xp25_ASAP7_75t_L g1895 ( 
.A(n_1878),
.B(n_1865),
.C(n_1867),
.D(n_1864),
.Y(n_1895)
);

OAI21xp5_ASAP7_75t_SL g1896 ( 
.A1(n_1881),
.A2(n_1864),
.B(n_1821),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1880),
.Y(n_1897)
);

NOR2xp33_ASAP7_75t_L g1898 ( 
.A(n_1879),
.B(n_1825),
.Y(n_1898)
);

OAI21xp5_ASAP7_75t_SL g1899 ( 
.A1(n_1895),
.A2(n_1880),
.B(n_1882),
.Y(n_1899)
);

NOR3xp33_ASAP7_75t_L g1900 ( 
.A(n_1891),
.B(n_1889),
.C(n_1888),
.Y(n_1900)
);

A2O1A1Ixp33_ASAP7_75t_L g1901 ( 
.A1(n_1896),
.A2(n_1885),
.B(n_1884),
.C(n_1868),
.Y(n_1901)
);

AOI22xp5_ASAP7_75t_L g1902 ( 
.A1(n_1897),
.A2(n_1821),
.B1(n_1723),
.B2(n_1720),
.Y(n_1902)
);

INVxp67_ASAP7_75t_L g1903 ( 
.A(n_1898),
.Y(n_1903)
);

NOR2x1_ASAP7_75t_L g1904 ( 
.A(n_1894),
.B(n_1759),
.Y(n_1904)
);

AOI221xp5_ASAP7_75t_L g1905 ( 
.A1(n_1900),
.A2(n_1892),
.B1(n_1887),
.B2(n_1893),
.C(n_1890),
.Y(n_1905)
);

AOI22xp33_ASAP7_75t_L g1906 ( 
.A1(n_1903),
.A2(n_1893),
.B1(n_1649),
.B2(n_1720),
.Y(n_1906)
);

NAND3xp33_ASAP7_75t_SL g1907 ( 
.A(n_1901),
.B(n_1772),
.C(n_1761),
.Y(n_1907)
);

INVx1_ASAP7_75t_L g1908 ( 
.A(n_1904),
.Y(n_1908)
);

AOI221xp5_ASAP7_75t_L g1909 ( 
.A1(n_1899),
.A2(n_1781),
.B1(n_1779),
.B2(n_1772),
.C(n_1720),
.Y(n_1909)
);

NOR2xp33_ASAP7_75t_L g1910 ( 
.A(n_1902),
.B(n_1779),
.Y(n_1910)
);

OAI21xp33_ASAP7_75t_L g1911 ( 
.A1(n_1899),
.A2(n_1781),
.B(n_1723),
.Y(n_1911)
);

AND2x4_ASAP7_75t_L g1912 ( 
.A(n_1908),
.B(n_1720),
.Y(n_1912)
);

NOR4xp25_ASAP7_75t_L g1913 ( 
.A(n_1907),
.B(n_1746),
.C(n_1745),
.D(n_1722),
.Y(n_1913)
);

BUFx2_ASAP7_75t_L g1914 ( 
.A(n_1905),
.Y(n_1914)
);

OAI322xp33_ASAP7_75t_L g1915 ( 
.A1(n_1910),
.A2(n_1700),
.A3(n_1745),
.B1(n_1746),
.B2(n_1744),
.C1(n_1722),
.C2(n_1731),
.Y(n_1915)
);

NOR2x1p5_ASAP7_75t_L g1916 ( 
.A(n_1909),
.B(n_1574),
.Y(n_1916)
);

AOI22xp5_ASAP7_75t_L g1917 ( 
.A1(n_1911),
.A2(n_1723),
.B1(n_1574),
.B2(n_1718),
.Y(n_1917)
);

NAND3xp33_ASAP7_75t_SL g1918 ( 
.A(n_1914),
.B(n_1906),
.C(n_1579),
.Y(n_1918)
);

NOR2x1_ASAP7_75t_L g1919 ( 
.A(n_1912),
.B(n_1574),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1916),
.Y(n_1920)
);

XNOR2xp5_ASAP7_75t_L g1921 ( 
.A(n_1918),
.B(n_1913),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1921),
.Y(n_1922)
);

OAI22x1_ASAP7_75t_L g1923 ( 
.A1(n_1922),
.A2(n_1920),
.B1(n_1919),
.B2(n_1917),
.Y(n_1923)
);

NAND2xp5_ASAP7_75t_L g1924 ( 
.A(n_1922),
.B(n_1915),
.Y(n_1924)
);

OAI22x1_ASAP7_75t_L g1925 ( 
.A1(n_1924),
.A2(n_1723),
.B1(n_1745),
.B2(n_1744),
.Y(n_1925)
);

OAI22xp5_ASAP7_75t_SL g1926 ( 
.A1(n_1923),
.A2(n_1565),
.B1(n_1579),
.B2(n_1571),
.Y(n_1926)
);

OAI221xp5_ASAP7_75t_SL g1927 ( 
.A1(n_1926),
.A2(n_1565),
.B1(n_1671),
.B2(n_1744),
.C(n_1746),
.Y(n_1927)
);

AOI22xp5_ASAP7_75t_L g1928 ( 
.A1(n_1925),
.A2(n_1565),
.B1(n_1729),
.B2(n_1734),
.Y(n_1928)
);

AO221x1_ASAP7_75t_L g1929 ( 
.A1(n_1927),
.A2(n_1722),
.B1(n_1731),
.B2(n_1742),
.C(n_1740),
.Y(n_1929)
);

OR2x6_ASAP7_75t_L g1930 ( 
.A(n_1929),
.B(n_1928),
.Y(n_1930)
);

OAI21xp5_ASAP7_75t_SL g1931 ( 
.A1(n_1930),
.A2(n_1562),
.B(n_1590),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_R g1932 ( 
.A1(n_1931),
.A2(n_1632),
.B1(n_1731),
.B2(n_1729),
.C(n_1734),
.Y(n_1932)
);

AOI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1558),
.B(n_1550),
.C(n_1571),
.Y(n_1933)
);


endmodule