module real_jpeg_14279_n_8 (n_5, n_4, n_0, n_1, n_2, n_6, n_7, n_3, n_8);

input n_5;
input n_4;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_8;

wire n_17;
wire n_43;
wire n_37;
wire n_21;
wire n_33;
wire n_35;
wire n_38;
wire n_50;
wire n_29;
wire n_49;
wire n_10;
wire n_31;
wire n_9;
wire n_52;
wire n_12;
wire n_24;
wire n_34;
wire n_28;
wire n_44;
wire n_46;
wire n_23;
wire n_51;
wire n_11;
wire n_14;
wire n_47;
wire n_45;
wire n_25;
wire n_42;
wire n_22;
wire n_18;
wire n_53;
wire n_36;
wire n_39;
wire n_40;
wire n_41;
wire n_26;
wire n_32;
wire n_20;
wire n_19;
wire n_48;
wire n_27;
wire n_30;
wire n_16;
wire n_15;
wire n_13;

BUFx2_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx4f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_2),
.A2(n_12),
.B1(n_13),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g19 ( 
.A1(n_3),
.A2(n_17),
.B1(n_20),
.B2(n_22),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_3),
.B(n_13),
.C(n_29),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g40 ( 
.A1(n_3),
.A2(n_16),
.B1(n_37),
.B2(n_41),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_5),
.A2(n_12),
.B1(n_13),
.B2(n_21),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_5),
.A2(n_21),
.B1(n_37),
.B2(n_41),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_6),
.A2(n_12),
.B1(n_13),
.B2(n_26),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx11_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

XOR2xp5_ASAP7_75t_L g8 ( 
.A(n_9),
.B(n_33),
.Y(n_8)
);

OAI21xp5_ASAP7_75t_L g9 ( 
.A1(n_10),
.A2(n_23),
.B(n_32),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_L g10 ( 
.A(n_11),
.B(n_19),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_15),
.Y(n_11)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_12),
.A2(n_13),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_13),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_13),
.B(n_17),
.Y(n_22)
);

INVx4_ASAP7_75t_L g13 ( 
.A(n_14),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_16),
.B(n_17),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_16),
.B(n_28),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_17),
.A2(n_20),
.B1(n_22),
.B2(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_18),
.A2(n_47),
.B1(n_48),
.B2(n_49),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_22),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_27),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_27),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g48 ( 
.A(n_25),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_29),
.A2(n_30),
.B1(n_37),
.B2(n_41),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_SL g29 ( 
.A(n_30),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_52),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_46),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_46),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_39),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_38),
.Y(n_36)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_37),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_42),
.B1(n_44),
.B2(n_45),
.Y(n_39)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);


endmodule