module real_jpeg_13612_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_201;
wire n_114;
wire n_49;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_249;
wire n_83;
wire n_286;
wire n_166;
wire n_221;
wire n_176;
wire n_215;
wire n_288;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_271;
wire n_47;
wire n_281;
wire n_131;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_173;
wire n_40;
wire n_105;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_267;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_290;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_219;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_222;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_258;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_150;
wire n_32;
wire n_20;
wire n_74;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_216;
wire n_244;
wire n_167;
wire n_128;
wire n_179;
wire n_202;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_256;
wire n_101;
wire n_274;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_273;
wire n_89;

BUFx2_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_3),
.A2(n_25),
.B1(n_29),
.B2(n_39),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_3),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_3),
.A2(n_35),
.B1(n_36),
.B2(n_39),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g160 ( 
.A1(n_3),
.A2(n_39),
.B1(n_48),
.B2(n_50),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_3),
.A2(n_39),
.B1(n_61),
.B2(n_64),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_4),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_5),
.A2(n_35),
.B1(n_36),
.B2(n_54),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g140 ( 
.A1(n_5),
.A2(n_48),
.B1(n_50),
.B2(n_54),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_5),
.A2(n_54),
.B1(n_61),
.B2(n_64),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_5),
.A2(n_25),
.B1(n_29),
.B2(n_54),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_6),
.A2(n_48),
.B1(n_50),
.B2(n_69),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_6),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_6),
.A2(n_61),
.B1(n_64),
.B2(n_69),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_6),
.A2(n_35),
.B1(n_36),
.B2(n_69),
.Y(n_217)
);

OAI22xp33_ASAP7_75t_SL g267 ( 
.A1(n_6),
.A2(n_25),
.B1(n_29),
.B2(n_69),
.Y(n_267)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_8),
.A2(n_61),
.B1(n_64),
.B2(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_8),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_8),
.A2(n_48),
.B1(n_50),
.B2(n_76),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_8),
.A2(n_35),
.B1(n_36),
.B2(n_76),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_8),
.A2(n_25),
.B1(n_29),
.B2(n_76),
.Y(n_286)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_10),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_24)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

O2A1O1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_10),
.A2(n_29),
.B(n_32),
.C(n_80),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_10),
.B(n_37),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_10),
.A2(n_28),
.B1(n_48),
.B2(n_50),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_10),
.A2(n_85),
.B1(n_114),
.B2(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_10),
.B(n_52),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_11),
.A2(n_61),
.B1(n_64),
.B2(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_11),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_11),
.A2(n_48),
.B1(n_50),
.B2(n_78),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_11),
.A2(n_35),
.B1(n_36),
.B2(n_78),
.Y(n_257)
);

BUFx8_ASAP7_75t_L g32 ( 
.A(n_12),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_13),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_13),
.A2(n_25),
.B1(n_29),
.B2(n_43),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_13),
.A2(n_43),
.B1(n_48),
.B2(n_50),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g165 ( 
.A1(n_13),
.A2(n_43),
.B1(n_61),
.B2(n_64),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_14),
.A2(n_48),
.B1(n_50),
.B2(n_66),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_14),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_14),
.A2(n_35),
.B1(n_36),
.B2(n_66),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_14),
.A2(n_61),
.B1(n_64),
.B2(n_66),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_14),
.A2(n_25),
.B1(n_29),
.B2(n_66),
.Y(n_244)
);

INVx11_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_271),
.Y(n_16)
);

AOI21xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_249),
.B(n_270),
.Y(n_17)
);

OAI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_222),
.B(n_248),
.Y(n_18)
);

O2A1O1Ixp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_123),
.B(n_201),
.C(n_221),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_96),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_21),
.B(n_96),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_70),
.C(n_83),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_22),
.B(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_40),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_23),
.B(n_41),
.C(n_55),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_23)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

INVx13_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp33_ASAP7_75t_L g80 ( 
.A1(n_28),
.A2(n_33),
.B(n_35),
.Y(n_80)
);

HAxp5_ASAP7_75t_SL g133 ( 
.A(n_28),
.B(n_36),
.CON(n_133),
.SN(n_133)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_28),
.B(n_59),
.C(n_64),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g171 ( 
.A(n_28),
.B(n_85),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_28),
.B(n_60),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_30),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_30),
.A2(n_37),
.B1(n_105),
.B2(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_30),
.B(n_267),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_34),
.Y(n_30)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_32),
.Y(n_33)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_34),
.A2(n_102),
.B1(n_103),
.B2(n_104),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g285 ( 
.A1(n_34),
.A2(n_286),
.B(n_287),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_35),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_51)
);

NOR3xp33_ASAP7_75t_L g134 ( 
.A(n_35),
.B(n_47),
.C(n_48),
.Y(n_134)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_37),
.B(n_244),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_37),
.B(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_38),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g40 ( 
.A(n_41),
.B(n_55),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_44),
.B1(n_52),
.B2(n_53),
.Y(n_41)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_42),
.Y(n_95)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_44),
.A2(n_52),
.B1(n_93),
.B2(n_133),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_L g215 ( 
.A1(n_44),
.A2(n_109),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_44),
.B(n_240),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_44),
.A2(n_52),
.B1(n_256),
.B2(n_257),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_51),
.Y(n_44)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_45),
.A2(n_92),
.B1(n_94),
.B2(n_95),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_45),
.B(n_217),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_45),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

OA22x2_ASAP7_75t_SL g45 ( 
.A1(n_46),
.A2(n_47),
.B1(n_48),
.B2(n_50),
.Y(n_45)
);

O2A1O1Ixp33_ASAP7_75t_SL g131 ( 
.A1(n_46),
.A2(n_50),
.B(n_132),
.C(n_134),
.Y(n_131)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_48),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_48),
.A2(n_50),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_50),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_109),
.Y(n_108)
);

CKINVDCx14_ASAP7_75t_R g107 ( 
.A(n_53),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_65),
.B(n_67),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_121),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_56),
.A2(n_140),
.B1(n_142),
.B2(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_56),
.A2(n_142),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_56),
.A2(n_142),
.B1(n_150),
.B2(n_160),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_56),
.A2(n_142),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_56),
.A2(n_67),
.B(n_210),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_56),
.A2(n_65),
.B(n_142),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_60),
.Y(n_56)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_64),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_60),
.B(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_60),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_60),
.Y(n_142)
);

CKINVDCx6p67_ASAP7_75t_R g64 ( 
.A(n_61),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_73),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_64),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_65),
.B(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_68),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_70),
.B(n_83),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_71),
.A2(n_79),
.B1(n_81),
.B2(n_82),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_77),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g86 ( 
.A(n_72),
.B(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_72),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_72),
.A2(n_117),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_72),
.A2(n_73),
.B1(n_164),
.B2(n_166),
.Y(n_163)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_73),
.B(n_136),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_75),
.A2(n_85),
.B(n_86),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_77),
.Y(n_115)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_79),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_79),
.B(n_81),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.C(n_91),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_84),
.A2(n_89),
.B1(n_90),
.B2(n_145),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_84),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_85),
.B(n_88),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_85),
.A2(n_114),
.B1(n_165),
.B2(n_173),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_85),
.A2(n_114),
.B(n_229),
.Y(n_228)
);

AND2x2_ASAP7_75t_L g207 ( 
.A(n_86),
.B(n_183),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_91),
.B(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

OAI21xp33_ASAP7_75t_L g280 ( 
.A1(n_94),
.A2(n_281),
.B(n_282),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_111),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_97),
.B(n_112),
.C(n_122),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_98),
.A2(n_99),
.B1(n_100),
.B2(n_110),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_98),
.Y(n_110)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_106),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_101),
.B(n_106),
.C(n_110),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_102),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_102),
.A2(n_265),
.B(n_266),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_122),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_118),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_113),
.B(n_118),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g113 ( 
.A1(n_114),
.A2(n_115),
.B(n_116),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_114),
.A2(n_167),
.B(n_183),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g209 ( 
.A(n_119),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_120),
.B(n_141),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_196),
.B(n_200),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_151),
.B(n_195),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_146),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_146),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_143),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_130),
.B(n_137),
.C(n_143),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_131),
.B(n_135),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g132 ( 
.A(n_133),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_136),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_138),
.A2(n_139),
.B(n_141),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.C(n_149),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_192),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_148),
.B(n_149),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_190),
.B(n_194),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_179),
.B(n_189),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_168),
.B(n_178),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_155),
.B(n_163),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_156),
.A2(n_158),
.B1(n_161),
.B2(n_162),
.Y(n_155)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_156),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_158),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_158),
.B(n_161),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_169),
.A2(n_174),
.B(n_177),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_172),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_175),
.B(n_176),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_180),
.B(n_181),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_184),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_182),
.B(n_185),
.C(n_188),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_185),
.A2(n_186),
.B1(n_187),
.B2(n_188),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_187),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_191),
.B(n_193),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_191),
.B(n_193),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_199),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_220),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_220),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_204),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_203),
.B(n_205),
.C(n_212),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_212),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_208),
.B2(n_211),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_211),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_207),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_208),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_213),
.B(n_215),
.C(n_218),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.Y(n_214)
);

INVxp33_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_217),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_219),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_224),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_247),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_232),
.B1(n_245),
.B2(n_246),
.Y(n_225)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_226),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_226),
.B(n_246),
.C(n_247),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_228),
.B1(n_230),
.B2(n_231),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_227),
.A2(n_228),
.B1(n_263),
.B2(n_264),
.Y(n_262)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_228),
.B(n_230),
.Y(n_261)
);

AOI21xp33_ASAP7_75t_L g275 ( 
.A1(n_228),
.A2(n_261),
.B(n_263),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_232),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_236),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_233),
.B(n_237),
.C(n_241),
.Y(n_252)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_238),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g265 ( 
.A(n_244),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_269),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_250),
.B(n_269),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_268),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_254),
.C(n_260),
.Y(n_273)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_253),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_260),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_258),
.B(n_259),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_255),
.B(n_258),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g274 ( 
.A(n_259),
.B(n_275),
.CI(n_276),
.CON(n_274),
.SN(n_274)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_289),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_274),
.Y(n_290)
);

BUFx24_ASAP7_75t_SL g292 ( 
.A(n_274),
.Y(n_292)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_278),
.B1(n_285),
.B2(n_288),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_283),
.B2(n_284),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_285),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);


endmodule