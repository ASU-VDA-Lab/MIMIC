module fake_ariane_1640_n_1464 (n_295, n_170, n_190, n_160, n_64, n_180, n_119, n_124, n_307, n_294, n_197, n_176, n_34, n_172, n_183, n_299, n_12, n_133, n_66, n_205, n_71, n_109, n_245, n_96, n_319, n_49, n_20, n_283, n_50, n_187, n_318, n_103, n_244, n_226, n_220, n_261, n_36, n_189, n_72, n_286, n_57, n_117, n_139, n_85, n_130, n_214, n_2, n_32, n_138, n_162, n_264, n_137, n_122, n_198, n_232, n_52, n_73, n_77, n_15, n_23, n_87, n_279, n_207, n_41, n_140, n_151, n_28, n_146, n_230, n_270, n_194, n_154, n_142, n_285, n_186, n_202, n_145, n_193, n_59, n_315, n_311, n_239, n_35, n_272, n_54, n_8, n_167, n_90, n_38, n_47, n_153, n_18, n_269, n_75, n_158, n_69, n_259, n_95, n_143, n_152, n_120, n_169, n_106, n_173, n_242, n_309, n_320, n_115, n_267, n_291, n_62, n_210, n_200, n_166, n_253, n_218, n_79, n_3, n_271, n_247, n_91, n_240, n_128, n_224, n_44, n_82, n_31, n_222, n_256, n_227, n_48, n_188, n_323, n_11, n_129, n_126, n_282, n_277, n_248, n_301, n_293, n_228, n_276, n_93, n_108, n_303, n_168, n_81, n_1, n_206, n_238, n_136, n_192, n_300, n_14, n_163, n_88, n_141, n_104, n_314, n_16, n_273, n_305, n_312, n_233, n_56, n_60, n_221, n_321, n_86, n_89, n_149, n_237, n_175, n_74, n_19, n_40, n_181, n_53, n_260, n_310, n_236, n_281, n_24, n_7, n_209, n_262, n_17, n_225, n_235, n_297, n_290, n_46, n_84, n_199, n_107, n_217, n_178, n_42, n_308, n_201, n_70, n_10, n_287, n_302, n_6, n_94, n_284, n_4, n_249, n_37, n_58, n_65, n_123, n_212, n_278, n_255, n_257, n_148, n_135, n_171, n_61, n_102, n_182, n_316, n_196, n_125, n_43, n_13, n_27, n_254, n_219, n_55, n_231, n_234, n_280, n_215, n_252, n_161, n_298, n_68, n_78, n_63, n_99, n_216, n_5, n_223, n_25, n_83, n_288, n_179, n_195, n_213, n_110, n_304, n_67, n_306, n_313, n_92, n_203, n_150, n_98, n_113, n_114, n_33, n_111, n_21, n_274, n_296, n_265, n_208, n_156, n_292, n_174, n_275, n_100, n_132, n_147, n_204, n_51, n_76, n_26, n_246, n_0, n_159, n_105, n_30, n_131, n_263, n_229, n_250, n_165, n_144, n_317, n_101, n_243, n_134, n_185, n_289, n_9, n_112, n_45, n_268, n_266, n_164, n_157, n_184, n_177, n_258, n_118, n_121, n_22, n_241, n_29, n_191, n_80, n_211, n_97, n_322, n_251, n_116, n_39, n_155, n_127, n_1464);

input n_295;
input n_170;
input n_190;
input n_160;
input n_64;
input n_180;
input n_119;
input n_124;
input n_307;
input n_294;
input n_197;
input n_176;
input n_34;
input n_172;
input n_183;
input n_299;
input n_12;
input n_133;
input n_66;
input n_205;
input n_71;
input n_109;
input n_245;
input n_96;
input n_319;
input n_49;
input n_20;
input n_283;
input n_50;
input n_187;
input n_318;
input n_103;
input n_244;
input n_226;
input n_220;
input n_261;
input n_36;
input n_189;
input n_72;
input n_286;
input n_57;
input n_117;
input n_139;
input n_85;
input n_130;
input n_214;
input n_2;
input n_32;
input n_138;
input n_162;
input n_264;
input n_137;
input n_122;
input n_198;
input n_232;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_87;
input n_279;
input n_207;
input n_41;
input n_140;
input n_151;
input n_28;
input n_146;
input n_230;
input n_270;
input n_194;
input n_154;
input n_142;
input n_285;
input n_186;
input n_202;
input n_145;
input n_193;
input n_59;
input n_315;
input n_311;
input n_239;
input n_35;
input n_272;
input n_54;
input n_8;
input n_167;
input n_90;
input n_38;
input n_47;
input n_153;
input n_18;
input n_269;
input n_75;
input n_158;
input n_69;
input n_259;
input n_95;
input n_143;
input n_152;
input n_120;
input n_169;
input n_106;
input n_173;
input n_242;
input n_309;
input n_320;
input n_115;
input n_267;
input n_291;
input n_62;
input n_210;
input n_200;
input n_166;
input n_253;
input n_218;
input n_79;
input n_3;
input n_271;
input n_247;
input n_91;
input n_240;
input n_128;
input n_224;
input n_44;
input n_82;
input n_31;
input n_222;
input n_256;
input n_227;
input n_48;
input n_188;
input n_323;
input n_11;
input n_129;
input n_126;
input n_282;
input n_277;
input n_248;
input n_301;
input n_293;
input n_228;
input n_276;
input n_93;
input n_108;
input n_303;
input n_168;
input n_81;
input n_1;
input n_206;
input n_238;
input n_136;
input n_192;
input n_300;
input n_14;
input n_163;
input n_88;
input n_141;
input n_104;
input n_314;
input n_16;
input n_273;
input n_305;
input n_312;
input n_233;
input n_56;
input n_60;
input n_221;
input n_321;
input n_86;
input n_89;
input n_149;
input n_237;
input n_175;
input n_74;
input n_19;
input n_40;
input n_181;
input n_53;
input n_260;
input n_310;
input n_236;
input n_281;
input n_24;
input n_7;
input n_209;
input n_262;
input n_17;
input n_225;
input n_235;
input n_297;
input n_290;
input n_46;
input n_84;
input n_199;
input n_107;
input n_217;
input n_178;
input n_42;
input n_308;
input n_201;
input n_70;
input n_10;
input n_287;
input n_302;
input n_6;
input n_94;
input n_284;
input n_4;
input n_249;
input n_37;
input n_58;
input n_65;
input n_123;
input n_212;
input n_278;
input n_255;
input n_257;
input n_148;
input n_135;
input n_171;
input n_61;
input n_102;
input n_182;
input n_316;
input n_196;
input n_125;
input n_43;
input n_13;
input n_27;
input n_254;
input n_219;
input n_55;
input n_231;
input n_234;
input n_280;
input n_215;
input n_252;
input n_161;
input n_298;
input n_68;
input n_78;
input n_63;
input n_99;
input n_216;
input n_5;
input n_223;
input n_25;
input n_83;
input n_288;
input n_179;
input n_195;
input n_213;
input n_110;
input n_304;
input n_67;
input n_306;
input n_313;
input n_92;
input n_203;
input n_150;
input n_98;
input n_113;
input n_114;
input n_33;
input n_111;
input n_21;
input n_274;
input n_296;
input n_265;
input n_208;
input n_156;
input n_292;
input n_174;
input n_275;
input n_100;
input n_132;
input n_147;
input n_204;
input n_51;
input n_76;
input n_26;
input n_246;
input n_0;
input n_159;
input n_105;
input n_30;
input n_131;
input n_263;
input n_229;
input n_250;
input n_165;
input n_144;
input n_317;
input n_101;
input n_243;
input n_134;
input n_185;
input n_289;
input n_9;
input n_112;
input n_45;
input n_268;
input n_266;
input n_164;
input n_157;
input n_184;
input n_177;
input n_258;
input n_118;
input n_121;
input n_22;
input n_241;
input n_29;
input n_191;
input n_80;
input n_211;
input n_97;
input n_322;
input n_251;
input n_116;
input n_39;
input n_155;
input n_127;

output n_1464;

wire n_913;
wire n_589;
wire n_1174;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_1463;
wire n_1238;
wire n_817;
wire n_924;
wire n_781;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_764;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1366;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_520;
wire n_870;
wire n_1453;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_338;
wire n_995;
wire n_1184;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_402;
wire n_1277;
wire n_829;
wire n_1062;
wire n_339;
wire n_738;
wire n_672;
wire n_740;
wire n_1283;
wire n_1018;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_989;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1276;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1195;
wire n_518;
wire n_1207;
wire n_786;
wire n_1404;
wire n_868;
wire n_1314;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1085;
wire n_432;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_587;
wire n_693;
wire n_863;
wire n_1254;
wire n_929;
wire n_352;
wire n_899;
wire n_611;
wire n_1295;
wire n_365;
wire n_1013;
wire n_334;
wire n_661;
wire n_533;
wire n_438;
wire n_440;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_490;
wire n_1461;
wire n_1391;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_676;
wire n_680;
wire n_380;
wire n_1432;
wire n_1108;
wire n_355;
wire n_851;
wire n_444;
wire n_1351;
wire n_1274;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_366;
wire n_762;
wire n_1253;
wire n_555;
wire n_804;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1026;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_619;
wire n_437;
wire n_337;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_1079;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1343;
wire n_563;
wire n_990;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_964;
wire n_382;
wire n_489;
wire n_974;
wire n_506;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1209;
wire n_1020;
wire n_646;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1455;
wire n_836;
wire n_1279;
wire n_564;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_713;
wire n_1255;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_1095;
wire n_370;
wire n_706;
wire n_1401;
wire n_1419;
wire n_776;
wire n_424;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_441;
wire n_1032;
wire n_1217;
wire n_637;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_905;
wire n_720;
wire n_926;
wire n_1163;
wire n_1384;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_487;
wire n_1456;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1287;
wire n_405;
wire n_1414;
wire n_1134;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_529;
wire n_502;
wire n_1304;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1061;
wire n_326;
wire n_681;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_1015;
wire n_545;
wire n_1377;
wire n_1162;
wire n_536;
wire n_325;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_442;
wire n_777;
wire n_1080;
wire n_920;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1371;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1218;
wire n_861;
wire n_1431;
wire n_877;
wire n_1119;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_735;
wire n_1005;
wire n_527;
wire n_1294;
wire n_888;
wire n_845;
wire n_1297;
wire n_551;
wire n_417;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_769;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_1075;
wire n_454;
wire n_1331;
wire n_1227;
wire n_655;
wire n_403;
wire n_1007;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_430;
wire n_1206;
wire n_722;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_521;
wire n_873;
wire n_1301;
wire n_1243;
wire n_1400;
wire n_342;
wire n_358;
wire n_608;
wire n_1037;
wire n_1329;
wire n_1257;
wire n_1078;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_1449;
wire n_687;
wire n_797;
wire n_480;
wire n_1327;
wire n_642;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_592;
wire n_854;
wire n_1318;
wire n_393;
wire n_474;
wire n_805;
wire n_1072;
wire n_695;
wire n_1305;
wire n_730;
wire n_386;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_640;
wire n_463;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_878;
wire n_771;
wire n_1321;
wire n_752;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_806;
wire n_1350;
wire n_649;
wire n_374;
wire n_1352;
wire n_643;
wire n_1441;
wire n_682;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_979;
wire n_897;
wire n_949;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1448;
wire n_1009;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1438;
wire n_597;
wire n_1047;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_1090;
wire n_1367;
wire n_928;
wire n_1153;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1192;
wire n_894;
wire n_1380;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_328;
wire n_368;
wire n_467;
wire n_1422;
wire n_644;
wire n_1197;
wire n_497;
wire n_1165;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1440;
wire n_1370;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1403;
wire n_1065;
wire n_453;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_593;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1040;
wire n_674;
wire n_1158;
wire n_1444;
wire n_820;
wire n_872;
wire n_1157;
wire n_848;
wire n_629;
wire n_532;
wire n_763;
wire n_540;
wire n_692;
wire n_984;
wire n_750;
wire n_834;
wire n_800;
wire n_395;
wire n_621;
wire n_1014;
wire n_724;
wire n_1427;
wire n_493;
wire n_1311;
wire n_1100;
wire n_585;
wire n_875;
wire n_827;
wire n_697;
wire n_622;
wire n_1335;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_739;
wire n_1028;
wire n_1221;
wire n_530;
wire n_792;
wire n_1262;
wire n_580;
wire n_494;
wire n_434;
wire n_975;
wire n_394;
wire n_923;
wire n_1124;
wire n_1381;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1407;
wire n_1204;
wire n_994;
wire n_1360;
wire n_973;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1054;
wire n_508;
wire n_353;
wire n_1361;
wire n_1057;
wire n_1011;
wire n_978;
wire n_828;
wire n_1411;
wire n_1359;
wire n_558;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1008;
wire n_332;
wire n_581;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1385;
wire n_541;
wire n_499;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1458;
wire n_679;
wire n_663;
wire n_443;
wire n_1412;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_391;
wire n_940;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1093;
wire n_1285;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1452;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_816;
wire n_1322;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1099;
wire n_839;
wire n_759;
wire n_567;
wire n_369;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_550;
wire n_1315;
wire n_997;
wire n_635;
wire n_694;
wire n_1320;
wire n_1113;
wire n_1152;
wire n_921;
wire n_1236;
wire n_1265;
wire n_671;
wire n_1409;
wire n_1148;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1289;
wire n_459;
wire n_1136;
wire n_458;
wire n_1190;
wire n_1144;
wire n_383;
wire n_838;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_709;
wire n_809;
wire n_881;
wire n_1019;
wire n_662;
wire n_641;
wire n_910;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_1114;
wire n_1325;
wire n_708;
wire n_1223;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_450;
wire n_896;
wire n_902;
wire n_1031;
wire n_853;
wire n_716;
wire n_1337;
wire n_774;
wire n_933;
wire n_596;
wire n_954;
wire n_1168;
wire n_1310;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_1229;
wire n_415;
wire n_1280;
wire n_544;
wire n_1186;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1126;
wire n_938;
wire n_1328;
wire n_895;
wire n_583;
wire n_1302;
wire n_1000;
wire n_626;
wire n_378;
wire n_946;
wire n_757;
wire n_375;
wire n_1146;
wire n_1203;
wire n_998;
wire n_472;
wire n_937;
wire n_1375;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_496;
wire n_866;
wire n_925;
wire n_1313;
wire n_1001;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1051;
wire n_719;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_548;
wire n_523;
wire n_457;
wire n_1299;
wire n_782;
wire n_364;
wire n_431;
wire n_1228;
wire n_1244;
wire n_411;
wire n_484;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1233;
wire n_893;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1374;
wire n_1451;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_157),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_185),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_217),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_300),
.Y(n_327)
);

INVx1_ASAP7_75t_SL g328 ( 
.A(n_60),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_226),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_280),
.Y(n_330)
);

BUFx3_ASAP7_75t_L g331 ( 
.A(n_204),
.Y(n_331)
);

CKINVDCx14_ASAP7_75t_R g332 ( 
.A(n_139),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_230),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_252),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g335 ( 
.A(n_261),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_133),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_170),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_315),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_264),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_90),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_207),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_307),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_253),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_1),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_266),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_16),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_2),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_59),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_249),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_110),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_158),
.Y(n_352)
);

BUFx10_ASAP7_75t_L g353 ( 
.A(n_254),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_114),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_182),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_242),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_269),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_120),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_12),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_285),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_184),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_135),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_165),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_299),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_257),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_199),
.Y(n_366)
);

INVx1_ASAP7_75t_SL g367 ( 
.A(n_308),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_37),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_236),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_316),
.Y(n_370)
);

INVx2_ASAP7_75t_SL g371 ( 
.A(n_245),
.Y(n_371)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_231),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_241),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g374 ( 
.A(n_247),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_183),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_128),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_221),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_26),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_235),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_132),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_39),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_234),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_80),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_116),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_60),
.Y(n_385)
);

BUFx10_ASAP7_75t_L g386 ( 
.A(n_98),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_258),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_13),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_203),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_295),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_136),
.Y(n_391)
);

CKINVDCx5p33_ASAP7_75t_R g392 ( 
.A(n_54),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_15),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_276),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_58),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_152),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_304),
.Y(n_397)
);

INVx4_ASAP7_75t_R g398 ( 
.A(n_191),
.Y(n_398)
);

BUFx2_ASAP7_75t_SL g399 ( 
.A(n_206),
.Y(n_399)
);

INVx2_ASAP7_75t_SL g400 ( 
.A(n_259),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_61),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_6),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_215),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g405 ( 
.A(n_84),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_176),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_298),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_92),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_220),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_313),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_63),
.Y(n_411)
);

BUFx6f_ASAP7_75t_L g412 ( 
.A(n_115),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_15),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_127),
.Y(n_414)
);

CKINVDCx20_ASAP7_75t_R g415 ( 
.A(n_237),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_51),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_95),
.Y(n_417)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_150),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_192),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_273),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_129),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_160),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_162),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_48),
.Y(n_424)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_45),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_188),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_303),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_119),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_88),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_229),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_82),
.Y(n_431)
);

INVxp67_ASAP7_75t_SL g432 ( 
.A(n_250),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_214),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_1),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_218),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_64),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_123),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_272),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_18),
.Y(n_439)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_16),
.Y(n_440)
);

CKINVDCx5p33_ASAP7_75t_R g441 ( 
.A(n_36),
.Y(n_441)
);

BUFx3_ASAP7_75t_L g442 ( 
.A(n_301),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_140),
.Y(n_443)
);

CKINVDCx20_ASAP7_75t_R g444 ( 
.A(n_251),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g445 ( 
.A(n_198),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_96),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_25),
.Y(n_447)
);

CKINVDCx16_ASAP7_75t_R g448 ( 
.A(n_200),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_244),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_111),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_144),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_122),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_51),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_256),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_209),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_8),
.Y(n_456)
);

INVx1_ASAP7_75t_SL g457 ( 
.A(n_163),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_105),
.Y(n_458)
);

CKINVDCx5p33_ASAP7_75t_R g459 ( 
.A(n_145),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_118),
.Y(n_460)
);

CKINVDCx5p33_ASAP7_75t_R g461 ( 
.A(n_156),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_34),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_108),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_149),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_196),
.Y(n_465)
);

INVxp67_ASAP7_75t_L g466 ( 
.A(n_177),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_155),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_0),
.Y(n_468)
);

BUFx3_ASAP7_75t_L g469 ( 
.A(n_97),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_143),
.Y(n_470)
);

BUFx5_ASAP7_75t_L g471 ( 
.A(n_255),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_102),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_34),
.Y(n_473)
);

INVx1_ASAP7_75t_SL g474 ( 
.A(n_239),
.Y(n_474)
);

CKINVDCx20_ASAP7_75t_R g475 ( 
.A(n_282),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_317),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_31),
.Y(n_477)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_211),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_74),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_29),
.Y(n_480)
);

BUFx6f_ASAP7_75t_L g481 ( 
.A(n_106),
.Y(n_481)
);

CKINVDCx20_ASAP7_75t_R g482 ( 
.A(n_297),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_59),
.Y(n_483)
);

CKINVDCx5p33_ASAP7_75t_R g484 ( 
.A(n_213),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_284),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_77),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_302),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_79),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_85),
.Y(n_489)
);

BUFx3_ASAP7_75t_L g490 ( 
.A(n_305),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_291),
.Y(n_491)
);

CKINVDCx5p33_ASAP7_75t_R g492 ( 
.A(n_194),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_270),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_197),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_142),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_322),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_195),
.Y(n_497)
);

CKINVDCx5p33_ASAP7_75t_R g498 ( 
.A(n_289),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_73),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_223),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_275),
.Y(n_501)
);

CKINVDCx5p33_ASAP7_75t_R g502 ( 
.A(n_306),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_312),
.Y(n_503)
);

INVx1_ASAP7_75t_SL g504 ( 
.A(n_168),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_210),
.Y(n_505)
);

BUFx2_ASAP7_75t_SL g506 ( 
.A(n_225),
.Y(n_506)
);

BUFx2_ASAP7_75t_L g507 ( 
.A(n_190),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_26),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_24),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_19),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_202),
.Y(n_511)
);

CKINVDCx5p33_ASAP7_75t_R g512 ( 
.A(n_201),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g513 ( 
.A(n_20),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_405),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_329),
.B(n_0),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_425),
.B(n_2),
.Y(n_516)
);

INVx5_ASAP7_75t_L g517 ( 
.A(n_333),
.Y(n_517)
);

BUFx6f_ASAP7_75t_L g518 ( 
.A(n_333),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_330),
.B(n_3),
.Y(n_519)
);

BUFx12f_ASAP7_75t_L g520 ( 
.A(n_353),
.Y(n_520)
);

INVx5_ASAP7_75t_L g521 ( 
.A(n_333),
.Y(n_521)
);

INVx2_ASAP7_75t_SL g522 ( 
.A(n_402),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_SL g523 ( 
.A(n_372),
.B(n_67),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_SL g524 ( 
.A(n_448),
.B(n_353),
.Y(n_524)
);

INVxp33_ASAP7_75t_SL g525 ( 
.A(n_344),
.Y(n_525)
);

BUFx8_ASAP7_75t_SL g526 ( 
.A(n_513),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_424),
.B(n_3),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_333),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_331),
.B(n_4),
.Y(n_529)
);

HB1xp67_ASAP7_75t_L g530 ( 
.A(n_425),
.Y(n_530)
);

AND2x2_ASAP7_75t_L g531 ( 
.A(n_332),
.B(n_4),
.Y(n_531)
);

INVx5_ASAP7_75t_L g532 ( 
.A(n_412),
.Y(n_532)
);

BUFx3_ASAP7_75t_L g533 ( 
.A(n_331),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_343),
.B(n_345),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_477),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_350),
.B(n_5),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_347),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_442),
.B(n_5),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_332),
.B(n_6),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_412),
.Y(n_540)
);

INVx5_ASAP7_75t_L g541 ( 
.A(n_412),
.Y(n_541)
);

INVx5_ASAP7_75t_L g542 ( 
.A(n_412),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_442),
.B(n_469),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_477),
.Y(n_544)
);

INVx5_ASAP7_75t_L g545 ( 
.A(n_481),
.Y(n_545)
);

HB1xp67_ASAP7_75t_L g546 ( 
.A(n_348),
.Y(n_546)
);

INVx3_ASAP7_75t_L g547 ( 
.A(n_477),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_469),
.B(n_7),
.Y(n_548)
);

BUFx6f_ASAP7_75t_L g549 ( 
.A(n_481),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_481),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_355),
.B(n_7),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_SL g552 ( 
.A(n_353),
.B(n_8),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_477),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_361),
.B(n_9),
.Y(n_554)
);

CKINVDCx5p33_ASAP7_75t_R g555 ( 
.A(n_334),
.Y(n_555)
);

INVx3_ASAP7_75t_L g556 ( 
.A(n_386),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_490),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_386),
.Y(n_558)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_363),
.B(n_9),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_490),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_378),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_365),
.B(n_10),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_375),
.B(n_10),
.Y(n_563)
);

INVx4_ASAP7_75t_L g564 ( 
.A(n_481),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_386),
.Y(n_565)
);

AND2x4_ASAP7_75t_L g566 ( 
.A(n_388),
.B(n_11),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_395),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_328),
.B(n_11),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_377),
.B(n_12),
.Y(n_569)
);

BUFx6f_ASAP7_75t_L g570 ( 
.A(n_486),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_486),
.Y(n_571)
);

INVx5_ASAP7_75t_L g572 ( 
.A(n_486),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_440),
.B(n_13),
.Y(n_573)
);

BUFx6f_ASAP7_75t_L g574 ( 
.A(n_486),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_389),
.B(n_14),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_418),
.Y(n_576)
);

HB1xp67_ASAP7_75t_L g577 ( 
.A(n_411),
.Y(n_577)
);

AND2x4_ASAP7_75t_L g578 ( 
.A(n_413),
.B(n_14),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_394),
.B(n_17),
.Y(n_579)
);

BUFx12f_ASAP7_75t_L g580 ( 
.A(n_346),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_408),
.B(n_17),
.Y(n_581)
);

BUFx3_ASAP7_75t_L g582 ( 
.A(n_409),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_359),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_419),
.B(n_18),
.Y(n_584)
);

INVx5_ASAP7_75t_L g585 ( 
.A(n_371),
.Y(n_585)
);

BUFx8_ASAP7_75t_SL g586 ( 
.A(n_513),
.Y(n_586)
);

BUFx6f_ASAP7_75t_L g587 ( 
.A(n_404),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_421),
.B(n_19),
.Y(n_588)
);

INVx4_ASAP7_75t_L g589 ( 
.A(n_324),
.Y(n_589)
);

BUFx6f_ASAP7_75t_L g590 ( 
.A(n_404),
.Y(n_590)
);

BUFx6f_ASAP7_75t_L g591 ( 
.A(n_417),
.Y(n_591)
);

INVx5_ASAP7_75t_L g592 ( 
.A(n_400),
.Y(n_592)
);

BUFx12f_ASAP7_75t_L g593 ( 
.A(n_368),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_416),
.B(n_20),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_417),
.Y(n_595)
);

NAND2xp5_ASAP7_75t_L g596 ( 
.A(n_435),
.B(n_21),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_L g597 ( 
.A(n_437),
.B(n_21),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_438),
.B(n_22),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_434),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_436),
.B(n_439),
.Y(n_600)
);

HB1xp67_ASAP7_75t_L g601 ( 
.A(n_453),
.Y(n_601)
);

AND2x4_ASAP7_75t_L g602 ( 
.A(n_473),
.B(n_22),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_458),
.B(n_23),
.Y(n_603)
);

AND2x2_ASAP7_75t_L g604 ( 
.A(n_480),
.B(n_23),
.Y(n_604)
);

AND2x4_ASAP7_75t_L g605 ( 
.A(n_509),
.B(n_24),
.Y(n_605)
);

AND2x2_ASAP7_75t_L g606 ( 
.A(n_381),
.B(n_25),
.Y(n_606)
);

INVx2_ASAP7_75t_L g607 ( 
.A(n_418),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_460),
.B(n_27),
.Y(n_608)
);

BUFx6f_ASAP7_75t_L g609 ( 
.A(n_431),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_418),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_431),
.Y(n_611)
);

BUFx6f_ASAP7_75t_L g612 ( 
.A(n_452),
.Y(n_612)
);

BUFx8_ASAP7_75t_SL g613 ( 
.A(n_335),
.Y(n_613)
);

BUFx12f_ASAP7_75t_L g614 ( 
.A(n_385),
.Y(n_614)
);

BUFx3_ASAP7_75t_L g615 ( 
.A(n_489),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_494),
.B(n_27),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_452),
.Y(n_617)
);

INVx5_ASAP7_75t_L g618 ( 
.A(n_423),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_496),
.B(n_28),
.Y(n_619)
);

BUFx6f_ASAP7_75t_L g620 ( 
.A(n_497),
.Y(n_620)
);

BUFx3_ASAP7_75t_L g621 ( 
.A(n_499),
.Y(n_621)
);

BUFx6f_ASAP7_75t_L g622 ( 
.A(n_497),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_418),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_503),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_505),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_398),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_392),
.Y(n_627)
);

BUFx8_ASAP7_75t_SL g628 ( 
.A(n_357),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_524),
.A2(n_410),
.B1(n_415),
.B2(n_370),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_587),
.Y(n_630)
);

AOI22xp5_ASAP7_75t_L g631 ( 
.A1(n_531),
.A2(n_539),
.B1(n_514),
.B2(n_516),
.Y(n_631)
);

INVx8_ASAP7_75t_L g632 ( 
.A(n_520),
.Y(n_632)
);

AND2x2_ASAP7_75t_L g633 ( 
.A(n_530),
.B(n_393),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_547),
.Y(n_634)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_537),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_547),
.Y(n_636)
);

BUFx6f_ASAP7_75t_SL g637 ( 
.A(n_558),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_SL g638 ( 
.A(n_523),
.B(n_426),
.Y(n_638)
);

AO22x2_ASAP7_75t_L g639 ( 
.A1(n_552),
.A2(n_367),
.B1(n_445),
.B2(n_374),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_564),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_SL g641 ( 
.A1(n_555),
.A2(n_472),
.B1(n_475),
.B2(n_444),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_561),
.Y(n_642)
);

INVx2_ASAP7_75t_SL g643 ( 
.A(n_556),
.Y(n_643)
);

OAI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_552),
.A2(n_401),
.B1(n_447),
.B2(n_441),
.Y(n_644)
);

OAI22xp5_ASAP7_75t_SL g645 ( 
.A1(n_530),
.A2(n_482),
.B1(n_456),
.B2(n_468),
.Y(n_645)
);

AND2x2_ASAP7_75t_SL g646 ( 
.A(n_516),
.B(n_399),
.Y(n_646)
);

OAI22xp33_ASAP7_75t_L g647 ( 
.A1(n_522),
.A2(n_483),
.B1(n_508),
.B2(n_462),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_556),
.B(n_358),
.Y(n_648)
);

INVx2_ASAP7_75t_SL g649 ( 
.A(n_565),
.Y(n_649)
);

AND2x2_ASAP7_75t_SL g650 ( 
.A(n_529),
.B(n_506),
.Y(n_650)
);

AOI22xp5_ASAP7_75t_L g651 ( 
.A1(n_525),
.A2(n_510),
.B1(n_457),
.B2(n_504),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_543),
.B(n_583),
.Y(n_652)
);

AOI22xp5_ASAP7_75t_L g653 ( 
.A1(n_568),
.A2(n_573),
.B1(n_606),
.B2(n_529),
.Y(n_653)
);

AO22x2_ASAP7_75t_L g654 ( 
.A1(n_527),
.A2(n_538),
.B1(n_578),
.B2(n_566),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_613),
.Y(n_655)
);

OAI22xp33_ASAP7_75t_L g656 ( 
.A1(n_534),
.A2(n_474),
.B1(n_478),
.B2(n_466),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_533),
.B(n_325),
.Y(n_657)
);

OAI22xp33_ASAP7_75t_L g658 ( 
.A1(n_546),
.A2(n_432),
.B1(n_327),
.B2(n_336),
.Y(n_658)
);

OAI22xp33_ASAP7_75t_L g659 ( 
.A1(n_546),
.A2(n_337),
.B1(n_338),
.B2(n_326),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_587),
.Y(n_660)
);

AO22x2_ASAP7_75t_L g661 ( 
.A1(n_527),
.A2(n_30),
.B1(n_28),
.B2(n_29),
.Y(n_661)
);

OAI22xp5_ASAP7_75t_SL g662 ( 
.A1(n_580),
.A2(n_340),
.B1(n_341),
.B2(n_339),
.Y(n_662)
);

AOI22xp5_ASAP7_75t_L g663 ( 
.A1(n_538),
.A2(n_349),
.B1(n_351),
.B2(n_342),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_535),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_587),
.Y(n_665)
);

AO22x2_ASAP7_75t_L g666 ( 
.A1(n_566),
.A2(n_32),
.B1(n_30),
.B2(n_31),
.Y(n_666)
);

AND2x4_ASAP7_75t_SL g667 ( 
.A(n_627),
.B(n_589),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_533),
.B(n_352),
.Y(n_668)
);

AND2x2_ASAP7_75t_L g669 ( 
.A(n_560),
.B(n_354),
.Y(n_669)
);

OAI22xp5_ASAP7_75t_L g670 ( 
.A1(n_578),
.A2(n_360),
.B1(n_362),
.B2(n_356),
.Y(n_670)
);

AO22x2_ASAP7_75t_L g671 ( 
.A1(n_602),
.A2(n_35),
.B1(n_32),
.B2(n_33),
.Y(n_671)
);

AND2x2_ASAP7_75t_SL g672 ( 
.A(n_548),
.B(n_602),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_587),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_SL g674 ( 
.A1(n_515),
.A2(n_554),
.B1(n_559),
.B2(n_519),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_560),
.B(n_364),
.Y(n_675)
);

AO22x2_ASAP7_75t_L g676 ( 
.A1(n_605),
.A2(n_36),
.B1(n_33),
.B2(n_35),
.Y(n_676)
);

CKINVDCx5p33_ASAP7_75t_R g677 ( 
.A(n_613),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_627),
.B(n_366),
.Y(n_678)
);

OAI22xp5_ASAP7_75t_SL g679 ( 
.A1(n_593),
.A2(n_373),
.B1(n_376),
.B2(n_369),
.Y(n_679)
);

OAI22xp33_ASAP7_75t_L g680 ( 
.A1(n_577),
.A2(n_380),
.B1(n_382),
.B2(n_379),
.Y(n_680)
);

AO22x2_ASAP7_75t_L g681 ( 
.A1(n_605),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_626),
.B(n_383),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_535),
.Y(n_683)
);

AOI22xp5_ASAP7_75t_L g684 ( 
.A1(n_614),
.A2(n_512),
.B1(n_511),
.B2(n_502),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_544),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_626),
.B(n_384),
.Y(n_686)
);

OAI22xp5_ASAP7_75t_SL g687 ( 
.A1(n_577),
.A2(n_501),
.B1(n_500),
.B2(n_498),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_626),
.B(n_387),
.Y(n_688)
);

INVx8_ASAP7_75t_L g689 ( 
.A(n_626),
.Y(n_689)
);

OAI22xp5_ASAP7_75t_L g690 ( 
.A1(n_562),
.A2(n_495),
.B1(n_493),
.B2(n_492),
.Y(n_690)
);

AOI22xp5_ASAP7_75t_SL g691 ( 
.A1(n_526),
.A2(n_491),
.B1(n_488),
.B2(n_487),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_590),
.Y(n_692)
);

OAI22xp33_ASAP7_75t_SL g693 ( 
.A1(n_563),
.A2(n_485),
.B1(n_484),
.B2(n_479),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g694 ( 
.A(n_589),
.B(n_390),
.Y(n_694)
);

OAI22xp5_ASAP7_75t_SL g695 ( 
.A1(n_601),
.A2(n_476),
.B1(n_470),
.B2(n_467),
.Y(n_695)
);

OAI22xp33_ASAP7_75t_L g696 ( 
.A1(n_601),
.A2(n_465),
.B1(n_396),
.B2(n_397),
.Y(n_696)
);

AOI22xp5_ASAP7_75t_L g697 ( 
.A1(n_536),
.A2(n_433),
.B1(n_464),
.B2(n_463),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_544),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_553),
.Y(n_699)
);

OR2x2_ASAP7_75t_L g700 ( 
.A(n_567),
.B(n_38),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_582),
.B(n_391),
.Y(n_701)
);

AND2x2_ASAP7_75t_L g702 ( 
.A(n_600),
.B(n_403),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_567),
.B(n_40),
.Y(n_703)
);

OAI22xp33_ASAP7_75t_R g704 ( 
.A1(n_536),
.A2(n_40),
.B1(n_41),
.B2(n_42),
.Y(n_704)
);

AND2x2_ASAP7_75t_L g705 ( 
.A(n_582),
.B(n_406),
.Y(n_705)
);

OAI22xp33_ASAP7_75t_L g706 ( 
.A1(n_569),
.A2(n_407),
.B1(n_414),
.B2(n_420),
.Y(n_706)
);

INVx2_ASAP7_75t_L g707 ( 
.A(n_553),
.Y(n_707)
);

AOI22xp5_ASAP7_75t_L g708 ( 
.A1(n_551),
.A2(n_446),
.B1(n_461),
.B2(n_459),
.Y(n_708)
);

AO22x2_ASAP7_75t_L g709 ( 
.A1(n_594),
.A2(n_41),
.B1(n_42),
.B2(n_43),
.Y(n_709)
);

OAI22xp5_ASAP7_75t_SL g710 ( 
.A1(n_551),
.A2(n_422),
.B1(n_427),
.B2(n_428),
.Y(n_710)
);

OR2x6_ASAP7_75t_L g711 ( 
.A(n_599),
.B(n_604),
.Y(n_711)
);

OAI22xp33_ASAP7_75t_SL g712 ( 
.A1(n_579),
.A2(n_429),
.B1(n_430),
.B2(n_443),
.Y(n_712)
);

AO22x2_ASAP7_75t_L g713 ( 
.A1(n_624),
.A2(n_43),
.B1(n_44),
.B2(n_45),
.Y(n_713)
);

OAI22xp33_ASAP7_75t_SL g714 ( 
.A1(n_581),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.Y(n_714)
);

AOI22xp5_ASAP7_75t_L g715 ( 
.A1(n_575),
.A2(n_455),
.B1(n_454),
.B2(n_471),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_564),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_575),
.A2(n_471),
.B1(n_418),
.B2(n_47),
.Y(n_717)
);

BUFx3_ASAP7_75t_L g718 ( 
.A(n_632),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_635),
.Y(n_719)
);

HB1xp67_ASAP7_75t_L g720 ( 
.A(n_652),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_642),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_716),
.Y(n_722)
);

AND2x2_ASAP7_75t_L g723 ( 
.A(n_702),
.B(n_615),
.Y(n_723)
);

NAND2x1p5_ASAP7_75t_L g724 ( 
.A(n_650),
.B(n_615),
.Y(n_724)
);

AND2x2_ASAP7_75t_L g725 ( 
.A(n_633),
.B(n_621),
.Y(n_725)
);

NAND2xp33_ASAP7_75t_SL g726 ( 
.A(n_637),
.B(n_584),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_634),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_636),
.Y(n_728)
);

NAND2x1p5_ASAP7_75t_L g729 ( 
.A(n_672),
.B(n_621),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_630),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_701),
.B(n_625),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_630),
.Y(n_732)
);

INVx1_ASAP7_75t_SL g733 ( 
.A(n_701),
.Y(n_733)
);

AND2x2_ASAP7_75t_L g734 ( 
.A(n_654),
.B(n_625),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_692),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_692),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_640),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_L g738 ( 
.A(n_640),
.B(n_576),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_660),
.Y(n_739)
);

XOR2x2_ASAP7_75t_L g740 ( 
.A(n_641),
.B(n_526),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_643),
.B(n_585),
.Y(n_741)
);

CKINVDCx20_ASAP7_75t_R g742 ( 
.A(n_655),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_665),
.Y(n_743)
);

AND2x6_ASAP7_75t_L g744 ( 
.A(n_717),
.B(n_557),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_654),
.B(n_557),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_673),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_664),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_711),
.B(n_599),
.Y(n_748)
);

INVx1_ASAP7_75t_L g749 ( 
.A(n_683),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_685),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_698),
.Y(n_751)
);

NOR2xp33_ASAP7_75t_SL g752 ( 
.A(n_638),
.B(n_588),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_674),
.B(n_576),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_699),
.Y(n_754)
);

INVx1_ASAP7_75t_L g755 ( 
.A(n_707),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_648),
.B(n_585),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_678),
.B(n_585),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_705),
.B(n_588),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_700),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_657),
.Y(n_760)
);

AND2x6_ASAP7_75t_L g761 ( 
.A(n_653),
.B(n_607),
.Y(n_761)
);

INVxp33_ASAP7_75t_SL g762 ( 
.A(n_677),
.Y(n_762)
);

INVx2_ASAP7_75t_L g763 ( 
.A(n_668),
.Y(n_763)
);

OAI21xp5_ASAP7_75t_L g764 ( 
.A1(n_715),
.A2(n_597),
.B(n_596),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_689),
.Y(n_765)
);

NOR2xp67_ASAP7_75t_L g766 ( 
.A(n_649),
.B(n_585),
.Y(n_766)
);

INVx1_ASAP7_75t_L g767 ( 
.A(n_669),
.Y(n_767)
);

NAND2x1p5_ASAP7_75t_L g768 ( 
.A(n_646),
.B(n_590),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_675),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_711),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_682),
.A2(n_610),
.B(n_607),
.Y(n_771)
);

CKINVDCx20_ASAP7_75t_R g772 ( 
.A(n_629),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_686),
.A2(n_623),
.B(n_610),
.Y(n_773)
);

INVxp67_ASAP7_75t_L g774 ( 
.A(n_694),
.Y(n_774)
);

AND2x2_ASAP7_75t_L g775 ( 
.A(n_631),
.B(n_616),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_703),
.Y(n_776)
);

NOR2xp67_ASAP7_75t_L g777 ( 
.A(n_684),
.B(n_592),
.Y(n_777)
);

INVx2_ASAP7_75t_L g778 ( 
.A(n_667),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_703),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_713),
.Y(n_780)
);

OR2x2_ASAP7_75t_L g781 ( 
.A(n_632),
.B(n_651),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_661),
.Y(n_782)
);

NOR2xp33_ASAP7_75t_L g783 ( 
.A(n_670),
.B(n_592),
.Y(n_783)
);

OAI21xp5_ASAP7_75t_L g784 ( 
.A1(n_697),
.A2(n_603),
.B(n_598),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_713),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_L g786 ( 
.A(n_689),
.B(n_623),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_688),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_661),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_708),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_666),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_666),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_659),
.B(n_592),
.Y(n_792)
);

AND2x2_ASAP7_75t_L g793 ( 
.A(n_691),
.B(n_616),
.Y(n_793)
);

OR2x2_ASAP7_75t_L g794 ( 
.A(n_645),
.B(n_608),
.Y(n_794)
);

CKINVDCx20_ASAP7_75t_R g795 ( 
.A(n_662),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_671),
.Y(n_796)
);

XOR2xp5_ASAP7_75t_L g797 ( 
.A(n_679),
.B(n_628),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_671),
.Y(n_798)
);

AOI21xp5_ASAP7_75t_L g799 ( 
.A1(n_690),
.A2(n_619),
.B(n_591),
.Y(n_799)
);

XOR2xp5_ASAP7_75t_L g800 ( 
.A(n_687),
.B(n_695),
.Y(n_800)
);

OAI21xp5_ASAP7_75t_L g801 ( 
.A1(n_663),
.A2(n_706),
.B(n_656),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_676),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_676),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_680),
.B(n_592),
.Y(n_804)
);

XNOR2xp5_ASAP7_75t_L g805 ( 
.A(n_639),
.B(n_628),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_681),
.Y(n_806)
);

HB1xp67_ASAP7_75t_L g807 ( 
.A(n_733),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_774),
.B(n_639),
.Y(n_808)
);

BUFx6f_ASAP7_75t_L g809 ( 
.A(n_765),
.Y(n_809)
);

OAI21xp5_ASAP7_75t_L g810 ( 
.A1(n_753),
.A2(n_696),
.B(n_693),
.Y(n_810)
);

INVx2_ASAP7_75t_SL g811 ( 
.A(n_733),
.Y(n_811)
);

AND2x2_ASAP7_75t_L g812 ( 
.A(n_734),
.B(n_745),
.Y(n_812)
);

AND2x2_ASAP7_75t_L g813 ( 
.A(n_775),
.B(n_681),
.Y(n_813)
);

BUFx3_ASAP7_75t_L g814 ( 
.A(n_768),
.Y(n_814)
);

INVxp67_ASAP7_75t_L g815 ( 
.A(n_718),
.Y(n_815)
);

BUFx3_ASAP7_75t_L g816 ( 
.A(n_768),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_738),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_774),
.B(n_758),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_725),
.B(n_731),
.Y(n_819)
);

BUFx6f_ASAP7_75t_L g820 ( 
.A(n_765),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_729),
.B(n_709),
.Y(n_821)
);

AND2x2_ASAP7_75t_L g822 ( 
.A(n_729),
.B(n_709),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_738),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_753),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_761),
.B(n_658),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_761),
.B(n_644),
.Y(n_826)
);

AND2x2_ASAP7_75t_L g827 ( 
.A(n_724),
.B(n_590),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_730),
.Y(n_828)
);

INVx2_ASAP7_75t_SL g829 ( 
.A(n_723),
.Y(n_829)
);

AND2x2_ASAP7_75t_SL g830 ( 
.A(n_752),
.B(n_704),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_789),
.B(n_801),
.Y(n_831)
);

OAI21xp5_ASAP7_75t_L g832 ( 
.A1(n_771),
.A2(n_714),
.B(n_712),
.Y(n_832)
);

AND2x2_ASAP7_75t_L g833 ( 
.A(n_724),
.B(n_590),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_732),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_720),
.B(n_591),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_720),
.B(n_591),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_748),
.B(n_591),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_735),
.Y(n_838)
);

NOR2xp33_ASAP7_75t_L g839 ( 
.A(n_752),
.B(n_710),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_748),
.B(n_595),
.Y(n_840)
);

AND2x2_ASAP7_75t_L g841 ( 
.A(n_759),
.B(n_595),
.Y(n_841)
);

BUFx5_ASAP7_75t_L g842 ( 
.A(n_761),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_736),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_761),
.B(n_719),
.Y(n_844)
);

AND2x2_ASAP7_75t_L g845 ( 
.A(n_782),
.B(n_595),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_761),
.B(n_647),
.Y(n_846)
);

INVx2_ASAP7_75t_L g847 ( 
.A(n_747),
.Y(n_847)
);

INVx1_ASAP7_75t_SL g848 ( 
.A(n_742),
.Y(n_848)
);

AND2x2_ASAP7_75t_L g849 ( 
.A(n_782),
.B(n_595),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_762),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_737),
.Y(n_851)
);

INVx2_ASAP7_75t_L g852 ( 
.A(n_749),
.Y(n_852)
);

NAND2xp5_ASAP7_75t_L g853 ( 
.A(n_721),
.B(n_618),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_722),
.B(n_618),
.Y(n_854)
);

AND2x2_ASAP7_75t_L g855 ( 
.A(n_798),
.B(n_609),
.Y(n_855)
);

AND2x2_ASAP7_75t_SL g856 ( 
.A(n_790),
.B(n_704),
.Y(n_856)
);

INVx1_ASAP7_75t_L g857 ( 
.A(n_750),
.Y(n_857)
);

OAI21x1_ASAP7_75t_L g858 ( 
.A1(n_771),
.A2(n_471),
.B(n_418),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_751),
.Y(n_859)
);

INVx1_ASAP7_75t_L g860 ( 
.A(n_754),
.Y(n_860)
);

AND2x2_ASAP7_75t_L g861 ( 
.A(n_788),
.B(n_609),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_765),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_L g863 ( 
.A(n_744),
.B(n_618),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_801),
.B(n_618),
.Y(n_864)
);

INVx3_ASAP7_75t_L g865 ( 
.A(n_739),
.Y(n_865)
);

AND2x2_ASAP7_75t_L g866 ( 
.A(n_763),
.B(n_791),
.Y(n_866)
);

AND2x2_ASAP7_75t_L g867 ( 
.A(n_796),
.B(n_609),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_R g868 ( 
.A(n_726),
.B(n_586),
.Y(n_868)
);

INVxp67_ASAP7_75t_L g869 ( 
.A(n_781),
.Y(n_869)
);

NAND2x1p5_ASAP7_75t_L g870 ( 
.A(n_802),
.B(n_609),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_803),
.B(n_806),
.Y(n_871)
);

INVx4_ASAP7_75t_L g872 ( 
.A(n_744),
.Y(n_872)
);

AND2x2_ASAP7_75t_L g873 ( 
.A(n_784),
.B(n_611),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_755),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_784),
.B(n_611),
.Y(n_875)
);

AND2x2_ASAP7_75t_L g876 ( 
.A(n_760),
.B(n_611),
.Y(n_876)
);

HB1xp67_ASAP7_75t_L g877 ( 
.A(n_778),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_767),
.B(n_611),
.Y(n_878)
);

AND2x2_ASAP7_75t_L g879 ( 
.A(n_769),
.B(n_612),
.Y(n_879)
);

AND2x2_ASAP7_75t_L g880 ( 
.A(n_780),
.B(n_612),
.Y(n_880)
);

AND2x4_ASAP7_75t_L g881 ( 
.A(n_785),
.B(n_612),
.Y(n_881)
);

AND2x2_ASAP7_75t_L g882 ( 
.A(n_793),
.B(n_612),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_744),
.B(n_617),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_743),
.Y(n_884)
);

INVx3_ASAP7_75t_SL g885 ( 
.A(n_795),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_764),
.B(n_617),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_764),
.B(n_617),
.Y(n_887)
);

AND2x2_ASAP7_75t_L g888 ( 
.A(n_794),
.B(n_617),
.Y(n_888)
);

AND2x2_ASAP7_75t_L g889 ( 
.A(n_727),
.B(n_620),
.Y(n_889)
);

BUFx6f_ASAP7_75t_L g890 ( 
.A(n_746),
.Y(n_890)
);

AND2x4_ASAP7_75t_L g891 ( 
.A(n_776),
.B(n_620),
.Y(n_891)
);

INVx3_ASAP7_75t_L g892 ( 
.A(n_787),
.Y(n_892)
);

AND2x2_ASAP7_75t_SL g893 ( 
.A(n_804),
.B(n_620),
.Y(n_893)
);

INVx3_ASAP7_75t_L g894 ( 
.A(n_728),
.Y(n_894)
);

AND2x2_ASAP7_75t_L g895 ( 
.A(n_779),
.B(n_620),
.Y(n_895)
);

AND2x2_ASAP7_75t_L g896 ( 
.A(n_770),
.B(n_622),
.Y(n_896)
);

AND2x2_ASAP7_75t_L g897 ( 
.A(n_783),
.B(n_622),
.Y(n_897)
);

INVx1_ASAP7_75t_SL g898 ( 
.A(n_772),
.Y(n_898)
);

INVx4_ASAP7_75t_L g899 ( 
.A(n_744),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_744),
.B(n_622),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_SL g901 ( 
.A(n_757),
.B(n_622),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_786),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_756),
.B(n_741),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_777),
.B(n_471),
.Y(n_904)
);

BUFx2_ASAP7_75t_L g905 ( 
.A(n_807),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_828),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_SL g907 ( 
.A(n_848),
.B(n_586),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_818),
.B(n_792),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_SL g909 ( 
.A(n_850),
.B(n_800),
.Y(n_909)
);

INVx3_ASAP7_75t_L g910 ( 
.A(n_809),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_888),
.B(n_786),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_888),
.B(n_799),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_819),
.B(n_740),
.Y(n_913)
);

INVx2_ASAP7_75t_L g914 ( 
.A(n_852),
.Y(n_914)
);

NOR2x1_ASAP7_75t_L g915 ( 
.A(n_862),
.B(n_766),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_839),
.B(n_799),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_830),
.B(n_805),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_831),
.B(n_773),
.Y(n_918)
);

NAND2xp5_ASAP7_75t_L g919 ( 
.A(n_882),
.B(n_773),
.Y(n_919)
);

INVx4_ASAP7_75t_L g920 ( 
.A(n_809),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_855),
.Y(n_921)
);

BUFx6f_ASAP7_75t_L g922 ( 
.A(n_809),
.Y(n_922)
);

OR2x6_ASAP7_75t_L g923 ( 
.A(n_811),
.B(n_797),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_811),
.B(n_518),
.Y(n_924)
);

AND2x6_ASAP7_75t_L g925 ( 
.A(n_814),
.B(n_518),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_855),
.Y(n_926)
);

NAND2x1p5_ASAP7_75t_L g927 ( 
.A(n_862),
.B(n_517),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_850),
.Y(n_928)
);

INVx1_ASAP7_75t_L g929 ( 
.A(n_828),
.Y(n_929)
);

OAI21x1_ASAP7_75t_L g930 ( 
.A1(n_858),
.A2(n_471),
.B(n_69),
.Y(n_930)
);

NAND2x1p5_ASAP7_75t_L g931 ( 
.A(n_862),
.B(n_517),
.Y(n_931)
);

NOR2xp33_ASAP7_75t_SL g932 ( 
.A(n_830),
.B(n_471),
.Y(n_932)
);

INVx3_ASAP7_75t_L g933 ( 
.A(n_809),
.Y(n_933)
);

INVx1_ASAP7_75t_L g934 ( 
.A(n_834),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_815),
.B(n_68),
.Y(n_935)
);

CKINVDCx5p33_ASAP7_75t_R g936 ( 
.A(n_868),
.Y(n_936)
);

AND2x2_ASAP7_75t_L g937 ( 
.A(n_819),
.B(n_44),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_852),
.Y(n_938)
);

BUFx2_ASAP7_75t_L g939 ( 
.A(n_882),
.Y(n_939)
);

AND2x4_ASAP7_75t_L g940 ( 
.A(n_871),
.B(n_46),
.Y(n_940)
);

HB1xp67_ASAP7_75t_L g941 ( 
.A(n_829),
.Y(n_941)
);

AND2x2_ASAP7_75t_SL g942 ( 
.A(n_830),
.B(n_856),
.Y(n_942)
);

AND2x2_ASAP7_75t_L g943 ( 
.A(n_812),
.B(n_46),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_809),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_834),
.Y(n_945)
);

AND2x2_ASAP7_75t_L g946 ( 
.A(n_812),
.B(n_47),
.Y(n_946)
);

AND2x6_ASAP7_75t_L g947 ( 
.A(n_814),
.B(n_518),
.Y(n_947)
);

CKINVDCx20_ASAP7_75t_R g948 ( 
.A(n_885),
.Y(n_948)
);

INVx1_ASAP7_75t_L g949 ( 
.A(n_838),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_871),
.B(n_48),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_813),
.B(n_49),
.Y(n_951)
);

NOR2x1_ASAP7_75t_L g952 ( 
.A(n_872),
.B(n_518),
.Y(n_952)
);

INVx4_ASAP7_75t_L g953 ( 
.A(n_820),
.Y(n_953)
);

INVxp67_ASAP7_75t_L g954 ( 
.A(n_837),
.Y(n_954)
);

HB1xp67_ASAP7_75t_L g955 ( 
.A(n_829),
.Y(n_955)
);

BUFx4f_ASAP7_75t_L g956 ( 
.A(n_820),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_838),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_845),
.Y(n_958)
);

CKINVDCx20_ASAP7_75t_R g959 ( 
.A(n_885),
.Y(n_959)
);

OR2x2_ASAP7_75t_L g960 ( 
.A(n_898),
.B(n_49),
.Y(n_960)
);

NOR2x1_ASAP7_75t_SL g961 ( 
.A(n_872),
.B(n_528),
.Y(n_961)
);

INVx6_ASAP7_75t_SL g962 ( 
.A(n_891),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_843),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_845),
.Y(n_964)
);

INVx6_ASAP7_75t_L g965 ( 
.A(n_820),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_849),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_849),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_869),
.B(n_50),
.Y(n_968)
);

AND2x2_ASAP7_75t_L g969 ( 
.A(n_813),
.B(n_50),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_874),
.Y(n_970)
);

INVx2_ASAP7_75t_SL g971 ( 
.A(n_820),
.Y(n_971)
);

BUFx5_ASAP7_75t_L g972 ( 
.A(n_814),
.Y(n_972)
);

INVx5_ASAP7_75t_L g973 ( 
.A(n_820),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_846),
.B(n_517),
.Y(n_974)
);

OR2x6_ASAP7_75t_L g975 ( 
.A(n_821),
.B(n_528),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_824),
.B(n_52),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_866),
.B(n_52),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_824),
.B(n_53),
.Y(n_978)
);

AND2x4_ASAP7_75t_L g979 ( 
.A(n_866),
.B(n_872),
.Y(n_979)
);

HB1xp67_ASAP7_75t_L g980 ( 
.A(n_837),
.Y(n_980)
);

NAND2x1p5_ASAP7_75t_L g981 ( 
.A(n_816),
.B(n_517),
.Y(n_981)
);

INVx4_ASAP7_75t_L g982 ( 
.A(n_872),
.Y(n_982)
);

AND2x4_ASAP7_75t_L g983 ( 
.A(n_899),
.B(n_53),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_914),
.Y(n_984)
);

INVx4_ASAP7_75t_L g985 ( 
.A(n_956),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_906),
.Y(n_986)
);

INVx4_ASAP7_75t_L g987 ( 
.A(n_956),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_906),
.Y(n_988)
);

BUFx3_ASAP7_75t_L g989 ( 
.A(n_973),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_973),
.Y(n_990)
);

HB1xp67_ASAP7_75t_L g991 ( 
.A(n_905),
.Y(n_991)
);

INVx5_ASAP7_75t_SL g992 ( 
.A(n_983),
.Y(n_992)
);

CKINVDCx16_ASAP7_75t_R g993 ( 
.A(n_907),
.Y(n_993)
);

INVx1_ASAP7_75t_L g994 ( 
.A(n_929),
.Y(n_994)
);

AND2x2_ASAP7_75t_L g995 ( 
.A(n_942),
.B(n_856),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_938),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_929),
.Y(n_997)
);

BUFx2_ASAP7_75t_L g998 ( 
.A(n_928),
.Y(n_998)
);

BUFx2_ASAP7_75t_L g999 ( 
.A(n_948),
.Y(n_999)
);

BUFx2_ASAP7_75t_SL g1000 ( 
.A(n_959),
.Y(n_1000)
);

BUFx12f_ASAP7_75t_L g1001 ( 
.A(n_936),
.Y(n_1001)
);

BUFx12f_ASAP7_75t_L g1002 ( 
.A(n_960),
.Y(n_1002)
);

CKINVDCx20_ASAP7_75t_R g1003 ( 
.A(n_913),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_934),
.Y(n_1004)
);

BUFx12f_ASAP7_75t_L g1005 ( 
.A(n_968),
.Y(n_1005)
);

BUFx6f_ASAP7_75t_L g1006 ( 
.A(n_973),
.Y(n_1006)
);

INVx3_ASAP7_75t_L g1007 ( 
.A(n_982),
.Y(n_1007)
);

AND2x2_ASAP7_75t_L g1008 ( 
.A(n_909),
.B(n_856),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_964),
.B(n_835),
.Y(n_1009)
);

BUFx12f_ASAP7_75t_L g1010 ( 
.A(n_923),
.Y(n_1010)
);

BUFx2_ASAP7_75t_R g1011 ( 
.A(n_916),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_982),
.Y(n_1012)
);

AND2x2_ASAP7_75t_L g1013 ( 
.A(n_977),
.B(n_821),
.Y(n_1013)
);

INVx1_ASAP7_75t_SL g1014 ( 
.A(n_940),
.Y(n_1014)
);

BUFx12f_ASAP7_75t_L g1015 ( 
.A(n_923),
.Y(n_1015)
);

BUFx10_ASAP7_75t_L g1016 ( 
.A(n_983),
.Y(n_1016)
);

INVxp67_ASAP7_75t_SL g1017 ( 
.A(n_979),
.Y(n_1017)
);

INVx1_ASAP7_75t_SL g1018 ( 
.A(n_940),
.Y(n_1018)
);

INVx3_ASAP7_75t_L g1019 ( 
.A(n_922),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_962),
.Y(n_1020)
);

INVx4_ASAP7_75t_L g1021 ( 
.A(n_979),
.Y(n_1021)
);

CKINVDCx20_ASAP7_75t_R g1022 ( 
.A(n_917),
.Y(n_1022)
);

BUFx24_ASAP7_75t_L g1023 ( 
.A(n_950),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_932),
.B(n_825),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_934),
.Y(n_1025)
);

CKINVDCx5p33_ASAP7_75t_R g1026 ( 
.A(n_941),
.Y(n_1026)
);

INVx1_ASAP7_75t_SL g1027 ( 
.A(n_950),
.Y(n_1027)
);

INVx4_ASAP7_75t_L g1028 ( 
.A(n_922),
.Y(n_1028)
);

BUFx12f_ASAP7_75t_L g1029 ( 
.A(n_977),
.Y(n_1029)
);

CKINVDCx20_ASAP7_75t_R g1030 ( 
.A(n_955),
.Y(n_1030)
);

INVx1_ASAP7_75t_L g1031 ( 
.A(n_945),
.Y(n_1031)
);

INVx3_ASAP7_75t_L g1032 ( 
.A(n_922),
.Y(n_1032)
);

BUFx6f_ASAP7_75t_L g1033 ( 
.A(n_965),
.Y(n_1033)
);

INVx5_ASAP7_75t_L g1034 ( 
.A(n_925),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_970),
.Y(n_1035)
);

BUFx2_ASAP7_75t_SL g1036 ( 
.A(n_925),
.Y(n_1036)
);

INVx2_ASAP7_75t_SL g1037 ( 
.A(n_965),
.Y(n_1037)
);

AND2x4_ASAP7_75t_L g1038 ( 
.A(n_939),
.B(n_899),
.Y(n_1038)
);

INVxp67_ASAP7_75t_SL g1039 ( 
.A(n_958),
.Y(n_1039)
);

AND2x2_ASAP7_75t_L g1040 ( 
.A(n_966),
.B(n_899),
.Y(n_1040)
);

BUFx5_ASAP7_75t_L g1041 ( 
.A(n_925),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_972),
.Y(n_1042)
);

OR2x2_ASAP7_75t_L g1043 ( 
.A(n_975),
.B(n_808),
.Y(n_1043)
);

BUFx4_ASAP7_75t_SL g1044 ( 
.A(n_975),
.Y(n_1044)
);

NOR2x1_ASAP7_75t_L g1045 ( 
.A(n_920),
.B(n_899),
.Y(n_1045)
);

CKINVDCx20_ASAP7_75t_R g1046 ( 
.A(n_951),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_945),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_967),
.B(n_835),
.Y(n_1048)
);

INVx3_ASAP7_75t_L g1049 ( 
.A(n_920),
.Y(n_1049)
);

INVx2_ASAP7_75t_SL g1050 ( 
.A(n_1001),
.Y(n_1050)
);

INVx2_ASAP7_75t_SL g1051 ( 
.A(n_1001),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_986),
.Y(n_1052)
);

OAI22xp33_ASAP7_75t_L g1053 ( 
.A1(n_1023),
.A2(n_1018),
.B1(n_1027),
.B2(n_1014),
.Y(n_1053)
);

BUFx2_ASAP7_75t_SL g1054 ( 
.A(n_1030),
.Y(n_1054)
);

CKINVDCx20_ASAP7_75t_R g1055 ( 
.A(n_993),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_1024),
.B(n_949),
.Y(n_1056)
);

INVx1_ASAP7_75t_L g1057 ( 
.A(n_988),
.Y(n_1057)
);

INVx5_ASAP7_75t_SL g1058 ( 
.A(n_1006),
.Y(n_1058)
);

AOI22xp33_ASAP7_75t_L g1059 ( 
.A1(n_1024),
.A2(n_893),
.B1(n_885),
.B2(n_810),
.Y(n_1059)
);

BUFx3_ASAP7_75t_L g1060 ( 
.A(n_998),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_1008),
.A2(n_893),
.B1(n_826),
.B2(n_822),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_991),
.B(n_969),
.Y(n_1062)
);

OAI22xp33_ASAP7_75t_L g1063 ( 
.A1(n_1023),
.A2(n_908),
.B1(n_954),
.B2(n_980),
.Y(n_1063)
);

BUFx3_ASAP7_75t_L g1064 ( 
.A(n_1030),
.Y(n_1064)
);

AOI22xp33_ASAP7_75t_SL g1065 ( 
.A1(n_995),
.A2(n_822),
.B1(n_893),
.B2(n_842),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_994),
.Y(n_1066)
);

AOI22xp33_ASAP7_75t_L g1067 ( 
.A1(n_1002),
.A2(n_1046),
.B1(n_1003),
.B2(n_1015),
.Y(n_1067)
);

BUFx10_ASAP7_75t_L g1068 ( 
.A(n_1026),
.Y(n_1068)
);

OR2x2_ASAP7_75t_L g1069 ( 
.A(n_1013),
.B(n_1026),
.Y(n_1069)
);

INVx1_ASAP7_75t_L g1070 ( 
.A(n_997),
.Y(n_1070)
);

BUFx8_ASAP7_75t_L g1071 ( 
.A(n_999),
.Y(n_1071)
);

AOI22xp33_ASAP7_75t_L g1072 ( 
.A1(n_1002),
.A2(n_842),
.B1(n_874),
.B2(n_827),
.Y(n_1072)
);

AOI22xp33_ASAP7_75t_L g1073 ( 
.A1(n_1046),
.A2(n_842),
.B1(n_827),
.B2(n_833),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_984),
.Y(n_1074)
);

AOI22xp33_ASAP7_75t_L g1075 ( 
.A1(n_1003),
.A2(n_842),
.B1(n_833),
.B2(n_877),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_1004),
.Y(n_1076)
);

INVx1_ASAP7_75t_SL g1077 ( 
.A(n_1044),
.Y(n_1077)
);

AOI22xp33_ASAP7_75t_SL g1078 ( 
.A1(n_1029),
.A2(n_1022),
.B1(n_1010),
.B2(n_1015),
.Y(n_1078)
);

CKINVDCx20_ASAP7_75t_R g1079 ( 
.A(n_1022),
.Y(n_1079)
);

AOI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_1017),
.A2(n_1029),
.B1(n_1038),
.B2(n_1005),
.Y(n_1080)
);

INVxp67_ASAP7_75t_SL g1081 ( 
.A(n_1047),
.Y(n_1081)
);

INVx2_ASAP7_75t_SL g1082 ( 
.A(n_1010),
.Y(n_1082)
);

INVx6_ASAP7_75t_L g1083 ( 
.A(n_1016),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1025),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_1000),
.Y(n_1085)
);

OAI21xp5_ASAP7_75t_SL g1086 ( 
.A1(n_1011),
.A2(n_937),
.B(n_943),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_1031),
.Y(n_1087)
);

AOI22xp33_ASAP7_75t_L g1088 ( 
.A1(n_1005),
.A2(n_842),
.B1(n_844),
.B2(n_892),
.Y(n_1088)
);

INVx2_ASAP7_75t_L g1089 ( 
.A(n_984),
.Y(n_1089)
);

INVx6_ASAP7_75t_L g1090 ( 
.A(n_1016),
.Y(n_1090)
);

BUFx3_ASAP7_75t_L g1091 ( 
.A(n_1020),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_1047),
.Y(n_1092)
);

INVx3_ASAP7_75t_L g1093 ( 
.A(n_985),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_996),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_996),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_1038),
.A2(n_842),
.B1(n_892),
.B2(n_847),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_992),
.B(n_946),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_1035),
.Y(n_1098)
);

BUFx6f_ASAP7_75t_L g1099 ( 
.A(n_1006),
.Y(n_1099)
);

AOI22xp5_ASAP7_75t_L g1100 ( 
.A1(n_1038),
.A2(n_842),
.B1(n_957),
.B2(n_949),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_1035),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_1039),
.Y(n_1102)
);

BUFx12f_ASAP7_75t_L g1103 ( 
.A(n_1006),
.Y(n_1103)
);

CKINVDCx11_ASAP7_75t_R g1104 ( 
.A(n_1016),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_985),
.B(n_953),
.Y(n_1105)
);

INVx4_ASAP7_75t_L g1106 ( 
.A(n_985),
.Y(n_1106)
);

NAND2xp5_ASAP7_75t_L g1107 ( 
.A(n_1040),
.B(n_957),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_1048),
.Y(n_1108)
);

AOI22xp33_ASAP7_75t_L g1109 ( 
.A1(n_1043),
.A2(n_842),
.B1(n_892),
.B2(n_847),
.Y(n_1109)
);

AOI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1021),
.A2(n_842),
.B1(n_963),
.B2(n_840),
.Y(n_1110)
);

AOI22xp5_ASAP7_75t_L g1111 ( 
.A1(n_1021),
.A2(n_963),
.B1(n_840),
.B2(n_926),
.Y(n_1111)
);

AOI22xp33_ASAP7_75t_L g1112 ( 
.A1(n_1040),
.A2(n_892),
.B1(n_847),
.B2(n_836),
.Y(n_1112)
);

AOI22xp33_ASAP7_75t_SL g1113 ( 
.A1(n_992),
.A2(n_978),
.B1(n_976),
.B2(n_875),
.Y(n_1113)
);

BUFx4f_ASAP7_75t_SL g1114 ( 
.A(n_1033),
.Y(n_1114)
);

BUFx3_ASAP7_75t_L g1115 ( 
.A(n_1033),
.Y(n_1115)
);

AOI22xp33_ASAP7_75t_SL g1116 ( 
.A1(n_992),
.A2(n_1034),
.B1(n_1036),
.B2(n_875),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_1052),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_1069),
.B(n_1062),
.Y(n_1118)
);

AOI22xp33_ASAP7_75t_SL g1119 ( 
.A1(n_1059),
.A2(n_897),
.B1(n_1034),
.B2(n_832),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_1054),
.B(n_836),
.Y(n_1120)
);

INVx4_ASAP7_75t_L g1121 ( 
.A(n_1114),
.Y(n_1121)
);

AOI22xp33_ASAP7_75t_L g1122 ( 
.A1(n_1065),
.A2(n_864),
.B1(n_1009),
.B2(n_921),
.Y(n_1122)
);

CKINVDCx20_ASAP7_75t_R g1123 ( 
.A(n_1079),
.Y(n_1123)
);

AOI22xp33_ASAP7_75t_L g1124 ( 
.A1(n_1065),
.A2(n_884),
.B1(n_878),
.B2(n_879),
.Y(n_1124)
);

CKINVDCx6p67_ASAP7_75t_R g1125 ( 
.A(n_1077),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_1061),
.A2(n_884),
.B1(n_878),
.B2(n_879),
.Y(n_1126)
);

BUFx12f_ASAP7_75t_L g1127 ( 
.A(n_1068),
.Y(n_1127)
);

OAI22xp5_ASAP7_75t_L g1128 ( 
.A1(n_1111),
.A2(n_1086),
.B1(n_1113),
.B2(n_1056),
.Y(n_1128)
);

OAI22xp5_ASAP7_75t_L g1129 ( 
.A1(n_1086),
.A2(n_1021),
.B1(n_903),
.B2(n_911),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1064),
.B(n_891),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_1102),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1108),
.B(n_876),
.Y(n_1132)
);

AOI22xp33_ASAP7_75t_L g1133 ( 
.A1(n_1113),
.A2(n_876),
.B1(n_857),
.B2(n_860),
.Y(n_1133)
);

AOI22xp33_ASAP7_75t_L g1134 ( 
.A1(n_1063),
.A2(n_857),
.B1(n_860),
.B2(n_859),
.Y(n_1134)
);

OAI22xp33_ASAP7_75t_L g1135 ( 
.A1(n_1080),
.A2(n_912),
.B1(n_1034),
.B2(n_987),
.Y(n_1135)
);

BUFx2_ASAP7_75t_L g1136 ( 
.A(n_1060),
.Y(n_1136)
);

OAI21xp33_ASAP7_75t_L g1137 ( 
.A1(n_1056),
.A2(n_841),
.B(n_873),
.Y(n_1137)
);

AND2x2_ASAP7_75t_L g1138 ( 
.A(n_1097),
.B(n_891),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_1057),
.Y(n_1139)
);

AOI22xp33_ASAP7_75t_L g1140 ( 
.A1(n_1078),
.A2(n_859),
.B1(n_881),
.B2(n_897),
.Y(n_1140)
);

HB1xp67_ASAP7_75t_L g1141 ( 
.A(n_1066),
.Y(n_1141)
);

OAI22xp33_ASAP7_75t_L g1142 ( 
.A1(n_1077),
.A2(n_1034),
.B1(n_987),
.B2(n_962),
.Y(n_1142)
);

AOI22xp33_ASAP7_75t_L g1143 ( 
.A1(n_1078),
.A2(n_881),
.B1(n_843),
.B2(n_873),
.Y(n_1143)
);

AOI22xp33_ASAP7_75t_SL g1144 ( 
.A1(n_1055),
.A2(n_1034),
.B1(n_886),
.B2(n_887),
.Y(n_1144)
);

OAI22xp5_ASAP7_75t_L g1145 ( 
.A1(n_1073),
.A2(n_865),
.B1(n_851),
.B2(n_987),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_1070),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1076),
.Y(n_1147)
);

INVx2_ASAP7_75t_L g1148 ( 
.A(n_1092),
.Y(n_1148)
);

AOI22xp33_ASAP7_75t_L g1149 ( 
.A1(n_1053),
.A2(n_881),
.B1(n_880),
.B2(n_890),
.Y(n_1149)
);

CKINVDCx11_ASAP7_75t_R g1150 ( 
.A(n_1068),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1084),
.Y(n_1151)
);

OAI222xp33_ASAP7_75t_L g1152 ( 
.A1(n_1075),
.A2(n_924),
.B1(n_883),
.B2(n_900),
.C1(n_851),
.C2(n_881),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_1085),
.Y(n_1153)
);

INVx3_ASAP7_75t_L g1154 ( 
.A(n_1099),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1087),
.Y(n_1155)
);

AND2x2_ASAP7_75t_L g1156 ( 
.A(n_1115),
.B(n_1067),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_SL g1157 ( 
.A1(n_1116),
.A2(n_887),
.B(n_886),
.Y(n_1157)
);

AOI22xp33_ASAP7_75t_L g1158 ( 
.A1(n_1072),
.A2(n_880),
.B1(n_890),
.B2(n_896),
.Y(n_1158)
);

HB1xp67_ASAP7_75t_SL g1159 ( 
.A(n_1071),
.Y(n_1159)
);

INVx3_ASAP7_75t_L g1160 ( 
.A(n_1099),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_1107),
.B(n_1081),
.Y(n_1161)
);

CKINVDCx8_ASAP7_75t_R g1162 ( 
.A(n_1099),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1107),
.A2(n_890),
.B1(n_896),
.B2(n_902),
.Y(n_1163)
);

OAI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1100),
.A2(n_924),
.B1(n_935),
.B2(n_816),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1074),
.Y(n_1165)
);

CKINVDCx5p33_ASAP7_75t_R g1166 ( 
.A(n_1071),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_1089),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1093),
.B(n_989),
.Y(n_1168)
);

BUFx4f_ASAP7_75t_SL g1169 ( 
.A(n_1103),
.Y(n_1169)
);

INVx4_ASAP7_75t_L g1170 ( 
.A(n_1104),
.Y(n_1170)
);

AOI222xp33_ASAP7_75t_L g1171 ( 
.A1(n_1081),
.A2(n_867),
.B1(n_861),
.B2(n_895),
.C1(n_891),
.C2(n_841),
.Y(n_1171)
);

INVx2_ASAP7_75t_L g1172 ( 
.A(n_1095),
.Y(n_1172)
);

AND2x2_ASAP7_75t_L g1173 ( 
.A(n_1082),
.B(n_895),
.Y(n_1173)
);

OAI22xp5_ASAP7_75t_L g1174 ( 
.A1(n_1110),
.A2(n_865),
.B1(n_817),
.B2(n_823),
.Y(n_1174)
);

OAI22xp5_ASAP7_75t_L g1175 ( 
.A1(n_1112),
.A2(n_865),
.B1(n_817),
.B2(n_823),
.Y(n_1175)
);

BUFx3_ASAP7_75t_L g1176 ( 
.A(n_1083),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_1094),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1058),
.B(n_1033),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1106),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1098),
.A2(n_890),
.B1(n_902),
.B2(n_867),
.Y(n_1180)
);

CKINVDCx6p67_ASAP7_75t_R g1181 ( 
.A(n_1091),
.Y(n_1181)
);

AOI22xp5_ASAP7_75t_L g1182 ( 
.A1(n_1083),
.A2(n_861),
.B1(n_816),
.B2(n_915),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_1090),
.Y(n_1183)
);

AOI22xp33_ASAP7_75t_L g1184 ( 
.A1(n_1101),
.A2(n_890),
.B1(n_919),
.B2(n_974),
.Y(n_1184)
);

CKINVDCx11_ASAP7_75t_R g1185 ( 
.A(n_1106),
.Y(n_1185)
);

AOI22xp5_ASAP7_75t_L g1186 ( 
.A1(n_1128),
.A2(n_1116),
.B1(n_1050),
.B2(n_1051),
.Y(n_1186)
);

AOI22xp33_ASAP7_75t_SL g1187 ( 
.A1(n_1129),
.A2(n_1090),
.B1(n_1041),
.B2(n_1058),
.Y(n_1187)
);

AOI22xp33_ASAP7_75t_L g1188 ( 
.A1(n_1119),
.A2(n_894),
.B1(n_1088),
.B2(n_865),
.Y(n_1188)
);

AOI22xp33_ASAP7_75t_L g1189 ( 
.A1(n_1124),
.A2(n_894),
.B1(n_1109),
.B2(n_889),
.Y(n_1189)
);

NAND2xp5_ASAP7_75t_L g1190 ( 
.A(n_1141),
.B(n_1058),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_1131),
.B(n_1093),
.Y(n_1191)
);

AOI22xp5_ASAP7_75t_L g1192 ( 
.A1(n_1143),
.A2(n_1096),
.B1(n_1037),
.B2(n_863),
.Y(n_1192)
);

AOI22xp33_ASAP7_75t_L g1193 ( 
.A1(n_1124),
.A2(n_894),
.B1(n_889),
.B2(n_918),
.Y(n_1193)
);

OAI22xp5_ASAP7_75t_L g1194 ( 
.A1(n_1133),
.A2(n_1007),
.B1(n_1012),
.B2(n_1105),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_L g1195 ( 
.A1(n_1156),
.A2(n_901),
.B1(n_972),
.B2(n_904),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1118),
.B(n_1019),
.Y(n_1196)
);

OAI221xp5_ASAP7_75t_L g1197 ( 
.A1(n_1133),
.A2(n_853),
.B1(n_894),
.B2(n_854),
.C(n_1037),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1117),
.Y(n_1198)
);

OAI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1134),
.A2(n_1007),
.B1(n_1012),
.B2(n_1105),
.Y(n_1199)
);

AOI22xp33_ASAP7_75t_SL g1200 ( 
.A1(n_1120),
.A2(n_1041),
.B1(n_972),
.B2(n_925),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1139),
.Y(n_1201)
);

AOI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_1143),
.A2(n_947),
.B1(n_972),
.B2(n_1041),
.Y(n_1202)
);

AOI22xp33_ASAP7_75t_L g1203 ( 
.A1(n_1137),
.A2(n_972),
.B1(n_947),
.B2(n_952),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1134),
.A2(n_947),
.B1(n_1041),
.B2(n_870),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1144),
.A2(n_947),
.B1(n_1041),
.B2(n_870),
.Y(n_1205)
);

AOI22xp5_ASAP7_75t_L g1206 ( 
.A1(n_1140),
.A2(n_1157),
.B1(n_1171),
.B2(n_1122),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_SL g1207 ( 
.A1(n_1132),
.A2(n_1041),
.B1(n_930),
.B2(n_961),
.Y(n_1207)
);

OAI222xp33_ASAP7_75t_L g1208 ( 
.A1(n_1122),
.A2(n_870),
.B1(n_981),
.B2(n_1028),
.C1(n_1032),
.C2(n_1019),
.Y(n_1208)
);

INVxp67_ASAP7_75t_L g1209 ( 
.A(n_1136),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1126),
.A2(n_1041),
.B1(n_1045),
.B2(n_989),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1126),
.A2(n_990),
.B1(n_1033),
.B2(n_933),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1149),
.A2(n_990),
.B1(n_933),
.B2(n_944),
.Y(n_1212)
);

INVx2_ASAP7_75t_SL g1213 ( 
.A(n_1181),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1146),
.B(n_1019),
.Y(n_1214)
);

AOI22xp33_ASAP7_75t_L g1215 ( 
.A1(n_1149),
.A2(n_944),
.B1(n_910),
.B2(n_1032),
.Y(n_1215)
);

OAI222xp33_ASAP7_75t_L g1216 ( 
.A1(n_1140),
.A2(n_1028),
.B1(n_1032),
.B2(n_1042),
.C1(n_1049),
.C2(n_971),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_SL g1217 ( 
.A1(n_1138),
.A2(n_961),
.B1(n_858),
.B2(n_1006),
.Y(n_1217)
);

AOI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1173),
.A2(n_910),
.B1(n_1042),
.B2(n_1049),
.Y(n_1218)
);

AOI22xp33_ASAP7_75t_L g1219 ( 
.A1(n_1163),
.A2(n_953),
.B1(n_1042),
.B2(n_1049),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_SL g1220 ( 
.A1(n_1161),
.A2(n_1028),
.B(n_931),
.Y(n_1220)
);

OAI222xp33_ASAP7_75t_L g1221 ( 
.A1(n_1182),
.A2(n_1177),
.B1(n_1172),
.B2(n_1167),
.C1(n_1165),
.C2(n_1155),
.Y(n_1221)
);

AOI22xp33_ASAP7_75t_L g1222 ( 
.A1(n_1130),
.A2(n_1012),
.B1(n_1007),
.B2(n_927),
.Y(n_1222)
);

CKINVDCx11_ASAP7_75t_R g1223 ( 
.A(n_1123),
.Y(n_1223)
);

OAI22xp5_ASAP7_75t_L g1224 ( 
.A1(n_1159),
.A2(n_54),
.B1(n_55),
.B2(n_56),
.Y(n_1224)
);

NAND3xp33_ASAP7_75t_SL g1225 ( 
.A(n_1166),
.B(n_55),
.C(n_56),
.Y(n_1225)
);

NAND3xp33_ASAP7_75t_L g1226 ( 
.A(n_1147),
.B(n_540),
.C(n_528),
.Y(n_1226)
);

AOI22xp33_ASAP7_75t_L g1227 ( 
.A1(n_1148),
.A2(n_528),
.B1(n_571),
.B2(n_570),
.Y(n_1227)
);

OAI221xp5_ASAP7_75t_L g1228 ( 
.A1(n_1163),
.A2(n_57),
.B1(n_58),
.B2(n_61),
.C(n_62),
.Y(n_1228)
);

AOI22xp33_ASAP7_75t_SL g1229 ( 
.A1(n_1151),
.A2(n_574),
.B1(n_540),
.B2(n_571),
.Y(n_1229)
);

OAI222xp33_ASAP7_75t_L g1230 ( 
.A1(n_1165),
.A2(n_57),
.B1(n_62),
.B2(n_63),
.C1(n_64),
.C2(n_65),
.Y(n_1230)
);

AOI22xp33_ASAP7_75t_L g1231 ( 
.A1(n_1180),
.A2(n_1158),
.B1(n_1175),
.B2(n_1164),
.Y(n_1231)
);

AND2x2_ASAP7_75t_L g1232 ( 
.A(n_1183),
.B(n_65),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1176),
.B(n_66),
.Y(n_1233)
);

OAI21xp33_ASAP7_75t_L g1234 ( 
.A1(n_1174),
.A2(n_66),
.B(n_574),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1148),
.B(n_540),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1145),
.A2(n_574),
.B1(n_540),
.B2(n_571),
.Y(n_1236)
);

AOI22xp33_ASAP7_75t_L g1237 ( 
.A1(n_1180),
.A2(n_574),
.B1(n_549),
.B2(n_571),
.Y(n_1237)
);

AND2x2_ASAP7_75t_L g1238 ( 
.A(n_1176),
.B(n_70),
.Y(n_1238)
);

AOI22xp33_ASAP7_75t_L g1239 ( 
.A1(n_1158),
.A2(n_549),
.B1(n_570),
.B2(n_550),
.Y(n_1239)
);

OAI22xp5_ASAP7_75t_L g1240 ( 
.A1(n_1125),
.A2(n_549),
.B1(n_570),
.B2(n_550),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1167),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_SL g1242 ( 
.A1(n_1170),
.A2(n_549),
.B1(n_570),
.B2(n_550),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1154),
.B(n_71),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1170),
.A2(n_550),
.B1(n_572),
.B2(n_545),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1135),
.A2(n_572),
.B1(n_545),
.B2(n_542),
.Y(n_1245)
);

OAI22xp5_ASAP7_75t_L g1246 ( 
.A1(n_1169),
.A2(n_572),
.B1(n_545),
.B2(n_542),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1184),
.A2(n_572),
.B(n_545),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1172),
.Y(n_1248)
);

NAND2xp5_ASAP7_75t_L g1249 ( 
.A(n_1168),
.B(n_1154),
.Y(n_1249)
);

OAI22xp5_ASAP7_75t_L g1250 ( 
.A1(n_1169),
.A2(n_1121),
.B1(n_1127),
.B2(n_1179),
.Y(n_1250)
);

OAI222xp33_ASAP7_75t_L g1251 ( 
.A1(n_1142),
.A2(n_1184),
.B1(n_1162),
.B2(n_1178),
.C1(n_1121),
.C2(n_1160),
.Y(n_1251)
);

AOI22xp33_ASAP7_75t_L g1252 ( 
.A1(n_1127),
.A2(n_542),
.B1(n_541),
.B2(n_532),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1209),
.B(n_1160),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1198),
.B(n_1168),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_L g1255 ( 
.A1(n_1206),
.A2(n_1150),
.B1(n_1185),
.B2(n_1153),
.Y(n_1255)
);

NAND2xp5_ASAP7_75t_L g1256 ( 
.A(n_1201),
.B(n_1179),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1186),
.B(n_1179),
.Y(n_1257)
);

NAND3xp33_ASAP7_75t_L g1258 ( 
.A(n_1228),
.B(n_1179),
.C(n_542),
.Y(n_1258)
);

NAND2xp33_ASAP7_75t_L g1259 ( 
.A(n_1234),
.B(n_1250),
.Y(n_1259)
);

AND2x2_ASAP7_75t_L g1260 ( 
.A(n_1196),
.B(n_72),
.Y(n_1260)
);

AND2x2_ASAP7_75t_L g1261 ( 
.A(n_1190),
.B(n_75),
.Y(n_1261)
);

NOR3xp33_ASAP7_75t_L g1262 ( 
.A(n_1225),
.B(n_1152),
.C(n_78),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1221),
.A2(n_76),
.B(n_81),
.Y(n_1263)
);

OAI21xp33_ASAP7_75t_L g1264 ( 
.A1(n_1224),
.A2(n_83),
.B(n_86),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1191),
.B(n_87),
.Y(n_1265)
);

NOR3xp33_ASAP7_75t_L g1266 ( 
.A(n_1230),
.B(n_89),
.C(n_91),
.Y(n_1266)
);

NAND4xp25_ASAP7_75t_L g1267 ( 
.A(n_1232),
.B(n_93),
.C(n_94),
.D(n_99),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1233),
.B(n_100),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1241),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_L g1270 ( 
.A(n_1214),
.B(n_101),
.Y(n_1270)
);

OAI22xp5_ASAP7_75t_L g1271 ( 
.A1(n_1231),
.A2(n_541),
.B1(n_532),
.B2(n_521),
.Y(n_1271)
);

OAI22xp5_ASAP7_75t_L g1272 ( 
.A1(n_1231),
.A2(n_541),
.B1(n_532),
.B2(n_521),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1249),
.B(n_103),
.Y(n_1273)
);

NAND3xp33_ASAP7_75t_L g1274 ( 
.A(n_1244),
.B(n_541),
.C(n_532),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1188),
.A2(n_521),
.B1(n_107),
.B2(n_109),
.Y(n_1275)
);

NAND2xp5_ASAP7_75t_L g1276 ( 
.A(n_1187),
.B(n_104),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1213),
.B(n_112),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_SL g1278 ( 
.A(n_1217),
.B(n_521),
.Y(n_1278)
);

OAI22xp5_ASAP7_75t_L g1279 ( 
.A1(n_1188),
.A2(n_1193),
.B1(n_1218),
.B2(n_1211),
.Y(n_1279)
);

OAI221xp5_ASAP7_75t_L g1280 ( 
.A1(n_1193),
.A2(n_113),
.B1(n_117),
.B2(n_121),
.C(n_124),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1238),
.B(n_125),
.Y(n_1281)
);

NAND3xp33_ASAP7_75t_L g1282 ( 
.A(n_1244),
.B(n_126),
.C(n_130),
.Y(n_1282)
);

NAND2xp5_ASAP7_75t_L g1283 ( 
.A(n_1220),
.B(n_323),
.Y(n_1283)
);

NAND2xp5_ASAP7_75t_L g1284 ( 
.A(n_1235),
.B(n_131),
.Y(n_1284)
);

OAI221xp5_ASAP7_75t_L g1285 ( 
.A1(n_1197),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.C(n_141),
.Y(n_1285)
);

AND2x2_ASAP7_75t_L g1286 ( 
.A(n_1243),
.B(n_320),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1189),
.A2(n_146),
.B1(n_147),
.B2(n_148),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1189),
.A2(n_1202),
.B1(n_1212),
.B2(n_1215),
.Y(n_1288)
);

NAND3xp33_ASAP7_75t_L g1289 ( 
.A(n_1194),
.B(n_151),
.C(n_153),
.Y(n_1289)
);

AND2x2_ASAP7_75t_L g1290 ( 
.A(n_1223),
.B(n_319),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1199),
.B(n_154),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_L g1292 ( 
.A(n_1248),
.B(n_314),
.Y(n_1292)
);

NOR3xp33_ASAP7_75t_L g1293 ( 
.A(n_1251),
.B(n_159),
.C(n_161),
.Y(n_1293)
);

AOI22xp33_ASAP7_75t_L g1294 ( 
.A1(n_1239),
.A2(n_164),
.B1(n_166),
.B2(n_167),
.Y(n_1294)
);

OAI221xp5_ASAP7_75t_L g1295 ( 
.A1(n_1222),
.A2(n_169),
.B1(n_171),
.B2(n_172),
.C(n_173),
.Y(n_1295)
);

AND2x2_ASAP7_75t_L g1296 ( 
.A(n_1219),
.B(n_311),
.Y(n_1296)
);

NOR3xp33_ASAP7_75t_SL g1297 ( 
.A(n_1216),
.B(n_174),
.C(n_175),
.Y(n_1297)
);

OAI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1210),
.A2(n_178),
.B1(n_179),
.B2(n_180),
.Y(n_1298)
);

NAND3xp33_ASAP7_75t_L g1299 ( 
.A(n_1195),
.B(n_181),
.C(n_186),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1219),
.B(n_310),
.Y(n_1300)
);

AOI211xp5_ASAP7_75t_L g1301 ( 
.A1(n_1208),
.A2(n_187),
.B(n_189),
.C(n_193),
.Y(n_1301)
);

NAND2xp5_ASAP7_75t_L g1302 ( 
.A(n_1192),
.B(n_309),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1263),
.B(n_1278),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1269),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1254),
.B(n_1207),
.Y(n_1305)
);

AND2x2_ASAP7_75t_L g1306 ( 
.A(n_1256),
.B(n_1245),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1290),
.B(n_1246),
.Y(n_1307)
);

NAND3xp33_ASAP7_75t_L g1308 ( 
.A(n_1259),
.B(n_1245),
.C(n_1239),
.Y(n_1308)
);

NOR2xp33_ASAP7_75t_L g1309 ( 
.A(n_1253),
.B(n_1200),
.Y(n_1309)
);

AND2x2_ASAP7_75t_L g1310 ( 
.A(n_1278),
.B(n_1261),
.Y(n_1310)
);

NAND4xp75_ASAP7_75t_L g1311 ( 
.A(n_1257),
.B(n_1247),
.C(n_1205),
.D(n_1204),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1292),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1260),
.B(n_1203),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1257),
.B(n_1236),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1266),
.A2(n_1240),
.B1(n_1237),
.B2(n_1226),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1263),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1263),
.Y(n_1317)
);

AO21x2_ASAP7_75t_L g1318 ( 
.A1(n_1302),
.A2(n_1229),
.B(n_1227),
.Y(n_1318)
);

NAND4xp75_ASAP7_75t_L g1319 ( 
.A(n_1297),
.B(n_1252),
.C(n_1242),
.D(n_1237),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1259),
.B(n_205),
.C(n_208),
.Y(n_1320)
);

NOR2xp33_ASAP7_75t_L g1321 ( 
.A(n_1267),
.B(n_212),
.Y(n_1321)
);

AND4x1_ASAP7_75t_L g1322 ( 
.A(n_1255),
.B(n_216),
.C(n_219),
.D(n_222),
.Y(n_1322)
);

NAND3xp33_ASAP7_75t_L g1323 ( 
.A(n_1262),
.B(n_224),
.C(n_227),
.Y(n_1323)
);

NOR2xp33_ASAP7_75t_L g1324 ( 
.A(n_1277),
.B(n_228),
.Y(n_1324)
);

INVx2_ASAP7_75t_L g1325 ( 
.A(n_1270),
.Y(n_1325)
);

AND2x2_ASAP7_75t_L g1326 ( 
.A(n_1255),
.B(n_232),
.Y(n_1326)
);

INVx2_ASAP7_75t_SL g1327 ( 
.A(n_1265),
.Y(n_1327)
);

NOR3xp33_ASAP7_75t_L g1328 ( 
.A(n_1258),
.B(n_233),
.C(n_238),
.Y(n_1328)
);

OA21x2_ASAP7_75t_L g1329 ( 
.A1(n_1291),
.A2(n_240),
.B(n_243),
.Y(n_1329)
);

AO21x2_ASAP7_75t_L g1330 ( 
.A1(n_1293),
.A2(n_246),
.B(n_248),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_L g1331 ( 
.A(n_1268),
.B(n_260),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_L g1332 ( 
.A(n_1297),
.B(n_262),
.C(n_263),
.Y(n_1332)
);

HB1xp67_ASAP7_75t_L g1333 ( 
.A(n_1304),
.Y(n_1333)
);

AND2x2_ASAP7_75t_L g1334 ( 
.A(n_1327),
.B(n_1300),
.Y(n_1334)
);

NAND4xp75_ASAP7_75t_SL g1335 ( 
.A(n_1329),
.B(n_1296),
.C(n_1286),
.D(n_1264),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1327),
.B(n_1273),
.Y(n_1336)
);

NAND4xp75_ASAP7_75t_SL g1337 ( 
.A(n_1329),
.B(n_1301),
.C(n_1289),
.D(n_1285),
.Y(n_1337)
);

NOR2x1_ASAP7_75t_L g1338 ( 
.A(n_1325),
.B(n_1283),
.Y(n_1338)
);

OR2x2_ASAP7_75t_L g1339 ( 
.A(n_1304),
.B(n_1279),
.Y(n_1339)
);

INVxp67_ASAP7_75t_SL g1340 ( 
.A(n_1325),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1312),
.Y(n_1341)
);

OA22x2_ASAP7_75t_L g1342 ( 
.A1(n_1310),
.A2(n_1288),
.B1(n_1271),
.B2(n_1272),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1312),
.B(n_1276),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1306),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1306),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1310),
.B(n_1281),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1309),
.B(n_1284),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1305),
.Y(n_1348)
);

INVx3_ASAP7_75t_L g1349 ( 
.A(n_1316),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1317),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1317),
.B(n_1299),
.Y(n_1351)
);

INVxp67_ASAP7_75t_SL g1352 ( 
.A(n_1303),
.Y(n_1352)
);

HB1xp67_ASAP7_75t_L g1353 ( 
.A(n_1316),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1344),
.B(n_1307),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1345),
.B(n_1303),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1341),
.Y(n_1356)
);

INVx1_ASAP7_75t_SL g1357 ( 
.A(n_1346),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1339),
.Y(n_1358)
);

XNOR2xp5_ASAP7_75t_L g1359 ( 
.A(n_1335),
.B(n_1322),
.Y(n_1359)
);

XOR2x2_ASAP7_75t_L g1360 ( 
.A(n_1342),
.B(n_1337),
.Y(n_1360)
);

XNOR2xp5_ASAP7_75t_L g1361 ( 
.A(n_1342),
.B(n_1322),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1339),
.Y(n_1362)
);

INVx1_ASAP7_75t_SL g1363 ( 
.A(n_1346),
.Y(n_1363)
);

INVx1_ASAP7_75t_SL g1364 ( 
.A(n_1334),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1350),
.Y(n_1365)
);

INVx2_ASAP7_75t_L g1366 ( 
.A(n_1349),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1342),
.A2(n_1308),
.B1(n_1330),
.B2(n_1320),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1356),
.Y(n_1368)
);

NAND2xp5_ASAP7_75t_L g1369 ( 
.A(n_1357),
.B(n_1350),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1361),
.A2(n_1347),
.B1(n_1330),
.B2(n_1348),
.Y(n_1370)
);

INVx2_ASAP7_75t_SL g1371 ( 
.A(n_1363),
.Y(n_1371)
);

INVx2_ASAP7_75t_L g1372 ( 
.A(n_1365),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1360),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1364),
.Y(n_1374)
);

AO22x2_ASAP7_75t_L g1375 ( 
.A1(n_1358),
.A2(n_1351),
.B1(n_1352),
.B2(n_1343),
.Y(n_1375)
);

OAI22x1_ASAP7_75t_L g1376 ( 
.A1(n_1361),
.A2(n_1334),
.B1(n_1303),
.B2(n_1338),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1362),
.Y(n_1377)
);

INVxp67_ASAP7_75t_L g1378 ( 
.A(n_1360),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1354),
.Y(n_1379)
);

BUFx3_ASAP7_75t_L g1380 ( 
.A(n_1359),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1355),
.Y(n_1381)
);

XOR2x2_ASAP7_75t_L g1382 ( 
.A(n_1367),
.B(n_1311),
.Y(n_1382)
);

OAI22xp5_ASAP7_75t_L g1383 ( 
.A1(n_1366),
.A2(n_1351),
.B1(n_1320),
.B2(n_1308),
.Y(n_1383)
);

INVx3_ASAP7_75t_L g1384 ( 
.A(n_1366),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1360),
.Y(n_1385)
);

OAI322xp33_ASAP7_75t_L g1386 ( 
.A1(n_1378),
.A2(n_1383),
.A3(n_1373),
.B1(n_1385),
.B2(n_1370),
.C1(n_1379),
.C2(n_1377),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_1368),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1372),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1369),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1369),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1374),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1378),
.A2(n_1332),
.B1(n_1330),
.B2(n_1319),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1384),
.Y(n_1393)
);

INVx3_ASAP7_75t_L g1394 ( 
.A(n_1384),
.Y(n_1394)
);

INVx1_ASAP7_75t_L g1395 ( 
.A(n_1371),
.Y(n_1395)
);

AOI322xp5_ASAP7_75t_L g1396 ( 
.A1(n_1373),
.A2(n_1385),
.A3(n_1380),
.B1(n_1382),
.B2(n_1375),
.C1(n_1353),
.C2(n_1383),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1387),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1388),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1394),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1389),
.Y(n_1400)
);

INVx2_ASAP7_75t_SL g1401 ( 
.A(n_1395),
.Y(n_1401)
);

OA22x2_ASAP7_75t_L g1402 ( 
.A1(n_1392),
.A2(n_1376),
.B1(n_1381),
.B2(n_1375),
.Y(n_1402)
);

OAI322xp33_ASAP7_75t_L g1403 ( 
.A1(n_1390),
.A2(n_1375),
.A3(n_1321),
.B1(n_1349),
.B2(n_1336),
.C1(n_1326),
.C2(n_1323),
.Y(n_1403)
);

AOI221xp5_ASAP7_75t_L g1404 ( 
.A1(n_1386),
.A2(n_1380),
.B1(n_1349),
.B2(n_1332),
.C(n_1326),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1391),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1393),
.Y(n_1406)
);

OAI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1402),
.A2(n_1392),
.B1(n_1396),
.B2(n_1394),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1397),
.Y(n_1408)
);

AOI22xp5_ASAP7_75t_L g1409 ( 
.A1(n_1404),
.A2(n_1329),
.B1(n_1311),
.B2(n_1331),
.Y(n_1409)
);

INVxp67_ASAP7_75t_SL g1410 ( 
.A(n_1401),
.Y(n_1410)
);

INVx2_ASAP7_75t_L g1411 ( 
.A(n_1399),
.Y(n_1411)
);

HB1xp67_ASAP7_75t_L g1412 ( 
.A(n_1397),
.Y(n_1412)
);

AOI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1405),
.A2(n_1329),
.B1(n_1319),
.B2(n_1313),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1410),
.B(n_1406),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1412),
.Y(n_1415)
);

AO22x2_ASAP7_75t_L g1416 ( 
.A1(n_1408),
.A2(n_1398),
.B1(n_1400),
.B2(n_1403),
.Y(n_1416)
);

AO22x2_ASAP7_75t_L g1417 ( 
.A1(n_1411),
.A2(n_1328),
.B1(n_1287),
.B2(n_1314),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1407),
.Y(n_1418)
);

INVx2_ASAP7_75t_SL g1419 ( 
.A(n_1409),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1413),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1412),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_1415),
.Y(n_1422)
);

AOI22xp5_ASAP7_75t_L g1423 ( 
.A1(n_1416),
.A2(n_1324),
.B1(n_1313),
.B2(n_1314),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1421),
.B(n_1333),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1414),
.Y(n_1425)
);

INVxp67_ASAP7_75t_L g1426 ( 
.A(n_1419),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1417),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1416),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1428),
.Y(n_1429)
);

NOR2x1p5_ASAP7_75t_L g1430 ( 
.A(n_1425),
.B(n_1418),
.Y(n_1430)
);

AOI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1423),
.A2(n_1417),
.B(n_1420),
.Y(n_1431)
);

NOR2x1_ASAP7_75t_L g1432 ( 
.A(n_1422),
.B(n_1280),
.Y(n_1432)
);

OAI22x1_ASAP7_75t_L g1433 ( 
.A1(n_1426),
.A2(n_1340),
.B1(n_1282),
.B2(n_1274),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1429),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1430),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1432),
.Y(n_1436)
);

INVx1_ASAP7_75t_L g1437 ( 
.A(n_1431),
.Y(n_1437)
);

AOI22xp5_ASAP7_75t_L g1438 ( 
.A1(n_1433),
.A2(n_1427),
.B1(n_1424),
.B2(n_1275),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1429),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1429),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1429),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1435),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1435),
.Y(n_1443)
);

OAI22xp5_ASAP7_75t_L g1444 ( 
.A1(n_1434),
.A2(n_1424),
.B1(n_1275),
.B2(n_1315),
.Y(n_1444)
);

OAI22xp5_ASAP7_75t_L g1445 ( 
.A1(n_1439),
.A2(n_1295),
.B1(n_1294),
.B2(n_1298),
.Y(n_1445)
);

OAI22xp5_ASAP7_75t_SL g1446 ( 
.A1(n_1436),
.A2(n_1294),
.B1(n_1318),
.B2(n_268),
.Y(n_1446)
);

AO22x2_ASAP7_75t_L g1447 ( 
.A1(n_1437),
.A2(n_1318),
.B1(n_267),
.B2(n_271),
.Y(n_1447)
);

INVx1_ASAP7_75t_L g1448 ( 
.A(n_1442),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1443),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1444),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1446),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1447),
.Y(n_1452)
);

OAI22xp5_ASAP7_75t_SL g1453 ( 
.A1(n_1448),
.A2(n_1441),
.B1(n_1440),
.B2(n_1438),
.Y(n_1453)
);

AOI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1449),
.A2(n_1445),
.B1(n_1318),
.B2(n_277),
.Y(n_1454)
);

OAI22xp5_ASAP7_75t_L g1455 ( 
.A1(n_1451),
.A2(n_1450),
.B1(n_1452),
.B2(n_278),
.Y(n_1455)
);

AOI22xp5_ASAP7_75t_L g1456 ( 
.A1(n_1448),
.A2(n_265),
.B1(n_274),
.B2(n_279),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1453),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1455),
.Y(n_1458)
);

INVx1_ASAP7_75t_L g1459 ( 
.A(n_1454),
.Y(n_1459)
);

AOI22xp5_ASAP7_75t_SL g1460 ( 
.A1(n_1457),
.A2(n_1456),
.B1(n_283),
.B2(n_286),
.Y(n_1460)
);

OAI22xp33_ASAP7_75t_L g1461 ( 
.A1(n_1458),
.A2(n_281),
.B1(n_287),
.B2(n_288),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1460),
.Y(n_1462)
);

AOI221xp5_ASAP7_75t_L g1463 ( 
.A1(n_1462),
.A2(n_1459),
.B1(n_1461),
.B2(n_293),
.C(n_294),
.Y(n_1463)
);

AOI211xp5_ASAP7_75t_L g1464 ( 
.A1(n_1463),
.A2(n_290),
.B(n_292),
.C(n_296),
.Y(n_1464)
);


endmodule