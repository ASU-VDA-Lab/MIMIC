module fake_jpeg_3050_n_584 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_584);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_584;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx2_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_18),
.Y(n_22)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_6),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_7),
.B(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_7),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

BUFx16f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_1),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g43 ( 
.A(n_6),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_18),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_0),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_9),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_8),
.Y(n_52)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_6),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_9),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_13),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_29),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_57),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_50),
.Y(n_58)
);

INVx4_ASAP7_75t_SL g139 ( 
.A(n_58),
.Y(n_139)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_55),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_59),
.Y(n_146)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_60),
.Y(n_144)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_61),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_62),
.B(n_63),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_40),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_40),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_64),
.B(n_84),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_20),
.B(n_10),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_65),
.B(n_69),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_66),
.Y(n_142)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_20),
.Y(n_67)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_67),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_55),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g152 ( 
.A(n_68),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_28),
.B(n_8),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_70),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_0),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_71),
.B(n_72),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_34),
.B(n_8),
.Y(n_72)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g160 ( 
.A(n_73),
.Y(n_160)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_28),
.Y(n_74)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_74),
.Y(n_141)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_33),
.Y(n_75)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_75),
.Y(n_153)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

INVx1_ASAP7_75t_SL g77 ( 
.A(n_50),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_77),
.B(n_125),
.Y(n_209)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_78),
.Y(n_145)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx5_ASAP7_75t_L g184 ( 
.A(n_79),
.Y(n_184)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_56),
.Y(n_80)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_34),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_81),
.B(n_85),
.Y(n_182)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_41),
.Y(n_82)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_82),
.Y(n_137)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_55),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g192 ( 
.A(n_83),
.Y(n_192)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_11),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_33),
.B(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_24),
.Y(n_86)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_86),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_46),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_87),
.B(n_113),
.Y(n_161)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_36),
.Y(n_88)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_88),
.Y(n_180)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_56),
.Y(n_89)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_89),
.Y(n_129)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g198 ( 
.A(n_90),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_46),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_91),
.B(n_123),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_36),
.B(n_44),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_92),
.B(n_95),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_39),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_93),
.Y(n_212)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_44),
.Y(n_94)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_94),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_34),
.B(n_51),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_96),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_19),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_97),
.B(n_101),
.Y(n_190)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_99),
.Y(n_143)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_27),
.Y(n_100)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_100),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_27),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_19),
.B(n_11),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_102),
.B(n_111),
.Y(n_197)
);

INVx11_ASAP7_75t_L g103 ( 
.A(n_30),
.Y(n_103)
);

INVx11_ASAP7_75t_L g200 ( 
.A(n_103),
.Y(n_200)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_30),
.Y(n_104)
);

INVx5_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_27),
.Y(n_105)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_105),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

INVx6_ASAP7_75t_L g150 ( 
.A(n_106),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g107 ( 
.A(n_37),
.Y(n_107)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_107),
.Y(n_163)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_39),
.Y(n_108)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_108),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_37),
.Y(n_109)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_52),
.Y(n_110)
);

INVx5_ASAP7_75t_L g214 ( 
.A(n_110),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_37),
.B(n_1),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_26),
.B(n_11),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_112),
.B(n_121),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_21),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_52),
.Y(n_114)
);

INVx6_ASAP7_75t_L g155 ( 
.A(n_114),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_52),
.Y(n_115)
);

INVx6_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_116),
.Y(n_154)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_30),
.Y(n_117)
);

INVx11_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_21),
.Y(n_118)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_52),
.Y(n_119)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_21),
.Y(n_120)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_120),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_26),
.B(n_12),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_21),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_122),
.B(n_124),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_31),
.B(n_12),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_22),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_23),
.B(n_22),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_22),
.Y(n_126)
);

INVx4_ASAP7_75t_L g186 ( 
.A(n_126),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_48),
.Y(n_127)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_127),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g128 ( 
.A1(n_125),
.A2(n_43),
.B1(n_35),
.B2(n_32),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_128),
.A2(n_135),
.B1(n_140),
.B2(n_167),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_91),
.A2(n_43),
.B1(n_23),
.B2(n_49),
.Y(n_133)
);

OA22x2_ASAP7_75t_L g225 ( 
.A1(n_133),
.A2(n_147),
.B1(n_157),
.B2(n_162),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_71),
.A2(n_31),
.B1(n_47),
.B2(n_45),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_98),
.A2(n_32),
.B1(n_35),
.B2(n_49),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_58),
.A2(n_49),
.B1(n_77),
.B2(n_48),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_120),
.A2(n_48),
.B1(n_47),
.B2(n_54),
.Y(n_157)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_81),
.B(n_45),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_159),
.B(n_16),
.Y(n_251)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_103),
.A2(n_48),
.B1(n_54),
.B2(n_42),
.Y(n_162)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_166),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_101),
.A2(n_111),
.B1(n_100),
.B2(n_105),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g169 ( 
.A1(n_117),
.A2(n_48),
.B1(n_42),
.B2(n_53),
.Y(n_169)
);

OA22x2_ASAP7_75t_L g243 ( 
.A1(n_169),
.A2(n_188),
.B1(n_202),
.B2(n_218),
.Y(n_243)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_116),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g254 ( 
.A(n_171),
.Y(n_254)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_73),
.Y(n_172)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_172),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_84),
.A2(n_126),
.B1(n_86),
.B2(n_119),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_174),
.A2(n_187),
.B1(n_2),
.B2(n_5),
.Y(n_249)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_79),
.Y(n_176)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_176),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_108),
.A2(n_66),
.B1(n_57),
.B2(n_115),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_178),
.A2(n_219),
.B1(n_124),
.B2(n_113),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_61),
.B(n_53),
.C(n_50),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_181),
.B(n_4),
.C(n_5),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_76),
.A2(n_38),
.B1(n_25),
.B2(n_53),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_78),
.A2(n_38),
.B1(n_25),
.B2(n_3),
.Y(n_188)
);

INVx4_ASAP7_75t_L g195 ( 
.A(n_104),
.Y(n_195)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_82),
.Y(n_196)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_196),
.Y(n_221)
);

BUFx2_ASAP7_75t_SL g199 ( 
.A(n_127),
.Y(n_199)
);

INVx3_ASAP7_75t_L g237 ( 
.A(n_199),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_80),
.A2(n_38),
.B1(n_25),
.B2(n_3),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_67),
.B(n_17),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_203),
.B(n_205),
.Y(n_248)
);

INVx4_ASAP7_75t_L g204 ( 
.A(n_59),
.Y(n_204)
);

INVx3_ASAP7_75t_L g239 ( 
.A(n_204),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_74),
.B(n_94),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_75),
.B(n_17),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_208),
.B(n_210),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_88),
.B(n_7),
.Y(n_210)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_89),
.Y(n_211)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx3_ASAP7_75t_L g213 ( 
.A(n_68),
.Y(n_213)
);

BUFx12f_ASAP7_75t_L g267 ( 
.A(n_213),
.Y(n_267)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_83),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_215),
.Y(n_282)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_118),
.Y(n_216)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

AOI22xp33_ASAP7_75t_SL g218 ( 
.A1(n_110),
.A2(n_5),
.B1(n_15),
.B2(n_3),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_70),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g289 ( 
.A(n_219),
.B(n_212),
.Y(n_289)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_220),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_156),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_222),
.B(n_224),
.Y(n_326)
);

INVx5_ASAP7_75t_L g223 ( 
.A(n_152),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g342 ( 
.A(n_223),
.Y(n_342)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_131),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_209),
.A2(n_110),
.B1(n_90),
.B2(n_106),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g319 ( 
.A(n_226),
.Y(n_319)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_227),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_SL g230 ( 
.A1(n_209),
.A2(n_114),
.B1(n_99),
.B2(n_93),
.Y(n_230)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_230),
.Y(n_334)
);

OR2x2_ASAP7_75t_SL g231 ( 
.A(n_197),
.B(n_109),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g310 ( 
.A(n_231),
.Y(n_310)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_207),
.Y(n_232)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_232),
.Y(n_303)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_173),
.Y(n_233)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_233),
.Y(n_322)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_153),
.Y(n_234)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_234),
.Y(n_306)
);

OR2x4_ASAP7_75t_L g235 ( 
.A(n_159),
.B(n_107),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_235),
.B(n_247),
.Y(n_304)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_138),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

INVx11_ASAP7_75t_L g238 ( 
.A(n_139),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g335 ( 
.A(n_238),
.Y(n_335)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_158),
.A2(n_13),
.B(n_16),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_240),
.A2(n_235),
.B(n_247),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_190),
.B(n_1),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_241),
.B(n_256),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_139),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_242),
.B(n_250),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_128),
.A2(n_96),
.B1(n_2),
.B2(n_1),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_244),
.A2(n_297),
.B1(n_245),
.B2(n_232),
.Y(n_311)
);

BUFx4f_ASAP7_75t_L g246 ( 
.A(n_186),
.Y(n_246)
);

INVx2_ASAP7_75t_L g323 ( 
.A(n_246),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_249),
.A2(n_260),
.B1(n_265),
.B2(n_266),
.Y(n_341)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_161),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g353 ( 
.A(n_251),
.B(n_264),
.Y(n_353)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_138),
.Y(n_253)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_253),
.Y(n_314)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_183),
.Y(n_255)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_255),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_177),
.B(n_2),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g257 ( 
.A1(n_164),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_257)
);

OAI22xp33_ASAP7_75t_SL g320 ( 
.A1(n_257),
.A2(n_263),
.B1(n_293),
.B2(n_230),
.Y(n_320)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_142),
.Y(n_258)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_258),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_182),
.B(n_2),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_259),
.B(n_271),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_180),
.A2(n_14),
.B1(n_15),
.B2(n_201),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_185),
.B(n_14),
.C(n_151),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_261),
.B(n_288),
.C(n_231),
.Y(n_307)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_170),
.A2(n_14),
.B1(n_140),
.B2(n_132),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_168),
.B(n_217),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g265 ( 
.A1(n_194),
.A2(n_145),
.B1(n_148),
.B2(n_215),
.Y(n_265)
);

AOI22xp33_ASAP7_75t_SL g266 ( 
.A1(n_152),
.A2(n_192),
.B1(n_133),
.B2(n_211),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g268 ( 
.A1(n_192),
.A2(n_129),
.B1(n_204),
.B2(n_154),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_268),
.A2(n_286),
.B1(n_238),
.B2(n_246),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_144),
.B(n_134),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_269),
.B(n_275),
.Y(n_313)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_175),
.Y(n_270)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_270),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_136),
.B(n_137),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_129),
.B(n_186),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_273),
.B(n_295),
.Y(n_347)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_143),
.Y(n_274)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_274),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_146),
.B(n_184),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_195),
.Y(n_276)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_276),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_157),
.B(n_189),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_277),
.B(n_280),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_146),
.B(n_193),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_278),
.B(n_285),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g279 ( 
.A(n_130),
.B(n_165),
.Y(n_279)
);

AND2x2_ASAP7_75t_L g327 ( 
.A(n_279),
.B(n_287),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_143),
.B(n_189),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_281),
.Y(n_332)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_142),
.Y(n_283)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_283),
.Y(n_339)
);

AO22x1_ASAP7_75t_SL g284 ( 
.A1(n_130),
.A2(n_165),
.B1(n_163),
.B2(n_212),
.Y(n_284)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_284),
.Y(n_349)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_191),
.Y(n_285)
);

AOI22xp33_ASAP7_75t_SL g286 ( 
.A1(n_188),
.A2(n_202),
.B1(n_160),
.B2(n_163),
.Y(n_286)
);

AND2x2_ASAP7_75t_L g287 ( 
.A(n_214),
.B(n_150),
.Y(n_287)
);

OR2x2_ASAP7_75t_SL g288 ( 
.A(n_218),
.B(n_147),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_289),
.B(n_290),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_150),
.B(n_155),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_149),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_291),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_155),
.B(n_149),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_292),
.B(n_272),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g293 ( 
.A1(n_198),
.A2(n_200),
.B1(n_206),
.B2(n_162),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_198),
.B(n_200),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_256),
.B(n_169),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_300),
.B(n_301),
.C(n_328),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_241),
.B(n_206),
.Y(n_301)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_307),
.B(n_320),
.Y(n_357)
);

HAxp5_ASAP7_75t_SL g395 ( 
.A(n_308),
.B(n_352),
.CON(n_395),
.SN(n_395)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_311),
.A2(n_337),
.B1(n_340),
.B2(n_343),
.Y(n_361)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_261),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_244),
.A2(n_277),
.B1(n_297),
.B2(n_280),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_329),
.A2(n_350),
.B1(n_272),
.B2(n_254),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_252),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g358 ( 
.A(n_333),
.B(n_351),
.Y(n_358)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_288),
.A2(n_225),
.B(n_243),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g373 ( 
.A1(n_336),
.A2(n_337),
.B(n_300),
.Y(n_373)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_243),
.A2(n_225),
.B1(n_274),
.B2(n_255),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_221),
.B(n_228),
.C(n_279),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_338),
.B(n_346),
.C(n_352),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_243),
.A2(n_225),
.B1(n_233),
.B2(n_287),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_243),
.A2(n_225),
.B1(n_287),
.B2(n_258),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g370 ( 
.A(n_344),
.B(n_345),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_248),
.B(n_240),
.Y(n_345)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_221),
.B(n_279),
.Y(n_346)
);

OAI22xp33_ASAP7_75t_SL g377 ( 
.A1(n_348),
.A2(n_237),
.B1(n_267),
.B2(n_341),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_228),
.A2(n_284),
.B1(n_272),
.B2(n_246),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_294),
.B(n_229),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_296),
.B(n_262),
.C(n_239),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_355),
.A2(n_366),
.B1(n_369),
.B2(n_379),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g356 ( 
.A(n_351),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g398 ( 
.A(n_356),
.B(n_359),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_312),
.B(n_294),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_340),
.A2(n_223),
.B1(n_284),
.B2(n_229),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_360),
.A2(n_368),
.B(n_373),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_312),
.B(n_254),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_362),
.B(n_375),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_254),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_363),
.B(n_372),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_311),
.A2(n_236),
.B1(n_291),
.B2(n_253),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_364),
.A2(n_380),
.B1(n_393),
.B2(n_335),
.Y(n_409)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_305),
.Y(n_365)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_365),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_336),
.A2(n_329),
.B1(n_349),
.B2(n_310),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_343),
.A2(n_282),
.B1(n_239),
.B2(n_262),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_349),
.A2(n_283),
.B1(n_296),
.B2(n_282),
.Y(n_369)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_328),
.B(n_237),
.C(n_267),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_371),
.B(n_381),
.C(n_384),
.Y(n_407)
);

CKINVDCx16_ASAP7_75t_R g372 ( 
.A(n_327),
.Y(n_372)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_303),
.Y(n_374)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_374),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_309),
.B(n_267),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_303),
.Y(n_376)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_377),
.Y(n_412)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_321),
.Y(n_378)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_378),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_334),
.A2(n_304),
.B1(n_308),
.B2(n_333),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_334),
.A2(n_304),
.B1(n_347),
.B2(n_307),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_304),
.B(n_309),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_316),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

OAI21xp5_ASAP7_75t_SL g383 ( 
.A1(n_347),
.A2(n_319),
.B(n_324),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g403 ( 
.A1(n_383),
.A2(n_335),
.B(n_330),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_301),
.B(n_346),
.C(n_298),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_299),
.B(n_326),
.Y(n_385)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_385),
.B(n_386),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_SL g386 ( 
.A(n_353),
.B(n_299),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_326),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_387),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g388 ( 
.A(n_316),
.Y(n_388)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_388),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_298),
.B(n_313),
.Y(n_389)
);

NOR2x1_ASAP7_75t_L g415 ( 
.A(n_389),
.B(n_391),
.Y(n_415)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_325),
.Y(n_390)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_390),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_338),
.B(n_327),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_SL g392 ( 
.A1(n_319),
.A2(n_350),
.B1(n_306),
.B2(n_302),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_315),
.B1(n_322),
.B2(n_323),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_302),
.A2(n_306),
.B1(n_331),
.B2(n_325),
.Y(n_393)
);

INVx4_ASAP7_75t_L g394 ( 
.A(n_342),
.Y(n_394)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_394),
.Y(n_431)
);

OAI22x1_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_330),
.B1(n_332),
.B2(n_315),
.Y(n_408)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_396),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_353),
.B(n_318),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_354),
.C(n_381),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_403),
.B(n_394),
.Y(n_456)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_408),
.B(n_433),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g449 ( 
.A1(n_409),
.A2(n_413),
.B1(n_430),
.B2(n_424),
.Y(n_449)
);

OAI22xp33_ASAP7_75t_L g410 ( 
.A1(n_361),
.A2(n_331),
.B1(n_317),
.B2(n_339),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g447 ( 
.A1(n_410),
.A2(n_411),
.B1(n_369),
.B2(n_355),
.Y(n_447)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_361),
.A2(n_314),
.B1(n_317),
.B2(n_339),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_L g413 ( 
.A1(n_364),
.A2(n_314),
.B1(n_316),
.B2(n_332),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_SL g443 ( 
.A1(n_414),
.A2(n_426),
.B1(n_432),
.B2(n_406),
.Y(n_443)
);

FAx1_ASAP7_75t_SL g416 ( 
.A(n_354),
.B(n_322),
.CI(n_342),
.CON(n_416),
.SN(n_416)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_416),
.B(n_426),
.Y(n_454)
);

AOI22xp5_ASAP7_75t_L g417 ( 
.A1(n_366),
.A2(n_323),
.B1(n_373),
.B2(n_379),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g442 ( 
.A1(n_417),
.A2(n_363),
.B1(n_387),
.B2(n_397),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_418),
.B(n_358),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g421 ( 
.A1(n_383),
.A2(n_359),
.B(n_362),
.Y(n_421)
);

OAI21xp5_ASAP7_75t_L g451 ( 
.A1(n_421),
.A2(n_422),
.B(n_417),
.Y(n_451)
);

OAI21xp5_ASAP7_75t_L g422 ( 
.A1(n_357),
.A2(n_356),
.B(n_380),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_384),
.B(n_367),
.C(n_391),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_425),
.B(n_429),
.C(n_357),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g426 ( 
.A(n_393),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_367),
.B(n_371),
.C(n_372),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_360),
.A2(n_358),
.B1(n_389),
.B2(n_368),
.Y(n_430)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_374),
.Y(n_432)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_432),
.Y(n_437)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_434),
.B(n_435),
.C(n_436),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_425),
.B(n_429),
.C(n_407),
.Y(n_436)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_406),
.Y(n_438)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_438),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_418),
.B(n_357),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_428),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g440 ( 
.A(n_399),
.B(n_375),
.Y(n_440)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_440),
.Y(n_480)
);

CKINVDCx14_ASAP7_75t_R g441 ( 
.A(n_423),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g483 ( 
.A1(n_441),
.A2(n_447),
.B1(n_449),
.B2(n_455),
.Y(n_483)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_442),
.A2(n_451),
.B1(n_464),
.B2(n_434),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_443),
.A2(n_456),
.B1(n_412),
.B2(n_428),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_407),
.B(n_363),
.C(n_370),
.Y(n_444)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_444),
.B(n_461),
.C(n_465),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_399),
.B(n_376),
.Y(n_445)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_445),
.Y(n_478)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_419),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_398),
.B(n_396),
.Y(n_448)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_448),
.Y(n_481)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_419),
.Y(n_450)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_450),
.Y(n_485)
);

INVxp67_ASAP7_75t_L g473 ( 
.A(n_451),
.Y(n_473)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_424),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_404),
.Y(n_453)
);

INVx1_ASAP7_75t_SL g490 ( 
.A(n_453),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_400),
.A2(n_392),
.B1(n_390),
.B2(n_388),
.Y(n_455)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_404),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_458),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g458 ( 
.A(n_398),
.B(n_382),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_405),
.B(n_382),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_459),
.B(n_462),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g460 ( 
.A1(n_400),
.A2(n_388),
.B1(n_422),
.B2(n_411),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_431),
.B1(n_402),
.B2(n_427),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g461 ( 
.A(n_415),
.B(n_433),
.C(n_405),
.Y(n_461)
);

CKINVDCx20_ASAP7_75t_R g462 ( 
.A(n_423),
.Y(n_462)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_463),
.A2(n_412),
.B(n_414),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_421),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_464),
.Y(n_472)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_433),
.B(n_416),
.C(n_403),
.Y(n_465)
);

FAx1_ASAP7_75t_SL g466 ( 
.A(n_461),
.B(n_416),
.CI(n_408),
.CON(n_466),
.SN(n_466)
);

A2O1A1Ixp33_ASAP7_75t_L g511 ( 
.A1(n_466),
.A2(n_473),
.B(n_471),
.C(n_481),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_467),
.A2(n_470),
.B1(n_484),
.B2(n_486),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_469),
.B(n_474),
.C(n_487),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g474 ( 
.A(n_439),
.B(n_401),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_436),
.B(n_401),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g498 ( 
.A(n_475),
.B(n_476),
.Y(n_498)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_435),
.B(n_420),
.Y(n_476)
);

NOR3xp33_ASAP7_75t_L g515 ( 
.A(n_482),
.B(n_469),
.C(n_466),
.Y(n_515)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_460),
.A2(n_410),
.B1(n_420),
.B2(n_402),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_444),
.B(n_431),
.C(n_427),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_465),
.B(n_442),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_488),
.B(n_459),
.C(n_445),
.Y(n_502)
);

OAI22xp5_ASAP7_75t_SL g489 ( 
.A1(n_455),
.A2(n_402),
.B1(n_462),
.B2(n_447),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_489),
.B(n_458),
.Y(n_504)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_463),
.B(n_454),
.Y(n_491)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_491),
.B(n_457),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_473),
.A2(n_482),
.B(n_472),
.Y(n_493)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_493),
.Y(n_533)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_492),
.Y(n_494)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_494),
.Y(n_517)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_492),
.Y(n_495)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_495),
.Y(n_518)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_480),
.Y(n_496)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_475),
.B(n_454),
.Y(n_500)
);

CKINVDCx14_ASAP7_75t_R g516 ( 
.A(n_500),
.Y(n_516)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_466),
.B(n_440),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_501),
.B(n_506),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g530 ( 
.A(n_502),
.B(n_468),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_476),
.B(n_448),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g525 ( 
.A(n_503),
.B(n_507),
.Y(n_525)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_504),
.Y(n_521)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_470),
.A2(n_437),
.B1(n_438),
.B2(n_446),
.Y(n_505)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_505),
.Y(n_529)
);

OAI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_481),
.A2(n_437),
.B1(n_450),
.B2(n_452),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_487),
.B(n_453),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_478),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g527 ( 
.A(n_508),
.B(n_509),
.Y(n_527)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_478),
.Y(n_509)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_510),
.B(n_474),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_511),
.B(n_512),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_490),
.Y(n_512)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_467),
.A2(n_491),
.B(n_477),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g522 ( 
.A(n_513),
.B(n_514),
.Y(n_522)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_479),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_488),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_523),
.A2(n_511),
.B(n_501),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g524 ( 
.A1(n_499),
.A2(n_495),
.B1(n_494),
.B2(n_504),
.Y(n_524)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_524),
.A2(n_489),
.B1(n_510),
.B2(n_497),
.Y(n_546)
);

XNOR2xp5_ASAP7_75t_L g541 ( 
.A(n_526),
.B(n_530),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g528 ( 
.A(n_502),
.B(n_468),
.Y(n_528)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_528),
.B(n_532),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_498),
.B(n_496),
.Y(n_532)
);

OAI22xp5_ASAP7_75t_SL g535 ( 
.A1(n_519),
.A2(n_493),
.B1(n_509),
.B2(n_508),
.Y(n_535)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_535),
.A2(n_540),
.B1(n_543),
.B2(n_546),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_527),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g552 ( 
.A(n_536),
.B(n_522),
.Y(n_552)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_527),
.Y(n_537)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_537),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g538 ( 
.A(n_520),
.B(n_506),
.Y(n_538)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

XOR2xp5_ASAP7_75t_L g539 ( 
.A(n_526),
.B(n_497),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g558 ( 
.A(n_539),
.B(n_548),
.Y(n_558)
);

OAI22xp5_ASAP7_75t_SL g540 ( 
.A1(n_519),
.A2(n_513),
.B1(n_484),
.B2(n_512),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_520),
.B(n_490),
.Y(n_542)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_542),
.A2(n_544),
.B(n_545),
.Y(n_554)
);

INVx1_ASAP7_75t_L g543 ( 
.A(n_524),
.Y(n_543)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_533),
.A2(n_505),
.B(n_483),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_530),
.B(n_498),
.C(n_471),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_547),
.B(n_525),
.Y(n_560)
);

XNOR2xp5_ASAP7_75t_L g548 ( 
.A(n_525),
.B(n_514),
.Y(n_548)
);

BUFx24_ASAP7_75t_SL g549 ( 
.A(n_544),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_549),
.B(n_551),
.Y(n_563)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_548),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g567 ( 
.A(n_552),
.B(n_555),
.Y(n_567)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_547),
.B(n_529),
.C(n_533),
.Y(n_555)
);

AOI21xp5_ASAP7_75t_L g556 ( 
.A1(n_534),
.A2(n_531),
.B(n_516),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g569 ( 
.A(n_556),
.B(n_557),
.Y(n_569)
);

XOR2xp5_ASAP7_75t_L g557 ( 
.A(n_546),
.B(n_531),
.Y(n_557)
);

NAND2xp5_ASAP7_75t_SL g565 ( 
.A(n_560),
.B(n_541),
.Y(n_565)
);

AO21x1_ASAP7_75t_L g561 ( 
.A1(n_554),
.A2(n_537),
.B(n_517),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_561),
.B(n_562),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g562 ( 
.A(n_558),
.B(n_539),
.C(n_541),
.Y(n_562)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_550),
.B(n_543),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_564),
.B(n_565),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_555),
.B(n_557),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_566),
.B(n_568),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_553),
.B(n_540),
.C(n_535),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_569),
.B(n_550),
.C(n_529),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g577 ( 
.A1(n_572),
.A2(n_575),
.B(n_561),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_567),
.B(n_559),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_574),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_L g575 ( 
.A1(n_564),
.A2(n_518),
.B1(n_517),
.B2(n_545),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_577),
.B(n_578),
.Y(n_580)
);

NOR3xp33_ASAP7_75t_L g578 ( 
.A(n_570),
.B(n_563),
.C(n_518),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_576),
.A2(n_573),
.B(n_571),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g581 ( 
.A1(n_579),
.A2(n_580),
.B(n_542),
.Y(n_581)
);

OAI21xp33_ASAP7_75t_L g582 ( 
.A1(n_581),
.A2(n_572),
.B(n_538),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g583 ( 
.A(n_582),
.B(n_521),
.C(n_485),
.Y(n_583)
);

BUFx24_ASAP7_75t_SL g584 ( 
.A(n_583),
.Y(n_584)
);


endmodule