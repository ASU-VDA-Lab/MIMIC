module fake_jpeg_1677_n_143 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_143);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_143;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_12),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_10),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_11),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_14),
.B(n_13),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_30),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g46 ( 
.A(n_31),
.B(n_32),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_15),
.B(n_0),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_21),
.Y(n_35)
);

CKINVDCx16_ASAP7_75t_R g59 ( 
.A(n_35),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_SL g36 ( 
.A(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_14),
.B(n_9),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_39),
.B(n_43),
.Y(n_48)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_27),
.Y(n_40)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_28),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_3),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_2),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_29),
.B(n_3),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_24),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g72 ( 
.A1(n_51),
.A2(n_57),
.B(n_64),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_30),
.B(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_52),
.B(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_20),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_33),
.B(n_29),
.C(n_24),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_42),
.C(n_22),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_18),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_39),
.A2(n_22),
.B1(n_26),
.B2(n_20),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_58),
.A2(n_36),
.B1(n_23),
.B2(n_26),
.Y(n_68)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_32),
.B(n_19),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_66),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_48),
.A2(n_31),
.B1(n_43),
.B2(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_67),
.B(n_70),
.Y(n_100)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_68),
.B(n_76),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_48),
.A2(n_34),
.B1(n_37),
.B2(n_42),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_48),
.A2(n_34),
.B1(n_42),
.B2(n_22),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_73),
.B(n_74),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_66),
.A2(n_37),
.B1(n_17),
.B2(n_16),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_78),
.B(n_80),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_66),
.A2(n_17),
.B1(n_23),
.B2(n_19),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g95 ( 
.A1(n_79),
.A2(n_80),
.B(n_73),
.Y(n_95)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_46),
.B(n_16),
.Y(n_80)
);

INVx2_ASAP7_75t_R g82 ( 
.A(n_59),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_62),
.B(n_60),
.Y(n_96)
);

AOI32xp33_ASAP7_75t_L g83 ( 
.A1(n_63),
.A2(n_25),
.A3(n_10),
.B1(n_5),
.B2(n_4),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_83),
.B(n_56),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_25),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_60),
.C(n_56),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_45),
.A2(n_4),
.B1(n_5),
.B2(n_55),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_89),
.Y(n_104)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_90),
.B(n_92),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_84),
.Y(n_91)
);

NAND3xp33_ASAP7_75t_L g105 ( 
.A(n_91),
.B(n_97),
.C(n_77),
.Y(n_105)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g94 ( 
.A(n_67),
.B(n_63),
.C(n_65),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_74),
.C(n_85),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_95),
.B(n_99),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_82),
.Y(n_109)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_75),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_96),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_101),
.B(n_105),
.Y(n_114)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_88),
.B(n_81),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_102),
.B(n_110),
.C(n_108),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_87),
.A2(n_79),
.B1(n_81),
.B2(n_72),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_103),
.B(n_109),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_107),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_108),
.B(n_87),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_88),
.B(n_70),
.C(n_76),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_93),
.B(n_47),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_112),
.B(n_90),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_101),
.A2(n_88),
.B(n_100),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_113),
.A2(n_106),
.B(n_110),
.Y(n_127)
);

OAI22xp33_ASAP7_75t_R g116 ( 
.A1(n_111),
.A2(n_86),
.B1(n_94),
.B2(n_95),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_115),
.B(n_114),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_117),
.B(n_119),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_99),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_109),
.A2(n_100),
.B(n_86),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_120),
.A2(n_92),
.B(n_50),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.C(n_102),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_129),
.C(n_121),
.Y(n_130)
);

INVx11_ASAP7_75t_L g124 ( 
.A(n_118),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_124),
.A2(n_128),
.B(n_118),
.Y(n_133)
);

FAx1_ASAP7_75t_SL g131 ( 
.A(n_126),
.B(n_120),
.CI(n_115),
.CON(n_131),
.SN(n_131)
);

OAI21xp5_ASAP7_75t_SL g132 ( 
.A1(n_127),
.A2(n_115),
.B(n_113),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_54),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_130),
.B(n_132),
.C(n_134),
.Y(n_135)
);

AOI31xp33_ASAP7_75t_L g138 ( 
.A1(n_131),
.A2(n_128),
.A3(n_124),
.B(n_5),
.Y(n_138)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_133),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_123),
.B(n_54),
.C(n_61),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_132),
.B(n_125),
.C(n_129),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g140 ( 
.A(n_137),
.Y(n_140)
);

OAI31xp33_ASAP7_75t_L g139 ( 
.A1(n_138),
.A2(n_136),
.A3(n_4),
.B(n_135),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_139),
.B(n_49),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_140),
.B(n_49),
.C(n_139),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_141),
.B(n_142),
.Y(n_143)
);


endmodule