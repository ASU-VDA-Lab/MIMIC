module fake_aes_5998_n_24 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_0, n_24);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_0;
output n_24;
wire n_20;
wire n_23;
wire n_8;
wire n_22;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
INVx2_ASAP7_75t_L g8 ( .A(n_4), .Y(n_8) );
CKINVDCx5p33_ASAP7_75t_R g9 ( .A(n_0), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_1), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_2), .Y(n_11) );
INVx1_ASAP7_75t_L g12 ( .A(n_11), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_13), .B(n_9), .Y(n_14) );
OAI21x1_ASAP7_75t_L g15 ( .A1(n_12), .A2(n_10), .B(n_8), .Y(n_15) );
INVx1_ASAP7_75t_SL g16 ( .A(n_14), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_16), .B(n_15), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_16), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
NOR2x1_ASAP7_75t_L g20 ( .A(n_19), .B(n_17), .Y(n_20) );
HB1xp67_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
XOR2xp5_ASAP7_75t_L g22 ( .A(n_21), .B(n_3), .Y(n_22) );
NOR3x2_ASAP7_75t_L g23 ( .A(n_22), .B(n_5), .C(n_6), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_7), .Y(n_24) );
endmodule