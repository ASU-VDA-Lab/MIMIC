module real_jpeg_25238_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_201;
wire n_114;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_215;
wire n_176;
wire n_104;
wire n_194;
wire n_153;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_87;
wire n_197;
wire n_105;
wire n_40;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_126;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_162;
wire n_121;
wire n_106;
wire n_160;
wire n_211;
wire n_172;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_165;
wire n_134;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_210;
wire n_206;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_2),
.A2(n_23),
.B1(n_24),
.B2(n_25),
.Y(n_22)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_2),
.A2(n_25),
.B1(n_39),
.B2(n_42),
.Y(n_121)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_5),
.A2(n_23),
.B1(n_24),
.B2(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_5),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g38 ( 
.A1(n_6),
.A2(n_39),
.B1(n_41),
.B2(n_42),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_6),
.A2(n_41),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_6),
.A2(n_23),
.B1(n_24),
.B2(n_41),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_6),
.A2(n_41),
.B1(n_53),
.B2(n_55),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_7),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_8),
.A2(n_23),
.B1(n_24),
.B2(n_32),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_8),
.A2(n_32),
.B1(n_39),
.B2(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_8),
.A2(n_32),
.B1(n_58),
.B2(n_62),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_8),
.A2(n_32),
.B1(n_53),
.B2(n_55),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_52),
.C(n_55),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_8),
.B(n_51),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_8),
.B(n_39),
.C(n_70),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_8),
.B(n_24),
.C(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_8),
.B(n_152),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_8),
.B(n_85),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_8),
.B(n_104),
.Y(n_194)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_9),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_9),
.A2(n_52),
.B1(n_56),
.B2(n_58),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_11),
.Y(n_99)
);

XOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_124),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_123),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_105),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_16),
.B(n_105),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_76),
.C(n_86),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_17),
.A2(n_18),
.B1(n_76),
.B2(n_216),
.Y(n_215)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_20),
.B1(n_47),
.B2(n_48),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_19),
.B(n_49),
.C(n_66),
.Y(n_106)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_33),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_21),
.A2(n_33),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_21),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_26),
.B(n_27),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g78 ( 
.A1(n_22),
.A2(n_29),
.B1(n_79),
.B2(n_81),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g34 ( 
.A1(n_23),
.A2(n_24),
.B1(n_35),
.B2(n_36),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_24),
.B(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_24),
.B(n_184),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_26),
.B(n_29),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g152 ( 
.A(n_26),
.Y(n_152)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_28),
.A2(n_97),
.B(n_152),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_31),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_29),
.Y(n_96)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_31),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_33),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_33),
.A2(n_130),
.B1(n_178),
.B2(n_180),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_33),
.B(n_180),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_33),
.A2(n_111),
.B1(n_113),
.B2(n_130),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_33),
.B(n_111),
.C(n_201),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B(n_43),
.Y(n_33)
);

AND2x2_ASAP7_75t_L g45 ( 
.A(n_34),
.B(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_34),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_34),
.A2(n_43),
.B(n_121),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_34),
.B(n_135),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_L g46 ( 
.A1(n_35),
.A2(n_36),
.B1(n_39),
.B2(n_42),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_38),
.A2(n_44),
.B1(n_45),
.B2(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_39),
.Y(n_42)
);

OA22x2_ASAP7_75t_SL g72 ( 
.A1(n_39),
.A2(n_42),
.B1(n_70),
.B2(n_71),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_39),
.B(n_179),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_45),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_44),
.B(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_45),
.Y(n_135)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_65),
.B1(n_66),
.B2(n_75),
.Y(n_48)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_49),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_49),
.A2(n_75),
.B1(n_145),
.B2(n_146),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g49 ( 
.A1(n_50),
.A2(n_57),
.B(n_60),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_64),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_51),
.A2(n_61),
.B1(n_63),
.B2(n_88),
.Y(n_87)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_55),
.B2(n_56),
.Y(n_51)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_SL g55 ( 
.A(n_53),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_53),
.A2(n_55),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_55),
.B(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_57),
.Y(n_88)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_58),
.Y(n_59)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_58),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_63),
.Y(n_60)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g66 ( 
.A1(n_67),
.A2(n_72),
.B(n_73),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_68),
.A2(n_74),
.B1(n_102),
.B2(n_104),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_68),
.B(n_74),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_72),
.Y(n_68)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_70),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_72),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_72),
.A2(n_103),
.B(n_112),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_113),
.C(n_133),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g216 ( 
.A(n_76),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_78),
.B(n_83),
.Y(n_109)
);

INVx5_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_81),
.B(n_117),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_83),
.A2(n_84),
.B1(n_194),
.B2(n_195),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_83),
.A2(n_84),
.B1(n_163),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_84),
.B(n_157),
.C(n_163),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_84),
.B(n_95),
.C(n_194),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_86),
.B(n_215),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_89),
.C(n_101),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_87),
.A2(n_111),
.B1(n_113),
.B2(n_114),
.Y(n_110)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_87),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_101),
.B1(n_114),
.B2(n_140),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_89),
.B(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_94),
.A2(n_95),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_95),
.B(n_186),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_95),
.B(n_186),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_98),
.B2(n_100),
.Y(n_95)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_100),
.B(n_118),
.Y(n_168)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_101),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_150),
.C(n_151),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_140),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_115),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_113),
.B1(n_133),
.B2(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_116),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_115)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_116),
.Y(n_122)
);

INVxp33_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_153),
.B(n_212),
.C(n_217),
.Y(n_124)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_142),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_126),
.B(n_142),
.Y(n_211)
);

AOI22xp33_ASAP7_75t_SL g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_138),
.B2(n_141),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_132),
.B1(n_136),
.B2(n_137),
.Y(n_128)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_129),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_129),
.B(n_137),
.C(n_141),
.Y(n_213)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_132),
.Y(n_137)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_138),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_148),
.C(n_149),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_143),
.A2(n_144),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_148),
.B(n_149),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_150),
.A2(n_151),
.B1(n_161),
.B2(n_162),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_150),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_151),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g182 ( 
.A(n_151),
.B(n_183),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_211),
.Y(n_153)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_172),
.B(n_210),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_169),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_156),
.B(n_169),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_157),
.A2(n_158),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_162),
.B(n_177),
.Y(n_188)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_163),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_167),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_164),
.A2(n_165),
.B1(n_167),
.B2(n_168),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_173),
.A2(n_203),
.B(n_209),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g173 ( 
.A1(n_174),
.A2(n_197),
.B(n_202),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_189),
.B(n_196),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_176),
.A2(n_181),
.B(n_188),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_178),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_185),
.B(n_187),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_190),
.B(n_191),
.Y(n_196)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_194),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_198),
.B(n_199),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_198),
.B(n_199),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_205),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_204),
.B(n_205),
.Y(n_209)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_206),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_213),
.B(n_214),
.Y(n_217)
);


endmodule