module real_aes_2386_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_678;
wire n_548;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_119;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_554;
wire n_475;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g217 ( .A(n_0), .B(n_160), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_1), .A2(n_142), .B(n_193), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g462 ( .A1(n_2), .A2(n_463), .B1(n_468), .B2(n_813), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_3), .B(n_112), .Y(n_111) );
AOI22xp5_ASAP7_75t_L g126 ( .A1(n_4), .A2(n_11), .B1(n_127), .B2(n_128), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g128 ( .A(n_4), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g206 ( .A(n_5), .B(n_150), .Y(n_206) );
INVx1_ASAP7_75t_L g147 ( .A(n_6), .Y(n_147) );
NAND2xp5_ASAP7_75t_L g170 ( .A(n_7), .B(n_150), .Y(n_170) );
AOI22xp5_ASAP7_75t_L g121 ( .A1(n_8), .A2(n_122), .B1(n_446), .B2(n_447), .Y(n_121) );
INVxp67_ASAP7_75t_L g447 ( .A(n_8), .Y(n_447) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_8), .B(n_137), .Y(n_504) );
INVx1_ASAP7_75t_L g532 ( .A(n_9), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g112 ( .A(n_10), .Y(n_112) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_11), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g547 ( .A(n_12), .Y(n_547) );
NAND2xp33_ASAP7_75t_L g187 ( .A(n_13), .B(n_154), .Y(n_187) );
INVx2_ASAP7_75t_L g139 ( .A(n_14), .Y(n_139) );
AOI221x1_ASAP7_75t_L g229 ( .A1(n_15), .A2(n_29), .B1(n_142), .B2(n_160), .C(n_230), .Y(n_229) );
CKINVDCx16_ASAP7_75t_R g113 ( .A(n_16), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_17), .B(n_160), .Y(n_183) );
AO21x2_ASAP7_75t_L g180 ( .A1(n_18), .A2(n_181), .B(n_182), .Y(n_180) );
INVx1_ASAP7_75t_L g513 ( .A(n_19), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_20), .B(n_173), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_21), .B(n_150), .Y(n_149) );
AO21x1_ASAP7_75t_L g201 ( .A1(n_22), .A2(n_160), .B(n_202), .Y(n_201) );
INVx1_ASAP7_75t_L g109 ( .A(n_23), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_24), .B(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g511 ( .A(n_25), .Y(n_511) );
INVx1_ASAP7_75t_SL g497 ( .A(n_26), .Y(n_497) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_27), .Y(n_822) );
NAND2xp5_ASAP7_75t_SL g591 ( .A(n_28), .B(n_161), .Y(n_591) );
NAND2x1_ASAP7_75t_L g215 ( .A(n_30), .B(n_150), .Y(n_215) );
AOI33xp33_ASAP7_75t_L g559 ( .A1(n_31), .A2(n_56), .A3(n_487), .B1(n_494), .B2(n_560), .B3(n_561), .Y(n_559) );
NAND2x1_ASAP7_75t_L g169 ( .A(n_32), .B(n_154), .Y(n_169) );
INVx1_ASAP7_75t_L g541 ( .A(n_33), .Y(n_541) );
OR2x2_ASAP7_75t_L g138 ( .A(n_34), .B(n_90), .Y(n_138) );
OA21x2_ASAP7_75t_L g178 ( .A1(n_34), .A2(n_90), .B(n_139), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g484 ( .A(n_35), .B(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_36), .B(n_154), .Y(n_195) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_37), .B(n_150), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_38), .B(n_154), .Y(n_205) );
AOI21xp5_ASAP7_75t_L g247 ( .A1(n_39), .A2(n_142), .B(n_248), .Y(n_247) );
AND2x2_ASAP7_75t_L g143 ( .A(n_40), .B(n_144), .Y(n_143) );
AND2x2_ASAP7_75t_L g158 ( .A(n_40), .B(n_147), .Y(n_158) );
INVx1_ASAP7_75t_L g493 ( .A(n_40), .Y(n_493) );
NOR3xp33_ASAP7_75t_L g110 ( .A(n_41), .B(n_111), .C(n_113), .Y(n_110) );
OR2x6_ASAP7_75t_L g452 ( .A(n_41), .B(n_453), .Y(n_452) );
XNOR2xp5_ASAP7_75t_L g464 ( .A(n_42), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_43), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g251 ( .A(n_44), .B(n_160), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_45), .B(n_485), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g584 ( .A1(n_46), .A2(n_137), .B1(n_177), .B2(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_47), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_48), .B(n_161), .Y(n_499) );
CKINVDCx20_ASAP7_75t_R g163 ( .A(n_49), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_50), .B(n_154), .Y(n_249) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_51), .B(n_181), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_52), .B(n_161), .Y(n_533) );
AOI21xp5_ASAP7_75t_L g167 ( .A1(n_53), .A2(n_142), .B(n_168), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g588 ( .A(n_54), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_55), .B(n_154), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_57), .B(n_161), .Y(n_571) );
INVx1_ASAP7_75t_L g146 ( .A(n_58), .Y(n_146) );
INVx1_ASAP7_75t_L g156 ( .A(n_58), .Y(n_156) );
AND2x2_ASAP7_75t_L g572 ( .A(n_59), .B(n_173), .Y(n_572) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_60), .A2(n_77), .B1(n_485), .B2(n_491), .C(n_531), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_61), .B(n_485), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_62), .B(n_150), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_63), .B(n_177), .Y(n_549) );
AOI21xp5_ASAP7_75t_SL g521 ( .A1(n_64), .A2(n_491), .B(n_522), .Y(n_521) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_65), .A2(n_142), .B(n_214), .Y(n_213) );
INVx1_ASAP7_75t_L g507 ( .A(n_66), .Y(n_507) );
AO21x1_ASAP7_75t_L g203 ( .A1(n_67), .A2(n_142), .B(n_204), .Y(n_203) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_68), .B(n_160), .Y(n_191) );
INVx1_ASAP7_75t_L g570 ( .A(n_69), .Y(n_570) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_70), .B(n_160), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_71), .A2(n_491), .B(n_569), .Y(n_568) );
AND2x2_ASAP7_75t_L g252 ( .A(n_72), .B(n_174), .Y(n_252) );
INVx1_ASAP7_75t_L g144 ( .A(n_73), .Y(n_144) );
INVx1_ASAP7_75t_L g152 ( .A(n_73), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_74), .A2(n_100), .B1(n_466), .B2(n_467), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g466 ( .A(n_74), .Y(n_466) );
AND2x2_ASAP7_75t_L g175 ( .A(n_75), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_76), .B(n_485), .Y(n_562) );
AND2x2_ASAP7_75t_L g500 ( .A(n_78), .B(n_176), .Y(n_500) );
INVx1_ASAP7_75t_L g508 ( .A(n_79), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_80), .A2(n_491), .B(n_496), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g589 ( .A1(n_81), .A2(n_491), .B(n_554), .C(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g108 ( .A(n_82), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g159 ( .A(n_83), .B(n_160), .Y(n_159) );
AND2x2_ASAP7_75t_L g189 ( .A(n_84), .B(n_176), .Y(n_189) );
AND2x2_ASAP7_75t_SL g519 ( .A(n_85), .B(n_176), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g556 ( .A1(n_86), .A2(n_491), .B1(n_557), .B2(n_558), .Y(n_556) );
OAI22xp5_ASAP7_75t_SL g123 ( .A1(n_87), .A2(n_124), .B1(n_125), .B2(n_126), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_87), .Y(n_124) );
XNOR2xp5_ASAP7_75t_L g463 ( .A(n_88), .B(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g202 ( .A(n_89), .B(n_137), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_91), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g219 ( .A(n_92), .B(n_176), .Y(n_219) );
INVx1_ASAP7_75t_L g523 ( .A(n_93), .Y(n_523) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_94), .B(n_150), .Y(n_250) );
AOI21xp5_ASAP7_75t_L g141 ( .A1(n_95), .A2(n_142), .B(n_148), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_96), .B(n_154), .Y(n_231) );
AND2x2_ASAP7_75t_L g563 ( .A(n_97), .B(n_176), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g194 ( .A(n_98), .B(n_150), .Y(n_194) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_99), .A2(n_539), .B(n_540), .C(n_542), .Y(n_538) );
CKINVDCx20_ASAP7_75t_R g467 ( .A(n_100), .Y(n_467) );
BUFx2_ASAP7_75t_L g119 ( .A(n_101), .Y(n_119) );
BUFx2_ASAP7_75t_SL g460 ( .A(n_101), .Y(n_460) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_102), .A2(n_142), .B(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_103), .B(n_161), .Y(n_524) );
AOI21xp33_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_114), .B(n_821), .Y(n_104) );
BUFx2_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
INVx3_ASAP7_75t_SL g825 ( .A(n_106), .Y(n_825) );
AND2x2_ASAP7_75t_SL g106 ( .A(n_107), .B(n_110), .Y(n_106) );
NOR2xp33_ASAP7_75t_L g107 ( .A(n_108), .B(n_109), .Y(n_107) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_108), .B(n_109), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_113), .B(n_451), .Y(n_450) );
AND2x6_ASAP7_75t_SL g472 ( .A(n_113), .B(n_452), .Y(n_472) );
OR2x6_ASAP7_75t_SL g475 ( .A(n_113), .B(n_451), .Y(n_475) );
OR2x2_ASAP7_75t_L g814 ( .A(n_113), .B(n_452), .Y(n_814) );
OA22x2_ASAP7_75t_L g114 ( .A1(n_115), .A2(n_120), .B1(n_457), .B2(n_461), .Y(n_114) );
INVx1_ASAP7_75t_SL g115 ( .A(n_116), .Y(n_115) );
BUFx3_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
OAI21xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_448), .B(n_454), .Y(n_120) );
INVx1_ASAP7_75t_L g446 ( .A(n_122), .Y(n_446) );
XNOR2x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_129), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g468 ( .A1(n_129), .A2(n_469), .B1(n_473), .B2(n_476), .Y(n_468) );
INVx2_ASAP7_75t_L g818 ( .A(n_129), .Y(n_818) );
OR2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_344), .Y(n_129) );
NAND3xp33_ASAP7_75t_SL g130 ( .A(n_131), .B(n_256), .C(n_311), .Y(n_130) );
AOI221xp5_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_196), .B1(n_220), .B2(n_224), .C(n_234), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_179), .Y(n_132) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_133), .B(n_223), .Y(n_222) );
INVx2_ASAP7_75t_L g255 ( .A(n_133), .Y(n_255) );
AND2x2_ASAP7_75t_L g300 ( .A(n_133), .B(n_237), .Y(n_300) );
AND2x4_ASAP7_75t_L g133 ( .A(n_134), .B(n_164), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx2_ASAP7_75t_L g288 ( .A(n_135), .Y(n_288) );
INVx1_ASAP7_75t_L g298 ( .A(n_135), .Y(n_298) );
AO21x2_ASAP7_75t_L g135 ( .A1(n_136), .A2(n_140), .B(n_162), .Y(n_135) );
NOR2xp33_ASAP7_75t_L g162 ( .A(n_136), .B(n_163), .Y(n_162) );
AO21x2_ASAP7_75t_L g262 ( .A1(n_136), .A2(n_140), .B(n_162), .Y(n_262) );
INVx1_ASAP7_75t_SL g136 ( .A(n_137), .Y(n_136) );
AOI21xp5_ASAP7_75t_L g182 ( .A1(n_137), .A2(n_183), .B(n_184), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_137), .B(n_208), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g515 ( .A(n_137), .B(n_157), .Y(n_515) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_137), .A2(n_521), .B(n_525), .Y(n_520) );
AND2x4_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
AND2x2_ASAP7_75t_SL g174 ( .A(n_138), .B(n_139), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_141), .B(n_159), .Y(n_140) );
AND2x6_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
BUFx3_ASAP7_75t_L g489 ( .A(n_143), .Y(n_489) );
AND2x6_ASAP7_75t_L g154 ( .A(n_144), .B(n_155), .Y(n_154) );
INVx2_ASAP7_75t_L g495 ( .A(n_144), .Y(n_495) );
AND2x4_ASAP7_75t_L g491 ( .A(n_145), .B(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g145 ( .A(n_146), .B(n_147), .Y(n_145) );
AND2x4_ASAP7_75t_L g150 ( .A(n_146), .B(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g487 ( .A(n_146), .Y(n_487) );
HB1xp67_ASAP7_75t_L g488 ( .A(n_147), .Y(n_488) );
AOI21xp5_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_153), .B(n_157), .Y(n_148) );
INVxp67_ASAP7_75t_L g514 ( .A(n_150), .Y(n_514) );
AND2x4_ASAP7_75t_L g161 ( .A(n_151), .B(n_155), .Y(n_161) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVxp67_ASAP7_75t_L g512 ( .A(n_154), .Y(n_512) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AOI21xp5_ASAP7_75t_L g168 ( .A1(n_157), .A2(n_169), .B(n_170), .Y(n_168) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_157), .A2(n_186), .B(n_187), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g193 ( .A1(n_157), .A2(n_194), .B(n_195), .Y(n_193) );
AOI21xp5_ASAP7_75t_L g204 ( .A1(n_157), .A2(n_205), .B(n_206), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_157), .A2(n_215), .B(n_216), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_157), .A2(n_231), .B(n_232), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_157), .A2(n_249), .B(n_250), .Y(n_248) );
O2A1O1Ixp33_ASAP7_75t_SL g496 ( .A1(n_157), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
O2A1O1Ixp33_ASAP7_75t_L g522 ( .A1(n_157), .A2(n_498), .B(n_523), .C(n_524), .Y(n_522) );
O2A1O1Ixp33_ASAP7_75t_SL g531 ( .A1(n_157), .A2(n_498), .B(n_532), .C(n_533), .Y(n_531) );
INVx1_ASAP7_75t_L g557 ( .A(n_157), .Y(n_557) );
O2A1O1Ixp33_ASAP7_75t_L g569 ( .A1(n_157), .A2(n_498), .B(n_570), .C(n_571), .Y(n_569) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_157), .A2(n_591), .B(n_592), .Y(n_590) );
INVx5_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
AND2x4_ASAP7_75t_L g160 ( .A(n_158), .B(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_158), .Y(n_542) );
INVx1_ASAP7_75t_L g509 ( .A(n_161), .Y(n_509) );
OR2x2_ASAP7_75t_L g277 ( .A(n_164), .B(n_180), .Y(n_277) );
NAND2x1p5_ASAP7_75t_L g308 ( .A(n_164), .B(n_223), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_164), .B(n_188), .Y(n_321) );
INVx2_ASAP7_75t_L g330 ( .A(n_164), .Y(n_330) );
AND2x2_ASAP7_75t_L g351 ( .A(n_164), .B(n_352), .Y(n_351) );
AND2x2_ASAP7_75t_L g435 ( .A(n_164), .B(n_254), .Y(n_435) );
INVx4_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
AND2x2_ASAP7_75t_L g263 ( .A(n_165), .B(n_188), .Y(n_263) );
AND2x2_ASAP7_75t_L g396 ( .A(n_165), .B(n_223), .Y(n_396) );
HB1xp67_ASAP7_75t_L g422 ( .A(n_165), .Y(n_422) );
AO21x2_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_172), .B(n_175), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_167), .B(n_171), .Y(n_166) );
AO21x2_ASAP7_75t_L g482 ( .A1(n_172), .A2(n_483), .B(n_500), .Y(n_482) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_173), .A2(n_191), .B(n_192), .Y(n_190) );
OA21x2_ASAP7_75t_L g228 ( .A1(n_173), .A2(n_229), .B(n_233), .Y(n_228) );
OA21x2_ASAP7_75t_L g240 ( .A1(n_173), .A2(n_229), .B(n_233), .Y(n_240) );
BUFx6f_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
INVx3_ASAP7_75t_L g218 ( .A(n_176), .Y(n_218) );
OAI22xp5_ASAP7_75t_L g537 ( .A1(n_176), .A2(n_218), .B1(n_538), .B2(n_543), .Y(n_537) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_177), .B(n_546), .Y(n_545) );
INVx3_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
BUFx4f_ASAP7_75t_L g181 ( .A(n_178), .Y(n_181) );
AND2x4_ASAP7_75t_L g350 ( .A(n_179), .B(n_351), .Y(n_350) );
AOI321xp33_ASAP7_75t_L g364 ( .A1(n_179), .A2(n_293), .A3(n_294), .B1(n_326), .B2(n_365), .C(n_368), .Y(n_364) );
AND2x2_ASAP7_75t_L g179 ( .A(n_180), .B(n_188), .Y(n_179) );
BUFx3_ASAP7_75t_L g221 ( .A(n_180), .Y(n_221) );
INVx2_ASAP7_75t_L g254 ( .A(n_180), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_180), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g287 ( .A(n_180), .B(n_288), .Y(n_287) );
INVx1_ASAP7_75t_L g320 ( .A(n_180), .Y(n_320) );
OA21x2_ASAP7_75t_L g529 ( .A1(n_181), .A2(n_530), .B(n_534), .Y(n_529) );
INVx2_ASAP7_75t_SL g554 ( .A(n_181), .Y(n_554) );
INVx5_ASAP7_75t_L g223 ( .A(n_188), .Y(n_223) );
NOR2x1_ASAP7_75t_SL g272 ( .A(n_188), .B(n_262), .Y(n_272) );
BUFx2_ASAP7_75t_L g367 ( .A(n_188), .Y(n_367) );
OR2x6_ASAP7_75t_L g188 ( .A(n_189), .B(n_190), .Y(n_188) );
INVxp67_ASAP7_75t_L g196 ( .A(n_197), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_209), .Y(n_197) );
NOR2xp33_ASAP7_75t_SL g265 ( .A(n_198), .B(n_266), .Y(n_265) );
NOR4xp25_ASAP7_75t_L g368 ( .A(n_198), .B(n_362), .C(n_366), .D(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g406 ( .A(n_198), .Y(n_406) );
AND2x2_ASAP7_75t_L g440 ( .A(n_198), .B(n_380), .Y(n_440) );
BUFx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx2_ASAP7_75t_L g241 ( .A(n_199), .Y(n_241) );
INVx2_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
INVx2_ASAP7_75t_L g295 ( .A(n_200), .Y(n_295) );
OAI21x1_ASAP7_75t_SL g200 ( .A1(n_201), .A2(n_203), .B(n_207), .Y(n_200) );
INVx1_ASAP7_75t_L g208 ( .A(n_202), .Y(n_208) );
AOI33xp33_ASAP7_75t_L g436 ( .A1(n_209), .A2(n_238), .A3(n_269), .B1(n_285), .B2(n_391), .B3(n_437), .Y(n_436) );
INVx1_ASAP7_75t_SL g209 ( .A(n_210), .Y(n_209) );
AND2x2_ASAP7_75t_L g226 ( .A(n_210), .B(n_227), .Y(n_226) );
AND2x4_ASAP7_75t_L g236 ( .A(n_210), .B(n_237), .Y(n_236) );
BUFx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
INVx2_ASAP7_75t_L g243 ( .A(n_211), .Y(n_243) );
INVxp67_ASAP7_75t_L g324 ( .A(n_211), .Y(n_324) );
AND2x2_ASAP7_75t_L g380 ( .A(n_211), .B(n_245), .Y(n_380) );
AO21x2_ASAP7_75t_L g211 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_211) );
AO21x2_ASAP7_75t_L g284 ( .A1(n_212), .A2(n_218), .B(n_219), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g212 ( .A(n_213), .B(n_217), .Y(n_212) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_218), .A2(n_246), .B(n_252), .Y(n_245) );
AO21x2_ASAP7_75t_L g281 ( .A1(n_218), .A2(n_246), .B(n_252), .Y(n_281) );
AO21x2_ASAP7_75t_L g565 ( .A1(n_218), .A2(n_566), .B(n_572), .Y(n_565) );
AO21x2_ASAP7_75t_L g603 ( .A1(n_218), .A2(n_566), .B(n_572), .Y(n_603) );
AOI21xp5_ASAP7_75t_L g401 ( .A1(n_220), .A2(n_402), .B(n_403), .Y(n_401) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_222), .Y(n_220) );
AND2x2_ASAP7_75t_L g389 ( .A(n_221), .B(n_263), .Y(n_389) );
AND3x2_ASAP7_75t_L g391 ( .A(n_221), .B(n_275), .C(n_330), .Y(n_391) );
INVx3_ASAP7_75t_SL g343 ( .A(n_222), .Y(n_343) );
INVx4_ASAP7_75t_L g237 ( .A(n_223), .Y(n_237) );
AND2x2_ASAP7_75t_L g275 ( .A(n_223), .B(n_262), .Y(n_275) );
INVxp67_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
BUFx2_ASAP7_75t_L g269 ( .A(n_227), .Y(n_269) );
AND2x4_ASAP7_75t_L g294 ( .A(n_227), .B(n_295), .Y(n_294) );
AND2x2_ASAP7_75t_L g357 ( .A(n_227), .B(n_245), .Y(n_357) );
INVx2_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx2_ASAP7_75t_L g327 ( .A(n_228), .Y(n_327) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_228), .Y(n_349) );
O2A1O1Ixp33_ASAP7_75t_R g234 ( .A1(n_235), .A2(n_238), .B(n_242), .C(n_253), .Y(n_234) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_236), .Y(n_235) );
AND2x2_ASAP7_75t_L g286 ( .A(n_237), .B(n_287), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_237), .B(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_237), .B(n_254), .Y(n_415) );
INVx1_ASAP7_75t_SL g238 ( .A(n_239), .Y(n_238) );
AND2x2_ASAP7_75t_L g397 ( .A(n_239), .B(n_387), .Y(n_397) );
AND2x2_ASAP7_75t_SL g239 ( .A(n_240), .B(n_241), .Y(n_239) );
AND2x2_ASAP7_75t_L g244 ( .A(n_240), .B(n_245), .Y(n_244) );
AND2x2_ASAP7_75t_L g266 ( .A(n_240), .B(n_267), .Y(n_266) );
AND2x2_ASAP7_75t_L g282 ( .A(n_240), .B(n_283), .Y(n_282) );
AND2x4_ASAP7_75t_L g315 ( .A(n_240), .B(n_295), .Y(n_315) );
AND2x4_ASAP7_75t_L g280 ( .A(n_241), .B(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g304 ( .A(n_241), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g342 ( .A(n_241), .B(n_267), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_243), .B(n_244), .Y(n_242) );
AND2x2_ASAP7_75t_L g270 ( .A(n_243), .B(n_267), .Y(n_270) );
AND2x2_ASAP7_75t_L g285 ( .A(n_243), .B(n_245), .Y(n_285) );
BUFx2_ASAP7_75t_L g341 ( .A(n_243), .Y(n_341) );
AND2x2_ASAP7_75t_L g355 ( .A(n_243), .B(n_266), .Y(n_355) );
INVx2_ASAP7_75t_L g267 ( .A(n_245), .Y(n_267) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_247), .B(n_251), .Y(n_246) );
OAI22xp33_ASAP7_75t_L g303 ( .A1(n_253), .A2(n_304), .B1(n_306), .B2(n_310), .Y(n_303) );
INVx2_ASAP7_75t_SL g334 ( .A(n_253), .Y(n_334) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
AND2x2_ASAP7_75t_L g309 ( .A(n_254), .B(n_262), .Y(n_309) );
INVx1_ASAP7_75t_L g416 ( .A(n_255), .Y(n_416) );
NOR3xp33_ASAP7_75t_L g256 ( .A(n_257), .B(n_289), .C(n_303), .Y(n_256) );
OAI221xp5_ASAP7_75t_SL g257 ( .A1(n_258), .A2(n_264), .B1(n_268), .B2(n_271), .C(n_273), .Y(n_257) );
INVx1_ASAP7_75t_SL g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_263), .Y(n_259) );
INVxp67_ASAP7_75t_SL g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g317 ( .A(n_261), .Y(n_317) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_261), .Y(n_445) );
INVx1_ASAP7_75t_L g408 ( .A(n_263), .Y(n_408) );
AND2x2_ASAP7_75t_SL g418 ( .A(n_263), .B(n_287), .Y(n_418) );
INVxp67_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_267), .B(n_295), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
OR2x2_ASAP7_75t_L g301 ( .A(n_269), .B(n_302), .Y(n_301) );
INVx1_ASAP7_75t_L g379 ( .A(n_269), .Y(n_379) );
AND2x2_ASAP7_75t_L g314 ( .A(n_270), .B(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g360 ( .A(n_272), .B(n_320), .Y(n_360) );
AND2x2_ASAP7_75t_L g437 ( .A(n_272), .B(n_435), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g273 ( .A1(n_274), .A2(n_278), .B1(n_285), .B2(n_286), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
INVx2_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g296 ( .A(n_277), .B(n_297), .Y(n_296) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_282), .Y(n_279) );
INVx2_ASAP7_75t_L g302 ( .A(n_280), .Y(n_302) );
AND2x4_ASAP7_75t_L g326 ( .A(n_280), .B(n_327), .Y(n_326) );
OAI21xp33_ASAP7_75t_SL g356 ( .A1(n_280), .A2(n_357), .B(n_358), .Y(n_356) );
AND2x2_ASAP7_75t_L g383 ( .A(n_280), .B(n_341), .Y(n_383) );
INVx2_ASAP7_75t_L g305 ( .A(n_281), .Y(n_305) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_281), .Y(n_338) );
INVx1_ASAP7_75t_SL g362 ( .A(n_282), .Y(n_362) );
INVx1_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
BUFx2_ASAP7_75t_L g293 ( .A(n_284), .Y(n_293) );
AND2x4_ASAP7_75t_SL g387 ( .A(n_284), .B(n_305), .Y(n_387) );
AND2x2_ASAP7_75t_L g384 ( .A(n_287), .B(n_330), .Y(n_384) );
AND2x2_ASAP7_75t_L g410 ( .A(n_287), .B(n_396), .Y(n_410) );
HB1xp67_ASAP7_75t_L g332 ( .A(n_288), .Y(n_332) );
INVx1_ASAP7_75t_L g352 ( .A(n_288), .Y(n_352) );
OAI22xp33_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_296), .B1(n_299), .B2(n_301), .Y(n_289) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_294), .Y(n_291) );
INVx2_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g310 ( .A(n_294), .B(n_305), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_294), .B(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g433 ( .A(n_294), .Y(n_433) );
INVx2_ASAP7_75t_SL g358 ( .A(n_296), .Y(n_358) );
AND2x2_ASAP7_75t_L g370 ( .A(n_298), .B(n_330), .Y(n_370) );
INVx2_ASAP7_75t_L g376 ( .A(n_298), .Y(n_376) );
INVxp33_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
INVx2_ASAP7_75t_L g335 ( .A(n_301), .Y(n_335) );
NOR2xp33_ASAP7_75t_L g361 ( .A(n_304), .B(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx1_ASAP7_75t_L g354 ( .A(n_306), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_309), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_307), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g365 ( .A(n_309), .B(n_366), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_309), .A2(n_439), .B1(n_440), .B2(n_441), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g311 ( .A(n_312), .B(n_333), .C(n_336), .Y(n_311) );
OAI221xp5_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_316), .B1(n_318), .B2(n_322), .C(n_325), .Y(n_312) );
INVx1_ASAP7_75t_SL g313 ( .A(n_314), .Y(n_313) );
INVx1_ASAP7_75t_SL g431 ( .A(n_316), .Y(n_431) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g400 ( .A(n_317), .B(n_366), .Y(n_400) );
OR2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
AND2x2_ASAP7_75t_L g331 ( .A(n_320), .B(n_332), .Y(n_331) );
INVx1_ASAP7_75t_L g402 ( .A(n_322), .Y(n_402) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g399 ( .A(n_323), .Y(n_399) );
INVx1_ASAP7_75t_L g405 ( .A(n_324), .Y(n_405) );
OR2x2_ASAP7_75t_L g428 ( .A(n_324), .B(n_429), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_328), .Y(n_325) );
INVx1_ASAP7_75t_SL g337 ( .A(n_327), .Y(n_337) );
AND2x2_ASAP7_75t_L g407 ( .A(n_327), .B(n_387), .Y(n_407) );
AND2x2_ASAP7_75t_SL g439 ( .A(n_327), .B(n_340), .Y(n_439) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx1_ASAP7_75t_L g444 ( .A(n_330), .Y(n_444) );
INVx1_ASAP7_75t_L g394 ( .A(n_332), .Y(n_394) );
AND2x2_ASAP7_75t_L g333 ( .A(n_334), .B(n_335), .Y(n_333) );
O2A1O1Ixp33_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_338), .B(n_339), .C(n_343), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_337), .B(n_387), .Y(n_411) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_340), .B(n_391), .Y(n_390) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_342), .Y(n_340) );
AND2x2_ASAP7_75t_L g348 ( .A(n_342), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g429 ( .A(n_342), .Y(n_429) );
NAND4xp75_ASAP7_75t_L g344 ( .A(n_345), .B(n_401), .C(n_417), .D(n_438), .Y(n_344) );
NOR3x1_ASAP7_75t_L g345 ( .A(n_346), .B(n_363), .C(n_385), .Y(n_345) );
NAND4xp75_ASAP7_75t_L g346 ( .A(n_347), .B(n_353), .C(n_356), .D(n_359), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g347 ( .A(n_348), .B(n_350), .Y(n_347) );
AND2x2_ASAP7_75t_L g398 ( .A(n_349), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g423 ( .A(n_350), .Y(n_423) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_SL g412 ( .A(n_355), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_364), .B(n_371), .Y(n_363) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g430 ( .A(n_367), .B(n_431), .Y(n_430) );
INVx1_ASAP7_75t_SL g369 ( .A(n_370), .Y(n_369) );
AOI21xp5_ASAP7_75t_L g371 ( .A1(n_372), .A2(n_377), .B(n_381), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI322xp33_ASAP7_75t_L g403 ( .A1(n_375), .A2(n_404), .A3(n_408), .B1(n_409), .B2(n_411), .C1(n_412), .C2(n_413), .Y(n_403) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_376), .B(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_380), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_379), .B(n_426), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_380), .B(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_383), .B(n_384), .Y(n_382) );
OAI211xp5_ASAP7_75t_L g385 ( .A1(n_386), .A2(n_388), .B(n_390), .C(n_392), .Y(n_385) );
INVx1_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_397), .B1(n_398), .B2(n_400), .Y(n_392) );
NOR2xp33_ASAP7_75t_SL g393 ( .A(n_394), .B(n_395), .Y(n_393) );
INVx2_ASAP7_75t_SL g395 ( .A(n_396), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B(n_407), .Y(n_404) );
INVxp67_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_410), .B(n_443), .Y(n_442) );
NAND2xp5_ASAP7_75t_SL g413 ( .A(n_414), .B(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g420 ( .A(n_415), .B(n_421), .Y(n_420) );
O2A1O1Ixp5_ASAP7_75t_L g417 ( .A1(n_418), .A2(n_419), .B(n_424), .C(n_427), .Y(n_417) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_420), .B(n_423), .Y(n_419) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
OAI221xp5_ASAP7_75t_SL g427 ( .A1(n_428), .A2(n_430), .B1(n_432), .B2(n_434), .C(n_436), .Y(n_427) );
INVxp67_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g443 ( .A(n_444), .B(n_445), .Y(n_443) );
INVx2_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx2_ASAP7_75t_L g456 ( .A(n_450), .Y(n_456) );
CKINVDCx5p33_ASAP7_75t_R g451 ( .A(n_452), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g457 ( .A(n_454), .B(n_458), .Y(n_457) );
INVx1_ASAP7_75t_SL g455 ( .A(n_456), .Y(n_455) );
CKINVDCx11_ASAP7_75t_R g458 ( .A(n_459), .Y(n_458) );
CKINVDCx8_ASAP7_75t_R g459 ( .A(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_462), .B(n_815), .Y(n_461) );
INVx1_ASAP7_75t_L g816 ( .A(n_463), .Y(n_816) );
CKINVDCx6p67_ASAP7_75t_R g469 ( .A(n_470), .Y(n_469) );
INVx4_ASAP7_75t_SL g819 ( .A(n_470), .Y(n_819) );
INVx3_ASAP7_75t_SL g470 ( .A(n_471), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
CKINVDCx11_ASAP7_75t_R g474 ( .A(n_475), .Y(n_474) );
OAI22x1_ASAP7_75t_L g817 ( .A1(n_475), .A2(n_818), .B1(n_819), .B2(n_820), .Y(n_817) );
INVx1_ASAP7_75t_L g820 ( .A(n_476), .Y(n_820) );
OR3x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_678), .C(n_749), .Y(n_476) );
NAND3x1_ASAP7_75t_SL g477 ( .A(n_478), .B(n_605), .C(n_627), .Y(n_477) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_595), .Y(n_478) );
AOI22xp33_ASAP7_75t_SL g479 ( .A1(n_480), .A2(n_526), .B1(n_573), .B2(n_577), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_480), .A2(n_781), .B1(n_782), .B2(n_784), .Y(n_780) );
AND2x2_ASAP7_75t_L g480 ( .A(n_481), .B(n_501), .Y(n_480) );
AND2x2_ASAP7_75t_L g596 ( .A(n_481), .B(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_SL g662 ( .A(n_481), .B(n_643), .Y(n_662) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g580 ( .A(n_482), .Y(n_580) );
AND2x2_ASAP7_75t_L g630 ( .A(n_482), .B(n_503), .Y(n_630) );
INVx1_ASAP7_75t_L g669 ( .A(n_482), .Y(n_669) );
OR2x2_ASAP7_75t_L g706 ( .A(n_482), .B(n_518), .Y(n_706) );
HB1xp67_ASAP7_75t_L g718 ( .A(n_482), .Y(n_718) );
HB1xp67_ASAP7_75t_L g742 ( .A(n_482), .Y(n_742) );
AND2x2_ASAP7_75t_L g799 ( .A(n_482), .B(n_626), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_490), .Y(n_483) );
INVx1_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
AND2x4_ASAP7_75t_L g485 ( .A(n_486), .B(n_489), .Y(n_485) );
INVx1_ASAP7_75t_L g586 ( .A(n_486), .Y(n_586) );
AND2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
OR2x6_ASAP7_75t_L g498 ( .A(n_487), .B(n_495), .Y(n_498) );
INVxp33_ASAP7_75t_L g560 ( .A(n_487), .Y(n_560) );
INVx1_ASAP7_75t_L g587 ( .A(n_489), .Y(n_587) );
INVxp67_ASAP7_75t_L g548 ( .A(n_491), .Y(n_548) );
NOR2x1p5_ASAP7_75t_L g492 ( .A(n_493), .B(n_494), .Y(n_492) );
INVx1_ASAP7_75t_L g561 ( .A(n_494), .Y(n_561) );
INVx3_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g506 ( .A1(n_498), .A2(n_507), .B1(n_508), .B2(n_509), .Y(n_506) );
INVxp67_ASAP7_75t_L g539 ( .A(n_498), .Y(n_539) );
INVx2_ASAP7_75t_L g593 ( .A(n_498), .Y(n_593) );
NOR2x1_ASAP7_75t_L g501 ( .A(n_502), .B(n_516), .Y(n_501) );
INVx1_ASAP7_75t_L g674 ( .A(n_502), .Y(n_674) );
AND2x2_ASAP7_75t_L g700 ( .A(n_502), .B(n_518), .Y(n_700) );
NAND2x1_ASAP7_75t_L g716 ( .A(n_502), .B(n_717), .Y(n_716) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AND2x2_ASAP7_75t_L g597 ( .A(n_503), .B(n_583), .Y(n_597) );
INVx3_ASAP7_75t_L g626 ( .A(n_503), .Y(n_626) );
NOR2x1_ASAP7_75t_SL g745 ( .A(n_503), .B(n_518), .Y(n_745) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
OAI21xp5_ASAP7_75t_L g505 ( .A1(n_506), .A2(n_510), .B(n_515), .Y(n_505) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_509), .B(n_541), .Y(n_540) );
OAI22xp5_ASAP7_75t_L g510 ( .A1(n_511), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_510) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_516), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g624 ( .A(n_517), .B(n_625), .Y(n_624) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
INVx4_ASAP7_75t_L g594 ( .A(n_518), .Y(n_594) );
BUFx6f_ASAP7_75t_L g639 ( .A(n_518), .Y(n_639) );
AND2x2_ASAP7_75t_L g711 ( .A(n_518), .B(n_583), .Y(n_711) );
AND2x4_ASAP7_75t_L g728 ( .A(n_518), .B(n_672), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g775 ( .A(n_518), .B(n_670), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_518), .B(n_579), .Y(n_804) );
OR2x6_ASAP7_75t_L g518 ( .A(n_519), .B(n_520), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g733 ( .A1(n_526), .A2(n_621), .B1(n_692), .B2(n_734), .Y(n_733) );
AND2x2_ASAP7_75t_L g526 ( .A(n_527), .B(n_551), .Y(n_526) );
INVx2_ASAP7_75t_L g694 ( .A(n_527), .Y(n_694) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_535), .Y(n_527) );
BUFx3_ASAP7_75t_L g684 ( .A(n_528), .Y(n_684) );
INVx1_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_529), .B(n_553), .Y(n_576) );
INVx2_ASAP7_75t_L g600 ( .A(n_529), .Y(n_600) );
INVx1_ASAP7_75t_L g612 ( .A(n_529), .Y(n_612) );
AND2x4_ASAP7_75t_L g619 ( .A(n_529), .B(n_620), .Y(n_619) );
AND2x2_ASAP7_75t_L g636 ( .A(n_529), .B(n_536), .Y(n_636) );
HB1xp67_ASAP7_75t_L g650 ( .A(n_529), .Y(n_650) );
INVxp67_ASAP7_75t_L g658 ( .A(n_529), .Y(n_658) );
AND2x2_ASAP7_75t_L g687 ( .A(n_535), .B(n_603), .Y(n_687) );
AND2x2_ASAP7_75t_L g703 ( .A(n_535), .B(n_604), .Y(n_703) );
NOR2xp67_ASAP7_75t_L g790 ( .A(n_535), .B(n_603), .Y(n_790) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
AND2x4_ASAP7_75t_L g599 ( .A(n_536), .B(n_600), .Y(n_599) );
INVx1_ASAP7_75t_L g610 ( .A(n_536), .Y(n_610) );
INVx1_ASAP7_75t_L g623 ( .A(n_536), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_536), .B(n_565), .Y(n_660) );
OR2x2_ASAP7_75t_L g536 ( .A(n_537), .B(n_544), .Y(n_536) );
OAI22xp5_ASAP7_75t_L g544 ( .A1(n_545), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_544) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g783 ( .A(n_551), .Y(n_783) );
AND2x4_ASAP7_75t_L g551 ( .A(n_552), .B(n_564), .Y(n_551) );
AND2x2_ASAP7_75t_L g657 ( .A(n_552), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g686 ( .A(n_552), .Y(n_686) );
AND2x2_ASAP7_75t_L g788 ( .A(n_552), .B(n_603), .Y(n_788) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_553), .B(n_565), .Y(n_648) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_555), .B(n_563), .Y(n_553) );
AO21x2_ASAP7_75t_L g604 ( .A1(n_554), .A2(n_555), .B(n_563), .Y(n_604) );
NAND2xp5_ASAP7_75t_SL g555 ( .A(n_556), .B(n_562), .Y(n_555) );
INVx1_ASAP7_75t_L g558 ( .A(n_559), .Y(n_558) );
INVx3_ASAP7_75t_L g574 ( .A(n_564), .Y(n_574) );
NAND2x1p5_ASAP7_75t_L g763 ( .A(n_564), .B(n_684), .Y(n_763) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_565), .Y(n_677) );
AND2x2_ASAP7_75t_L g704 ( .A(n_565), .B(n_650), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_567), .B(n_568), .Y(n_566) );
AND2x2_ASAP7_75t_L g573 ( .A(n_574), .B(n_575), .Y(n_573) );
AND2x2_ASAP7_75t_L g618 ( .A(n_574), .B(n_619), .Y(n_618) );
INVx1_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
AND2x2_ASAP7_75t_L g722 ( .A(n_574), .B(n_599), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_574), .B(n_742), .Y(n_747) );
AND2x2_ASAP7_75t_L g757 ( .A(n_574), .B(n_636), .Y(n_757) );
OR2x2_ASAP7_75t_L g794 ( .A(n_574), .B(n_694), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_575), .B(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g754 ( .A(n_575), .B(n_610), .Y(n_754) );
AND2x2_ASAP7_75t_L g770 ( .A(n_575), .B(n_771), .Y(n_770) );
INVx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
OR2x2_ASAP7_75t_L g764 ( .A(n_576), .B(n_660), .Y(n_764) );
AND2x2_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .Y(n_577) );
INVx1_ASAP7_75t_L g646 ( .A(n_578), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_578), .B(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g744 ( .A(n_578), .B(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_578), .B(n_625), .Y(n_769) );
INVx3_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
HB1xp67_ASAP7_75t_L g616 ( .A(n_579), .Y(n_616) );
INVx2_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
HB1xp67_ASAP7_75t_L g725 ( .A(n_580), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g631 ( .A1(n_581), .A2(n_614), .B1(n_632), .B2(n_635), .Y(n_631) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_581), .B(n_716), .Y(n_715) );
INVx2_ASAP7_75t_SL g748 ( .A(n_581), .Y(n_748) );
AND2x4_ASAP7_75t_SL g581 ( .A(n_582), .B(n_594), .Y(n_581) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
AND2x4_ASAP7_75t_L g625 ( .A(n_583), .B(n_626), .Y(n_625) );
INVx2_ASAP7_75t_L g645 ( .A(n_583), .Y(n_645) );
INVx1_ASAP7_75t_L g672 ( .A(n_583), .Y(n_672) );
AND2x2_ASAP7_75t_L g583 ( .A(n_584), .B(n_589), .Y(n_583) );
NOR3xp33_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .C(n_588), .Y(n_585) );
HB1xp67_ASAP7_75t_L g614 ( .A(n_594), .Y(n_614) );
AND2x4_ASAP7_75t_L g671 ( .A(n_594), .B(n_672), .Y(n_671) );
NOR2x1_ASAP7_75t_L g732 ( .A(n_594), .B(n_701), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_596), .B(n_598), .Y(n_595) );
AND2x2_ASAP7_75t_L g696 ( .A(n_596), .B(n_639), .Y(n_696) );
OAI21xp5_ASAP7_75t_L g776 ( .A1(n_596), .A2(n_777), .B(n_778), .Y(n_776) );
INVx2_ASAP7_75t_L g654 ( .A(n_597), .Y(n_654) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_598), .A2(n_708), .B1(n_712), .B2(n_715), .Y(n_707) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
HB1xp67_ASAP7_75t_L g665 ( .A(n_599), .Y(n_665) );
AND2x2_ASAP7_75t_L g675 ( .A(n_599), .B(n_676), .Y(n_675) );
INVx3_ASAP7_75t_L g714 ( .A(n_599), .Y(n_714) );
NAND2x1_ASAP7_75t_SL g739 ( .A(n_599), .B(n_608), .Y(n_739) );
AND2x2_ASAP7_75t_L g635 ( .A(n_601), .B(n_636), .Y(n_635) );
AND2x4_ASAP7_75t_L g601 ( .A(n_602), .B(n_604), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_603), .Y(n_602) );
NOR2x1_ASAP7_75t_L g611 ( .A(n_603), .B(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g608 ( .A(n_604), .Y(n_608) );
INVx2_ASAP7_75t_L g620 ( .A(n_604), .Y(n_620) );
AOI21xp5_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_613), .B(n_617), .Y(n_605) );
INVx1_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_609), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_608), .B(n_802), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_609), .A2(n_698), .B1(n_702), .B2(n_705), .Y(n_697) );
AND2x2_ASAP7_75t_L g609 ( .A(n_610), .B(n_611), .Y(n_609) );
BUFx2_ASAP7_75t_L g802 ( .A(n_610), .Y(n_802) );
INVx1_ASAP7_75t_SL g809 ( .A(n_610), .Y(n_809) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_611), .Y(n_772) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_614), .B(n_615), .Y(n_613) );
HB1xp67_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
OA21x2_ASAP7_75t_L g617 ( .A1(n_618), .A2(n_621), .B(n_624), .Y(n_617) );
AND2x2_ASAP7_75t_L g621 ( .A(n_619), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g663 ( .A(n_619), .B(n_659), .Y(n_663) );
AND2x2_ASAP7_75t_L g778 ( .A(n_619), .B(n_676), .Y(n_778) );
AND2x2_ASAP7_75t_L g781 ( .A(n_619), .B(n_687), .Y(n_781) );
AND2x4_ASAP7_75t_L g789 ( .A(n_619), .B(n_790), .Y(n_789) );
OAI21xp33_ASAP7_75t_L g743 ( .A1(n_621), .A2(n_744), .B(n_746), .Y(n_743) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
INVx1_ASAP7_75t_L g771 ( .A(n_623), .Y(n_771) );
AND2x2_ASAP7_75t_L g787 ( .A(n_623), .B(n_788), .Y(n_787) );
INVx4_ASAP7_75t_L g701 ( .A(n_625), .Y(n_701) );
INVx1_ASAP7_75t_L g670 ( .A(n_626), .Y(n_670) );
AND2x2_ASAP7_75t_L g692 ( .A(n_626), .B(n_645), .Y(n_692) );
NOR2x1_ASAP7_75t_L g627 ( .A(n_628), .B(n_651), .Y(n_627) );
OAI21xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_631), .B(n_637), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g638 ( .A(n_630), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_SL g791 ( .A(n_630), .B(n_643), .Y(n_791) );
AND2x2_ASAP7_75t_L g812 ( .A(n_630), .B(n_728), .Y(n_812) );
INVx1_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx2_ASAP7_75t_L g738 ( .A(n_635), .Y(n_738) );
OAI21xp5_ASAP7_75t_SL g637 ( .A1(n_638), .A2(n_640), .B(n_647), .Y(n_637) );
OR2x6_ASAP7_75t_L g690 ( .A(n_639), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_642), .B(n_646), .Y(n_641) );
INVx2_ASAP7_75t_SL g642 ( .A(n_643), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_648), .B(n_649), .Y(n_647) );
OR2x2_ASAP7_75t_L g713 ( .A(n_648), .B(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g810 ( .A(n_648), .Y(n_810) );
NOR2xp33_ASAP7_75t_L g782 ( .A(n_649), .B(n_783), .Y(n_782) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_664), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_661), .B2(n_663), .Y(n_652) );
OR2x2_ASAP7_75t_L g724 ( .A(n_654), .B(n_725), .Y(n_724) );
INVx3_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_656), .Y(n_681) );
NAND2x1p5_ASAP7_75t_L g656 ( .A(n_657), .B(n_659), .Y(n_656) );
INVx1_ASAP7_75t_L g730 ( .A(n_659), .Y(n_730) );
INVx2_ASAP7_75t_SL g659 ( .A(n_660), .Y(n_659) );
INVxp67_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_666), .B1(n_673), .B2(n_675), .Y(n_664) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_668), .B(n_671), .Y(n_667) );
AND2x4_ASAP7_75t_SL g668 ( .A(n_669), .B(n_670), .Y(n_668) );
AND2x2_ASAP7_75t_L g673 ( .A(n_671), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g734 ( .A(n_674), .B(n_728), .Y(n_734) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g678 ( .A(n_679), .B(n_719), .Y(n_678) );
NOR2xp67_ASAP7_75t_L g679 ( .A(n_680), .B(n_693), .Y(n_679) );
AOI21xp33_ASAP7_75t_SL g680 ( .A1(n_681), .A2(n_682), .B(n_688), .Y(n_680) );
OR2x2_ASAP7_75t_L g682 ( .A(n_683), .B(n_685), .Y(n_682) );
INVx3_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
NAND2x1p5_ASAP7_75t_L g685 ( .A(n_686), .B(n_687), .Y(n_685) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
OAI22xp33_ASAP7_75t_SL g758 ( .A1(n_690), .A2(n_759), .B1(n_761), .B2(n_764), .Y(n_758) );
NOR2x1_ASAP7_75t_L g705 ( .A(n_691), .B(n_706), .Y(n_705) );
INVx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
AND2x2_ASAP7_75t_L g741 ( .A(n_692), .B(n_742), .Y(n_741) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_695), .B(n_697), .C(n_707), .Y(n_693) );
INVx2_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
NAND2xp33_ASAP7_75t_SL g698 ( .A(n_699), .B(n_701), .Y(n_698) );
INVxp33_ASAP7_75t_L g699 ( .A(n_700), .Y(n_699) );
INVx2_ASAP7_75t_L g710 ( .A(n_701), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g721 ( .A1(n_702), .A2(n_722), .B1(n_723), .B2(n_726), .C(n_729), .Y(n_721) );
AND2x4_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g762 ( .A(n_703), .Y(n_762) );
INVx2_ASAP7_75t_SL g760 ( .A(n_706), .Y(n_760) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_710), .B(n_711), .Y(n_709) );
NAND2x1_ASAP7_75t_L g759 ( .A(n_710), .B(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g756 ( .A(n_716), .Y(n_756) );
INVx1_ASAP7_75t_L g785 ( .A(n_717), .Y(n_785) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
NOR2x1_ASAP7_75t_L g719 ( .A(n_720), .B(n_735), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_721), .B(n_733), .Y(n_720) );
INVx1_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx1_ASAP7_75t_L g774 ( .A(n_725), .Y(n_774) );
INVx1_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
AND2x2_ASAP7_75t_L g795 ( .A(n_728), .B(n_796), .Y(n_795) );
INVx2_ASAP7_75t_L g800 ( .A(n_728), .Y(n_800) );
NOR2xp33_ASAP7_75t_L g729 ( .A(n_730), .B(n_731), .Y(n_729) );
INVxp33_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
BUFx2_ASAP7_75t_L g753 ( .A(n_732), .Y(n_753) );
OAI21xp5_ASAP7_75t_SL g735 ( .A1(n_736), .A2(n_740), .B(n_743), .Y(n_735) );
INVxp67_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_738), .B(n_739), .Y(n_737) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
BUFx2_ASAP7_75t_L g796 ( .A(n_742), .Y(n_796) );
AND2x2_ASAP7_75t_L g784 ( .A(n_745), .B(n_785), .Y(n_784) );
NOR2xp33_ASAP7_75t_R g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND3xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_765), .C(n_792), .Y(n_749) );
NOR2xp33_ASAP7_75t_L g750 ( .A(n_751), .B(n_758), .Y(n_750) );
NAND2xp5_ASAP7_75t_SL g751 ( .A(n_752), .B(n_755), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_753), .B(n_754), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
OR2x2_ASAP7_75t_L g761 ( .A(n_762), .B(n_763), .Y(n_761) );
NOR2xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_779), .Y(n_765) );
NAND2xp5_ASAP7_75t_SL g766 ( .A(n_767), .B(n_776), .Y(n_766) );
AOI22xp33_ASAP7_75t_SL g767 ( .A1(n_768), .A2(n_770), .B1(n_772), .B2(n_773), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
NOR2x1_ASAP7_75t_L g773 ( .A(n_774), .B(n_775), .Y(n_773) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_775), .Y(n_777) );
NAND2xp5_ASAP7_75t_SL g779 ( .A(n_780), .B(n_786), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g786 ( .A1(n_787), .A2(n_789), .B(n_791), .Y(n_786) );
INVx1_ASAP7_75t_L g805 ( .A(n_789), .Y(n_805) );
AOI211xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_795), .B(n_797), .C(n_806), .Y(n_792) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g797 ( .A1(n_798), .A2(n_801), .B1(n_803), .B2(n_805), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_799), .B(n_800), .Y(n_798) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
NOR2xp33_ASAP7_75t_L g806 ( .A(n_807), .B(n_811), .Y(n_806) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
INVxp67_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_816), .B(n_817), .Y(n_815) );
NOR2xp33_ASAP7_75t_L g821 ( .A(n_822), .B(n_823), .Y(n_821) );
HB1xp67_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx2_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
endmodule