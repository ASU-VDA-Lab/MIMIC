module fake_jpeg_11345_n_40 (n_3, n_2, n_1, n_0, n_4, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

AND2x2_ASAP7_75t_SL g6 ( 
.A(n_4),
.B(n_0),
.Y(n_6)
);

NOR2xp33_ASAP7_75t_L g7 ( 
.A(n_0),
.B(n_1),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_2),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

BUFx12f_ASAP7_75t_L g10 ( 
.A(n_4),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx2_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g13 ( 
.A(n_6),
.B(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_13),
.Y(n_20)
);

INVx2_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx3_ASAP7_75t_SL g15 ( 
.A(n_11),
.Y(n_15)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_15),
.A2(n_16),
.B1(n_10),
.B2(n_6),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

AND2x6_ASAP7_75t_L g19 ( 
.A(n_17),
.B(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_18),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_19),
.B(n_7),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_22),
.B(n_14),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g28 ( 
.A(n_23),
.B(n_20),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx5p33_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_23),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_29),
.B(n_25),
.Y(n_32)
);

OAI21xp5_ASAP7_75t_SL g35 ( 
.A1(n_32),
.A2(n_34),
.B(n_30),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g36 ( 
.A(n_33),
.B(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.C(n_29),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_37),
.B(n_15),
.C(n_12),
.Y(n_38)
);

AOI322xp5_ASAP7_75t_L g39 ( 
.A1(n_38),
.A2(n_3),
.A3(n_5),
.B1(n_10),
.B2(n_16),
.C1(n_17),
.C2(n_25),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_39),
.B(n_3),
.Y(n_40)
);


endmodule