module fake_ariane_623_n_872 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_187, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_188, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_186, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_872);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_187;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_188;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_186;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_872;

wire n_295;
wire n_356;
wire n_556;
wire n_190;
wire n_698;
wire n_695;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_830;
wire n_691;
wire n_404;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_836;
wire n_541;
wire n_499;
wire n_789;
wire n_788;
wire n_850;
wire n_771;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_421;
wire n_245;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_525;
wire n_806;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_817;
wire n_244;
wire n_643;
wire n_679;
wire n_226;
wire n_781;
wire n_261;
wire n_220;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_819;
wire n_286;
wire n_443;
wire n_586;
wire n_864;
wire n_686;
wire n_605;
wire n_776;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_826;
wire n_524;
wire n_391;
wire n_349;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_807;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_802;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_870;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_790;
wire n_857;
wire n_363;
wire n_720;
wire n_354;
wire n_813;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_338;
wire n_285;
wire n_473;
wire n_801;
wire n_202;
wire n_193;
wire n_761;
wire n_733;
wire n_818;
wire n_500;
wire n_754;
wire n_336;
wire n_779;
wire n_665;
wire n_731;
wire n_871;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_829;
wire n_668;
wire n_339;
wire n_758;
wire n_738;
wire n_833;
wire n_672;
wire n_487;
wire n_740;
wire n_422;
wire n_648;
wire n_784;
wire n_269;
wire n_597;
wire n_816;
wire n_855;
wire n_259;
wire n_835;
wire n_808;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_814;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_858;
wire n_242;
wire n_645;
wire n_309;
wire n_320;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_822;
wire n_344;
wire n_381;
wire n_795;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_840;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_253;
wire n_561;
wire n_770;
wire n_218;
wire n_821;
wire n_839;
wire n_271;
wire n_507;
wire n_465;
wire n_486;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_825;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_787;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_786;
wire n_510;
wire n_831;
wire n_256;
wire n_868;
wire n_326;
wire n_681;
wire n_778;
wire n_227;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_689;
wire n_694;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_727;
wire n_699;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_823;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_859;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_863;
wire n_303;
wire n_671;
wire n_442;
wire n_777;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_843;
wire n_511;
wire n_611;
wire n_365;
wire n_238;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_775;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_869;
wire n_846;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_844;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_838;
wire n_237;
wire n_780;
wire n_861;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_810;
wire n_723;
wire n_658;
wire n_616;
wire n_617;
wire n_630;
wire n_705;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_809;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_772;
wire n_747;
wire n_847;
wire n_371;
wire n_845;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_865;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_860;
wire n_249;
wire n_534;
wire n_355;
wire n_212;
wire n_444;
wire n_609;
wire n_278;
wire n_851;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_842;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_519;
wire n_384;
wire n_468;
wire n_853;
wire n_526;
wire n_716;
wire n_742;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_798;
wire n_769;
wire n_820;
wire n_577;
wire n_407;
wire n_774;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_832;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_848;
wire n_804;
wire n_280;
wire n_215;
wire n_252;
wire n_629;
wire n_664;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_794;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_768;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_834;
wire n_389;
wire n_800;
wire n_657;
wire n_513;
wire n_837;
wire n_288;
wire n_812;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_862;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_785;
wire n_827;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_292;
wire n_793;
wire n_852;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_866;
wire n_246;
wire n_517;
wire n_530;
wire n_792;
wire n_824;
wire n_428;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_773;
wire n_317;
wire n_867;
wire n_243;
wire n_803;
wire n_329;
wire n_718;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_815;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_632;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_782;
wire n_856;
wire n_425;
wire n_431;
wire n_811;
wire n_508;
wire n_624;
wire n_791;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_849;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_797;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_828;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_799;
wire n_558;
wire n_592;
wire n_397;
wire n_841;
wire n_854;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_573;
wire n_796;
wire n_805;
wire n_531;
wire n_783;
wire n_675;

INVx1_ASAP7_75t_L g189 ( 
.A(n_169),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_25),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_52),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_108),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_50),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_13),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_3),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_80),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_24),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_26),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_103),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_137),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_36),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_116),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_178),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_40),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_119),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_43),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_84),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_148),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_57),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_167),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_12),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_145),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_16),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_186),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_65),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g216 ( 
.A(n_21),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g217 ( 
.A(n_9),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_133),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_11),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_20),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_66),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_123),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_9),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_106),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g225 ( 
.A(n_156),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_183),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_138),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_49),
.Y(n_229)
);

INVx2_ASAP7_75t_SL g230 ( 
.A(n_126),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_158),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_67),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_111),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

INVx1_ASAP7_75t_SL g236 ( 
.A(n_55),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_51),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_157),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_69),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_151),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_94),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_7),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_44),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_64),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_144),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_68),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_17),
.Y(n_247)
);

INVx2_ASAP7_75t_SL g248 ( 
.A(n_110),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_47),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_1),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_86),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_173),
.Y(n_252)
);

BUFx3_ASAP7_75t_L g253 ( 
.A(n_98),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_93),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_81),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_135),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_46),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_166),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_146),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_59),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_96),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_15),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_31),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_5),
.Y(n_264)
);

HB1xp67_ASAP7_75t_L g265 ( 
.A(n_8),
.Y(n_265)
);

BUFx12f_ASAP7_75t_L g266 ( 
.A(n_217),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

BUFx3_ASAP7_75t_L g268 ( 
.A(n_225),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_223),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_216),
.Y(n_270)
);

OAI21x1_ASAP7_75t_L g271 ( 
.A1(n_196),
.A2(n_23),
.B(n_22),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_192),
.B(n_0),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_189),
.B(n_202),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_225),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_217),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g277 ( 
.A(n_253),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_204),
.B(n_0),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g279 ( 
.A(n_216),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_212),
.Y(n_280)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

INVx4_ASAP7_75t_L g282 ( 
.A(n_216),
.Y(n_282)
);

AOI22x1_ASAP7_75t_SL g283 ( 
.A1(n_214),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_283)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_253),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_232),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g286 ( 
.A(n_216),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_233),
.B(n_2),
.Y(n_287)
);

BUFx2_ASAP7_75t_L g288 ( 
.A(n_194),
.Y(n_288)
);

OA21x2_ASAP7_75t_L g289 ( 
.A1(n_240),
.A2(n_4),
.B(n_5),
.Y(n_289)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_243),
.A2(n_255),
.B(n_251),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

BUFx8_ASAP7_75t_L g292 ( 
.A(n_230),
.Y(n_292)
);

BUFx6f_ASAP7_75t_L g293 ( 
.A(n_235),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_256),
.B(n_4),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_259),
.B(n_6),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g296 ( 
.A(n_235),
.Y(n_296)
);

BUFx8_ASAP7_75t_SL g297 ( 
.A(n_229),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_195),
.Y(n_298)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_196),
.Y(n_299)
);

BUFx2_ASAP7_75t_L g300 ( 
.A(n_211),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_235),
.Y(n_301)
);

BUFx2_ASAP7_75t_L g302 ( 
.A(n_213),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_237),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_219),
.Y(n_304)
);

BUFx8_ASAP7_75t_SL g305 ( 
.A(n_239),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_242),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_237),
.Y(n_307)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_209),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_248),
.Y(n_309)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_190),
.Y(n_310)
);

AND2x4_ASAP7_75t_L g311 ( 
.A(n_197),
.B(n_6),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_247),
.Y(n_312)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_262),
.B(n_7),
.Y(n_313)
);

HB1xp67_ASAP7_75t_L g314 ( 
.A(n_191),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_236),
.Y(n_315)
);

BUFx8_ASAP7_75t_L g316 ( 
.A(n_193),
.Y(n_316)
);

OA21x2_ASAP7_75t_L g317 ( 
.A1(n_198),
.A2(n_8),
.B(n_10),
.Y(n_317)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_272),
.C(n_311),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_297),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_282),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_297),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_269),
.Y(n_322)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_268),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_305),
.Y(n_324)
);

NAND2xp33_ASAP7_75t_R g325 ( 
.A(n_288),
.B(n_199),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_305),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_316),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_315),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_R g329 ( 
.A(n_298),
.B(n_200),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_274),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_R g332 ( 
.A(n_304),
.B(n_263),
.Y(n_332)
);

CKINVDCx20_ASAP7_75t_R g333 ( 
.A(n_316),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_314),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_266),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_303),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_266),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_310),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_281),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_R g340 ( 
.A(n_312),
.B(n_201),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_R g342 ( 
.A(n_315),
.B(n_261),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_310),
.Y(n_343)
);

INVx3_ASAP7_75t_L g344 ( 
.A(n_268),
.Y(n_344)
);

BUFx2_ASAP7_75t_L g345 ( 
.A(n_288),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_310),
.B(n_203),
.Y(n_346)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_270),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_300),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_300),
.Y(n_350)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_283),
.B(n_10),
.Y(n_351)
);

AOI21x1_ASAP7_75t_L g352 ( 
.A1(n_290),
.A2(n_206),
.B(n_205),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_302),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_302),
.Y(n_354)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_207),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_R g356 ( 
.A(n_277),
.B(n_260),
.Y(n_356)
);

NAND2xp33_ASAP7_75t_R g357 ( 
.A(n_317),
.B(n_208),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_275),
.Y(n_358)
);

NOR2xp67_ASAP7_75t_L g359 ( 
.A(n_282),
.B(n_210),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_277),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_292),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_275),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_284),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_292),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_292),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_285),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_285),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_284),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_282),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_308),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_R g371 ( 
.A(n_280),
.B(n_215),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_347),
.B(n_267),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_336),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_319),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_328),
.B(n_309),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_328),
.B(n_311),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_348),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_341),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_362),
.Y(n_380)
);

INVx3_ASAP7_75t_L g381 ( 
.A(n_323),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_338),
.B(n_307),
.Y(n_382)
);

INVx2_ASAP7_75t_SL g383 ( 
.A(n_366),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_323),
.B(n_309),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_344),
.B(n_311),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_363),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_367),
.B(n_313),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_320),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_343),
.B(n_307),
.Y(n_389)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_344),
.B(n_308),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_342),
.B(n_313),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_368),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_369),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_346),
.B(n_308),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_360),
.B(n_276),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g397 ( 
.A(n_318),
.B(n_308),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_322),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_355),
.B(n_299),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_330),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_371),
.B(n_278),
.Y(n_401)
);

INVxp67_ASAP7_75t_SL g402 ( 
.A(n_359),
.Y(n_402)
);

BUFx3_ASAP7_75t_L g403 ( 
.A(n_339),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_348),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_329),
.B(n_299),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_352),
.B(n_287),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_332),
.B(n_299),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_348),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g409 ( 
.A(n_345),
.B(n_290),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_340),
.B(n_290),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_371),
.B(n_356),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_348),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_361),
.B(n_294),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_334),
.Y(n_414)
);

INVx2_ASAP7_75t_L g415 ( 
.A(n_350),
.Y(n_415)
);

AO221x1_ASAP7_75t_L g416 ( 
.A1(n_357),
.A2(n_317),
.B1(n_289),
.B2(n_270),
.C(n_286),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_353),
.B(n_295),
.Y(n_417)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_364),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_354),
.Y(n_419)
);

AND2x2_ASAP7_75t_L g420 ( 
.A(n_365),
.B(n_317),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_331),
.B(n_218),
.Y(n_421)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_325),
.A2(n_246),
.B1(n_221),
.B2(n_222),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_335),
.B(n_289),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_349),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_337),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_SL g426 ( 
.A(n_325),
.B(n_220),
.Y(n_426)
);

INVx1_ASAP7_75t_SL g427 ( 
.A(n_321),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_327),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_333),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_324),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_351),
.B(n_224),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_357),
.B(n_270),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_326),
.B(n_226),
.Y(n_433)
);

BUFx2_ASAP7_75t_R g434 ( 
.A(n_319),
.Y(n_434)
);

NAND2xp33_ASAP7_75t_L g435 ( 
.A(n_338),
.B(n_227),
.Y(n_435)
);

NOR3xp33_ASAP7_75t_L g436 ( 
.A(n_318),
.B(n_271),
.C(n_231),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_328),
.B(n_228),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_348),
.Y(n_438)
);

A2O1A1Ixp33_ASAP7_75t_L g439 ( 
.A1(n_385),
.A2(n_271),
.B(n_234),
.C(n_257),
.Y(n_439)
);

AOI22xp33_ASAP7_75t_L g440 ( 
.A1(n_416),
.A2(n_289),
.B1(n_270),
.B2(n_286),
.Y(n_440)
);

NOR2x2_ASAP7_75t_L g441 ( 
.A(n_415),
.B(n_11),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_385),
.B(n_238),
.Y(n_442)
);

INVx5_ASAP7_75t_L g443 ( 
.A(n_378),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g444 ( 
.A(n_409),
.B(n_241),
.Y(n_444)
);

INVx3_ASAP7_75t_L g445 ( 
.A(n_381),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_393),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_SL g447 ( 
.A(n_383),
.B(n_244),
.Y(n_447)
);

OR2x6_ASAP7_75t_L g448 ( 
.A(n_403),
.B(n_286),
.Y(n_448)
);

AND2x6_ASAP7_75t_SL g449 ( 
.A(n_431),
.B(n_12),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_398),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_411),
.B(n_245),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_374),
.Y(n_452)
);

INVx2_ASAP7_75t_SL g453 ( 
.A(n_414),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_375),
.Y(n_454)
);

OAI21xp5_ASAP7_75t_L g455 ( 
.A1(n_406),
.A2(n_252),
.B(n_249),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_382),
.B(n_13),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_379),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_388),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_376),
.B(n_254),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g460 ( 
.A(n_427),
.Y(n_460)
);

INVx2_ASAP7_75t_SL g461 ( 
.A(n_372),
.Y(n_461)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_400),
.Y(n_462)
);

NOR2x2_ASAP7_75t_L g463 ( 
.A(n_424),
.B(n_14),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_436),
.A2(n_286),
.B1(n_296),
.B2(n_293),
.Y(n_464)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_436),
.A2(n_301),
.B1(n_296),
.B2(n_293),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_376),
.B(n_258),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_373),
.Y(n_467)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_395),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_389),
.B(n_279),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_406),
.A2(n_301),
.B(n_296),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_377),
.A2(n_437),
.B1(n_397),
.B2(n_401),
.Y(n_471)
);

AND2x2_ASAP7_75t_L g472 ( 
.A(n_419),
.B(n_14),
.Y(n_472)
);

AND2x2_ASAP7_75t_L g473 ( 
.A(n_417),
.B(n_15),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_381),
.B(n_16),
.Y(n_474)
);

INVx3_ASAP7_75t_L g475 ( 
.A(n_438),
.Y(n_475)
);

NAND2xp5_ASAP7_75t_SL g476 ( 
.A(n_422),
.B(n_279),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_397),
.A2(n_301),
.B1(n_296),
.B2(n_293),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_437),
.B(n_279),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_405),
.B(n_279),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_407),
.B(n_279),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_418),
.B(n_291),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_R g483 ( 
.A(n_430),
.B(n_27),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_399),
.B(n_291),
.Y(n_484)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_423),
.A2(n_402),
.B1(n_420),
.B2(n_391),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_418),
.B(n_291),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_386),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_392),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_384),
.B(n_291),
.Y(n_489)
);

BUFx6f_ASAP7_75t_L g490 ( 
.A(n_378),
.Y(n_490)
);

CKINVDCx5p33_ASAP7_75t_R g491 ( 
.A(n_434),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_408),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_384),
.B(n_291),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_418),
.B(n_293),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_390),
.Y(n_495)
);

INVx2_ASAP7_75t_L g496 ( 
.A(n_404),
.Y(n_496)
);

INVx2_ASAP7_75t_L g497 ( 
.A(n_412),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_402),
.B(n_293),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_418),
.B(n_296),
.Y(n_499)
);

NAND2xp33_ASAP7_75t_L g500 ( 
.A(n_410),
.B(n_301),
.Y(n_500)
);

AND2x2_ASAP7_75t_L g501 ( 
.A(n_431),
.B(n_17),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_390),
.B(n_301),
.Y(n_502)
);

INVx1_ASAP7_75t_SL g503 ( 
.A(n_428),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_394),
.B(n_18),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_378),
.Y(n_505)
);

BUFx12f_ASAP7_75t_L g506 ( 
.A(n_378),
.Y(n_506)
);

O2A1O1Ixp33_ASAP7_75t_L g507 ( 
.A1(n_387),
.A2(n_18),
.B(n_19),
.C(n_28),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_425),
.B(n_29),
.Y(n_508)
);

BUFx3_ASAP7_75t_L g509 ( 
.A(n_429),
.Y(n_509)
);

A2O1A1Ixp33_ASAP7_75t_L g510 ( 
.A1(n_455),
.A2(n_394),
.B(n_426),
.C(n_435),
.Y(n_510)
);

OAI21xp33_ASAP7_75t_L g511 ( 
.A1(n_456),
.A2(n_413),
.B(n_433),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_501),
.B(n_396),
.Y(n_512)
);

INVx1_ASAP7_75t_SL g513 ( 
.A(n_460),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_471),
.B(n_421),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_442),
.A2(n_432),
.B1(n_438),
.B2(n_19),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_450),
.B(n_473),
.Y(n_516)
);

AOI21xp5_ASAP7_75t_L g517 ( 
.A1(n_478),
.A2(n_438),
.B(n_32),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_456),
.B(n_438),
.Y(n_518)
);

OAI21xp33_ASAP7_75t_L g519 ( 
.A1(n_474),
.A2(n_30),
.B(n_33),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_467),
.Y(n_520)
);

AOI21xp5_ASAP7_75t_L g521 ( 
.A1(n_495),
.A2(n_34),
.B(n_35),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_479),
.B(n_37),
.Y(n_522)
);

BUFx4f_ASAP7_75t_L g523 ( 
.A(n_448),
.Y(n_523)
);

AOI221xp5_ASAP7_75t_L g524 ( 
.A1(n_461),
.A2(n_472),
.B1(n_487),
.B2(n_488),
.C(n_507),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_446),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g526 ( 
.A1(n_459),
.A2(n_38),
.B(n_39),
.Y(n_526)
);

AOI21xp33_ASAP7_75t_L g527 ( 
.A1(n_444),
.A2(n_41),
.B(n_42),
.Y(n_527)
);

O2A1O1Ixp33_ASAP7_75t_SL g528 ( 
.A1(n_451),
.A2(n_45),
.B(n_48),
.C(n_53),
.Y(n_528)
);

CKINVDCx6p67_ASAP7_75t_R g529 ( 
.A(n_454),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g530 ( 
.A1(n_466),
.A2(n_54),
.B(n_56),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_SL g531 ( 
.A(n_453),
.B(n_58),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_506),
.Y(n_532)
);

INVx1_ASAP7_75t_SL g533 ( 
.A(n_503),
.Y(n_533)
);

NAND2xp5_ASAP7_75t_SL g534 ( 
.A(n_485),
.B(n_60),
.Y(n_534)
);

AOI21xp5_ASAP7_75t_L g535 ( 
.A1(n_469),
.A2(n_61),
.B(n_62),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_462),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_SL g537 ( 
.A(n_508),
.B(n_63),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_504),
.A2(n_70),
.B(n_71),
.Y(n_538)
);

INVx4_ASAP7_75t_L g539 ( 
.A(n_448),
.Y(n_539)
);

OR2x6_ASAP7_75t_L g540 ( 
.A(n_448),
.B(n_72),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_L g541 ( 
.A1(n_445),
.A2(n_474),
.B1(n_475),
.B2(n_465),
.Y(n_541)
);

BUFx6f_ASAP7_75t_L g542 ( 
.A(n_490),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_452),
.Y(n_543)
);

INVx3_ASAP7_75t_L g544 ( 
.A(n_509),
.Y(n_544)
);

OAI22xp5_ASAP7_75t_L g545 ( 
.A1(n_445),
.A2(n_73),
.B1(n_74),
.B2(n_75),
.Y(n_545)
);

A2O1A1Ixp33_ASAP7_75t_L g546 ( 
.A1(n_507),
.A2(n_76),
.B(n_77),
.C(n_78),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_457),
.Y(n_547)
);

BUFx6f_ASAP7_75t_L g548 ( 
.A(n_490),
.Y(n_548)
);

AOI21xp5_ASAP7_75t_L g549 ( 
.A1(n_470),
.A2(n_79),
.B(n_82),
.Y(n_549)
);

O2A1O1Ixp5_ASAP7_75t_L g550 ( 
.A1(n_439),
.A2(n_83),
.B(n_85),
.C(n_87),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_491),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g552 ( 
.A(n_447),
.B(n_188),
.Y(n_552)
);

BUFx6f_ASAP7_75t_SL g553 ( 
.A(n_463),
.Y(n_553)
);

O2A1O1Ixp33_ASAP7_75t_L g554 ( 
.A1(n_458),
.A2(n_88),
.B(n_89),
.C(n_90),
.Y(n_554)
);

NAND2xp5_ASAP7_75t_L g555 ( 
.A(n_468),
.B(n_91),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_483),
.Y(n_556)
);

INVx4_ASAP7_75t_L g557 ( 
.A(n_443),
.Y(n_557)
);

OAI22x1_ASAP7_75t_L g558 ( 
.A1(n_441),
.A2(n_92),
.B1(n_95),
.B2(n_97),
.Y(n_558)
);

AND2x6_ASAP7_75t_L g559 ( 
.A(n_475),
.B(n_99),
.Y(n_559)
);

BUFx12f_ASAP7_75t_L g560 ( 
.A(n_449),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_496),
.Y(n_561)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_470),
.A2(n_100),
.B(n_101),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_484),
.A2(n_102),
.B(n_104),
.Y(n_563)
);

INVx2_ASAP7_75t_SL g564 ( 
.A(n_508),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_490),
.Y(n_565)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_498),
.A2(n_105),
.B(n_107),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_497),
.Y(n_567)
);

OAI22xp5_ASAP7_75t_L g568 ( 
.A1(n_465),
.A2(n_109),
.B1(n_112),
.B2(n_113),
.Y(n_568)
);

A2O1A1Ixp33_ASAP7_75t_L g569 ( 
.A1(n_464),
.A2(n_114),
.B(n_115),
.C(n_117),
.Y(n_569)
);

OR2x6_ASAP7_75t_L g570 ( 
.A(n_540),
.B(n_482),
.Y(n_570)
);

INVx2_ASAP7_75t_SL g571 ( 
.A(n_523),
.Y(n_571)
);

AOI22x1_ASAP7_75t_L g572 ( 
.A1(n_517),
.A2(n_505),
.B1(n_490),
.B2(n_492),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_529),
.Y(n_573)
);

INVx2_ASAP7_75t_L g574 ( 
.A(n_536),
.Y(n_574)
);

CKINVDCx20_ASAP7_75t_R g575 ( 
.A(n_551),
.Y(n_575)
);

OAI21x1_ASAP7_75t_L g576 ( 
.A1(n_550),
.A2(n_440),
.B(n_502),
.Y(n_576)
);

BUFx6f_ASAP7_75t_L g577 ( 
.A(n_542),
.Y(n_577)
);

CKINVDCx16_ASAP7_75t_R g578 ( 
.A(n_553),
.Y(n_578)
);

BUFx8_ASAP7_75t_SL g579 ( 
.A(n_560),
.Y(n_579)
);

AO21x2_ASAP7_75t_L g580 ( 
.A1(n_518),
.A2(n_500),
.B(n_476),
.Y(n_580)
);

AO21x2_ASAP7_75t_L g581 ( 
.A1(n_534),
.A2(n_481),
.B(n_480),
.Y(n_581)
);

AOI22xp5_ASAP7_75t_L g582 ( 
.A1(n_556),
.A2(n_499),
.B1(n_494),
.B2(n_486),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_549),
.A2(n_440),
.B(n_464),
.Y(n_583)
);

INVx3_ASAP7_75t_L g584 ( 
.A(n_542),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_543),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_562),
.A2(n_493),
.B(n_489),
.Y(n_586)
);

AO21x2_ASAP7_75t_L g587 ( 
.A1(n_510),
.A2(n_483),
.B(n_477),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_542),
.B(n_443),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_541),
.A2(n_477),
.B(n_443),
.Y(n_589)
);

BUFx12f_ASAP7_75t_L g590 ( 
.A(n_532),
.Y(n_590)
);

AO21x1_ASAP7_75t_L g591 ( 
.A1(n_515),
.A2(n_443),
.B(n_120),
.Y(n_591)
);

BUFx12f_ASAP7_75t_L g592 ( 
.A(n_540),
.Y(n_592)
);

BUFx3_ASAP7_75t_L g593 ( 
.A(n_544),
.Y(n_593)
);

AO21x2_ASAP7_75t_L g594 ( 
.A1(n_519),
.A2(n_118),
.B(n_121),
.Y(n_594)
);

INVx3_ASAP7_75t_L g595 ( 
.A(n_548),
.Y(n_595)
);

INVx5_ASAP7_75t_L g596 ( 
.A(n_559),
.Y(n_596)
);

INVx5_ASAP7_75t_SL g597 ( 
.A(n_548),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_516),
.B(n_122),
.Y(n_598)
);

NAND2x1p5_ASAP7_75t_L g599 ( 
.A(n_548),
.B(n_124),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_547),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_520),
.Y(n_601)
);

INVx3_ASAP7_75t_L g602 ( 
.A(n_559),
.Y(n_602)
);

OA21x2_ASAP7_75t_L g603 ( 
.A1(n_546),
.A2(n_125),
.B(n_127),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_513),
.Y(n_604)
);

AND2x2_ASAP7_75t_L g605 ( 
.A(n_525),
.B(n_128),
.Y(n_605)
);

AO21x2_ASAP7_75t_L g606 ( 
.A1(n_514),
.A2(n_130),
.B(n_131),
.Y(n_606)
);

OAI21x1_ASAP7_75t_SL g607 ( 
.A1(n_522),
.A2(n_132),
.B(n_134),
.Y(n_607)
);

INVx1_ASAP7_75t_SL g608 ( 
.A(n_533),
.Y(n_608)
);

AO21x2_ASAP7_75t_L g609 ( 
.A1(n_527),
.A2(n_136),
.B(n_139),
.Y(n_609)
);

AOI22x1_ASAP7_75t_L g610 ( 
.A1(n_526),
.A2(n_140),
.B1(n_141),
.B2(n_142),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_561),
.Y(n_611)
);

INVx2_ASAP7_75t_L g612 ( 
.A(n_567),
.Y(n_612)
);

OAI21xp5_ASAP7_75t_L g613 ( 
.A1(n_511),
.A2(n_143),
.B(n_147),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_565),
.Y(n_614)
);

OAI21x1_ASAP7_75t_L g615 ( 
.A1(n_530),
.A2(n_149),
.B(n_150),
.Y(n_615)
);

INVx2_ASAP7_75t_L g616 ( 
.A(n_555),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_539),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_557),
.Y(n_618)
);

AND2x4_ASAP7_75t_L g619 ( 
.A(n_564),
.B(n_512),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_559),
.Y(n_620)
);

OAI21x1_ASAP7_75t_L g621 ( 
.A1(n_572),
.A2(n_535),
.B(n_538),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_604),
.B(n_558),
.Y(n_622)
);

AOI22xp33_ASAP7_75t_SL g623 ( 
.A1(n_592),
.A2(n_568),
.B1(n_552),
.B2(n_559),
.Y(n_623)
);

OAI21xp5_ASAP7_75t_L g624 ( 
.A1(n_583),
.A2(n_524),
.B(n_521),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_612),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_593),
.Y(n_626)
);

INVx4_ASAP7_75t_L g627 ( 
.A(n_590),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_575),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_601),
.Y(n_629)
);

INVx6_ASAP7_75t_L g630 ( 
.A(n_590),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_612),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_611),
.Y(n_632)
);

AOI22xp33_ASAP7_75t_L g633 ( 
.A1(n_592),
.A2(n_537),
.B1(n_531),
.B2(n_545),
.Y(n_633)
);

OAI22xp5_ASAP7_75t_L g634 ( 
.A1(n_598),
.A2(n_569),
.B1(n_554),
.B2(n_566),
.Y(n_634)
);

AOI22xp33_ASAP7_75t_L g635 ( 
.A1(n_611),
.A2(n_563),
.B1(n_528),
.B2(n_154),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_574),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_574),
.Y(n_637)
);

OAI21x1_ASAP7_75t_L g638 ( 
.A1(n_586),
.A2(n_152),
.B(n_153),
.Y(n_638)
);

OAI22xp5_ASAP7_75t_L g639 ( 
.A1(n_598),
.A2(n_155),
.B1(n_160),
.B2(n_161),
.Y(n_639)
);

CKINVDCx6p67_ASAP7_75t_R g640 ( 
.A(n_578),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_596),
.B(n_162),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_585),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_585),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_SL g644 ( 
.A1(n_596),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_644)
);

AOI21xp33_ASAP7_75t_L g645 ( 
.A1(n_587),
.A2(n_168),
.B(n_170),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_600),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_600),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_605),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_575),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_597),
.Y(n_650)
);

OAI21x1_ASAP7_75t_L g651 ( 
.A1(n_586),
.A2(n_171),
.B(n_172),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_608),
.B(n_187),
.Y(n_652)
);

AOI21x1_ASAP7_75t_L g653 ( 
.A1(n_591),
.A2(n_174),
.B(n_175),
.Y(n_653)
);

OAI21x1_ASAP7_75t_L g654 ( 
.A1(n_576),
.A2(n_176),
.B(n_177),
.Y(n_654)
);

BUFx6f_ASAP7_75t_L g655 ( 
.A(n_577),
.Y(n_655)
);

INVx2_ASAP7_75t_L g656 ( 
.A(n_614),
.Y(n_656)
);

OR2x6_ASAP7_75t_L g657 ( 
.A(n_571),
.B(n_179),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_605),
.Y(n_658)
);

AOI21x1_ASAP7_75t_L g659 ( 
.A1(n_591),
.A2(n_180),
.B(n_181),
.Y(n_659)
);

BUFx10_ASAP7_75t_L g660 ( 
.A(n_571),
.Y(n_660)
);

NAND2x1p5_ASAP7_75t_L g661 ( 
.A(n_596),
.B(n_182),
.Y(n_661)
);

INVx1_ASAP7_75t_SL g662 ( 
.A(n_604),
.Y(n_662)
);

NOR2x1p5_ASAP7_75t_L g663 ( 
.A(n_640),
.B(n_573),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_629),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_628),
.Y(n_665)
);

INVx1_ASAP7_75t_L g666 ( 
.A(n_631),
.Y(n_666)
);

INVx3_ASAP7_75t_L g667 ( 
.A(n_655),
.Y(n_667)
);

INVx1_ASAP7_75t_L g668 ( 
.A(n_625),
.Y(n_668)
);

NAND2xp33_ASAP7_75t_R g669 ( 
.A(n_657),
.B(n_602),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_632),
.Y(n_670)
);

AND2x2_ASAP7_75t_L g671 ( 
.A(n_622),
.B(n_593),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_662),
.B(n_619),
.Y(n_672)
);

INVxp33_ASAP7_75t_L g673 ( 
.A(n_626),
.Y(n_673)
);

AND2x4_ASAP7_75t_L g674 ( 
.A(n_650),
.B(n_595),
.Y(n_674)
);

INVx1_ASAP7_75t_SL g675 ( 
.A(n_662),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_636),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_637),
.Y(n_677)
);

CKINVDCx11_ASAP7_75t_R g678 ( 
.A(n_660),
.Y(n_678)
);

OAI222xp33_ASAP7_75t_L g679 ( 
.A1(n_623),
.A2(n_596),
.B1(n_570),
.B2(n_602),
.C1(n_620),
.C2(n_599),
.Y(n_679)
);

OAI22xp5_ASAP7_75t_L g680 ( 
.A1(n_648),
.A2(n_596),
.B1(n_613),
.B2(n_602),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_649),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_658),
.B(n_614),
.Y(n_682)
);

BUFx3_ASAP7_75t_L g683 ( 
.A(n_630),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_642),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_643),
.Y(n_685)
);

BUFx12f_ASAP7_75t_L g686 ( 
.A(n_627),
.Y(n_686)
);

AO31x2_ASAP7_75t_L g687 ( 
.A1(n_634),
.A2(n_616),
.A3(n_639),
.B(n_647),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g688 ( 
.A(n_646),
.B(n_584),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_L g689 ( 
.A(n_657),
.B(n_619),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_656),
.Y(n_690)
);

CKINVDCx16_ASAP7_75t_R g691 ( 
.A(n_627),
.Y(n_691)
);

AND2x2_ASAP7_75t_L g692 ( 
.A(n_657),
.B(n_619),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_655),
.Y(n_693)
);

AOI22xp5_ASAP7_75t_L g694 ( 
.A1(n_639),
.A2(n_570),
.B1(n_587),
.B2(n_573),
.Y(n_694)
);

AND2x2_ASAP7_75t_L g695 ( 
.A(n_660),
.B(n_617),
.Y(n_695)
);

AND2x2_ASAP7_75t_L g696 ( 
.A(n_652),
.B(n_570),
.Y(n_696)
);

AND2x2_ASAP7_75t_L g697 ( 
.A(n_630),
.B(n_570),
.Y(n_697)
);

AND2x2_ASAP7_75t_L g698 ( 
.A(n_650),
.B(n_597),
.Y(n_698)
);

NAND3xp33_ASAP7_75t_SL g699 ( 
.A(n_633),
.B(n_582),
.C(n_599),
.Y(n_699)
);

CKINVDCx5p33_ASAP7_75t_R g700 ( 
.A(n_655),
.Y(n_700)
);

AND2x2_ASAP7_75t_L g701 ( 
.A(n_644),
.B(n_597),
.Y(n_701)
);

INVx1_ASAP7_75t_SL g702 ( 
.A(n_641),
.Y(n_702)
);

BUFx2_ASAP7_75t_SL g703 ( 
.A(n_634),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_641),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_624),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_L g706 ( 
.A(n_624),
.B(n_584),
.Y(n_706)
);

AOI22xp5_ASAP7_75t_L g707 ( 
.A1(n_645),
.A2(n_587),
.B1(n_594),
.B2(n_603),
.Y(n_707)
);

OR2x6_ASAP7_75t_L g708 ( 
.A(n_661),
.B(n_589),
.Y(n_708)
);

OR2x6_ASAP7_75t_L g709 ( 
.A(n_661),
.B(n_589),
.Y(n_709)
);

AOI221xp5_ASAP7_75t_L g710 ( 
.A1(n_645),
.A2(n_607),
.B1(n_594),
.B2(n_606),
.C(n_609),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_653),
.Y(n_711)
);

BUFx3_ASAP7_75t_L g712 ( 
.A(n_638),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_SL g713 ( 
.A(n_635),
.B(n_599),
.C(n_588),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_664),
.Y(n_714)
);

INVx1_ASAP7_75t_L g715 ( 
.A(n_666),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_670),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_684),
.Y(n_717)
);

BUFx6f_ASAP7_75t_L g718 ( 
.A(n_708),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_700),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_676),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_705),
.B(n_703),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_706),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_677),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_685),
.Y(n_724)
);

AOI221xp5_ASAP7_75t_SL g725 ( 
.A1(n_675),
.A2(n_584),
.B1(n_595),
.B2(n_577),
.C(n_659),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_668),
.Y(n_726)
);

INVx3_ASAP7_75t_L g727 ( 
.A(n_712),
.Y(n_727)
);

HB1xp67_ASAP7_75t_L g728 ( 
.A(n_682),
.Y(n_728)
);

AND2x2_ASAP7_75t_L g729 ( 
.A(n_706),
.B(n_606),
.Y(n_729)
);

AOI22xp33_ASAP7_75t_SL g730 ( 
.A1(n_689),
.A2(n_594),
.B1(n_609),
.B2(n_603),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_690),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_687),
.Y(n_732)
);

OR2x2_ASAP7_75t_L g733 ( 
.A(n_672),
.B(n_606),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_687),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_687),
.B(n_577),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_688),
.Y(n_736)
);

AND2x2_ASAP7_75t_L g737 ( 
.A(n_687),
.B(n_577),
.Y(n_737)
);

AO31x2_ASAP7_75t_L g738 ( 
.A1(n_680),
.A2(n_616),
.A3(n_603),
.B(n_609),
.Y(n_738)
);

INVx1_ASAP7_75t_L g739 ( 
.A(n_688),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_673),
.B(n_595),
.Y(n_740)
);

AND2x2_ASAP7_75t_L g741 ( 
.A(n_671),
.B(n_577),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_708),
.Y(n_742)
);

NOR2x1_ASAP7_75t_L g743 ( 
.A(n_663),
.B(n_580),
.Y(n_743)
);

CKINVDCx20_ASAP7_75t_R g744 ( 
.A(n_678),
.Y(n_744)
);

AND2x2_ASAP7_75t_L g745 ( 
.A(n_673),
.B(n_583),
.Y(n_745)
);

AND2x2_ASAP7_75t_L g746 ( 
.A(n_693),
.B(n_654),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_708),
.Y(n_747)
);

AND2x2_ASAP7_75t_L g748 ( 
.A(n_692),
.B(n_580),
.Y(n_748)
);

INVxp67_ASAP7_75t_L g749 ( 
.A(n_695),
.Y(n_749)
);

AND2x2_ASAP7_75t_L g750 ( 
.A(n_694),
.B(n_580),
.Y(n_750)
);

AND2x4_ASAP7_75t_L g751 ( 
.A(n_709),
.B(n_651),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_689),
.B(n_597),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_667),
.B(n_576),
.Y(n_753)
);

INVx4_ASAP7_75t_R g754 ( 
.A(n_719),
.Y(n_754)
);

AND2x2_ASAP7_75t_L g755 ( 
.A(n_721),
.B(n_691),
.Y(n_755)
);

HB1xp67_ASAP7_75t_L g756 ( 
.A(n_722),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_715),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_718),
.B(n_709),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_715),
.Y(n_759)
);

HB1xp67_ASAP7_75t_L g760 ( 
.A(n_722),
.Y(n_760)
);

INVx2_ASAP7_75t_SL g761 ( 
.A(n_727),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_716),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_721),
.B(n_697),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_728),
.B(n_667),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_741),
.B(n_683),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_716),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_736),
.B(n_696),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_741),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_720),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_714),
.Y(n_770)
);

NAND2xp5_ASAP7_75t_L g771 ( 
.A(n_739),
.B(n_704),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_720),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_717),
.Y(n_773)
);

AND2x4_ASAP7_75t_L g774 ( 
.A(n_718),
.B(n_709),
.Y(n_774)
);

NAND2x1p5_ASAP7_75t_L g775 ( 
.A(n_743),
.B(n_702),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_726),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_745),
.Y(n_777)
);

NOR3xp33_ASAP7_75t_L g778 ( 
.A(n_740),
.B(n_699),
.C(n_710),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_756),
.Y(n_779)
);

INVx2_ASAP7_75t_L g780 ( 
.A(n_769),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_768),
.B(n_749),
.Y(n_781)
);

NAND2x1_ASAP7_75t_SL g782 ( 
.A(n_756),
.B(n_735),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_755),
.B(n_719),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_760),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_777),
.B(n_745),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_769),
.Y(n_786)
);

NOR2x1_ASAP7_75t_L g787 ( 
.A(n_764),
.B(n_744),
.Y(n_787)
);

HB1xp67_ASAP7_75t_L g788 ( 
.A(n_777),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_761),
.B(n_737),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_772),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_760),
.B(n_744),
.Y(n_791)
);

INVx2_ASAP7_75t_SL g792 ( 
.A(n_754),
.Y(n_792)
);

HB1xp67_ASAP7_75t_L g793 ( 
.A(n_757),
.Y(n_793)
);

AND2x2_ASAP7_75t_L g794 ( 
.A(n_765),
.B(n_748),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_780),
.Y(n_795)
);

OAI22xp5_ASAP7_75t_L g796 ( 
.A1(n_791),
.A2(n_778),
.B1(n_730),
.B2(n_767),
.Y(n_796)
);

INVxp67_ASAP7_75t_L g797 ( 
.A(n_791),
.Y(n_797)
);

OA222x2_ASAP7_75t_L g798 ( 
.A1(n_782),
.A2(n_733),
.B1(n_771),
.B2(n_747),
.C1(n_742),
.C2(n_669),
.Y(n_798)
);

OAI22xp5_ASAP7_75t_L g799 ( 
.A1(n_787),
.A2(n_773),
.B1(n_770),
.B2(n_707),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_793),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_785),
.B(n_761),
.Y(n_801)
);

OR2x2_ASAP7_75t_L g802 ( 
.A(n_779),
.B(n_776),
.Y(n_802)
);

NAND4xp75_ASAP7_75t_L g803 ( 
.A(n_792),
.B(n_725),
.C(n_701),
.D(n_750),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_783),
.B(n_686),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_780),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_793),
.B(n_759),
.Y(n_806)
);

OAI221xp5_ASAP7_75t_SL g807 ( 
.A1(n_796),
.A2(n_781),
.B1(n_788),
.B2(n_734),
.C(n_710),
.Y(n_807)
);

AOI21xp33_ASAP7_75t_L g808 ( 
.A1(n_796),
.A2(n_784),
.B(n_669),
.Y(n_808)
);

AOI211xp5_ASAP7_75t_SL g809 ( 
.A1(n_799),
.A2(n_797),
.B(n_804),
.C(n_800),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_795),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_806),
.Y(n_811)
);

HB1xp67_ASAP7_75t_L g812 ( 
.A(n_811),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_810),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_809),
.B(n_788),
.Y(n_814)
);

NAND2x1_ASAP7_75t_SL g815 ( 
.A(n_808),
.B(n_789),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_813),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_812),
.B(n_665),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_814),
.B(n_807),
.Y(n_818)
);

AOI211x1_ASAP7_75t_L g819 ( 
.A1(n_818),
.A2(n_799),
.B(n_807),
.C(n_815),
.Y(n_819)
);

AOI211xp5_ASAP7_75t_L g820 ( 
.A1(n_817),
.A2(n_798),
.B(n_699),
.C(n_679),
.Y(n_820)
);

NOR4xp25_ASAP7_75t_L g821 ( 
.A(n_819),
.B(n_816),
.C(n_802),
.D(n_801),
.Y(n_821)
);

AOI211xp5_ASAP7_75t_L g822 ( 
.A1(n_820),
.A2(n_679),
.B(n_681),
.C(n_680),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_819),
.B(n_803),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_821),
.B(n_794),
.Y(n_824)
);

NOR2x1_ASAP7_75t_L g825 ( 
.A(n_823),
.B(n_579),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_822),
.B(n_789),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_823),
.Y(n_827)
);

NOR2x1_ASAP7_75t_L g828 ( 
.A(n_823),
.B(n_579),
.Y(n_828)
);

AND2x2_ASAP7_75t_L g829 ( 
.A(n_821),
.B(n_678),
.Y(n_829)
);

NOR2xp33_ASAP7_75t_L g830 ( 
.A(n_825),
.B(n_789),
.Y(n_830)
);

INVx1_ASAP7_75t_L g831 ( 
.A(n_827),
.Y(n_831)
);

NOR3xp33_ASAP7_75t_L g832 ( 
.A(n_828),
.B(n_618),
.C(n_713),
.Y(n_832)
);

NAND2x1p5_ASAP7_75t_L g833 ( 
.A(n_829),
.B(n_698),
.Y(n_833)
);

NAND5xp2_ASAP7_75t_L g834 ( 
.A(n_824),
.B(n_775),
.C(n_752),
.D(n_746),
.E(n_763),
.Y(n_834)
);

INVxp33_ASAP7_75t_SL g835 ( 
.A(n_826),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_827),
.Y(n_836)
);

AOI222xp33_ASAP7_75t_L g837 ( 
.A1(n_831),
.A2(n_734),
.B1(n_750),
.B2(n_713),
.C1(n_729),
.C2(n_732),
.Y(n_837)
);

BUFx6f_ASAP7_75t_L g838 ( 
.A(n_836),
.Y(n_838)
);

BUFx2_ASAP7_75t_L g839 ( 
.A(n_833),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_835),
.A2(n_830),
.B(n_834),
.Y(n_840)
);

AOI211xp5_ASAP7_75t_L g841 ( 
.A1(n_832),
.A2(n_746),
.B(n_751),
.C(n_727),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_831),
.B(n_805),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_831),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_838),
.Y(n_844)
);

INVx2_ASAP7_75t_SL g845 ( 
.A(n_838),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_842),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_843),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_839),
.A2(n_727),
.B1(n_775),
.B2(n_751),
.Y(n_848)
);

AOI22xp5_ASAP7_75t_L g849 ( 
.A1(n_840),
.A2(n_751),
.B1(n_674),
.B2(n_729),
.Y(n_849)
);

OA22x2_ASAP7_75t_L g850 ( 
.A1(n_841),
.A2(n_674),
.B1(n_711),
.B2(n_753),
.Y(n_850)
);

XNOR2xp5_ASAP7_75t_L g851 ( 
.A(n_837),
.B(n_588),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_838),
.Y(n_852)
);

OAI31xp33_ASAP7_75t_L g853 ( 
.A1(n_846),
.A2(n_618),
.A3(n_588),
.B(n_733),
.Y(n_853)
);

OAI22xp33_ASAP7_75t_L g854 ( 
.A1(n_849),
.A2(n_790),
.B1(n_786),
.B2(n_766),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_SL g855 ( 
.A1(n_847),
.A2(n_737),
.B1(n_735),
.B2(n_610),
.Y(n_855)
);

AOI211xp5_ASAP7_75t_L g856 ( 
.A1(n_844),
.A2(n_615),
.B(n_753),
.C(n_621),
.Y(n_856)
);

OAI22xp5_ASAP7_75t_L g857 ( 
.A1(n_852),
.A2(n_762),
.B1(n_732),
.B2(n_786),
.Y(n_857)
);

AOI31xp33_ASAP7_75t_L g858 ( 
.A1(n_845),
.A2(n_774),
.A3(n_758),
.B(n_742),
.Y(n_858)
);

OAI22xp33_ASAP7_75t_L g859 ( 
.A1(n_850),
.A2(n_790),
.B1(n_718),
.B2(n_731),
.Y(n_859)
);

AOI31xp33_ASAP7_75t_L g860 ( 
.A1(n_848),
.A2(n_851),
.A3(n_774),
.B(n_758),
.Y(n_860)
);

AOI31xp33_ASAP7_75t_L g861 ( 
.A1(n_845),
.A2(n_774),
.A3(n_758),
.B(n_747),
.Y(n_861)
);

OAI22xp5_ASAP7_75t_SL g862 ( 
.A1(n_855),
.A2(n_718),
.B1(n_724),
.B2(n_723),
.Y(n_862)
);

OAI22x1_ASAP7_75t_L g863 ( 
.A1(n_860),
.A2(n_772),
.B1(n_724),
.B2(n_723),
.Y(n_863)
);

XNOR2x1_ASAP7_75t_L g864 ( 
.A(n_859),
.B(n_615),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_857),
.Y(n_865)
);

HB1xp67_ASAP7_75t_L g866 ( 
.A(n_856),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_866),
.A2(n_861),
.B1(n_858),
.B2(n_854),
.Y(n_867)
);

XOR2xp5_ASAP7_75t_L g868 ( 
.A(n_865),
.B(n_853),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_867),
.A2(n_864),
.B1(n_862),
.B2(n_863),
.Y(n_869)
);

AOI22xp5_ASAP7_75t_L g870 ( 
.A1(n_869),
.A2(n_868),
.B1(n_748),
.B2(n_581),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_870),
.B(n_718),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_871),
.A2(n_581),
.B1(n_738),
.B2(n_184),
.Y(n_872)
);


endmodule