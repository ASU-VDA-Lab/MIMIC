module fake_jpeg_15864_n_189 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx4_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx2_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx4f_ASAP7_75t_SL g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_10),
.Y(n_23)
);

INVx5_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_19),
.B(n_2),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_31),
.B(n_33),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g33 ( 
.A(n_19),
.B(n_2),
.Y(n_33)
);

OR2x2_ASAP7_75t_L g34 ( 
.A(n_19),
.B(n_2),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_34),
.B(n_35),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_19),
.B(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_39),
.A2(n_24),
.B1(n_16),
.B2(n_29),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_34),
.B(n_18),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_43),
.B(n_45),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g70 ( 
.A(n_48),
.B(n_52),
.Y(n_70)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_50),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_34),
.B(n_16),
.Y(n_52)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_56),
.Y(n_61)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_38),
.A2(n_3),
.B(n_4),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g68 ( 
.A1(n_55),
.A2(n_18),
.B(n_29),
.C(n_25),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_33),
.B(n_30),
.Y(n_56)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_58),
.B(n_62),
.Y(n_84)
);

O2A1O1Ixp33_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_57),
.B(n_43),
.C(n_55),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_60),
.A2(n_74),
.B1(n_53),
.B2(n_22),
.Y(n_91)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_42),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g64 ( 
.A(n_45),
.B(n_27),
.C(n_23),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_64),
.A2(n_68),
.B(n_28),
.C(n_22),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_49),
.B(n_35),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_65),
.B(n_67),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_32),
.C(n_22),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_69),
.C(n_71),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_44),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_32),
.C(n_49),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g71 ( 
.A(n_51),
.B(n_37),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_54),
.B(n_27),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_72),
.B(n_75),
.Y(n_93)
);

A2O1A1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_41),
.A2(n_37),
.B(n_36),
.C(n_38),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_76),
.B(n_50),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_47),
.A2(n_16),
.B1(n_18),
.B2(n_20),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_77),
.A2(n_47),
.B1(n_20),
.B2(n_25),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_53),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_81),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_61),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_82),
.B(n_89),
.Y(n_105)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_71),
.Y(n_85)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_85),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_86),
.A2(n_90),
.B1(n_92),
.B2(n_94),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_36),
.C(n_22),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_87),
.B(n_91),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_88),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_41),
.B1(n_26),
.B2(n_30),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_63),
.A2(n_21),
.B1(n_4),
.B2(n_5),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_62),
.A2(n_28),
.B1(n_26),
.B2(n_23),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_95),
.B(n_98),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_70),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_96),
.A2(n_74),
.B(n_6),
.Y(n_108)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_68),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_81),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_100),
.B(n_104),
.Y(n_125)
);

MAJx2_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_60),
.C(n_73),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_83),
.C(n_82),
.Y(n_131)
);

CKINVDCx12_ASAP7_75t_R g103 ( 
.A(n_93),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_103),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_79),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_88),
.B(n_67),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_75),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_108),
.A2(n_117),
.B(n_87),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_84),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_109),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_95),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_89),
.A2(n_60),
.B(n_85),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

OA22x2_ASAP7_75t_L g121 ( 
.A1(n_108),
.A2(n_92),
.B1(n_80),
.B2(n_74),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_121),
.A2(n_111),
.B1(n_101),
.B2(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g138 ( 
.A1(n_124),
.A2(n_131),
.B(n_115),
.Y(n_138)
);

INVx2_ASAP7_75t_SL g126 ( 
.A(n_100),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_83),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_127),
.B(n_132),
.Y(n_136)
);

OA21x2_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_74),
.B(n_96),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_129),
.A2(n_78),
.B(n_97),
.Y(n_147)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_130),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_106),
.B(n_74),
.Y(n_132)
);

AO21x1_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_112),
.B(n_111),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_58),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_120),
.A2(n_118),
.B1(n_114),
.B2(n_115),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_119),
.B1(n_140),
.B2(n_141),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_147),
.C(n_142),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_139),
.B(n_141),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_125),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_145),
.B1(n_146),
.B2(n_126),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_102),
.B1(n_101),
.B2(n_59),
.Y(n_145)
);

CKINVDCx14_ASAP7_75t_R g146 ( 
.A(n_134),
.Y(n_146)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_147),
.Y(n_152)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_149),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g150 ( 
.A(n_144),
.B(n_128),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_150),
.B(n_153),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_136),
.B(n_127),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_154),
.C(n_158),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_136),
.A2(n_126),
.B1(n_132),
.B2(n_131),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_145),
.B(n_124),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_155),
.B(n_157),
.Y(n_168)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_160),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_138),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_162),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_154),
.B(n_139),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_148),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_163),
.B(n_156),
.Y(n_170)
);

OR2x2_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_143),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_164),
.B(n_140),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_170),
.B(n_172),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_171),
.A2(n_169),
.B1(n_166),
.B2(n_17),
.Y(n_179)
);

HB1xp67_ASAP7_75t_L g172 ( 
.A(n_164),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_165),
.B(n_133),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_174),
.C(n_168),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_133),
.Y(n_174)
);

AOI321xp33_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_153),
.A3(n_158),
.B1(n_129),
.B2(n_121),
.C(n_13),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_175),
.A2(n_121),
.B(n_8),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_176),
.B(n_179),
.Y(n_181)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_172),
.A2(n_166),
.A3(n_121),
.B1(n_59),
.B2(n_17),
.C1(n_15),
.C2(n_7),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_178),
.Y(n_182)
);

OAI321xp33_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_7),
.A3(n_9),
.B1(n_11),
.B2(n_13),
.C(n_14),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_183),
.A2(n_184),
.B(n_15),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_180),
.B(n_9),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_15),
.Y(n_185)
);

BUFx24_ASAP7_75t_SL g187 ( 
.A(n_185),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_187),
.B(n_186),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_188),
.B(n_181),
.Y(n_189)
);


endmodule