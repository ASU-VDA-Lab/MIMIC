module fake_netlist_1_4405_n_32 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
INVx1_ASAP7_75t_L g11 ( .A(n_4), .Y(n_11) );
INVx3_ASAP7_75t_L g12 ( .A(n_5), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_2), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx3_ASAP7_75t_L g15 ( .A(n_1), .Y(n_15) );
INVx2_ASAP7_75t_L g16 ( .A(n_15), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_15), .Y(n_17) );
NAND3xp33_ASAP7_75t_SL g18 ( .A(n_11), .B(n_0), .C(n_2), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
AOI22xp5_ASAP7_75t_L g20 ( .A1(n_18), .A2(n_15), .B1(n_14), .B2(n_13), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_20), .A2(n_17), .B1(n_14), .B2(n_13), .Y(n_21) );
NAND4xp25_ASAP7_75t_L g22 ( .A(n_19), .B(n_11), .C(n_16), .D(n_12), .Y(n_22) );
NAND2xp5_ASAP7_75t_L g23 ( .A(n_21), .B(n_12), .Y(n_23) );
NOR3xp33_ASAP7_75t_L g24 ( .A(n_22), .B(n_12), .C(n_3), .Y(n_24) );
NOR2x1_ASAP7_75t_L g25 ( .A(n_23), .B(n_0), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_24), .B(n_3), .Y(n_26) );
INVxp67_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
NOR2x1_ASAP7_75t_L g28 ( .A(n_25), .B(n_4), .Y(n_28) );
CKINVDCx5p33_ASAP7_75t_R g29 ( .A(n_27), .Y(n_29) );
OR2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_10), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
AOI222xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B1(n_7), .B2(n_8), .C1(n_9), .C2(n_6), .Y(n_32) );
endmodule