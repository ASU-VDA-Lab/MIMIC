module fake_jpeg_15835_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx6f_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

INVx3_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx6f_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

CKINVDCx14_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx3_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

INVx13_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_14),
.A2(n_15),
.B1(n_17),
.B2(n_12),
.Y(n_18)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_16),
.B(n_6),
.C(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_18),
.Y(n_24)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_15),
.B(n_8),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_21),
.C(n_16),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_20),
.A2(n_16),
.B1(n_0),
.B2(n_2),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_22),
.A2(n_21),
.B1(n_0),
.B2(n_4),
.Y(n_29)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_19),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g27 ( 
.A(n_25),
.B(n_26),
.Y(n_27)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

XNOR2xp5_ASAP7_75t_SL g30 ( 
.A(n_29),
.B(n_22),
.Y(n_30)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_32),
.C(n_28),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_24),
.Y(n_31)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_25),
.B(n_23),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_28),
.C(n_26),
.Y(n_35)
);

XOR2xp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_36),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_37),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_4),
.Y(n_39)
);


endmodule