module real_jpeg_5774_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_128;
wire n_202;
wire n_216;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_215;
wire n_286;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_420;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx8_ASAP7_75t_L g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_1),
.A2(n_80),
.B1(n_83),
.B2(n_84),
.Y(n_79)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_1),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_1),
.A2(n_117),
.B1(n_120),
.B2(n_121),
.Y(n_116)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_1),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_1),
.A2(n_121),
.B1(n_157),
.B2(n_159),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_1),
.A2(n_197),
.B1(n_199),
.B2(n_200),
.Y(n_196)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_1),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_2),
.A2(n_25),
.B1(n_43),
.B2(n_46),
.Y(n_42)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_46),
.B1(n_141),
.B2(n_143),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_2),
.A2(n_46),
.B1(n_189),
.B2(n_191),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_2),
.A2(n_46),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g258 ( 
.A1(n_2),
.A2(n_259),
.B(n_262),
.C(n_265),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_2),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_2),
.B(n_51),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_2),
.B(n_301),
.C(n_302),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_2),
.B(n_109),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g322 ( 
.A(n_2),
.B(n_74),
.C(n_323),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_2),
.B(n_27),
.Y(n_338)
);

OAI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_3),
.A2(n_74),
.B1(n_76),
.B2(n_77),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_3),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_3),
.A2(n_76),
.B1(n_111),
.B2(n_113),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_3),
.A2(n_76),
.B1(n_126),
.B2(n_128),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_3),
.A2(n_76),
.B1(n_170),
.B2(n_174),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_4),
.A2(n_22),
.B1(n_24),
.B2(n_25),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_4),
.A2(n_24),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_4),
.A2(n_24),
.B1(n_71),
.B2(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_4),
.A2(n_24),
.B1(n_269),
.B2(n_270),
.Y(n_268)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_5),
.Y(n_55)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_5),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_5),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g424 ( 
.A(n_6),
.Y(n_424)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_7),
.Y(n_93)
);

INVx8_ASAP7_75t_L g167 ( 
.A(n_8),
.Y(n_167)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_8),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_8),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_8),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_9),
.Y(n_261)
);

BUFx5_ASAP7_75t_L g264 ( 
.A(n_9),
.Y(n_264)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx3_ASAP7_75t_L g421 ( 
.A(n_11),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_12),
.Y(n_127)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_13),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_13),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_13),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_419),
.B(n_422),
.Y(n_14)
);

XNOR2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_415),
.Y(n_15)
);

AO21x2_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_130),
.B(n_414),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_124),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_18),
.B(n_124),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_115),
.C(n_122),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_19),
.B(n_411),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_48),
.C(n_78),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_20),
.A2(n_138),
.B1(n_139),
.B2(n_152),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_20),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_20),
.B(n_139),
.C(n_153),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_20),
.B(n_240),
.C(n_257),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_20),
.A2(n_152),
.B1(n_240),
.B2(n_339),
.Y(n_362)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_20),
.A2(n_152),
.B1(n_386),
.B2(n_387),
.Y(n_385)
);

OA22x2_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_26),
.B1(n_42),
.B2(n_47),
.Y(n_20)
);

OA22x2_ASAP7_75t_L g228 ( 
.A1(n_21),
.A2(n_26),
.B1(n_42),
.B2(n_47),
.Y(n_228)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g265 ( 
.A(n_25),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_26),
.A2(n_42),
.B1(n_47),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_26),
.A2(n_47),
.B1(n_116),
.B2(n_125),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_26),
.A2(n_42),
.B(n_47),
.Y(n_235)
);

AO21x1_ASAP7_75t_L g417 ( 
.A1(n_26),
.A2(n_47),
.B(n_125),
.Y(n_417)
);

OR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_35),
.Y(n_26)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g27 ( 
.A1(n_28),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_27)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_28),
.Y(n_147)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_29),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_29),
.Y(n_145)
);

INVx6_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_30),
.Y(n_85)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_30),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_30),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g151 ( 
.A(n_30),
.Y(n_151)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_38),
.B1(n_39),
.B2(n_40),
.Y(n_35)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_36),
.Y(n_119)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_37),
.Y(n_129)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g262 ( 
.A1(n_46),
.A2(n_141),
.B(n_263),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g387 ( 
.A1(n_48),
.A2(n_78),
.B1(n_388),
.B2(n_389),
.Y(n_387)
);

CKINVDCx14_ASAP7_75t_R g389 ( 
.A(n_48),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_48),
.B(n_228),
.C(n_391),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_48),
.A2(n_389),
.B1(n_391),
.B2(n_398),
.Y(n_397)
);

AND2x2_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_73),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_49),
.B(n_188),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_50),
.B(n_61),
.Y(n_49)
);

OA22x2_ASAP7_75t_L g181 ( 
.A1(n_50),
.A2(n_61),
.B1(n_182),
.B2(n_187),
.Y(n_181)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

NOR2x1_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_63),
.Y(n_62)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_51),
.A2(n_196),
.B(n_203),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_51),
.B(n_183),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_51),
.A2(n_62),
.B1(n_73),
.B2(n_196),
.Y(n_239)
);

AO22x1_ASAP7_75t_SL g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_56),
.B2(n_59),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_52),
.A2(n_64),
.B1(n_67),
.B2(n_70),
.Y(n_63)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_55),
.Y(n_159)
);

BUFx6f_ASAP7_75t_L g225 ( 
.A(n_55),
.Y(n_225)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_55),
.Y(n_272)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_57),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g158 ( 
.A(n_58),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_58),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_62),
.B(n_188),
.Y(n_204)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_66),
.Y(n_72)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_66),
.Y(n_106)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_66),
.Y(n_202)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g186 ( 
.A(n_72),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_72),
.Y(n_192)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_74),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_75),
.Y(n_190)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_78),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_86),
.B1(n_109),
.B2(n_110),
.Y(n_78)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_79),
.Y(n_392)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_85),
.Y(n_114)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_85),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_86),
.B(n_227),
.Y(n_393)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_87),
.B(n_101),
.Y(n_123)
);

OA22x2_ASAP7_75t_L g139 ( 
.A1(n_87),
.A2(n_101),
.B1(n_140),
.B2(n_146),
.Y(n_139)
);

OA22x2_ASAP7_75t_L g240 ( 
.A1(n_87),
.A2(n_101),
.B1(n_140),
.B2(n_146),
.Y(n_240)
);

NAND2x1_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_101),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g88 ( 
.A1(n_89),
.A2(n_94),
.B1(n_96),
.B2(n_99),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_92),
.Y(n_98)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_93),
.Y(n_104)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

INVx8_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx6_ASAP7_75t_L g323 ( 
.A(n_98),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_101),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_L g391 ( 
.A1(n_101),
.A2(n_392),
.B(n_393),
.Y(n_391)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_103),
.B1(n_105),
.B2(n_107),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_104),
.Y(n_108)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_110),
.B(n_123),
.Y(n_122)
);

INVx6_ASAP7_75t_SL g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g411 ( 
.A(n_115),
.B(n_122),
.Y(n_411)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_123),
.B(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_124),
.B(n_417),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g418 ( 
.A(n_124),
.B(n_417),
.Y(n_418)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_409),
.B(n_413),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_132),
.A2(n_380),
.B(n_406),
.Y(n_131)
);

OAI211xp5_ASAP7_75t_L g132 ( 
.A1(n_133),
.A2(n_276),
.B(n_374),
.C(n_379),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_245),
.Y(n_133)
);

A2O1A1Ixp33_ASAP7_75t_L g374 ( 
.A1(n_134),
.A2(n_245),
.B(n_375),
.C(n_378),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_229),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g379 ( 
.A(n_135),
.B(n_229),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_193),
.C(n_211),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_136),
.B(n_193),
.Y(n_247)
);

XNOR2x1_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_153),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_138),
.A2(n_139),
.B1(n_214),
.B2(n_295),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_138),
.B(n_295),
.C(n_316),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_138),
.A2(n_139),
.B1(n_349),
.B2(n_350),
.Y(n_348)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_139),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_139),
.B(n_228),
.C(n_349),
.Y(n_366)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_140),
.Y(n_227)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_151),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_180),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_154),
.A2(n_180),
.B1(n_181),
.B2(n_255),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_154),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_155),
.A2(n_160),
.B1(n_168),
.B2(n_177),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_156),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_156),
.A2(n_217),
.B(n_220),
.Y(n_216)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx6_ASAP7_75t_L g285 ( 
.A(n_159),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_160),
.B(n_207),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_160),
.B(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_161),
.A2(n_222),
.B1(n_268),
.B2(n_273),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_161),
.A2(n_218),
.B1(n_222),
.B2(n_268),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx3_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_167),
.Y(n_209)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_167),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_206),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g170 ( 
.A(n_171),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

BUFx5_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_174),
.Y(n_302)
);

INVx4_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_176),
.Y(n_223)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_180),
.A2(n_181),
.B1(n_309),
.B2(n_310),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_180),
.A2(n_181),
.B1(n_331),
.B2(n_332),
.Y(n_330)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_181),
.B(n_267),
.C(n_309),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_181),
.B(n_331),
.C(n_333),
.Y(n_344)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx4_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_189),
.Y(n_198)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_190),
.Y(n_189)
);

INVx11_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_195),
.B1(n_205),
.B2(n_210),
.Y(n_193)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_195),
.B(n_205),
.Y(n_236)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

BUFx3_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx4_ASAP7_75t_L g299 ( 
.A(n_202),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

AND2x2_ASAP7_75t_SL g214 ( 
.A(n_204),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_205),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_205),
.A2(n_210),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g400 ( 
.A1(n_205),
.A2(n_235),
.B(n_236),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_206),
.B(n_222),
.Y(n_324)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx8_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_211),
.B(n_247),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_226),
.C(n_228),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_213),
.B(n_251),
.Y(n_250)
);

NOR2xp67_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_216),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_214),
.A2(n_295),
.B1(n_296),
.B2(n_303),
.Y(n_294)
);

INVx2_ASAP7_75t_L g295 ( 
.A(n_214),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_L g364 ( 
.A1(n_214),
.A2(n_216),
.B1(n_295),
.B2(n_365),
.Y(n_364)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_216),
.Y(n_365)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_226),
.A2(n_228),
.B1(n_252),
.B2(n_253),
.Y(n_251)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_226),
.Y(n_253)
);

INVx2_ASAP7_75t_SL g252 ( 
.A(n_228),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_228),
.A2(n_252),
.B1(n_347),
.B2(n_348),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g383 ( 
.A1(n_228),
.A2(n_252),
.B1(n_384),
.B2(n_385),
.Y(n_383)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_228),
.A2(n_252),
.B1(n_396),
.B2(n_397),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_228),
.B(n_385),
.C(n_390),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_243),
.B2(n_244),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_237),
.B1(n_238),
.B2(n_242),
.Y(n_231)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_232),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g405 ( 
.A(n_237),
.B(n_242),
.C(n_244),
.Y(n_405)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_240),
.B(n_241),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_240),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_240),
.A2(n_335),
.B1(n_336),
.B2(n_339),
.Y(n_334)
);

CKINVDCx16_ASAP7_75t_R g339 ( 
.A(n_240),
.Y(n_339)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_241),
.Y(n_399)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_241),
.A2(n_395),
.B1(n_399),
.B2(n_404),
.Y(n_403)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_246),
.B(n_248),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_249),
.B(n_254),
.C(n_256),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_249),
.A2(n_250),
.B1(n_254),
.B2(n_373),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_254),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g371 ( 
.A(n_256),
.B(n_372),
.Y(n_371)
);

XOR2xp5_ASAP7_75t_L g361 ( 
.A(n_257),
.B(n_362),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_266),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_258),
.A2(n_266),
.B1(n_267),
.B2(n_356),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_258),
.Y(n_356)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx3_ASAP7_75t_SL g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_266),
.A2(n_267),
.B1(n_307),
.B2(n_308),
.Y(n_306)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_290),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_267),
.B(n_290),
.Y(n_291)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_358),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_278),
.A2(n_343),
.B(n_357),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_328),
.B(n_342),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_313),
.B(n_327),
.Y(n_279)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_281),
.A2(n_305),
.B(n_312),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_282),
.A2(n_292),
.B(n_304),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_283),
.A2(n_289),
.B(n_291),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_288),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_288),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_288),
.A2(n_293),
.B1(n_337),
.B2(n_338),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_294),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_293),
.B(n_337),
.C(n_339),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_303),
.Y(n_311)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_296),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_300),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx4_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_311),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_311),
.Y(n_312)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_309),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_315),
.Y(n_327)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_326),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_317),
.A2(n_318),
.B1(n_324),
.B2(n_325),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_317),
.B(n_325),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_319),
.B(n_322),
.Y(n_318)
);

INVx3_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx2_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_324),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_329),
.B(n_341),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_329),
.B(n_341),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_330),
.A2(n_333),
.B1(n_334),
.B2(n_340),
.Y(n_329)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_330),
.Y(n_340)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_331),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

CKINVDCx14_ASAP7_75t_R g337 ( 
.A(n_338),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_344),
.B(n_345),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_351),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_353),
.C(n_354),
.Y(n_367)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_349),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_352),
.A2(n_353),
.B1(n_354),
.B2(n_355),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

NOR2x1_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_368),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_360),
.B(n_367),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_360),
.B(n_367),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_363),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_361),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_366),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_364),
.B(n_366),
.C(n_370),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_368),
.A2(n_376),
.B(n_377),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_371),
.Y(n_368)
);

OR2x2_ASAP7_75t_L g377 ( 
.A(n_369),
.B(n_371),
.Y(n_377)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_381),
.B(n_401),
.Y(n_380)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_381),
.A2(n_407),
.B(n_408),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_394),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_382),
.B(n_394),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_390),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_391),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_399),
.C(n_400),
.Y(n_394)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_395),
.Y(n_404)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_400),
.B(n_403),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_402),
.B(n_405),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_405),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_412),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_410),
.B(n_412),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_418),
.Y(n_415)
);

BUFx4f_ASAP7_75t_SL g419 ( 
.A(n_420),
.Y(n_419)
);

INVx13_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

INVx5_ASAP7_75t_L g423 ( 
.A(n_421),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);


endmodule