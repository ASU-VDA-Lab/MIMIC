module fake_jpeg_18755_n_203 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_0),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

INVx6_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx16f_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_14),
.B(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_31),
.B(n_32),
.Y(n_53)
);

INVx6_ASAP7_75t_SL g32 ( 
.A(n_18),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_33),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_18),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_35),
.B(n_39),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_23),
.B(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_37),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_23),
.B(n_1),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_23),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_40),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

INVx2_ASAP7_75t_SL g41 ( 
.A(n_29),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_42),
.Y(n_56)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_29),
.B(n_2),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_43),
.A2(n_26),
.B1(n_16),
.B2(n_22),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_26),
.B1(n_16),
.B2(n_14),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_45),
.A2(n_51),
.B1(n_38),
.B2(n_40),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_43),
.Y(n_61)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_48),
.B(n_49),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_42),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_15),
.B1(n_21),
.B2(n_30),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_36),
.A2(n_22),
.B1(n_21),
.B2(n_28),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_52),
.A2(n_57),
.B1(n_40),
.B2(n_3),
.Y(n_83)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_32),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_54),
.B(n_27),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_43),
.A2(n_24),
.B1(n_28),
.B2(n_19),
.Y(n_57)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_60),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_61),
.A2(n_65),
.B1(n_78),
.B2(n_2),
.Y(n_99)
);

INVx13_ASAP7_75t_L g63 ( 
.A(n_54),
.Y(n_63)
);

INVx13_ASAP7_75t_L g107 ( 
.A(n_63),
.Y(n_107)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_44),
.A2(n_37),
.B1(n_36),
.B2(n_38),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_60),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_69),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_44),
.B(n_37),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_68),
.B(n_73),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_55),
.Y(n_69)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_70),
.Y(n_105)
);

OR2x4_ASAP7_75t_L g71 ( 
.A(n_46),
.B(n_41),
.Y(n_71)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_71),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_49),
.B(n_39),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_53),
.A2(n_29),
.B(n_35),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_76),
.A2(n_31),
.B(n_25),
.Y(n_101)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_40),
.B1(n_38),
.B2(n_35),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_80),
.Y(n_109)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_59),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_56),
.B(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_81),
.B(n_82),
.Y(n_110)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_50),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_83),
.A2(n_90),
.B1(n_24),
.B2(n_27),
.Y(n_96)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_84),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_48),
.A2(n_19),
.B1(n_30),
.B2(n_20),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_56),
.B(n_34),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_86),
.B(n_89),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_55),
.Y(n_87)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_59),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_50),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_47),
.A2(n_52),
.B1(n_25),
.B2(n_20),
.Y(n_90)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_89),
.A2(n_53),
.B(n_34),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_92),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_34),
.C(n_33),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_94),
.B(n_97),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_86),
.B1(n_81),
.B2(n_66),
.Y(n_119)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_65),
.B(n_61),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_99),
.B(n_83),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_77),
.B(n_59),
.C(n_27),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_100),
.B(n_74),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_73),
.B(n_3),
.Y(n_103)
);

CKINVDCx16_ASAP7_75t_R g114 ( 
.A(n_103),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_113),
.A2(n_119),
.B1(n_129),
.B2(n_103),
.Y(n_147)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_115),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_93),
.A2(n_84),
.B1(n_82),
.B2(n_71),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_116),
.A2(n_96),
.B1(n_102),
.B2(n_111),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_109),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_118),
.B(n_120),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_95),
.Y(n_120)
);

A2O1A1O1Ixp25_ASAP7_75t_L g121 ( 
.A1(n_93),
.A2(n_76),
.B(n_63),
.C(n_72),
.D(n_62),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_98),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_95),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_123),
.B(n_124),
.Y(n_133)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_125),
.B(n_127),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_108),
.B(n_72),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_128),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_97),
.B(n_62),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_13),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g132 ( 
.A(n_130),
.B(n_103),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_126),
.B(n_94),
.C(n_108),
.Y(n_131)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_131),
.B(n_139),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_132),
.B(n_147),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_136),
.A2(n_145),
.B1(n_115),
.B2(n_125),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_111),
.C(n_104),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_129),
.B(n_116),
.C(n_127),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_141),
.B(n_143),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_128),
.B(n_104),
.C(n_110),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_117),
.A2(n_92),
.B(n_102),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_144),
.A2(n_114),
.B(n_121),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_113),
.A2(n_99),
.B1(n_110),
.B2(n_106),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_112),
.B(n_100),
.C(n_101),
.Y(n_146)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_146),
.B(n_114),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_134),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_148),
.B(n_149),
.Y(n_169)
);

CKINVDCx14_ASAP7_75t_R g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_135),
.B(n_120),
.Y(n_151)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_151),
.Y(n_164)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_152),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_142),
.A2(n_112),
.B1(n_123),
.B2(n_119),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_153),
.A2(n_155),
.B1(n_161),
.B2(n_107),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_144),
.C(n_141),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_154),
.B(n_150),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_143),
.B(n_122),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_156),
.A2(n_132),
.B(n_138),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_158),
.B(n_146),
.C(n_139),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_160),
.A2(n_140),
.B1(n_136),
.B2(n_145),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_124),
.B1(n_70),
.B2(n_64),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_163),
.C(n_168),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_165),
.A2(n_170),
.B1(n_161),
.B2(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_166),
.B(n_167),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_107),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_148),
.A2(n_91),
.B1(n_105),
.B2(n_88),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_159),
.B(n_107),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_171),
.A2(n_154),
.B(n_157),
.Y(n_175)
);

BUFx2_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_174),
.A2(n_165),
.B1(n_91),
.B2(n_171),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_162),
.Y(n_182)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_169),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_176),
.A2(n_178),
.B1(n_179),
.B2(n_181),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_153),
.B(n_150),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_180),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_170),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_172),
.A2(n_4),
.B(n_5),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_182),
.B(n_185),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_183),
.B(n_184),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_173),
.B(n_168),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_88),
.B1(n_80),
.B2(n_91),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_186),
.B(n_4),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_174),
.B(n_88),
.C(n_6),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_4),
.C(n_7),
.Y(n_189)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_189),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_190),
.B(n_193),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_187),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_192),
.B(n_188),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g198 ( 
.A(n_196),
.B(n_191),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g197 ( 
.A1(n_194),
.A2(n_190),
.B(n_188),
.Y(n_197)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_197),
.A2(n_198),
.B(n_195),
.Y(n_199)
);

AOI322xp5_ASAP7_75t_L g200 ( 
.A1(n_199),
.A2(n_185),
.A3(n_182),
.B1(n_9),
.B2(n_10),
.C1(n_11),
.C2(n_8),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_200),
.B(n_7),
.C(n_8),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_9),
.C(n_10),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_10),
.Y(n_203)
);


endmodule