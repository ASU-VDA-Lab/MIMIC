module fake_aes_5778_n_536 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_536);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_536;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_119;
wire n_141;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_447;
wire n_171;
wire n_196;
wire n_192;
wire n_502;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_133;
wire n_149;
wire n_81;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_107;
wire n_403;
wire n_516;
wire n_254;
wire n_262;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_376;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_435;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_445;
wire n_398;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_418;
wire n_493;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g77 ( .A(n_24), .Y(n_77) );
CKINVDCx5p33_ASAP7_75t_R g78 ( .A(n_51), .Y(n_78) );
CKINVDCx20_ASAP7_75t_R g79 ( .A(n_7), .Y(n_79) );
CKINVDCx20_ASAP7_75t_R g80 ( .A(n_18), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_66), .Y(n_81) );
INVx1_ASAP7_75t_SL g82 ( .A(n_68), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_9), .Y(n_83) );
CKINVDCx20_ASAP7_75t_R g84 ( .A(n_67), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_34), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_1), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_21), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_45), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_15), .Y(n_89) );
BUFx3_ASAP7_75t_L g90 ( .A(n_16), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_50), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_38), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_20), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_25), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_28), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_39), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_2), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_65), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_42), .Y(n_99) );
INVxp67_ASAP7_75t_L g100 ( .A(n_40), .Y(n_100) );
CKINVDCx16_ASAP7_75t_R g101 ( .A(n_52), .Y(n_101) );
BUFx2_ASAP7_75t_L g102 ( .A(n_22), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_7), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_54), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_61), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_75), .Y(n_106) );
INVxp67_ASAP7_75t_SL g107 ( .A(n_73), .Y(n_107) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_55), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_49), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_12), .Y(n_110) );
HB1xp67_ASAP7_75t_L g111 ( .A(n_59), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_36), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_85), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_85), .Y(n_114) );
AND2x2_ASAP7_75t_L g115 ( .A(n_102), .B(n_0), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g117 ( .A(n_102), .B(n_0), .Y(n_117) );
OAI22x1_ASAP7_75t_SL g118 ( .A1(n_79), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_88), .Y(n_119) );
OA21x2_ASAP7_75t_L g120 ( .A1(n_77), .A2(n_35), .B(n_74), .Y(n_120) );
AND2x4_ASAP7_75t_L g121 ( .A(n_86), .B(n_3), .Y(n_121) );
INVx2_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
NOR2x1_ASAP7_75t_L g123 ( .A(n_93), .B(n_4), .Y(n_123) );
INVx3_ASAP7_75t_L g124 ( .A(n_97), .Y(n_124) );
AND2x4_ASAP7_75t_L g125 ( .A(n_86), .B(n_4), .Y(n_125) );
AND2x4_ASAP7_75t_L g126 ( .A(n_91), .B(n_5), .Y(n_126) );
HB1xp67_ASAP7_75t_L g127 ( .A(n_83), .Y(n_127) );
INVx2_ASAP7_75t_L g128 ( .A(n_91), .Y(n_128) );
BUFx8_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_90), .Y(n_130) );
INVx3_ASAP7_75t_L g131 ( .A(n_97), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_94), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_98), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_99), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_97), .Y(n_135) );
INVxp67_ASAP7_75t_SL g136 ( .A(n_115), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_115), .Y(n_137) );
NOR2x1p5_ASAP7_75t_L g138 ( .A(n_117), .B(n_78), .Y(n_138) );
INVx4_ASAP7_75t_L g139 ( .A(n_121), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g140 ( .A(n_113), .B(n_111), .Y(n_140) );
AOI22xp33_ASAP7_75t_L g141 ( .A1(n_121), .A2(n_110), .B1(n_89), .B2(n_103), .Y(n_141) );
INVx1_ASAP7_75t_SL g142 ( .A(n_115), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_116), .B(n_100), .Y(n_143) );
INVx4_ASAP7_75t_L g144 ( .A(n_121), .Y(n_144) );
NOR2xp33_ASAP7_75t_L g145 ( .A(n_116), .B(n_101), .Y(n_145) );
INVx2_ASAP7_75t_SL g146 ( .A(n_129), .Y(n_146) );
NAND2xp5_ASAP7_75t_SL g147 ( .A(n_129), .B(n_108), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_119), .B(n_112), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_122), .Y(n_149) );
NAND2xp5_ASAP7_75t_L g150 ( .A(n_113), .B(n_104), .Y(n_150) );
INVxp33_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_131), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_131), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_114), .B(n_109), .Y(n_154) );
INVx1_ASAP7_75t_SL g155 ( .A(n_127), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_122), .Y(n_156) );
AND3x2_ASAP7_75t_L g157 ( .A(n_127), .B(n_107), .C(n_84), .Y(n_157) );
INVx2_ASAP7_75t_SL g158 ( .A(n_129), .Y(n_158) );
NOR2xp33_ASAP7_75t_L g159 ( .A(n_119), .B(n_109), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_131), .Y(n_160) );
NAND2x1p5_ASAP7_75t_L g161 ( .A(n_155), .B(n_121), .Y(n_161) );
AND2x6_ASAP7_75t_L g162 ( .A(n_142), .B(n_121), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_155), .B(n_125), .Y(n_163) );
AOI221xp5_ASAP7_75t_L g164 ( .A1(n_136), .A2(n_114), .B1(n_134), .B2(n_133), .C(n_132), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_154), .B(n_129), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g166 ( .A(n_154), .B(n_129), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_139), .Y(n_167) );
NAND2xp33_ASAP7_75t_L g168 ( .A(n_146), .B(n_78), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_151), .B(n_134), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_142), .Y(n_170) );
AO22x1_ASAP7_75t_L g171 ( .A1(n_137), .A2(n_125), .B1(n_126), .B2(n_96), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_149), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_149), .Y(n_173) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_146), .B(n_158), .Y(n_174) );
BUFx6f_ASAP7_75t_L g175 ( .A(n_146), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_139), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_156), .Y(n_177) );
NAND2xp5_ASAP7_75t_SL g178 ( .A(n_158), .B(n_125), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_156), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_145), .B(n_133), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_139), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_158), .B(n_125), .Y(n_182) );
NAND2xp5_ASAP7_75t_SL g183 ( .A(n_139), .B(n_125), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g184 ( .A(n_140), .B(n_132), .Y(n_184) );
INVxp67_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
AOI22xp33_ASAP7_75t_SL g186 ( .A1(n_140), .A2(n_80), .B1(n_92), .B2(n_126), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_143), .B(n_126), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_138), .B(n_126), .Y(n_188) );
OAI22xp5_ASAP7_75t_L g189 ( .A1(n_141), .A2(n_126), .B1(n_123), .B2(n_130), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_144), .B(n_130), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_144), .B(n_130), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_138), .B(n_106), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_144), .B(n_106), .Y(n_193) );
BUFx12f_ASAP7_75t_L g194 ( .A(n_163), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_172), .Y(n_195) );
BUFx2_ASAP7_75t_L g196 ( .A(n_163), .Y(n_196) );
O2A1O1Ixp33_ASAP7_75t_L g197 ( .A1(n_189), .A2(n_147), .B(n_150), .C(n_148), .Y(n_197) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_161), .A2(n_144), .B1(n_150), .B2(n_95), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_185), .B(n_157), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g200 ( .A1(n_161), .A2(n_87), .B1(n_95), .B2(n_96), .Y(n_200) );
OAI21xp5_ASAP7_75t_L g201 ( .A1(n_183), .A2(n_120), .B(n_123), .Y(n_201) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_165), .B(n_87), .Y(n_202) );
INVx2_ASAP7_75t_SL g203 ( .A(n_169), .Y(n_203) );
AND2x2_ASAP7_75t_L g204 ( .A(n_184), .B(n_122), .Y(n_204) );
AOI21xp5_ASAP7_75t_L g205 ( .A1(n_178), .A2(n_120), .B(n_153), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_173), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_170), .B(n_128), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_177), .Y(n_208) );
BUFx4f_ASAP7_75t_L g209 ( .A(n_162), .Y(n_209) );
INVx4_ASAP7_75t_L g210 ( .A(n_162), .Y(n_210) );
NAND2x1p5_ASAP7_75t_L g211 ( .A(n_181), .B(n_120), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_179), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_164), .B(n_105), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g214 ( .A1(n_178), .A2(n_120), .B(n_153), .Y(n_214) );
INVx2_ASAP7_75t_L g215 ( .A(n_167), .Y(n_215) );
NAND3xp33_ASAP7_75t_SL g216 ( .A(n_186), .B(n_105), .C(n_82), .Y(n_216) );
AND2x4_ASAP7_75t_L g217 ( .A(n_176), .B(n_128), .Y(n_217) );
A2O1A1Ixp33_ASAP7_75t_L g218 ( .A1(n_180), .A2(n_128), .B(n_124), .C(n_131), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_171), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g220 ( .A1(n_182), .A2(n_174), .B(n_166), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_162), .B(n_97), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_192), .B(n_118), .Y(n_222) );
O2A1O1Ixp33_ASAP7_75t_L g223 ( .A1(n_188), .A2(n_124), .B(n_131), .C(n_135), .Y(n_223) );
O2A1O1Ixp33_ASAP7_75t_L g224 ( .A1(n_187), .A2(n_124), .B(n_135), .C(n_152), .Y(n_224) );
NOR2x1_ASAP7_75t_L g225 ( .A(n_193), .B(n_118), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_203), .Y(n_226) );
A2O1A1Ixp33_ASAP7_75t_L g227 ( .A1(n_197), .A2(n_182), .B(n_190), .C(n_191), .Y(n_227) );
OAI21xp5_ASAP7_75t_L g228 ( .A1(n_220), .A2(n_191), .B(n_190), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_205), .A2(n_174), .B(n_168), .Y(n_229) );
AOI21xp5_ASAP7_75t_L g230 ( .A1(n_214), .A2(n_175), .B(n_120), .Y(n_230) );
NAND2x1p5_ASAP7_75t_L g231 ( .A(n_210), .B(n_175), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_203), .B(n_162), .Y(n_232) );
AOI21xp5_ASAP7_75t_L g233 ( .A1(n_202), .A2(n_175), .B(n_152), .Y(n_233) );
OAI21x1_ASAP7_75t_L g234 ( .A1(n_211), .A2(n_201), .B(n_221), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_225), .B(n_162), .Y(n_235) );
INVx3_ASAP7_75t_L g236 ( .A(n_210), .Y(n_236) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_218), .A2(n_124), .B(n_135), .C(n_97), .Y(n_237) );
A2O1A1Ixp33_ASAP7_75t_L g238 ( .A1(n_218), .A2(n_135), .B(n_175), .C(n_153), .Y(n_238) );
OAI22x1_ASAP7_75t_L g239 ( .A1(n_219), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_202), .A2(n_160), .B(n_152), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_204), .Y(n_241) );
INVx2_ASAP7_75t_SL g242 ( .A(n_194), .Y(n_242) );
OAI21xp5_ASAP7_75t_L g243 ( .A1(n_215), .A2(n_160), .B(n_135), .Y(n_243) );
AOI21xp5_ASAP7_75t_L g244 ( .A1(n_198), .A2(n_160), .B(n_41), .Y(n_244) );
BUFx3_ASAP7_75t_L g245 ( .A(n_194), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_222), .B(n_6), .Y(n_246) );
OAI22xp33_ASAP7_75t_SL g247 ( .A1(n_219), .A2(n_8), .B1(n_9), .B2(n_10), .Y(n_247) );
INVx2_ASAP7_75t_SL g248 ( .A(n_209), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_204), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_207), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_195), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_241), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_230), .A2(n_211), .B(n_224), .Y(n_253) );
AO31x2_ASAP7_75t_L g254 ( .A1(n_237), .A2(n_238), .A3(n_229), .B(n_227), .Y(n_254) );
INVx5_ASAP7_75t_L g255 ( .A(n_236), .Y(n_255) );
OA21x2_ASAP7_75t_L g256 ( .A1(n_234), .A2(n_195), .B(n_206), .Y(n_256) );
INVx1_ASAP7_75t_SL g257 ( .A(n_245), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_236), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_249), .B(n_212), .Y(n_259) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_233), .A2(n_209), .B(n_206), .Y(n_260) );
AO31x2_ASAP7_75t_L g261 ( .A1(n_237), .A2(n_208), .A3(n_212), .B(n_210), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_232), .A2(n_199), .B1(n_216), .B2(n_200), .Y(n_262) );
OR2x6_ASAP7_75t_L g263 ( .A(n_248), .B(n_196), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_227), .A2(n_209), .B(n_208), .Y(n_264) );
AOI21xp33_ASAP7_75t_L g265 ( .A1(n_232), .A2(n_223), .B(n_207), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_251), .B(n_217), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_250), .B(n_213), .Y(n_267) );
INVx6_ASAP7_75t_L g268 ( .A(n_245), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_251), .Y(n_269) );
BUFx2_ASAP7_75t_L g270 ( .A(n_226), .Y(n_270) );
OAI21x1_ASAP7_75t_L g271 ( .A1(n_234), .A2(n_215), .B(n_217), .Y(n_271) );
AND2x4_ASAP7_75t_L g272 ( .A(n_248), .B(n_217), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_235), .Y(n_273) );
INVx2_ASAP7_75t_L g274 ( .A(n_256), .Y(n_274) );
INVx2_ASAP7_75t_SL g275 ( .A(n_255), .Y(n_275) );
AOI21xp5_ASAP7_75t_SL g276 ( .A1(n_256), .A2(n_239), .B(n_238), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_257), .B(n_242), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_269), .B(n_228), .Y(n_278) );
AND2x2_ASAP7_75t_L g279 ( .A(n_269), .B(n_236), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_259), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_256), .Y(n_281) );
INVx2_ASAP7_75t_L g282 ( .A(n_271), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_271), .Y(n_283) );
OA21x2_ASAP7_75t_L g284 ( .A1(n_253), .A2(n_244), .B(n_243), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_273), .A2(n_246), .B1(n_242), .B2(n_247), .Y(n_285) );
AND2x4_ASAP7_75t_L g286 ( .A(n_255), .B(n_240), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_254), .Y(n_287) );
AND2x2_ASAP7_75t_L g288 ( .A(n_259), .B(n_231), .Y(n_288) );
INVxp67_ASAP7_75t_SL g289 ( .A(n_266), .Y(n_289) );
OR2x2_ASAP7_75t_L g290 ( .A(n_252), .B(n_231), .Y(n_290) );
INVx3_ASAP7_75t_L g291 ( .A(n_255), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_268), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_254), .B(n_10), .Y(n_293) );
AND2x2_ASAP7_75t_L g294 ( .A(n_254), .B(n_11), .Y(n_294) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_261), .Y(n_295) );
AOI211xp5_ASAP7_75t_SL g296 ( .A1(n_276), .A2(n_262), .B(n_265), .C(n_264), .Y(n_296) );
AOI221xp5_ASAP7_75t_L g297 ( .A1(n_285), .A2(n_267), .B1(n_270), .B2(n_266), .C(n_272), .Y(n_297) );
AND2x2_ASAP7_75t_SL g298 ( .A(n_293), .B(n_270), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_293), .B(n_261), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_274), .Y(n_300) );
INVx2_ASAP7_75t_L g301 ( .A(n_274), .Y(n_301) );
OAI22xp5_ASAP7_75t_L g302 ( .A1(n_275), .A2(n_263), .B1(n_255), .B2(n_268), .Y(n_302) );
INVx2_ASAP7_75t_L g303 ( .A(n_274), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_281), .Y(n_304) );
INVx4_ASAP7_75t_L g305 ( .A(n_291), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_281), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_281), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_280), .B(n_268), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_293), .B(n_261), .Y(n_309) );
AND2x4_ASAP7_75t_L g310 ( .A(n_294), .B(n_261), .Y(n_310) );
OR2x2_ASAP7_75t_L g311 ( .A(n_280), .B(n_254), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_294), .B(n_258), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_294), .B(n_258), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_282), .Y(n_314) );
BUFx2_ASAP7_75t_L g315 ( .A(n_291), .Y(n_315) );
OR2x2_ASAP7_75t_L g316 ( .A(n_287), .B(n_263), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_282), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_287), .B(n_263), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_278), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_288), .B(n_258), .Y(n_320) );
INVx1_ASAP7_75t_L g321 ( .A(n_278), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_278), .Y(n_322) );
INVx2_ASAP7_75t_SL g323 ( .A(n_291), .Y(n_323) );
AND2x2_ASAP7_75t_L g324 ( .A(n_288), .B(n_258), .Y(n_324) );
AND2x2_ASAP7_75t_L g325 ( .A(n_288), .B(n_255), .Y(n_325) );
INVxp67_ASAP7_75t_L g326 ( .A(n_315), .Y(n_326) );
AND2x2_ASAP7_75t_L g327 ( .A(n_299), .B(n_287), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_319), .B(n_275), .Y(n_328) );
INVx2_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
NAND4xp25_ASAP7_75t_SL g330 ( .A(n_297), .B(n_292), .C(n_290), .D(n_277), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_299), .B(n_295), .Y(n_331) );
INVx2_ASAP7_75t_SL g332 ( .A(n_305), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_304), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g334 ( .A(n_308), .B(n_290), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_301), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_301), .Y(n_337) );
HB1xp67_ASAP7_75t_L g338 ( .A(n_315), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_307), .Y(n_339) );
INVx1_ASAP7_75t_SL g340 ( .A(n_325), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_309), .B(n_295), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_311), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_309), .B(n_283), .Y(n_344) );
INVx2_ASAP7_75t_SL g345 ( .A(n_305), .Y(n_345) );
AND3x1_ASAP7_75t_L g346 ( .A(n_296), .B(n_291), .C(n_275), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_319), .B(n_283), .Y(n_347) );
AND2x4_ASAP7_75t_L g348 ( .A(n_310), .B(n_283), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_321), .B(n_282), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_303), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_321), .B(n_289), .Y(n_352) );
AND2x2_ASAP7_75t_L g353 ( .A(n_322), .B(n_289), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g354 ( .A(n_322), .B(n_279), .Y(n_354) );
AND2x2_ASAP7_75t_L g355 ( .A(n_310), .B(n_279), .Y(n_355) );
NAND2xp33_ASAP7_75t_SL g356 ( .A(n_305), .B(n_279), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_320), .B(n_286), .Y(n_357) );
OR2x2_ASAP7_75t_L g358 ( .A(n_316), .B(n_318), .Y(n_358) );
OR2x2_ASAP7_75t_L g359 ( .A(n_316), .B(n_286), .Y(n_359) );
NOR4xp25_ASAP7_75t_SL g360 ( .A(n_305), .B(n_286), .C(n_12), .D(n_13), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_303), .Y(n_361) );
NOR3xp33_ASAP7_75t_SL g362 ( .A(n_302), .B(n_260), .C(n_13), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_310), .B(n_286), .Y(n_363) );
NOR2x1_ASAP7_75t_R g364 ( .A(n_310), .B(n_286), .Y(n_364) );
AND2x2_ASAP7_75t_L g365 ( .A(n_312), .B(n_284), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_320), .B(n_272), .Y(n_366) );
AOI22xp33_ASAP7_75t_L g367 ( .A1(n_298), .A2(n_272), .B1(n_263), .B2(n_284), .Y(n_367) );
AND2x4_ASAP7_75t_L g368 ( .A(n_312), .B(n_46), .Y(n_368) );
AND2x2_ASAP7_75t_L g369 ( .A(n_313), .B(n_284), .Y(n_369) );
INVx1_ASAP7_75t_SL g370 ( .A(n_340), .Y(n_370) );
OR2x2_ASAP7_75t_L g371 ( .A(n_358), .B(n_343), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_327), .B(n_313), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_333), .Y(n_373) );
INVxp67_ASAP7_75t_SL g374 ( .A(n_338), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_327), .B(n_303), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_343), .B(n_298), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_358), .B(n_306), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_333), .Y(n_378) );
AND2x2_ASAP7_75t_L g379 ( .A(n_344), .B(n_306), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_344), .B(n_306), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_349), .B(n_318), .Y(n_381) );
INVx1_ASAP7_75t_SL g382 ( .A(n_332), .Y(n_382) );
NAND2x1p5_ASAP7_75t_L g383 ( .A(n_346), .B(n_298), .Y(n_383) );
OR2x2_ASAP7_75t_L g384 ( .A(n_349), .B(n_300), .Y(n_384) );
OR2x2_ASAP7_75t_L g385 ( .A(n_331), .B(n_300), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_335), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_365), .B(n_324), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_365), .B(n_324), .Y(n_388) );
NOR2x1_ASAP7_75t_L g389 ( .A(n_330), .B(n_325), .Y(n_389) );
NAND2xp5_ASAP7_75t_L g390 ( .A(n_352), .B(n_323), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_369), .B(n_317), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_329), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_335), .Y(n_393) );
NOR2xp67_ASAP7_75t_L g394 ( .A(n_332), .B(n_323), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_369), .B(n_317), .Y(n_395) );
OR2x2_ASAP7_75t_L g396 ( .A(n_331), .B(n_341), .Y(n_396) );
INVx2_ASAP7_75t_L g397 ( .A(n_329), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_352), .B(n_317), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_339), .Y(n_399) );
HB1xp67_ASAP7_75t_L g400 ( .A(n_326), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_345), .Y(n_401) );
INVx2_ASAP7_75t_SL g402 ( .A(n_345), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_339), .Y(n_403) );
NAND2xp33_ASAP7_75t_SL g404 ( .A(n_362), .B(n_314), .Y(n_404) );
OR2x2_ASAP7_75t_L g405 ( .A(n_341), .B(n_314), .Y(n_405) );
AND2x2_ASAP7_75t_L g406 ( .A(n_355), .B(n_314), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g407 ( .A(n_334), .B(n_328), .Y(n_407) );
INVx2_ASAP7_75t_L g408 ( .A(n_329), .Y(n_408) );
INVxp67_ASAP7_75t_L g409 ( .A(n_346), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_342), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_355), .B(n_284), .Y(n_411) );
AND2x2_ASAP7_75t_L g412 ( .A(n_363), .B(n_353), .Y(n_412) );
INVx2_ASAP7_75t_SL g413 ( .A(n_361), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_363), .B(n_284), .Y(n_414) );
INVx2_ASAP7_75t_SL g415 ( .A(n_361), .Y(n_415) );
AND4x1_ASAP7_75t_L g416 ( .A(n_367), .B(n_11), .C(n_14), .D(n_15), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_353), .B(n_14), .Y(n_417) );
INVxp67_ASAP7_75t_L g418 ( .A(n_356), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_337), .Y(n_419) );
AND2x2_ASAP7_75t_L g420 ( .A(n_348), .B(n_17), .Y(n_420) );
INVx2_ASAP7_75t_SL g421 ( .A(n_337), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_371), .Y(n_422) );
NAND2xp33_ASAP7_75t_L g423 ( .A(n_383), .B(n_342), .Y(n_423) );
INVx1_ASAP7_75t_SL g424 ( .A(n_370), .Y(n_424) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_407), .B(n_366), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_412), .B(n_359), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_371), .B(n_347), .Y(n_427) );
INVx5_ASAP7_75t_L g428 ( .A(n_420), .Y(n_428) );
HB1xp67_ASAP7_75t_L g429 ( .A(n_413), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_412), .B(n_359), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_387), .B(n_388), .Y(n_431) );
NAND2x1p5_ASAP7_75t_L g432 ( .A(n_394), .B(n_368), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_413), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_373), .B(n_378), .Y(n_434) );
OR2x2_ASAP7_75t_L g435 ( .A(n_396), .B(n_357), .Y(n_435) );
NAND2x1_ASAP7_75t_L g436 ( .A(n_402), .B(n_368), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_396), .B(n_354), .Y(n_437) );
NAND2xp5_ASAP7_75t_L g438 ( .A(n_386), .B(n_350), .Y(n_438) );
NAND2xp33_ASAP7_75t_L g439 ( .A(n_383), .B(n_364), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_409), .B(n_364), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_393), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_399), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_403), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_415), .Y(n_444) );
INVxp33_ASAP7_75t_L g445 ( .A(n_383), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_410), .Y(n_446) );
A2O1A1Ixp33_ASAP7_75t_L g447 ( .A1(n_389), .A2(n_368), .B(n_348), .C(n_351), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_400), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_381), .Y(n_449) );
INVxp67_ASAP7_75t_SL g450 ( .A(n_401), .Y(n_450) );
AND2x2_ASAP7_75t_L g451 ( .A(n_387), .B(n_348), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_385), .B(n_351), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_391), .B(n_350), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_402), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_388), .B(n_348), .Y(n_455) );
AOI211xp5_ASAP7_75t_SL g456 ( .A1(n_418), .A2(n_417), .B(n_420), .C(n_374), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_381), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_385), .Y(n_458) );
INVx1_ASAP7_75t_SL g459 ( .A(n_382), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_405), .B(n_351), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_415), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_377), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g463 ( .A1(n_404), .A2(n_360), .B(n_368), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_391), .B(n_347), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_395), .B(n_337), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_451), .B(n_372), .Y(n_466) );
INVxp67_ASAP7_75t_L g467 ( .A(n_429), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_455), .B(n_372), .Y(n_468) );
AOI221xp5_ASAP7_75t_L g469 ( .A1(n_448), .A2(n_404), .B1(n_417), .B2(n_376), .C(n_414), .Y(n_469) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_445), .A2(n_405), .B1(n_390), .B2(n_377), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_422), .B(n_395), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_434), .Y(n_472) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_431), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_453), .B(n_375), .Y(n_474) );
NOR2x1_ASAP7_75t_L g475 ( .A(n_439), .B(n_384), .Y(n_475) );
NAND3xp33_ASAP7_75t_L g476 ( .A(n_456), .B(n_416), .C(n_360), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_434), .Y(n_477) );
AOI22xp5_ASAP7_75t_L g478 ( .A1(n_440), .A2(n_411), .B1(n_414), .B2(n_406), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_427), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_426), .B(n_406), .Y(n_480) );
OAI22xp5_ASAP7_75t_L g481 ( .A1(n_447), .A2(n_375), .B1(n_379), .B2(n_380), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_430), .B(n_411), .Y(n_482) );
OAI32xp33_ASAP7_75t_L g483 ( .A1(n_459), .A2(n_398), .A3(n_384), .B1(n_380), .B2(n_379), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_428), .B(n_421), .Y(n_484) );
INVx3_ASAP7_75t_L g485 ( .A(n_436), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_427), .Y(n_486) );
AOI222xp33_ASAP7_75t_L g487 ( .A1(n_423), .A2(n_421), .B1(n_419), .B2(n_408), .C1(n_397), .C2(n_392), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_438), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_450), .Y(n_489) );
OAI22xp5_ASAP7_75t_L g490 ( .A1(n_432), .A2(n_419), .B1(n_408), .B2(n_397), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g491 ( .A(n_424), .B(n_392), .Y(n_491) );
HB1xp67_ASAP7_75t_L g492 ( .A(n_433), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g493 ( .A(n_425), .B(n_336), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_438), .Y(n_494) );
AOI22xp5_ASAP7_75t_L g495 ( .A1(n_473), .A2(n_449), .B1(n_457), .B2(n_454), .Y(n_495) );
NOR2xp67_ASAP7_75t_L g496 ( .A(n_485), .B(n_428), .Y(n_496) );
OAI21xp33_ASAP7_75t_L g497 ( .A1(n_478), .A2(n_456), .B(n_462), .Y(n_497) );
CKINVDCx16_ASAP7_75t_R g498 ( .A(n_475), .Y(n_498) );
OAI211xp5_ASAP7_75t_SL g499 ( .A1(n_469), .A2(n_463), .B(n_461), .C(n_458), .Y(n_499) );
INVxp33_ASAP7_75t_L g500 ( .A(n_491), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_472), .Y(n_501) );
OR2x2_ASAP7_75t_L g502 ( .A(n_474), .B(n_464), .Y(n_502) );
OAI211xp5_ASAP7_75t_L g503 ( .A1(n_476), .A2(n_428), .B(n_444), .C(n_437), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_477), .Y(n_504) );
O2A1O1Ixp33_ASAP7_75t_L g505 ( .A1(n_489), .A2(n_443), .B(n_441), .C(n_446), .Y(n_505) );
AOI222xp33_ASAP7_75t_L g506 ( .A1(n_489), .A2(n_442), .B1(n_464), .B2(n_453), .C1(n_465), .C2(n_428), .Y(n_506) );
NAND4xp25_ASAP7_75t_SL g507 ( .A(n_487), .B(n_435), .C(n_452), .D(n_432), .Y(n_507) );
OAI221xp5_ASAP7_75t_L g508 ( .A1(n_485), .A2(n_460), .B1(n_336), .B2(n_26), .C(n_27), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_488), .Y(n_509) );
AOI21xp33_ASAP7_75t_L g510 ( .A1(n_467), .A2(n_19), .B(n_23), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_L g511 ( .A1(n_483), .A2(n_29), .B(n_30), .C(n_31), .Y(n_511) );
NOR2xp33_ASAP7_75t_L g512 ( .A(n_498), .B(n_467), .Y(n_512) );
XNOR2x1_ASAP7_75t_L g513 ( .A(n_495), .B(n_470), .Y(n_513) );
AOI222xp33_ASAP7_75t_L g514 ( .A1(n_497), .A2(n_499), .B1(n_503), .B2(n_500), .C1(n_504), .C2(n_501), .Y(n_514) );
AOI222xp33_ASAP7_75t_L g515 ( .A1(n_503), .A2(n_481), .B1(n_491), .B2(n_494), .C1(n_486), .C2(n_479), .Y(n_515) );
AOI32xp33_ASAP7_75t_L g516 ( .A1(n_507), .A2(n_490), .A3(n_493), .B1(n_466), .B2(n_468), .Y(n_516) );
INVxp33_ASAP7_75t_SL g517 ( .A(n_506), .Y(n_517) );
NAND3xp33_ASAP7_75t_L g518 ( .A(n_511), .B(n_492), .C(n_484), .Y(n_518) );
AOI221xp5_ASAP7_75t_L g519 ( .A1(n_505), .A2(n_492), .B1(n_471), .B2(n_482), .C(n_480), .Y(n_519) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_502), .B(n_32), .Y(n_520) );
NOR5xp2_ASAP7_75t_L g521 ( .A(n_518), .B(n_508), .C(n_509), .D(n_510), .E(n_496), .Y(n_521) );
NAND5xp2_ASAP7_75t_L g522 ( .A(n_514), .B(n_33), .C(n_37), .D(n_43), .E(n_44), .Y(n_522) );
AOI221xp5_ASAP7_75t_L g523 ( .A1(n_517), .A2(n_47), .B1(n_48), .B2(n_53), .C(n_56), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_512), .Y(n_524) );
AOI211xp5_ASAP7_75t_L g525 ( .A1(n_519), .A2(n_57), .B(n_58), .C(n_60), .Y(n_525) );
NOR3xp33_ASAP7_75t_L g526 ( .A(n_522), .B(n_516), .C(n_520), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_524), .Y(n_527) );
NAND5xp2_ASAP7_75t_L g528 ( .A(n_525), .B(n_515), .C(n_513), .D(n_64), .E(n_69), .Y(n_528) );
NAND3xp33_ASAP7_75t_L g529 ( .A(n_527), .B(n_521), .C(n_523), .Y(n_529) );
INVxp67_ASAP7_75t_SL g530 ( .A(n_526), .Y(n_530) );
INVx2_ASAP7_75t_L g531 ( .A(n_530), .Y(n_531) );
INVx2_ASAP7_75t_L g532 ( .A(n_531), .Y(n_532) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_532), .A2(n_529), .B1(n_528), .B2(n_70), .Y(n_533) );
INVx2_ASAP7_75t_SL g534 ( .A(n_533), .Y(n_534) );
OA21x2_ASAP7_75t_L g535 ( .A1(n_534), .A2(n_62), .B(n_63), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g536 ( .A1(n_535), .A2(n_71), .B1(n_72), .B2(n_76), .Y(n_536) );
endmodule