module real_jpeg_18495_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_475;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_502;
wire n_418;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_0),
.A2(n_19),
.B(n_501),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_0),
.B(n_502),
.Y(n_501)
);

AND2x2_ASAP7_75t_SL g36 ( 
.A(n_1),
.B(n_37),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_1),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_1),
.B(n_97),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_1),
.B(n_142),
.Y(n_141)
);

NAND2x1p5_ASAP7_75t_L g190 ( 
.A(n_1),
.B(n_191),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_1),
.B(n_138),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_1),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_1),
.B(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_2),
.Y(n_92)
);

BUFx3_ASAP7_75t_L g166 ( 
.A(n_2),
.Y(n_166)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_2),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_3),
.Y(n_66)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_3),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g392 ( 
.A(n_3),
.Y(n_392)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_4),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_4),
.A2(n_11),
.B1(n_116),
.B2(n_120),
.Y(n_115)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_4),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_4),
.B(n_56),
.Y(n_195)
);

AND2x2_ASAP7_75t_L g266 ( 
.A(n_4),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_4),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_4),
.B(n_457),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_4),
.B(n_499),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_5),
.B(n_44),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g63 ( 
.A(n_5),
.B(n_64),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_5),
.B(n_86),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_5),
.B(n_111),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_5),
.B(n_91),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g242 ( 
.A(n_5),
.B(n_243),
.Y(n_242)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_5),
.B(n_293),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_SL g459 ( 
.A(n_5),
.B(n_460),
.Y(n_459)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_6),
.Y(n_84)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_6),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g138 ( 
.A(n_6),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_6),
.Y(n_375)
);

INVxp33_ASAP7_75t_L g502 ( 
.A(n_7),
.Y(n_502)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_8),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_8),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g169 ( 
.A(n_8),
.Y(n_169)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_8),
.Y(n_269)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_8),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_9),
.B(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_SL g69 ( 
.A(n_9),
.B(n_70),
.Y(n_69)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_9),
.B(n_94),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_9),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_9),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_9),
.B(n_325),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_9),
.B(n_331),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_9),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_10),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_10),
.B(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_10),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_10),
.B(n_164),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_10),
.B(n_346),
.Y(n_345)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_10),
.B(n_392),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_10),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_SL g427 ( 
.A(n_10),
.B(n_428),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_11),
.B(n_33),
.Y(n_32)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_11),
.B(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_11),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_11),
.B(n_357),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_11),
.B(n_378),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_11),
.B(n_407),
.Y(n_406)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_12),
.Y(n_79)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_12),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_13),
.B(n_54),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g72 ( 
.A(n_13),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_13),
.B(n_84),
.Y(n_83)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_13),
.B(n_207),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g265 ( 
.A(n_13),
.B(n_91),
.Y(n_265)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_13),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_14),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_15),
.Y(n_88)
);

BUFx4f_ASAP7_75t_L g109 ( 
.A(n_15),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g334 ( 
.A(n_15),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_16),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_16),
.B(n_77),
.Y(n_147)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_16),
.B(n_171),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g350 ( 
.A(n_16),
.B(n_351),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_SL g388 ( 
.A(n_16),
.B(n_389),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_16),
.B(n_415),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_16),
.B(n_421),
.Y(n_420)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_17),
.Y(n_62)
);

BUFx8_ASAP7_75t_L g104 ( 
.A(n_17),
.Y(n_104)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_17),
.Y(n_220)
);

BUFx3_ASAP7_75t_L g283 ( 
.A(n_17),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_476),
.Y(n_19)
);

OAI21xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_443),
.B(n_475),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2x1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_437),
.Y(n_22)
);

NAND4xp25_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_225),
.C(n_308),
.D(n_313),
.Y(n_23)
);

NOR2x1_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_174),
.Y(n_24)
);

NOR2xp67_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_148),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g439 ( 
.A(n_26),
.B(n_148),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_99),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_27),
.B(n_100),
.C(n_125),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_67),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.Y(n_28)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_29),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_42),
.B2(n_43),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_36),
.B1(n_40),
.B2(n_41),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_32),
.B(n_41),
.C(n_42),
.Y(n_224)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_36),
.A2(n_41),
.B1(n_59),
.B2(n_128),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_37),
.Y(n_70)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_42),
.A2(n_43),
.B1(n_295),
.B2(n_299),
.Y(n_294)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g471 ( 
.A(n_43),
.B(n_292),
.C(n_299),
.Y(n_471)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_47),
.Y(n_179)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_58),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_49),
.A2(n_52),
.B1(n_53),
.B2(n_57),
.Y(n_48)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_49),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_L g199 ( 
.A1(n_49),
.A2(n_53),
.B(n_58),
.C(n_200),
.Y(n_199)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_51),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_52),
.B(n_57),
.Y(n_200)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_55),
.Y(n_417)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_59),
.B(n_61),
.C(n_63),
.Y(n_58)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_59),
.A2(n_63),
.B1(n_128),
.B2(n_129),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_59),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g466 ( 
.A1(n_59),
.A2(n_96),
.B1(n_128),
.B2(n_159),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_59),
.B(n_159),
.C(n_467),
.Y(n_487)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_61),
.B(n_127),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g491 ( 
.A(n_62),
.Y(n_491)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_63),
.Y(n_129)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_63),
.B(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_66),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_67),
.B(n_178),
.C(n_179),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_80),
.C(n_89),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_SL g152 ( 
.A(n_68),
.B(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_69),
.B(n_72),
.C(n_76),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_76),
.Y(n_71)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_80),
.A2(n_81),
.B1(n_89),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_82),
.A2(n_83),
.B1(n_85),
.B2(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g430 ( 
.A(n_84),
.Y(n_430)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_85),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_85),
.A2(n_161),
.B1(n_222),
.B2(n_223),
.Y(n_221)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_87),
.Y(n_142)
);

INVx2_ASAP7_75t_L g378 ( 
.A(n_87),
.Y(n_378)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g426 ( 
.A(n_88),
.Y(n_426)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_89),
.Y(n_154)
);

MAJx2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_93),
.C(n_96),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_90),
.A2(n_96),
.B1(n_158),
.B2(n_159),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_90),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_92),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_SL g156 ( 
.A(n_93),
.B(n_157),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g207 ( 
.A(n_95),
.Y(n_207)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_96),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_96),
.A2(n_141),
.B1(n_159),
.B2(n_259),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_96),
.B(n_259),
.C(n_302),
.Y(n_472)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_98),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_125),
.Y(n_99)
);

XOR2x2_ASAP7_75t_SL g100 ( 
.A(n_101),
.B(n_115),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_114),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_102),
.B(n_184),
.C(n_185),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_103),
.B(n_105),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_103),
.B(n_107),
.C(n_110),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B1(n_110),
.B2(n_113),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g113 ( 
.A(n_110),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_141),
.Y(n_140)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_112),
.Y(n_119)
);

XNOR2x1_ASAP7_75t_SL g322 ( 
.A(n_113),
.B(n_141),
.Y(n_322)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_114),
.Y(n_185)
);

AOI21xp5_ASAP7_75t_L g130 ( 
.A1(n_115),
.A2(n_131),
.B(n_134),
.Y(n_130)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_115),
.Y(n_184)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx4_ASAP7_75t_SL g408 ( 
.A(n_118),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_120),
.Y(n_133)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_122),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_123),
.Y(n_458)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_124),
.Y(n_173)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_124),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_124),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_130),
.C(n_139),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g150 ( 
.A(n_126),
.B(n_130),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_129),
.B(n_264),
.C(n_270),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_132),
.B(n_168),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_132),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_136),
.Y(n_134)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g149 ( 
.A(n_139),
.B(n_150),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_143),
.C(n_146),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g319 ( 
.A(n_140),
.B(n_320),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_141),
.A2(n_222),
.B1(n_223),
.B2(n_259),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_141),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_141),
.B(n_223),
.C(n_254),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_143),
.A2(n_144),
.B1(n_146),
.B2(n_147),
.Y(n_320)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_151),
.C(n_155),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_149),
.B(n_336),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_151),
.A2(n_152),
.B1(n_155),
.B2(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_155),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_160),
.C(n_162),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g317 ( 
.A(n_156),
.B(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_160),
.B(n_162),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_161),
.B(n_216),
.C(n_223),
.Y(n_261)
);

MAJx2_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.C(n_170),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g360 ( 
.A(n_163),
.B(n_170),
.Y(n_360)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_167),
.B(n_360),
.Y(n_359)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

OAI21x1_ASAP7_75t_SL g438 ( 
.A1(n_174),
.A2(n_439),
.B(n_440),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

OR2x2_ASAP7_75t_L g440 ( 
.A(n_175),
.B(n_176),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_180),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_177),
.B(n_181),
.C(n_204),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_203),
.B2(n_204),
.Y(n_180)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_183),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_199),
.B1(n_201),
.B2(n_202),
.Y(n_186)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_189),
.B1(n_197),
.B2(n_198),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_190),
.A2(n_194),
.B1(n_195),
.B2(n_196),
.Y(n_189)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_190),
.Y(n_196)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_196),
.C(n_198),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_SL g198 ( 
.A(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_199),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g250 ( 
.A(n_199),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_201),
.B(n_250),
.C(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_214),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_205),
.B(n_224),
.C(n_231),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_208),
.Y(n_205)
);

MAJx2_ASAP7_75t_L g245 ( 
.A(n_206),
.B(n_209),
.C(n_213),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_SL g208 ( 
.A(n_209),
.B(n_213),
.Y(n_208)
);

INVx4_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_211),
.Y(n_469)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_211),
.Y(n_499)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_212),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_SL g453 ( 
.A1(n_213),
.A2(n_454),
.B1(n_455),
.B2(n_456),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_213),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_213),
.B(n_455),
.C(n_459),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_224),
.Y(n_214)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_215),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_221),
.Y(n_215)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_218),
.Y(n_460)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_222),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g380 ( 
.A(n_222),
.B(n_330),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_223),
.B(n_330),
.Y(n_329)
);

A2O1A1O1Ixp25_ASAP7_75t_L g437 ( 
.A1(n_225),
.A2(n_308),
.B(n_438),
.C(n_441),
.D(n_442),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_271),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_226),
.B(n_271),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_248),
.C(n_252),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_227),
.A2(n_228),
.B1(n_252),
.B2(n_312),
.Y(n_311)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_230),
.B1(n_232),
.B2(n_247),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_233),
.C(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_232),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_235),
.B2(n_246),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g246 ( 
.A(n_235),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_245),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_241),
.B2(n_242),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_238),
.B(n_241),
.C(n_245),
.Y(n_278)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g496 ( 
.A1(n_241),
.A2(n_242),
.B1(n_497),
.B2(n_498),
.Y(n_496)
);

INVx2_ASAP7_75t_SL g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_242),
.B(n_281),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_242),
.B(n_286),
.C(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_249),
.B(n_311),
.Y(n_310)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_252),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_260),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_261),
.C(n_262),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_258),
.Y(n_253)
);

INVx4_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx4_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_270),
.Y(n_263)
);

INVx1_ASAP7_75t_SL g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_266),
.Y(n_270)
);

INVx6_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_272),
.B(n_274),
.C(n_474),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_274),
.B(n_288),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_276),
.B1(n_277),
.B2(n_287),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_275),
.B(n_278),
.C(n_279),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_277),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_SL g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

AO22x1_ASAP7_75t_SL g279 ( 
.A1(n_280),
.A2(n_284),
.B1(n_285),
.B2(n_286),
.Y(n_279)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_281),
.Y(n_463)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

INVx1_ASAP7_75t_SL g286 ( 
.A(n_284),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_288),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_289),
.B(n_300),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g449 ( 
.A(n_290),
.B(n_291),
.C(n_300),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_294),
.Y(n_291)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

INVx5_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx5_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_301),
.B(n_302),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_303),
.B(n_468),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g489 ( 
.A(n_303),
.B(n_490),
.Y(n_489)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_309),
.B(n_310),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_338),
.B(n_436),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_335),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_315),
.B(n_335),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.C(n_321),
.Y(n_315)
);

AOI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_316),
.A2(n_317),
.B1(n_362),
.B2(n_363),
.Y(n_361)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_319),
.B(n_321),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_323),
.C(n_329),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_322),
.A2(n_323),
.B1(n_324),
.B2(n_343),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_322),
.Y(n_343)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_SL g341 ( 
.A(n_329),
.B(n_342),
.Y(n_341)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

INVx3_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g405 ( 
.A(n_334),
.Y(n_405)
);

AOI21x1_ASAP7_75t_SL g338 ( 
.A1(n_339),
.A2(n_364),
.B(n_435),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_361),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g435 ( 
.A(n_340),
.B(n_361),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_344),
.C(n_359),
.Y(n_340)
);

XNOR2xp5_ASAP7_75t_L g381 ( 
.A(n_341),
.B(n_382),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_359),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_350),
.C(n_356),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_345),
.B(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_349),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_350),
.B(n_356),
.Y(n_369)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx2_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

BUFx3_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx3_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_363),
.Y(n_362)
);

OAI21x1_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_383),
.B(n_434),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_381),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_366),
.B(n_381),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.C(n_379),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_L g393 ( 
.A1(n_367),
.A2(n_368),
.B1(n_394),
.B2(n_396),
.Y(n_393)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g394 ( 
.A1(n_370),
.A2(n_379),
.B1(n_380),
.B2(n_395),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_370),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_376),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_372),
.B1(n_376),
.B2(n_377),
.Y(n_386)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_384),
.A2(n_397),
.B(n_433),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_393),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_SL g433 ( 
.A(n_385),
.B(n_393),
.Y(n_433)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.C(n_391),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_410),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g410 ( 
.A1(n_387),
.A2(n_388),
.B1(n_391),
.B2(n_411),
.Y(n_410)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_391),
.Y(n_411)
);

INVxp67_ASAP7_75t_SL g396 ( 
.A(n_394),
.Y(n_396)
);

OAI21xp5_ASAP7_75t_SL g397 ( 
.A1(n_398),
.A2(n_412),
.B(n_432),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_399),
.B(n_409),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g432 ( 
.A(n_399),
.B(n_409),
.Y(n_432)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_400),
.B(n_406),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_400),
.B(n_406),
.Y(n_418)
);

INVx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_408),
.Y(n_407)
);

AOI21xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_419),
.B(n_431),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_418),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_SL g431 ( 
.A(n_414),
.B(n_418),
.Y(n_431)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_427),
.Y(n_419)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_424),
.Y(n_423)
);

INVx3_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_429),
.Y(n_428)
);

INVx6_ASAP7_75t_L g429 ( 
.A(n_430),
.Y(n_429)
);

CKINVDCx14_ASAP7_75t_R g443 ( 
.A(n_444),
.Y(n_443)
);

OR2x2_ASAP7_75t_SL g444 ( 
.A(n_445),
.B(n_473),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_473),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_446),
.B(n_447),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_446),
.B(n_448),
.C(n_464),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g447 ( 
.A(n_448),
.B(n_464),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_450),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_449),
.B(n_451),
.C(n_462),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_462),
.Y(n_450)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_452),
.A2(n_453),
.B1(n_459),
.B2(n_461),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_453),
.Y(n_452)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_456),
.Y(n_455)
);

INVx8_ASAP7_75t_L g457 ( 
.A(n_458),
.Y(n_457)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_459),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_465),
.B(n_470),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_465),
.B(n_471),
.C(n_472),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g465 ( 
.A(n_466),
.B(n_467),
.Y(n_465)
);

INVx3_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_471),
.B(n_472),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_477),
.B(n_500),
.Y(n_476)
);

INVxp33_ASAP7_75t_L g477 ( 
.A(n_478),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_480),
.Y(n_478)
);

NOR2xp67_ASAP7_75t_SL g500 ( 
.A(n_479),
.B(n_480),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_481),
.B(n_482),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_484),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_485),
.A2(n_486),
.B1(n_493),
.B2(n_494),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_486),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_L g486 ( 
.A(n_487),
.B(n_488),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_489),
.B(n_492),
.Y(n_488)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_491),
.Y(n_490)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_SL g494 ( 
.A(n_495),
.B(n_496),
.Y(n_494)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_498),
.Y(n_497)
);


endmodule