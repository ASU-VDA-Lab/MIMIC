module fake_jpeg_2572_n_124 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_124);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_124;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

BUFx4f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_27),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_3),
.Y(n_45)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_3),
.Y(n_46)
);

BUFx12_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_47),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_38),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_45),
.Y(n_54)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_50),
.Y(n_58)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

NAND3xp33_ASAP7_75t_L g65 ( 
.A(n_54),
.B(n_46),
.C(n_1),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_52),
.A2(n_35),
.B1(n_44),
.B2(n_43),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_56),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_52),
.A2(n_46),
.B1(n_42),
.B2(n_41),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_37),
.C(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_35),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_59),
.B(n_64),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_40),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_70),
.Y(n_84)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_63),
.Y(n_66)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_66),
.Y(n_85)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_0),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_55),
.B(n_2),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_71),
.B(n_73),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_72),
.B(n_76),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_59),
.B(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_60),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_61),
.A2(n_37),
.B1(n_47),
.B2(n_6),
.Y(n_75)
);

OR2x2_ASAP7_75t_L g90 ( 
.A(n_75),
.B(n_4),
.Y(n_90)
);

INVx13_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_77),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_62),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_80),
.B(n_82),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_72),
.B(n_62),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_70),
.B(n_61),
.Y(n_83)
);

OAI32xp33_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_77),
.A3(n_21),
.B1(n_22),
.B2(n_33),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_66),
.A2(n_60),
.B1(n_57),
.B2(n_58),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_86),
.A2(n_89),
.B1(n_7),
.B2(n_8),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_58),
.B1(n_5),
.B2(n_7),
.Y(n_89)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_90),
.B(n_14),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_93),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_101),
.B1(n_90),
.B2(n_86),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_8),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_83),
.A2(n_9),
.B(n_10),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_95),
.Y(n_106)
);

NAND3xp33_ASAP7_75t_L g95 ( 
.A(n_81),
.B(n_9),
.C(n_10),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_84),
.B(n_12),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_96),
.B(n_98),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_87),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_99),
.B(n_100),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_15),
.Y(n_101)
);

BUFx24_ASAP7_75t_SL g104 ( 
.A(n_101),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_28),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_110),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_102),
.A2(n_89),
.B1(n_78),
.B2(n_20),
.Y(n_108)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_108),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_93),
.A2(n_17),
.B1(n_18),
.B2(n_23),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_100),
.C(n_26),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_114),
.B(n_116),
.C(n_109),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_107),
.B(n_25),
.Y(n_115)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_115),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_117),
.B(n_103),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g120 ( 
.A1(n_119),
.A2(n_118),
.B(n_113),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_112),
.C(n_106),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_121),
.A2(n_111),
.B(n_30),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_122),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_123),
.B(n_31),
.Y(n_124)
);


endmodule