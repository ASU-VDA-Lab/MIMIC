module fake_jpeg_3116_n_40 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_40);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_40;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_39;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

INVx2_ASAP7_75t_L g8 ( 
.A(n_3),
.Y(n_8)
);

INVx3_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_4),
.B(n_3),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_12),
.B(n_1),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_15),
.B(n_19),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g16 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g24 ( 
.A1(n_16),
.A2(n_18),
.B1(n_22),
.B2(n_10),
.Y(n_24)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_17),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g18 ( 
.A1(n_11),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_4),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_11),
.B(n_0),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_21),
.Y(n_29)
);

INVx13_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_9),
.A2(n_0),
.B(n_5),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g23 ( 
.A(n_20),
.B(n_7),
.C(n_10),
.Y(n_23)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_25),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_24),
.A2(n_28),
.B1(n_22),
.B2(n_21),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_17),
.B(n_13),
.C(n_14),
.Y(n_25)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_19),
.B(n_13),
.C(n_14),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_27),
.B(n_29),
.Y(n_35)
);

OAI22x1_ASAP7_75t_SL g28 ( 
.A1(n_22),
.A2(n_16),
.B1(n_18),
.B2(n_21),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_26),
.B(n_15),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_32),
.C(n_33),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_29),
.B(n_22),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_35),
.B(n_5),
.C(n_6),
.Y(n_37)
);

AOI21xp5_ASAP7_75t_SL g36 ( 
.A1(n_35),
.A2(n_28),
.B(n_30),
.Y(n_36)
);

AOI21xp5_ASAP7_75t_SL g39 ( 
.A1(n_36),
.A2(n_37),
.B(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_39),
.A2(n_33),
.B1(n_34),
.B2(n_31),
.Y(n_40)
);


endmodule