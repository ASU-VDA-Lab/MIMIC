module fake_jpeg_18622_n_264 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_264);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_264;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_12),
.B(n_2),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

INVx8_ASAP7_75t_SL g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_4),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx5_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_17),
.B(n_15),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_17),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_41),
.B(n_31),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_45),
.Y(n_48)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_45),
.B1(n_39),
.B2(n_44),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_49),
.A2(n_53),
.B1(n_57),
.B2(n_58),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_44),
.A2(n_21),
.B1(n_34),
.B2(n_33),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_63),
.B1(n_26),
.B2(n_46),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_40),
.Y(n_51)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_51),
.B(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_44),
.A2(n_21),
.B1(n_26),
.B2(n_18),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_36),
.B(n_35),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_54),
.A2(n_36),
.B(n_38),
.Y(n_87)
);

BUFx16f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_37),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_45),
.A2(n_16),
.B1(n_20),
.B2(n_23),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_59),
.B(n_41),
.Y(n_74)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_62),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_44),
.A2(n_45),
.B1(n_39),
.B2(n_43),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_40),
.B(n_28),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_33),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_42),
.A2(n_27),
.B1(n_31),
.B2(n_22),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_65),
.A2(n_69),
.B1(n_42),
.B2(n_43),
.Y(n_72)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_66),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_42),
.A2(n_27),
.B1(n_18),
.B2(n_22),
.Y(n_69)
);

NAND2xp33_ASAP7_75t_SL g70 ( 
.A(n_54),
.B(n_36),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_70),
.B(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_71),
.B(n_74),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_72),
.A2(n_95),
.B1(n_101),
.B2(n_87),
.Y(n_129)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_61),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g112 ( 
.A(n_73),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_52),
.A2(n_43),
.B1(n_42),
.B2(n_29),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_75),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_59),
.B(n_30),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_76),
.B(n_79),
.Y(n_133)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_78),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_30),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_80),
.B(n_102),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_47),
.B(n_29),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_81),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_48),
.Y(n_83)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

BUFx2_ASAP7_75t_SL g84 ( 
.A(n_55),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_84),
.Y(n_123)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_60),
.Y(n_86)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_86),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_88),
.B(n_91),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_51),
.A2(n_25),
.B(n_19),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_53),
.B(n_25),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_90),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_36),
.Y(n_91)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_67),
.Y(n_92)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_66),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_94),
.B(n_2),
.Y(n_139)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_97),
.Y(n_137)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_98),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_57),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g120 ( 
.A1(n_99),
.A2(n_100),
.B(n_105),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g100 ( 
.A1(n_54),
.A2(n_19),
.B(n_1),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_55),
.B(n_0),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_69),
.Y(n_102)
);

BUFx4f_ASAP7_75t_SL g103 ( 
.A(n_55),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_104),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_68),
.A2(n_35),
.B1(n_34),
.B2(n_33),
.Y(n_105)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_62),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_34),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_36),
.C(n_52),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_113),
.B(n_134),
.C(n_106),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_82),
.A2(n_67),
.B1(n_49),
.B2(n_46),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_117),
.A2(n_124),
.B1(n_128),
.B2(n_105),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_97),
.A2(n_67),
.B1(n_38),
.B2(n_46),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_36),
.B(n_52),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_126),
.A2(n_130),
.B(n_9),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_46),
.B1(n_61),
.B2(n_56),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_138),
.B1(n_94),
.B2(n_77),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_61),
.B1(n_56),
.B2(n_34),
.Y(n_128)
);

A2O1A1Ixp33_ASAP7_75t_SL g165 ( 
.A1(n_129),
.A2(n_15),
.B(n_12),
.C(n_13),
.Y(n_165)
);

OAI32xp33_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_56),
.A3(n_35),
.B1(n_33),
.B2(n_28),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_28),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_83),
.B(n_28),
.C(n_3),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g138 ( 
.A1(n_95),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_138)
);

AO22x1_ASAP7_75t_L g145 ( 
.A1(n_139),
.A2(n_88),
.B1(n_98),
.B2(n_85),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_156),
.Y(n_174)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_121),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_142),
.B(n_149),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_143),
.A2(n_145),
.B(n_160),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_90),
.B1(n_86),
.B2(n_77),
.Y(n_144)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_119),
.Y(n_146)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_146),
.Y(n_188)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_147),
.Y(n_171)
);

AO22x1_ASAP7_75t_L g148 ( 
.A1(n_118),
.A2(n_91),
.B1(n_107),
.B2(n_106),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_125),
.B(n_103),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_135),
.B(n_91),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_150),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_166),
.Y(n_168)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g153 ( 
.A(n_135),
.B(n_3),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_157),
.Y(n_178)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_154),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_118),
.A2(n_92),
.B1(n_73),
.B2(n_103),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_114),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_161),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_132),
.B(n_6),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_162),
.C(n_111),
.Y(n_169)
);

OAI32xp33_ASAP7_75t_L g160 ( 
.A1(n_110),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_108),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_111),
.B(n_93),
.C(n_11),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_133),
.B(n_93),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_163),
.B(n_108),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_164),
.A2(n_110),
.B(n_139),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_165),
.A2(n_116),
.B1(n_124),
.B2(n_137),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_114),
.B(n_15),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_180),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_169),
.B(n_179),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_151),
.B(n_113),
.C(n_115),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_181),
.C(n_185),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_115),
.Y(n_172)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_172),
.Y(n_196)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_173),
.A2(n_145),
.B(n_143),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_134),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_122),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_155),
.B(n_137),
.C(n_120),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_182),
.B(n_186),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_148),
.B(n_120),
.C(n_122),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_148),
.B(n_130),
.C(n_131),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_187),
.B(n_164),
.Y(n_194)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_171),
.Y(n_191)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_191),
.Y(n_209)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_193),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_194),
.B(n_178),
.C(n_130),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_175),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_195),
.B(n_198),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_167),
.B(n_145),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_181),
.A2(n_162),
.B1(n_165),
.B2(n_160),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_199),
.A2(n_123),
.B(n_188),
.Y(n_220)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_200),
.B(n_201),
.Y(n_216)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_189),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_202),
.B(n_203),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_175),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_183),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_204),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_184),
.A2(n_154),
.B1(n_116),
.B2(n_136),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_205),
.A2(n_207),
.B1(n_177),
.B2(n_159),
.Y(n_215)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_183),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_206),
.B(n_123),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_184),
.A2(n_174),
.B1(n_187),
.B2(n_185),
.Y(n_207)
);

OAI321xp33_ASAP7_75t_L g210 ( 
.A1(n_192),
.A2(n_176),
.A3(n_174),
.B1(n_165),
.B2(n_182),
.C(n_140),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_210),
.B(n_221),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_192),
.A2(n_170),
.B1(n_176),
.B2(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

AOI322xp5_ASAP7_75t_L g214 ( 
.A1(n_197),
.A2(n_178),
.A3(n_177),
.B1(n_173),
.B2(n_186),
.C1(n_165),
.C2(n_169),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_214),
.B(n_208),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_215),
.B(n_222),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_205),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_L g226 ( 
.A1(n_220),
.A2(n_199),
.B(n_206),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_207),
.A2(n_188),
.B1(n_128),
.B2(n_146),
.Y(n_222)
);

INVx4_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_223),
.A2(n_224),
.B(n_200),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_SL g224 ( 
.A1(n_198),
.A2(n_202),
.B(n_201),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_SL g225 ( 
.A(n_213),
.B(n_208),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_SL g246 ( 
.A(n_225),
.B(n_226),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_227),
.B(n_231),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_217),
.B(n_190),
.C(n_194),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_232),
.C(n_234),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_196),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_L g241 ( 
.A1(n_233),
.A2(n_212),
.B(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_215),
.B(n_191),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_219),
.B(n_193),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_235),
.B(n_237),
.C(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_222),
.B(n_224),
.C(n_216),
.Y(n_237)
);

AOI322xp5_ASAP7_75t_L g238 ( 
.A1(n_230),
.A2(n_210),
.A3(n_216),
.B1(n_211),
.B2(n_209),
.C1(n_221),
.C2(n_223),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g250 ( 
.A(n_238),
.B(n_245),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_236),
.A2(n_212),
.B1(n_218),
.B2(n_211),
.Y(n_240)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_240),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_241),
.A2(n_242),
.B(n_237),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_228),
.A2(n_209),
.B(n_109),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_243),
.B(n_229),
.Y(n_248)
);

NOR2xp67_ASAP7_75t_L g245 ( 
.A(n_225),
.B(n_109),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_243),
.B(n_235),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_247),
.B(n_249),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_251),
.C(n_239),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_239),
.B(n_234),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_250),
.A2(n_244),
.B(n_246),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_254),
.Y(n_257)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_247),
.B(n_246),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_256),
.A2(n_251),
.B(n_248),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_255),
.B(n_252),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_258),
.B(n_259),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_257),
.B(n_119),
.C(n_112),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_112),
.B(n_9),
.Y(n_262)
);

NAND3xp33_ASAP7_75t_SL g263 ( 
.A(n_262),
.B(n_14),
.C(n_260),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_263),
.B(n_14),
.Y(n_264)
);


endmodule