module real_aes_8724_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_635;
wire n_503;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_552;
wire n_602;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_713;
wire n_288;
wire n_404;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_354;
wire n_265;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_266;
wire n_183;
wire n_312;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_639;
wire n_546;
wire n_587;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_719;
wire n_473;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g262 ( .A1(n_0), .A2(n_263), .B(n_264), .C(n_267), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_1), .B(n_204), .Y(n_268) );
INVx1_ASAP7_75t_L g110 ( .A(n_2), .Y(n_110) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_3), .B(n_174), .Y(n_240) );
A2O1A1Ixp33_ASAP7_75t_L g453 ( .A1(n_4), .A2(n_144), .B(n_147), .C(n_454), .Y(n_453) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_5), .A2(n_164), .B(n_494), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g194 ( .A1(n_6), .A2(n_164), .B(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_7), .B(n_204), .Y(n_500) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_8), .A2(n_131), .B(n_184), .Y(n_183) );
AND2x6_ASAP7_75t_L g144 ( .A(n_9), .B(n_145), .Y(n_144) );
A2O1A1Ixp33_ASAP7_75t_L g146 ( .A1(n_10), .A2(n_144), .B(n_147), .C(n_150), .Y(n_146) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_11), .A2(n_45), .B1(n_118), .B2(n_119), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_11), .Y(n_118) );
INVx1_ASAP7_75t_L g107 ( .A(n_12), .Y(n_107) );
NOR2xp33_ASAP7_75t_L g442 ( .A(n_12), .B(n_41), .Y(n_442) );
INVx1_ASAP7_75t_L g470 ( .A(n_13), .Y(n_470) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_14), .B(n_154), .Y(n_456) );
INVx1_ASAP7_75t_L g136 ( .A(n_15), .Y(n_136) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_16), .B(n_174), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_17), .A2(n_152), .B(n_478), .C(n_480), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_18), .B(n_204), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_19), .B(n_228), .Y(n_513) );
A2O1A1Ixp33_ASAP7_75t_L g223 ( .A1(n_20), .A2(n_147), .B(n_191), .C(n_224), .Y(n_223) );
A2O1A1Ixp33_ASAP7_75t_L g486 ( .A1(n_21), .A2(n_156), .B(n_266), .C(n_487), .Y(n_486) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_22), .B(n_154), .Y(n_532) );
CKINVDCx20_ASAP7_75t_R g741 ( .A(n_23), .Y(n_741) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_24), .B(n_154), .Y(n_521) );
CKINVDCx16_ASAP7_75t_R g528 ( .A(n_25), .Y(n_528) );
INVx1_ASAP7_75t_L g520 ( .A(n_26), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g186 ( .A1(n_27), .A2(n_147), .B(n_187), .C(n_191), .Y(n_186) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_28), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g452 ( .A(n_29), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_30), .A2(n_102), .B1(n_115), .B2(n_744), .Y(n_101) );
INVx1_ASAP7_75t_L g511 ( .A(n_31), .Y(n_511) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_32), .A2(n_164), .B(n_260), .Y(n_259) );
INVx2_ASAP7_75t_L g142 ( .A(n_33), .Y(n_142) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_34), .A2(n_166), .B(n_177), .C(n_212), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g459 ( .A(n_35), .Y(n_459) );
A2O1A1Ixp33_ASAP7_75t_L g496 ( .A1(n_36), .A2(n_266), .B(n_497), .C(n_499), .Y(n_496) );
INVxp67_ASAP7_75t_L g512 ( .A(n_37), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g188 ( .A(n_38), .B(n_189), .Y(n_188) );
CKINVDCx14_ASAP7_75t_R g495 ( .A(n_39), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_40), .A2(n_147), .B(n_191), .C(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_41), .B(n_107), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_42), .A2(n_267), .B(n_468), .C(n_469), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_43), .B(n_222), .Y(n_221) );
CKINVDCx20_ASAP7_75t_R g159 ( .A(n_44), .Y(n_159) );
INVx1_ASAP7_75t_L g119 ( .A(n_45), .Y(n_119) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_46), .B(n_174), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g185 ( .A(n_47), .B(n_164), .Y(n_185) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_48), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g508 ( .A(n_49), .Y(n_508) );
A2O1A1Ixp33_ASAP7_75t_L g165 ( .A1(n_50), .A2(n_166), .B(n_168), .C(n_177), .Y(n_165) );
INVx1_ASAP7_75t_L g265 ( .A(n_51), .Y(n_265) );
INVx1_ASAP7_75t_L g169 ( .A(n_52), .Y(n_169) );
INVx1_ASAP7_75t_L g485 ( .A(n_53), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_54), .B(n_164), .Y(n_163) );
OAI22xp5_ASAP7_75t_SL g732 ( .A1(n_55), .A2(n_59), .B1(n_733), .B2(n_734), .Y(n_732) );
CKINVDCx20_ASAP7_75t_R g734 ( .A(n_55), .Y(n_734) );
CKINVDCx20_ASAP7_75t_R g719 ( .A(n_56), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g231 ( .A(n_57), .Y(n_231) );
CKINVDCx14_ASAP7_75t_R g466 ( .A(n_58), .Y(n_466) );
CKINVDCx20_ASAP7_75t_R g733 ( .A(n_59), .Y(n_733) );
INVx1_ASAP7_75t_L g145 ( .A(n_60), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_61), .B(n_164), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_62), .B(n_204), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_63), .A2(n_198), .B(n_200), .C(n_202), .Y(n_197) );
INVx1_ASAP7_75t_L g135 ( .A(n_64), .Y(n_135) );
INVx1_ASAP7_75t_SL g498 ( .A(n_65), .Y(n_498) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_66), .Y(n_727) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_67), .B(n_174), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_68), .B(n_204), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_69), .B(n_152), .Y(n_151) );
INVx1_ASAP7_75t_L g531 ( .A(n_70), .Y(n_531) );
CKINVDCx16_ASAP7_75t_R g261 ( .A(n_71), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_72), .B(n_171), .Y(n_225) );
A2O1A1Ixp33_ASAP7_75t_L g237 ( .A1(n_73), .A2(n_147), .B(n_177), .C(n_238), .Y(n_237) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_74), .Y(n_196) );
INVx1_ASAP7_75t_L g114 ( .A(n_75), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g464 ( .A1(n_76), .A2(n_164), .B(n_465), .Y(n_464) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_77), .Y(n_534) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_78), .A2(n_164), .B(n_475), .Y(n_474) );
AOI21xp5_ASAP7_75t_L g506 ( .A1(n_79), .A2(n_222), .B(n_507), .Y(n_506) );
INVx1_ASAP7_75t_L g476 ( .A(n_80), .Y(n_476) );
CKINVDCx16_ASAP7_75t_R g517 ( .A(n_81), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_82), .B(n_170), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g216 ( .A(n_83), .Y(n_216) );
AOI21xp5_ASAP7_75t_L g483 ( .A1(n_84), .A2(n_164), .B(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g479 ( .A(n_85), .Y(n_479) );
INVx2_ASAP7_75t_L g133 ( .A(n_86), .Y(n_133) );
INVx1_ASAP7_75t_L g455 ( .A(n_87), .Y(n_455) );
CKINVDCx20_ASAP7_75t_R g245 ( .A(n_88), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_89), .B(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g111 ( .A(n_90), .Y(n_111) );
OR2x2_ASAP7_75t_L g440 ( .A(n_90), .B(n_441), .Y(n_440) );
OR2x2_ASAP7_75t_L g737 ( .A(n_90), .B(n_724), .Y(n_737) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_91), .A2(n_147), .B(n_177), .C(n_530), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_92), .B(n_164), .Y(n_210) );
INVx1_ASAP7_75t_L g213 ( .A(n_93), .Y(n_213) );
INVxp67_ASAP7_75t_L g201 ( .A(n_94), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_95), .B(n_131), .Y(n_471) );
INVx2_ASAP7_75t_L g488 ( .A(n_96), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_97), .B(n_114), .Y(n_113) );
INVx1_ASAP7_75t_L g138 ( .A(n_98), .Y(n_138) );
INVx1_ASAP7_75t_L g239 ( .A(n_99), .Y(n_239) );
AND2x2_ASAP7_75t_L g180 ( .A(n_100), .B(n_179), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g102 ( .A(n_103), .Y(n_102) );
CKINVDCx16_ASAP7_75t_R g103 ( .A(n_104), .Y(n_103) );
INVx2_ASAP7_75t_L g746 ( .A(n_104), .Y(n_746) );
AND2x2_ASAP7_75t_L g104 ( .A(n_105), .B(n_108), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
CKINVDCx14_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
NAND3xp33_ASAP7_75t_SL g109 ( .A(n_110), .B(n_111), .C(n_112), .Y(n_109) );
AND2x2_ASAP7_75t_L g441 ( .A(n_110), .B(n_442), .Y(n_441) );
OR2x2_ASAP7_75t_L g711 ( .A(n_111), .B(n_441), .Y(n_711) );
NOR2x2_ASAP7_75t_L g723 ( .A(n_111), .B(n_724), .Y(n_723) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
AO221x1_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_725), .B1(n_728), .B2(n_738), .C(n_740), .Y(n_115) );
OAI222xp33_ASAP7_75t_SL g116 ( .A1(n_117), .A2(n_120), .B1(n_712), .B2(n_713), .C1(n_719), .C2(n_720), .Y(n_116) );
INVx1_ASAP7_75t_L g712 ( .A(n_117), .Y(n_712) );
INVxp67_ASAP7_75t_L g120 ( .A(n_121), .Y(n_120) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_122), .A2(n_438), .B1(n_443), .B2(n_709), .Y(n_121) );
INVx2_ASAP7_75t_L g716 ( .A(n_122), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g730 ( .A1(n_122), .A2(n_716), .B1(n_731), .B2(n_732), .Y(n_730) );
OR3x1_ASAP7_75t_L g122 ( .A(n_123), .B(n_336), .C(n_401), .Y(n_122) );
NAND4xp25_ASAP7_75t_SL g123 ( .A(n_124), .B(n_277), .C(n_303), .D(n_326), .Y(n_123) );
AOI221xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_205), .B1(n_246), .B2(n_253), .C(n_269), .Y(n_124) );
CKINVDCx14_ASAP7_75t_R g125 ( .A(n_126), .Y(n_125) );
OAI22xp5_ASAP7_75t_L g424 ( .A1(n_126), .A2(n_270), .B1(n_294), .B2(n_425), .Y(n_424) );
OR2x2_ASAP7_75t_L g126 ( .A(n_127), .B(n_181), .Y(n_126) );
INVx1_ASAP7_75t_SL g330 ( .A(n_127), .Y(n_330) );
OR2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_161), .Y(n_127) );
OR2x2_ASAP7_75t_L g251 ( .A(n_128), .B(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g272 ( .A(n_128), .B(n_182), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_128), .B(n_192), .Y(n_285) );
AND2x2_ASAP7_75t_L g302 ( .A(n_128), .B(n_161), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_128), .B(n_249), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_128), .B(n_301), .Y(n_413) );
NOR2xp33_ASAP7_75t_L g423 ( .A(n_128), .B(n_181), .Y(n_423) );
AOI211xp5_ASAP7_75t_SL g434 ( .A1(n_128), .A2(n_340), .B(n_435), .C(n_436), .Y(n_434) );
INVx5_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
NAND2xp5_ASAP7_75t_SL g306 ( .A(n_129), .B(n_182), .Y(n_306) );
AND2x2_ASAP7_75t_L g309 ( .A(n_129), .B(n_183), .Y(n_309) );
OR2x2_ASAP7_75t_L g354 ( .A(n_129), .B(n_182), .Y(n_354) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_129), .B(n_192), .Y(n_363) );
AO21x2_ASAP7_75t_L g129 ( .A1(n_130), .A2(n_137), .B(n_158), .Y(n_129) );
INVx3_ASAP7_75t_L g204 ( .A(n_130), .Y(n_204) );
NOR2xp33_ASAP7_75t_L g215 ( .A(n_130), .B(n_216), .Y(n_215) );
AO21x2_ASAP7_75t_L g235 ( .A1(n_130), .A2(n_236), .B(n_244), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_130), .B(n_245), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g458 ( .A(n_130), .B(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_130), .B(n_523), .Y(n_522) );
AO21x2_ASAP7_75t_L g526 ( .A1(n_130), .A2(n_527), .B(n_533), .Y(n_526) );
INVx4_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
AOI21xp5_ASAP7_75t_L g184 ( .A1(n_131), .A2(n_185), .B(n_186), .Y(n_184) );
HB1xp67_ASAP7_75t_L g193 ( .A(n_131), .Y(n_193) );
BUFx6f_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_134), .Y(n_132) );
AND2x2_ASAP7_75t_SL g179 ( .A(n_133), .B(n_134), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g134 ( .A(n_135), .B(n_136), .Y(n_134) );
OAI21xp5_ASAP7_75t_L g137 ( .A1(n_138), .A2(n_139), .B(n_146), .Y(n_137) );
OAI21xp5_ASAP7_75t_L g451 ( .A1(n_139), .A2(n_452), .B(n_453), .Y(n_451) );
O2A1O1Ixp33_ASAP7_75t_L g516 ( .A1(n_139), .A2(n_179), .B(n_517), .C(n_518), .Y(n_516) );
OAI21xp5_ASAP7_75t_L g527 ( .A1(n_139), .A2(n_528), .B(n_529), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g139 ( .A(n_140), .B(n_144), .Y(n_139) );
AND2x4_ASAP7_75t_L g164 ( .A(n_140), .B(n_144), .Y(n_164) );
AND2x2_ASAP7_75t_L g140 ( .A(n_141), .B(n_143), .Y(n_140) );
INVx1_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx1_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
INVx2_ASAP7_75t_L g148 ( .A(n_142), .Y(n_148) );
INVx1_ASAP7_75t_L g157 ( .A(n_142), .Y(n_157) );
INVx1_ASAP7_75t_L g149 ( .A(n_143), .Y(n_149) );
INVx3_ASAP7_75t_L g152 ( .A(n_143), .Y(n_152) );
BUFx6f_ASAP7_75t_L g154 ( .A(n_143), .Y(n_154) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_143), .Y(n_172) );
INVx1_ASAP7_75t_L g189 ( .A(n_143), .Y(n_189) );
INVx4_ASAP7_75t_SL g178 ( .A(n_144), .Y(n_178) );
BUFx3_ASAP7_75t_L g191 ( .A(n_144), .Y(n_191) );
INVx5_ASAP7_75t_L g167 ( .A(n_147), .Y(n_167) );
AND2x6_ASAP7_75t_L g147 ( .A(n_148), .B(n_149), .Y(n_147) );
BUFx3_ASAP7_75t_L g176 ( .A(n_148), .Y(n_176) );
BUFx6f_ASAP7_75t_L g242 ( .A(n_148), .Y(n_242) );
AOI21xp5_ASAP7_75t_L g150 ( .A1(n_151), .A2(n_153), .B(n_155), .Y(n_150) );
INVx5_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g469 ( .A(n_152), .B(n_470), .Y(n_469) );
INVx4_ASAP7_75t_L g266 ( .A(n_154), .Y(n_266) );
INVx2_ASAP7_75t_L g468 ( .A(n_154), .Y(n_468) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_155), .A2(n_188), .B(n_190), .Y(n_187) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
NOR2xp33_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
INVx2_ASAP7_75t_L g505 ( .A(n_160), .Y(n_505) );
INVx5_ASAP7_75t_SL g252 ( .A(n_161), .Y(n_252) );
AND2x2_ASAP7_75t_L g271 ( .A(n_161), .B(n_272), .Y(n_271) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_161), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g357 ( .A(n_161), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g389 ( .A(n_161), .B(n_192), .Y(n_389) );
OR2x2_ASAP7_75t_L g395 ( .A(n_161), .B(n_285), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_161), .B(n_345), .Y(n_404) );
OR2x6_ASAP7_75t_L g161 ( .A(n_162), .B(n_180), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g162 ( .A1(n_163), .A2(n_165), .B(n_179), .Y(n_162) );
BUFx2_ASAP7_75t_L g222 ( .A(n_164), .Y(n_222) );
INVx2_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
O2A1O1Ixp33_ASAP7_75t_L g195 ( .A1(n_167), .A2(n_178), .B(n_196), .C(n_197), .Y(n_195) );
O2A1O1Ixp33_ASAP7_75t_SL g260 ( .A1(n_167), .A2(n_178), .B(n_261), .C(n_262), .Y(n_260) );
O2A1O1Ixp33_ASAP7_75t_SL g465 ( .A1(n_167), .A2(n_178), .B(n_466), .C(n_467), .Y(n_465) );
O2A1O1Ixp33_ASAP7_75t_SL g475 ( .A1(n_167), .A2(n_178), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g484 ( .A1(n_167), .A2(n_178), .B(n_485), .C(n_486), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g494 ( .A1(n_167), .A2(n_178), .B(n_495), .C(n_496), .Y(n_494) );
O2A1O1Ixp33_ASAP7_75t_SL g507 ( .A1(n_167), .A2(n_178), .B(n_508), .C(n_509), .Y(n_507) );
O2A1O1Ixp33_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_173), .C(n_175), .Y(n_168) );
O2A1O1Ixp33_ASAP7_75t_L g212 ( .A1(n_170), .A2(n_175), .B(n_213), .C(n_214), .Y(n_212) );
O2A1O1Ixp5_ASAP7_75t_L g454 ( .A1(n_170), .A2(n_455), .B(n_456), .C(n_457), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_170), .A2(n_457), .B(n_531), .C(n_532), .Y(n_530) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx4_ASAP7_75t_L g199 ( .A(n_172), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_174), .B(n_201), .Y(n_200) );
INVx2_ASAP7_75t_L g263 ( .A(n_174), .Y(n_263) );
OAI22xp33_ASAP7_75t_L g510 ( .A1(n_174), .A2(n_199), .B1(n_511), .B2(n_512), .Y(n_510) );
O2A1O1Ixp33_ASAP7_75t_L g519 ( .A1(n_174), .A2(n_227), .B(n_520), .C(n_521), .Y(n_519) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_176), .Y(n_175) );
INVx2_ASAP7_75t_L g267 ( .A(n_176), .Y(n_267) );
INVx1_ASAP7_75t_L g480 ( .A(n_176), .Y(n_480) );
INVx1_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_179), .A2(n_210), .B(n_211), .Y(n_209) );
INVx2_ASAP7_75t_L g229 ( .A(n_179), .Y(n_229) );
INVx1_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
OA21x2_ASAP7_75t_L g463 ( .A1(n_179), .A2(n_464), .B(n_471), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g181 ( .A(n_182), .B(n_192), .Y(n_181) );
AND2x2_ASAP7_75t_L g286 ( .A(n_182), .B(n_252), .Y(n_286) );
INVx1_ASAP7_75t_SL g299 ( .A(n_182), .Y(n_299) );
OR2x2_ASAP7_75t_L g334 ( .A(n_182), .B(n_335), .Y(n_334) );
OR2x2_ASAP7_75t_L g340 ( .A(n_182), .B(n_192), .Y(n_340) );
AND2x2_ASAP7_75t_L g398 ( .A(n_182), .B(n_249), .Y(n_398) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_183), .B(n_252), .Y(n_325) );
INVx3_ASAP7_75t_L g249 ( .A(n_192), .Y(n_249) );
OR2x2_ASAP7_75t_L g291 ( .A(n_192), .B(n_252), .Y(n_291) );
AND2x2_ASAP7_75t_L g301 ( .A(n_192), .B(n_299), .Y(n_301) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_192), .Y(n_349) );
AND2x2_ASAP7_75t_L g358 ( .A(n_192), .B(n_272), .Y(n_358) );
OA21x2_ASAP7_75t_L g192 ( .A1(n_193), .A2(n_194), .B(n_203), .Y(n_192) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_193), .A2(n_474), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g482 ( .A1(n_193), .A2(n_483), .B(n_489), .Y(n_482) );
OA21x2_ASAP7_75t_L g492 ( .A1(n_193), .A2(n_493), .B(n_500), .Y(n_492) );
O2A1O1Ixp33_ASAP7_75t_L g238 ( .A1(n_198), .A2(n_239), .B(n_240), .C(n_241), .Y(n_238) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_199), .B(n_479), .Y(n_478) );
NOR2xp33_ASAP7_75t_L g487 ( .A(n_199), .B(n_488), .Y(n_487) );
INVx2_ASAP7_75t_L g227 ( .A(n_202), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g509 ( .A(n_202), .B(n_510), .Y(n_509) );
OA21x2_ASAP7_75t_L g258 ( .A1(n_204), .A2(n_259), .B(n_268), .Y(n_258) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_205), .A2(n_375), .B1(n_377), .B2(n_379), .C(n_382), .Y(n_374) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
OR2x2_ASAP7_75t_L g206 ( .A(n_207), .B(n_217), .Y(n_206) );
AND2x2_ASAP7_75t_L g348 ( .A(n_207), .B(n_329), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_207), .B(n_407), .Y(n_411) );
OR2x2_ASAP7_75t_L g432 ( .A(n_207), .B(n_433), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g436 ( .A(n_207), .B(n_437), .Y(n_436) );
BUFx2_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
INVx5_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
AND2x2_ASAP7_75t_L g356 ( .A(n_208), .B(n_219), .Y(n_356) );
AND2x2_ASAP7_75t_L g417 ( .A(n_208), .B(n_296), .Y(n_417) );
AND2x2_ASAP7_75t_L g430 ( .A(n_208), .B(n_249), .Y(n_430) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_215), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_218), .B(n_233), .Y(n_217) );
AND2x4_ASAP7_75t_L g256 ( .A(n_218), .B(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g275 ( .A(n_218), .B(n_276), .Y(n_275) );
INVx2_ASAP7_75t_L g282 ( .A(n_218), .Y(n_282) );
AND2x2_ASAP7_75t_L g351 ( .A(n_218), .B(n_329), .Y(n_351) );
AND2x2_ASAP7_75t_L g361 ( .A(n_218), .B(n_279), .Y(n_361) );
HB1xp67_ASAP7_75t_L g369 ( .A(n_218), .Y(n_369) );
AND2x2_ASAP7_75t_L g381 ( .A(n_218), .B(n_258), .Y(n_381) );
NOR2xp33_ASAP7_75t_L g385 ( .A(n_218), .B(n_313), .Y(n_385) );
AND2x2_ASAP7_75t_L g422 ( .A(n_218), .B(n_417), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_218), .B(n_296), .Y(n_433) );
OR2x2_ASAP7_75t_L g435 ( .A(n_218), .B(n_371), .Y(n_435) );
INVx5_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
AND2x2_ASAP7_75t_L g321 ( .A(n_219), .B(n_322), .Y(n_321) );
AND2x2_ASAP7_75t_L g331 ( .A(n_219), .B(n_276), .Y(n_331) );
AND2x2_ASAP7_75t_L g343 ( .A(n_219), .B(n_258), .Y(n_343) );
HB1xp67_ASAP7_75t_L g373 ( .A(n_219), .Y(n_373) );
AND2x4_ASAP7_75t_L g407 ( .A(n_219), .B(n_257), .Y(n_407) );
OR2x6_ASAP7_75t_L g219 ( .A(n_220), .B(n_230), .Y(n_219) );
AOI21xp5_ASAP7_75t_SL g220 ( .A1(n_221), .A2(n_223), .B(n_228), .Y(n_220) );
AOI21xp5_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_226), .B(n_227), .Y(n_224) );
INVx1_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g533 ( .A(n_229), .B(n_534), .Y(n_533) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_231), .B(n_232), .Y(n_230) );
AO21x2_ASAP7_75t_L g450 ( .A1(n_232), .A2(n_451), .B(n_458), .Y(n_450) );
BUFx2_ASAP7_75t_L g255 ( .A(n_233), .Y(n_255) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
INVx2_ASAP7_75t_L g296 ( .A(n_234), .Y(n_296) );
AND2x2_ASAP7_75t_L g329 ( .A(n_234), .B(n_258), .Y(n_329) );
INVx2_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AND2x2_ASAP7_75t_L g276 ( .A(n_235), .B(n_258), .Y(n_276) );
BUFx2_ASAP7_75t_L g322 ( .A(n_235), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
HB1xp67_ASAP7_75t_L g241 ( .A(n_242), .Y(n_241) );
INVx3_ASAP7_75t_L g499 ( .A(n_242), .Y(n_499) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_248), .B(n_330), .Y(n_409) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_249), .B(n_272), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_249), .B(n_252), .Y(n_311) );
AND2x2_ASAP7_75t_L g366 ( .A(n_249), .B(n_302), .Y(n_366) );
AOI221xp5_ASAP7_75t_SL g303 ( .A1(n_250), .A2(n_304), .B1(n_312), .B2(n_314), .C(n_318), .Y(n_303) );
INVx2_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g298 ( .A(n_251), .B(n_299), .Y(n_298) );
OR2x2_ASAP7_75t_L g339 ( .A(n_251), .B(n_340), .Y(n_339) );
OAI321xp33_ASAP7_75t_L g346 ( .A1(n_251), .A2(n_305), .A3(n_347), .B1(n_349), .B2(n_350), .C(n_352), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_252), .B(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_255), .B(n_256), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_255), .B(n_407), .Y(n_425) );
AND2x2_ASAP7_75t_L g312 ( .A(n_256), .B(n_313), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_256), .B(n_316), .Y(n_315) );
HB1xp67_ASAP7_75t_L g288 ( .A(n_257), .Y(n_288) );
AND2x2_ASAP7_75t_L g295 ( .A(n_257), .B(n_296), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g400 ( .A(n_257), .B(n_370), .Y(n_400) );
INVx1_ASAP7_75t_L g437 ( .A(n_257), .Y(n_437) );
INVx2_ASAP7_75t_L g257 ( .A(n_258), .Y(n_257) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
NOR2xp33_ASAP7_75t_L g497 ( .A(n_266), .B(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g457 ( .A(n_267), .Y(n_457) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_270), .A2(n_273), .B(n_274), .Y(n_269) );
INVx1_ASAP7_75t_SL g270 ( .A(n_271), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g429 ( .A1(n_271), .A2(n_381), .B(n_430), .C(n_431), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_272), .B(n_290), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_272), .B(n_310), .Y(n_376) );
INVx1_ASAP7_75t_SL g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g319 ( .A(n_276), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_276), .B(n_279), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g342 ( .A(n_276), .B(n_343), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_276), .B(n_361), .Y(n_360) );
AOI22xp33_ASAP7_75t_L g277 ( .A1(n_278), .A2(n_280), .B1(n_292), .B2(n_297), .Y(n_277) );
HB1xp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
OR2x2_ASAP7_75t_L g293 ( .A(n_279), .B(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g316 ( .A(n_279), .B(n_317), .Y(n_316) );
AND2x2_ASAP7_75t_L g328 ( .A(n_279), .B(n_329), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_279), .B(n_322), .Y(n_364) );
OR2x2_ASAP7_75t_L g371 ( .A(n_279), .B(n_296), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_279), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g421 ( .A(n_279), .B(n_407), .Y(n_421) );
OAI22xp33_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B1(n_287), .B2(n_289), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
AND2x2_ASAP7_75t_L g327 ( .A(n_282), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
OAI22xp33_ASAP7_75t_L g367 ( .A1(n_285), .A2(n_300), .B1(n_368), .B2(n_372), .Y(n_367) );
INVx1_ASAP7_75t_L g415 ( .A(n_286), .Y(n_415) );
INVx1_ASAP7_75t_L g287 ( .A(n_288), .Y(n_287) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_290), .A2(n_327), .B1(n_330), .B2(n_331), .C(n_332), .Y(n_326) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
OR2x2_ASAP7_75t_L g305 ( .A(n_291), .B(n_306), .Y(n_305) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_295), .B(n_361), .Y(n_393) );
HB1xp67_ASAP7_75t_L g313 ( .A(n_296), .Y(n_313) );
INVx1_ASAP7_75t_L g317 ( .A(n_296), .Y(n_317) );
NAND2xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_300), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g335 ( .A(n_302), .Y(n_335) );
AND2x2_ASAP7_75t_L g344 ( .A(n_302), .B(n_345), .Y(n_344) );
NAND2xp33_ASAP7_75t_L g304 ( .A(n_305), .B(n_307), .Y(n_304) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x4_ASAP7_75t_L g308 ( .A(n_309), .B(n_310), .Y(n_308) );
AND2x2_ASAP7_75t_L g388 ( .A(n_309), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
AOI221xp5_ASAP7_75t_L g337 ( .A1(n_312), .A2(n_338), .B1(n_341), .B2(n_344), .C(n_346), .Y(n_337) );
INVx1_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_316), .B(n_373), .Y(n_372) );
AOI21xp33_ASAP7_75t_SL g318 ( .A1(n_319), .A2(n_320), .B(n_323), .Y(n_318) );
INVx2_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
CKINVDCx16_ASAP7_75t_R g420 ( .A(n_323), .Y(n_420) );
OR2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
OR2x2_ASAP7_75t_L g362 ( .A(n_325), .B(n_363), .Y(n_362) );
INVx1_ASAP7_75t_SL g383 ( .A(n_328), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_328), .B(n_388), .Y(n_428) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_331), .B(n_353), .Y(n_352) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_333), .B(n_334), .Y(n_332) );
NAND4xp25_ASAP7_75t_L g336 ( .A(n_337), .B(n_355), .C(n_374), .D(n_387), .Y(n_336) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
INVx1_ASAP7_75t_SL g345 ( .A(n_340), .Y(n_345) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
OR2x2_ASAP7_75t_L g378 ( .A(n_349), .B(n_354), .Y(n_378) );
INVxp67_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
AOI211xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_357), .B(n_359), .C(n_367), .Y(n_355) );
AOI211xp5_ASAP7_75t_L g426 ( .A1(n_357), .A2(n_399), .B(n_427), .C(n_434), .Y(n_426) );
INVx1_ASAP7_75t_SL g386 ( .A(n_358), .Y(n_386) );
OAI22xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_362), .B1(n_364), .B2(n_365), .Y(n_359) );
INVx1_ASAP7_75t_L g390 ( .A(n_364), .Y(n_390) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_370), .B(n_407), .Y(n_406) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_370), .B(n_381), .Y(n_414) );
INVx2_ASAP7_75t_SL g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_SL g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g391 ( .A(n_381), .Y(n_391) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_383), .A2(n_384), .B(n_386), .Y(n_382) );
INVxp33_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
AOI322xp5_ASAP7_75t_L g387 ( .A1(n_388), .A2(n_390), .A3(n_391), .B1(n_392), .B2(n_394), .C1(n_396), .C2(n_399), .Y(n_387) );
INVxp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
NAND3xp33_ASAP7_75t_SL g401 ( .A(n_402), .B(n_419), .C(n_426), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_403), .A2(n_405), .B1(n_408), .B2(n_410), .C(n_412), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVx1_ASAP7_75t_SL g418 ( .A(n_407), .Y(n_418) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
INVxp67_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
OAI22xp33_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g419 ( .A1(n_420), .A2(n_421), .B1(n_422), .B2(n_423), .C(n_424), .Y(n_419) );
NAND2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_429), .Y(n_427) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g715 ( .A(n_439), .Y(n_715) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g724 ( .A(n_441), .Y(n_724) );
INVx2_ASAP7_75t_L g717 ( .A(n_443), .Y(n_717) );
OR2x2_ASAP7_75t_SL g443 ( .A(n_444), .B(n_664), .Y(n_443) );
NAND5xp2_ASAP7_75t_L g444 ( .A(n_445), .B(n_576), .C(n_614), .D(n_635), .E(n_652), .Y(n_444) );
NOR3xp33_ASAP7_75t_L g445 ( .A(n_446), .B(n_548), .C(n_569), .Y(n_445) );
OAI221xp5_ASAP7_75t_SL g446 ( .A1(n_447), .A2(n_490), .B1(n_514), .B2(n_535), .C(n_539), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_448), .B(n_460), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_449), .B(n_537), .Y(n_556) );
OR2x2_ASAP7_75t_L g583 ( .A(n_449), .B(n_473), .Y(n_583) );
AND2x2_ASAP7_75t_L g597 ( .A(n_449), .B(n_473), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g611 ( .A(n_449), .B(n_463), .Y(n_611) );
AND2x2_ASAP7_75t_L g649 ( .A(n_449), .B(n_613), .Y(n_649) );
AND2x2_ASAP7_75t_L g678 ( .A(n_449), .B(n_588), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_449), .B(n_560), .Y(n_695) );
INVx4_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
AND2x2_ASAP7_75t_L g575 ( .A(n_450), .B(n_472), .Y(n_575) );
BUFx3_ASAP7_75t_L g600 ( .A(n_450), .Y(n_600) );
AND2x2_ASAP7_75t_L g629 ( .A(n_450), .B(n_473), .Y(n_629) );
AND3x2_ASAP7_75t_L g642 ( .A(n_450), .B(n_643), .C(n_644), .Y(n_642) );
INVx1_ASAP7_75t_L g565 ( .A(n_460), .Y(n_565) );
AND2x2_ASAP7_75t_L g460 ( .A(n_461), .B(n_472), .Y(n_460) );
AOI32xp33_ASAP7_75t_L g620 ( .A1(n_461), .A2(n_572), .A3(n_621), .B1(n_624), .B2(n_625), .Y(n_620) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g547 ( .A(n_462), .B(n_472), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g618 ( .A(n_462), .B(n_575), .Y(n_618) );
AND2x2_ASAP7_75t_L g625 ( .A(n_462), .B(n_597), .Y(n_625) );
OR2x2_ASAP7_75t_L g631 ( .A(n_462), .B(n_632), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_462), .B(n_586), .Y(n_656) );
OR2x2_ASAP7_75t_L g674 ( .A(n_462), .B(n_502), .Y(n_674) );
BUFx3_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
AND2x2_ASAP7_75t_L g538 ( .A(n_463), .B(n_482), .Y(n_538) );
INVx2_ASAP7_75t_L g560 ( .A(n_463), .Y(n_560) );
OR2x2_ASAP7_75t_L g582 ( .A(n_463), .B(n_482), .Y(n_582) );
AND2x2_ASAP7_75t_L g587 ( .A(n_463), .B(n_588), .Y(n_587) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_463), .B(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g643 ( .A(n_463), .B(n_537), .Y(n_643) );
INVx1_ASAP7_75t_SL g694 ( .A(n_472), .Y(n_694) );
AND2x2_ASAP7_75t_L g472 ( .A(n_473), .B(n_482), .Y(n_472) );
INVx1_ASAP7_75t_SL g537 ( .A(n_473), .Y(n_537) );
HB1xp67_ASAP7_75t_L g586 ( .A(n_473), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_473), .B(n_623), .Y(n_622) );
NAND3xp33_ASAP7_75t_L g689 ( .A(n_473), .B(n_560), .C(n_678), .Y(n_689) );
INVx2_ASAP7_75t_L g588 ( .A(n_482), .Y(n_588) );
HB1xp67_ASAP7_75t_L g602 ( .A(n_482), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_501), .Y(n_490) );
INVx1_ASAP7_75t_L g624 ( .A(n_491), .Y(n_624) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
AND2x2_ASAP7_75t_L g542 ( .A(n_492), .B(n_525), .Y(n_542) );
INVx2_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
AND2x2_ASAP7_75t_L g564 ( .A(n_492), .B(n_526), .Y(n_564) );
AND2x2_ASAP7_75t_L g579 ( .A(n_492), .B(n_515), .Y(n_579) );
AND2x2_ASAP7_75t_L g591 ( .A(n_492), .B(n_563), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_501), .B(n_607), .Y(n_606) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_501), .B(n_564), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_501), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_501), .B(n_558), .Y(n_686) );
BUFx3_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
OR2x2_ASAP7_75t_L g524 ( .A(n_502), .B(n_525), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_502), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g568 ( .A(n_502), .B(n_515), .Y(n_568) );
AND2x2_ASAP7_75t_L g594 ( .A(n_502), .B(n_525), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_502), .B(n_634), .Y(n_633) );
OA21x2_ASAP7_75t_L g502 ( .A1(n_503), .A2(n_506), .B(n_513), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_504), .Y(n_503) );
AO21x2_ASAP7_75t_L g552 ( .A1(n_504), .A2(n_553), .B(n_554), .Y(n_552) );
INVx1_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
INVx1_ASAP7_75t_L g553 ( .A(n_506), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_513), .Y(n_554) );
OR2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_515), .B(n_545), .Y(n_544) );
AND2x4_ASAP7_75t_L g558 ( .A(n_515), .B(n_559), .Y(n_558) );
INVx3_ASAP7_75t_SL g563 ( .A(n_515), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_515), .B(n_550), .Y(n_616) );
OR2x2_ASAP7_75t_L g626 ( .A(n_515), .B(n_552), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_515), .B(n_594), .Y(n_654) );
OR2x2_ASAP7_75t_L g684 ( .A(n_515), .B(n_525), .Y(n_684) );
AND2x2_ASAP7_75t_L g688 ( .A(n_515), .B(n_526), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g701 ( .A(n_515), .B(n_564), .Y(n_701) );
AND2x2_ASAP7_75t_L g708 ( .A(n_515), .B(n_590), .Y(n_708) );
OR2x6_ASAP7_75t_L g515 ( .A(n_516), .B(n_522), .Y(n_515) );
INVx1_ASAP7_75t_SL g651 ( .A(n_524), .Y(n_651) );
AND2x2_ASAP7_75t_L g590 ( .A(n_525), .B(n_552), .Y(n_590) );
AND2x2_ASAP7_75t_L g604 ( .A(n_525), .B(n_559), .Y(n_604) );
AND2x2_ASAP7_75t_L g607 ( .A(n_525), .B(n_563), .Y(n_607) );
INVx1_ASAP7_75t_L g634 ( .A(n_525), .Y(n_634) );
INVx2_ASAP7_75t_SL g525 ( .A(n_526), .Y(n_525) );
BUFx2_ASAP7_75t_L g546 ( .A(n_526), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_536), .B(n_538), .Y(n_535) );
A2O1A1Ixp33_ASAP7_75t_L g705 ( .A1(n_536), .A2(n_582), .B(n_706), .C(n_707), .Y(n_705) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
AND2x2_ASAP7_75t_L g612 ( .A(n_537), .B(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_538), .B(n_555), .Y(n_570) );
AND2x2_ASAP7_75t_L g596 ( .A(n_538), .B(n_597), .Y(n_596) );
OAI21xp5_ASAP7_75t_SL g539 ( .A1(n_540), .A2(n_543), .B(n_547), .Y(n_539) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
NOR2xp33_ASAP7_75t_L g640 ( .A(n_541), .B(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g567 ( .A(n_542), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_542), .B(n_563), .Y(n_608) );
AND2x2_ASAP7_75t_L g699 ( .A(n_542), .B(n_550), .Y(n_699) );
INVxp67_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g572 ( .A(n_546), .B(n_559), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_546), .B(n_557), .Y(n_573) );
OAI322xp33_ASAP7_75t_L g548 ( .A1(n_549), .A2(n_556), .A3(n_557), .B1(n_560), .B2(n_561), .C1(n_565), .C2(n_566), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_555), .Y(n_549) );
AND2x2_ASAP7_75t_L g660 ( .A(n_550), .B(n_572), .Y(n_660) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_550), .B(n_624), .Y(n_706) );
INVx2_ASAP7_75t_L g550 ( .A(n_551), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g603 ( .A(n_552), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
OR2x2_ASAP7_75t_L g669 ( .A(n_556), .B(n_582), .Y(n_669) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_557), .B(n_651), .Y(n_650) );
INVx3_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_558), .B(n_590), .Y(n_647) );
AND2x2_ASAP7_75t_L g593 ( .A(n_559), .B(n_563), .Y(n_593) );
AND2x2_ASAP7_75t_L g601 ( .A(n_560), .B(n_602), .Y(n_601) );
A2O1A1Ixp33_ASAP7_75t_L g698 ( .A1(n_560), .A2(n_639), .B(n_699), .C(n_700), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g671 ( .A1(n_561), .A2(n_574), .B(n_672), .Y(n_671) );
INVx1_ASAP7_75t_SL g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_564), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_563), .B(n_590), .Y(n_630) );
AND2x2_ASAP7_75t_L g636 ( .A(n_563), .B(n_604), .Y(n_636) );
AND2x2_ASAP7_75t_L g670 ( .A(n_563), .B(n_572), .Y(n_670) );
NOR2xp33_ASAP7_75t_L g578 ( .A(n_564), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_SL g680 ( .A(n_564), .Y(n_680) );
INVx1_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
AOI22xp5_ASAP7_75t_L g595 ( .A1(n_568), .A2(n_596), .B1(n_598), .B2(n_603), .Y(n_595) );
OAI22xp5_ASAP7_75t_SL g569 ( .A1(n_570), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_569) );
OAI22xp33_ASAP7_75t_L g605 ( .A1(n_570), .A2(n_606), .B1(n_608), .B2(n_609), .Y(n_605) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_SL g574 ( .A(n_575), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g676 ( .A1(n_575), .A2(n_677), .B1(n_679), .B2(n_681), .C(n_685), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_580), .B(n_584), .C(n_605), .Y(n_576) );
INVxp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx1_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
OR2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
OR2x2_ASAP7_75t_L g646 ( .A(n_582), .B(n_599), .Y(n_646) );
INVx1_ASAP7_75t_L g697 ( .A(n_582), .Y(n_697) );
OAI221xp5_ASAP7_75t_L g584 ( .A1(n_583), .A2(n_585), .B1(n_589), .B2(n_592), .C(n_595), .Y(n_584) );
INVx2_ASAP7_75t_SL g639 ( .A(n_583), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_586), .B(n_587), .Y(n_585) );
INVx1_ASAP7_75t_L g704 ( .A(n_586), .Y(n_704) );
AND2x2_ASAP7_75t_L g628 ( .A(n_587), .B(n_629), .Y(n_628) );
INVx2_ASAP7_75t_L g613 ( .A(n_588), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_590), .B(n_591), .Y(n_589) );
INVx1_ASAP7_75t_L g675 ( .A(n_591), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_593), .B(n_594), .Y(n_592) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_601), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g700 ( .A(n_599), .B(n_701), .Y(n_700) );
CKINVDCx16_ASAP7_75t_R g599 ( .A(n_600), .Y(n_599) );
INVxp67_ASAP7_75t_L g644 ( .A(n_602), .Y(n_644) );
O2A1O1Ixp33_ASAP7_75t_L g614 ( .A1(n_603), .A2(n_615), .B(n_617), .C(n_619), .Y(n_614) );
INVx1_ASAP7_75t_L g692 ( .A(n_606), .Y(n_692) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
NOR2xp33_ASAP7_75t_L g667 ( .A(n_610), .B(n_668), .Y(n_667) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
INVx2_ASAP7_75t_L g623 ( .A(n_613), .Y(n_623) );
INVx1_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
OAI222xp33_ASAP7_75t_L g619 ( .A1(n_620), .A2(n_626), .B1(n_627), .B2(n_630), .C1(n_631), .C2(n_633), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_SL g659 ( .A(n_623), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g679 ( .A(n_626), .B(n_680), .Y(n_679) );
NAND2xp33_ASAP7_75t_SL g657 ( .A(n_627), .B(n_658), .Y(n_657) );
INVx1_ASAP7_75t_SL g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_SL g632 ( .A(n_629), .Y(n_632) );
AND2x2_ASAP7_75t_L g696 ( .A(n_629), .B(n_697), .Y(n_696) );
OR2x2_ASAP7_75t_L g662 ( .A(n_632), .B(n_659), .Y(n_662) );
INVx1_ASAP7_75t_L g691 ( .A(n_633), .Y(n_691) );
AOI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .B(n_640), .C(n_645), .Y(n_635) );
INVx1_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_639), .B(n_659), .Y(n_658) );
INVx2_ASAP7_75t_SL g641 ( .A(n_642), .Y(n_641) );
AOI322xp5_ASAP7_75t_L g690 ( .A1(n_642), .A2(n_670), .A3(n_675), .B1(n_691), .B2(n_692), .C1(n_693), .C2(n_696), .Y(n_690) );
AND2x2_ASAP7_75t_L g677 ( .A(n_643), .B(n_678), .Y(n_677) );
OAI22xp33_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_647), .B1(n_648), .B2(n_650), .Y(n_645) );
INVxp33_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_655), .B1(n_657), .B2(n_660), .C(n_661), .Y(n_652) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
NOR2xp33_ASAP7_75t_L g661 ( .A(n_662), .B(n_663), .Y(n_661) );
NAND5xp2_ASAP7_75t_L g664 ( .A(n_665), .B(n_676), .C(n_690), .D(n_698), .E(n_702), .Y(n_664) );
AOI21xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_670), .B(n_671), .Y(n_665) );
INVxp67_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_L g668 ( .A(n_669), .Y(n_668) );
INVxp33_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
A2O1A1Ixp33_ASAP7_75t_L g702 ( .A1(n_678), .A2(n_703), .B(n_704), .C(n_705), .Y(n_702) );
AOI31xp33_ASAP7_75t_L g685 ( .A1(n_680), .A2(n_686), .A3(n_687), .B(n_689), .Y(n_685) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g693 ( .A(n_694), .B(n_695), .Y(n_693) );
INVx1_ASAP7_75t_L g703 ( .A(n_701), .Y(n_703) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g718 ( .A(n_710), .Y(n_718) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVxp67_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI22x1_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B1(n_717), .B2(n_718), .Y(n_714) );
INVx1_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
BUFx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx2_ASAP7_75t_L g726 ( .A(n_727), .Y(n_726) );
INVx1_ASAP7_75t_L g739 ( .A(n_727), .Y(n_739) );
INVxp67_ASAP7_75t_L g728 ( .A(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_SL g729 ( .A(n_730), .B(n_735), .Y(n_729) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_SL g735 ( .A(n_736), .Y(n_735) );
INVx1_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
INVx1_ASAP7_75t_SL g743 ( .A(n_737), .Y(n_743) );
INVx1_ASAP7_75t_L g738 ( .A(n_739), .Y(n_738) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_741), .B(n_742), .Y(n_740) );
INVx1_ASAP7_75t_SL g742 ( .A(n_743), .Y(n_742) );
INVx1_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
endmodule