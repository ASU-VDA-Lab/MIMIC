module fake_jpeg_16965_n_82 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_82);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_82;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

INVx11_ASAP7_75t_SL g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_27),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx2_ASAP7_75t_SL g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_34),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_35),
.B(n_38),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_28),
.Y(n_36)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_1),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_43),
.B(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_2),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_41),
.B(n_32),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_49),
.B(n_51),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_3),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_33),
.Y(n_53)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_53),
.Y(n_63)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_54),
.B(n_57),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_33),
.C(n_31),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_55),
.B(n_12),
.C(n_13),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_46),
.B(n_3),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_56),
.B(n_59),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

OAI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_50),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_58),
.B(n_14),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_43),
.B(n_9),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_45),
.B(n_10),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_60),
.B(n_11),
.Y(n_62)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_64),
.B(n_66),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_65),
.A2(n_67),
.B1(n_70),
.B2(n_19),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_61),
.B(n_50),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_15),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_57),
.B(n_17),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g73 ( 
.A(n_69),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_73),
.Y(n_76)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_74),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g77 ( 
.A1(n_76),
.A2(n_71),
.B(n_63),
.Y(n_77)
);

FAx1_ASAP7_75t_SL g78 ( 
.A(n_77),
.B(n_73),
.CI(n_75),
.CON(n_78),
.SN(n_78)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_78),
.B(n_68),
.C(n_72),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_79),
.A2(n_78),
.B(n_75),
.Y(n_80)
);

AOI322xp5_ASAP7_75t_L g81 ( 
.A1(n_80),
.A2(n_20),
.A3(n_21),
.B1(n_22),
.B2(n_23),
.C1(n_24),
.C2(n_25),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_26),
.Y(n_82)
);


endmodule