module fake_jpeg_9903_n_278 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_175;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_96;

BUFx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx11_ASAP7_75t_SL g18 ( 
.A(n_0),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx16f_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx2_ASAP7_75t_L g30 ( 
.A(n_12),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_5),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_17),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_37),
.B(n_39),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_17),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_43),
.Y(n_58)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_44),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_43),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_45)
);

OAI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_45),
.A2(n_53),
.B1(n_57),
.B2(n_62),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_46)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_46),
.A2(n_52),
.B1(n_33),
.B2(n_32),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_22),
.B1(n_28),
.B2(n_19),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_47),
.A2(n_49),
.B1(n_55),
.B2(n_63),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_37),
.A2(n_26),
.B1(n_21),
.B2(n_31),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_39),
.A2(n_19),
.B1(n_31),
.B2(n_21),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_43),
.A2(n_39),
.B1(n_44),
.B2(n_41),
.Y(n_53)
);

AND2x2_ASAP7_75t_SL g54 ( 
.A(n_40),
.B(n_24),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_54),
.B(n_66),
.C(n_42),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_39),
.A2(n_26),
.B1(n_34),
.B2(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_40),
.B(n_30),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_54),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_34),
.B1(n_33),
.B2(n_32),
.Y(n_57)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_58),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_43),
.A2(n_33),
.B1(n_32),
.B2(n_23),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_40),
.A2(n_33),
.B1(n_32),
.B2(n_23),
.Y(n_63)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_24),
.C(n_17),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_53),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_67),
.B(n_71),
.Y(n_109)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_64),
.Y(n_68)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_68),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g118 ( 
.A(n_69),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g70 ( 
.A(n_49),
.B(n_38),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_70),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_51),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_36),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_72),
.B(n_73),
.Y(n_111)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_48),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_75),
.B(n_100),
.Y(n_107)
);

OAI22x1_ASAP7_75t_R g76 ( 
.A1(n_54),
.A2(n_42),
.B1(n_38),
.B2(n_41),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_76),
.B(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_36),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_77),
.B(n_78),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_61),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_79),
.Y(n_115)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVx1_ASAP7_75t_SL g125 ( 
.A(n_80),
.Y(n_125)
);

CKINVDCx6p67_ASAP7_75t_R g81 ( 
.A(n_59),
.Y(n_81)
);

INVx13_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_55),
.A2(n_44),
.B1(n_36),
.B2(n_41),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_82),
.A2(n_86),
.B1(n_96),
.B2(n_97),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_49),
.B(n_36),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_83),
.B(n_85),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_61),
.A2(n_38),
.B(n_35),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_84),
.B(n_101),
.Y(n_121)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_48),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g86 ( 
.A1(n_56),
.A2(n_44),
.B1(n_42),
.B2(n_23),
.Y(n_86)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_88),
.Y(n_106)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_64),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_89),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_52),
.B(n_30),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_55),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_92),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_41),
.Y(n_93)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_46),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_46),
.A2(n_42),
.B1(n_30),
.B2(n_27),
.Y(n_96)
);

OAI22x1_ASAP7_75t_L g97 ( 
.A1(n_45),
.A2(n_35),
.B1(n_30),
.B2(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_50),
.B(n_1),
.Y(n_98)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_98),
.Y(n_123)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_48),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_99),
.Y(n_126)
);

CKINVDCx14_ASAP7_75t_R g100 ( 
.A(n_57),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_63),
.A2(n_27),
.B1(n_25),
.B2(n_35),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_25),
.B1(n_24),
.B2(n_3),
.Y(n_102)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_102),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_75),
.B(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_108),
.B(n_116),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_54),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_74),
.B(n_66),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_119),
.B(n_129),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_66),
.Y(n_129)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_131),
.B(n_133),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_99),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_134),
.B(n_135),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_84),
.Y(n_135)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_109),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_136),
.B(n_137),
.Y(n_163)
);

A2O1A1O1Ixp25_ASAP7_75t_L g137 ( 
.A1(n_127),
.A2(n_70),
.B(n_76),
.C(n_97),
.D(n_79),
.Y(n_137)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_138),
.B(n_139),
.Y(n_170)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_117),
.Y(n_139)
);

INVx1_ASAP7_75t_SL g140 ( 
.A(n_122),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_141),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_127),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_110),
.B(n_73),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g175 ( 
.A(n_142),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_87),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_152),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_122),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_144),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_105),
.A2(n_129),
.B1(n_119),
.B2(n_112),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_145),
.A2(n_149),
.B1(n_155),
.B2(n_103),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_109),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_146),
.B(n_148),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_76),
.C(n_60),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_147),
.B(n_157),
.C(n_121),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_126),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_112),
.B1(n_104),
.B2(n_114),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_85),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_150),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_151),
.Y(n_169)
);

NOR3xp33_ASAP7_75t_SL g152 ( 
.A(n_114),
.B(n_81),
.C(n_60),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_126),
.Y(n_153)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_153),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_86),
.Y(n_154)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_154),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_104),
.A2(n_90),
.B1(n_96),
.B2(n_50),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_107),
.B(n_50),
.Y(n_156)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_107),
.B(n_47),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_103),
.A2(n_65),
.B1(n_88),
.B2(n_89),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_158),
.A2(n_106),
.B1(n_124),
.B2(n_65),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_115),
.A2(n_68),
.B1(n_71),
.B2(n_80),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_159),
.A2(n_120),
.B1(n_113),
.B2(n_122),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_132),
.A2(n_115),
.B(n_128),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_162),
.A2(n_168),
.B(n_184),
.Y(n_202)
);

NOR2x1_ASAP7_75t_L g164 ( 
.A(n_152),
.B(n_81),
.Y(n_164)
);

NOR2x1_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_183),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_165),
.B(n_174),
.C(n_143),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_166),
.A2(n_140),
.B1(n_137),
.B2(n_113),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_167),
.A2(n_173),
.B1(n_158),
.B2(n_155),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_L g168 ( 
.A1(n_136),
.A2(n_120),
.B(n_121),
.C(n_106),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_128),
.C(n_81),
.Y(n_174)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_156),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_178),
.B(n_180),
.Y(n_199)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g181 ( 
.A(n_132),
.B(n_130),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_181),
.B(n_162),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_128),
.B(n_120),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_24),
.B(n_18),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_186),
.A2(n_1),
.B(n_4),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_170),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_187),
.B(n_192),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_176),
.B(n_157),
.Y(n_188)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_188),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_190),
.B1(n_204),
.B2(n_164),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_182),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_191),
.B(n_193),
.Y(n_218)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_179),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_161),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_179),
.Y(n_194)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_194),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_195),
.B(n_200),
.C(n_201),
.Y(n_213)
);

NOR4xp25_ASAP7_75t_L g196 ( 
.A(n_163),
.B(n_16),
.C(n_15),
.D(n_138),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_177),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_185),
.B(n_113),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_171),
.B(n_16),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g219 ( 
.A(n_198),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_165),
.B(n_64),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_144),
.C(n_24),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_25),
.C(n_2),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_203),
.B(n_206),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_168),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_207),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_185),
.B(n_4),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_208),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_199),
.A2(n_167),
.B1(n_180),
.B2(n_172),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_210),
.A2(n_223),
.B1(n_173),
.B2(n_201),
.Y(n_231)
);

AOI221xp5_ASAP7_75t_L g228 ( 
.A1(n_211),
.A2(n_202),
.B1(n_186),
.B2(n_207),
.C(n_204),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_217),
.Y(n_239)
);

AO22x1_ASAP7_75t_SL g220 ( 
.A1(n_205),
.A2(n_177),
.B1(n_172),
.B2(n_178),
.Y(n_220)
);

BUFx2_ASAP7_75t_L g236 ( 
.A(n_220),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_206),
.B(n_184),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_221),
.B(n_200),
.C(n_175),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_189),
.A2(n_190),
.B1(n_202),
.B2(n_192),
.Y(n_223)
);

HB1xp67_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_224),
.B(n_226),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g227 ( 
.A(n_213),
.B(n_195),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_227),
.B(n_232),
.C(n_213),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_228),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_211),
.A2(n_169),
.B1(n_175),
.B2(n_171),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_229),
.A2(n_234),
.B1(n_235),
.B2(n_217),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_203),
.Y(n_230)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_230),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_231),
.B(n_238),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_220),
.A2(n_169),
.B1(n_160),
.B2(n_166),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_220),
.A2(n_160),
.B1(n_7),
.B2(n_8),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_215),
.B(n_6),
.Y(n_237)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_237),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_6),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_6),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_240),
.B(n_219),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g241 ( 
.A1(n_234),
.A2(n_209),
.B1(n_212),
.B2(n_223),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_241),
.A2(n_214),
.B1(n_216),
.B2(n_226),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_239),
.B(n_235),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_242),
.B(n_249),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_229),
.A2(n_212),
.B(n_210),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_243),
.A2(n_233),
.B(n_236),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_216),
.C(n_221),
.Y(n_256)
);

BUFx24_ASAP7_75t_SL g247 ( 
.A(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_250),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_244),
.B(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_252),
.B(n_250),
.Y(n_263)
);

FAx1_ASAP7_75t_SL g253 ( 
.A(n_243),
.B(n_236),
.CI(n_230),
.CON(n_253),
.SN(n_253)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_253),
.B(n_258),
.Y(n_262)
);

AOI21xp5_ASAP7_75t_L g264 ( 
.A1(n_254),
.A2(n_255),
.B(n_259),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_245),
.A2(n_251),
.B(n_246),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_256),
.B(n_248),
.C(n_8),
.Y(n_266)
);

OR2x2_ASAP7_75t_L g258 ( 
.A(n_242),
.B(n_222),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_256),
.B(n_257),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_263),
.C(n_266),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_253),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_265),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_266),
.B(n_260),
.C(n_259),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_269),
.B(n_9),
.C(n_10),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_262),
.A2(n_7),
.B(n_8),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_270),
.B(n_7),
.Y(n_271)
);

AOI322xp5_ASAP7_75t_L g275 ( 
.A1(n_271),
.A2(n_273),
.A3(n_9),
.B1(n_11),
.B2(n_13),
.C1(n_14),
.C2(n_219),
.Y(n_275)
);

AOI21xp33_ASAP7_75t_L g272 ( 
.A1(n_267),
.A2(n_264),
.B(n_261),
.Y(n_272)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_268),
.B(n_10),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_274),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_275),
.C(n_11),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);


endmodule