module real_jpeg_4048_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_203;
wire n_198;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_216;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_393;
wire n_221;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

AND2x2_ASAP7_75t_SL g70 ( 
.A(n_0),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_SL g84 ( 
.A(n_0),
.B(n_85),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_0),
.B(n_101),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_0),
.B(n_139),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_0),
.B(n_154),
.Y(n_153)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_1),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_1),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g262 ( 
.A(n_1),
.Y(n_262)
);

BUFx5_ASAP7_75t_L g314 ( 
.A(n_1),
.Y(n_314)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_1),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g343 ( 
.A(n_1),
.Y(n_343)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_2),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_2),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g160 ( 
.A(n_2),
.Y(n_160)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_2),
.Y(n_217)
);

INVx6_ASAP7_75t_L g283 ( 
.A(n_2),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_3),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_3),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_3),
.B(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_3),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_3),
.B(n_182),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_3),
.B(n_270),
.Y(n_269)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_3),
.B(n_292),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_3),
.B(n_226),
.Y(n_408)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_4),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g192 ( 
.A(n_4),
.Y(n_192)
);

BUFx5_ASAP7_75t_L g393 ( 
.A(n_4),
.Y(n_393)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_5),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_6),
.B(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_6),
.B(n_311),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_6),
.B(n_314),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_6),
.B(n_333),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g348 ( 
.A(n_6),
.B(n_120),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_6),
.B(n_58),
.Y(n_377)
);

AND2x2_ASAP7_75t_L g392 ( 
.A(n_6),
.B(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_7),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_7),
.Y(n_130)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_7),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g330 ( 
.A(n_7),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_8),
.Y(n_503)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_9),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_10),
.Y(n_140)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_10),
.Y(n_205)
);

BUFx3_ASAP7_75t_L g271 ( 
.A(n_10),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g191 ( 
.A(n_11),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_11),
.B(n_46),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_11),
.B(n_58),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_11),
.B(n_225),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_11),
.B(n_322),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_11),
.B(n_330),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_11),
.B(n_374),
.Y(n_373)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_11),
.B(n_399),
.Y(n_398)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_13),
.B(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_13),
.B(n_62),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_13),
.B(n_122),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_13),
.B(n_128),
.Y(n_127)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_13),
.B(n_203),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g224 ( 
.A(n_13),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_14),
.B(n_44),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_14),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_14),
.B(n_102),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_14),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_14),
.B(n_194),
.Y(n_193)
);

AND2x2_ASAP7_75t_SL g284 ( 
.A(n_14),
.B(n_285),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_14),
.B(n_226),
.Y(n_362)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_14),
.B(n_407),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_15),
.B(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_15),
.B(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_15),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g295 ( 
.A(n_15),
.B(n_58),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_15),
.B(n_324),
.Y(n_323)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_15),
.B(n_341),
.Y(n_340)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_15),
.B(n_290),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_16),
.B(n_216),
.Y(n_215)
);

NAND2x1p5_ASAP7_75t_L g266 ( 
.A(n_16),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_16),
.B(n_308),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_16),
.B(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_16),
.B(n_347),
.Y(n_346)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_16),
.B(n_379),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_16),
.B(n_389),
.Y(n_388)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_17),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_17),
.B(n_158),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_17),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_17),
.B(n_230),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_17),
.B(n_290),
.Y(n_289)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_17),
.B(n_343),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_17),
.B(n_365),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g400 ( 
.A(n_17),
.B(n_401),
.Y(n_400)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_19),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_19),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_19),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_19),
.B(n_228),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_19),
.B(n_262),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_498),
.B(n_501),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_173),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_172),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_107),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_25),
.B(n_107),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_90),
.B1(n_91),
.B2(n_106),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_26),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_60),
.C(n_74),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_27),
.A2(n_28),
.B1(n_169),
.B2(n_171),
.Y(n_168)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

XNOR2xp5_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_42),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_30),
.B(n_35),
.C(n_42),
.Y(n_105)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_34),
.Y(n_115)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_47),
.C(n_54),
.Y(n_42)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_43),
.B(n_143),
.Y(n_142)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_47),
.A2(n_48),
.B1(n_54),
.B2(n_55),
.Y(n_143)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

BUFx2_ASAP7_75t_L g198 ( 
.A(n_51),
.Y(n_198)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g274 ( 
.A(n_52),
.Y(n_274)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_53),
.Y(n_88)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_53),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_53),
.Y(n_187)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_53),
.Y(n_379)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g230 ( 
.A(n_59),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g391 ( 
.A(n_59),
.Y(n_391)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_60),
.A2(n_74),
.B1(n_75),
.B2(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_60),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_64),
.C(n_69),
.Y(n_60)
);

XNOR2xp5_ASAP7_75t_SL g164 ( 
.A(n_61),
.B(n_165),
.Y(n_164)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_64),
.A2(n_65),
.B1(n_138),
.B2(n_141),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_64),
.A2(n_65),
.B1(n_69),
.B2(n_70),
.Y(n_165)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_65),
.B(n_135),
.C(n_138),
.Y(n_166)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_68),
.Y(n_228)
);

INVx5_ASAP7_75t_L g294 ( 
.A(n_68),
.Y(n_294)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_68),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_69),
.A2(n_70),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_70),
.B(n_83),
.C(n_89),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_72),
.Y(n_124)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx5_ASAP7_75t_L g196 ( 
.A(n_72),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g290 ( 
.A(n_72),
.Y(n_290)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_73),
.Y(n_183)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_73),
.Y(n_334)
);

INVx3_ASAP7_75t_L g347 ( 
.A(n_73),
.Y(n_347)
);

BUFx3_ASAP7_75t_L g375 ( 
.A(n_73),
.Y(n_375)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_81),
.B1(n_82),
.B2(n_89),
.Y(n_75)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_76),
.Y(n_89)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_80),
.Y(n_79)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_80),
.Y(n_210)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_83),
.A2(n_84),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_105),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_97),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_94),
.B(n_96),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_104),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_103),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_163),
.C(n_168),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_108),
.A2(n_109),
.B1(n_481),
.B2(n_482),
.Y(n_480)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_142),
.C(n_144),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_SL g485 ( 
.A(n_110),
.B(n_486),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_125),
.C(n_134),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_111),
.A2(n_112),
.B1(n_125),
.B2(n_234),
.Y(n_233)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_116),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_113),
.B(n_117),
.C(n_121),
.Y(n_167)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_121),
.Y(n_116)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx11_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_125),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_127),
.C(n_131),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_126),
.B(n_131),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_127),
.B(n_246),
.Y(n_245)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g232 ( 
.A(n_134),
.B(n_233),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_137),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_138),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_147),
.C(n_152),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_138),
.A2(n_141),
.B1(n_152),
.B2(n_153),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_140),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g407 ( 
.A(n_140),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_142),
.A2(n_144),
.B1(n_145),
.B2(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_142),
.Y(n_487)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_156),
.C(n_161),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g239 ( 
.A(n_146),
.B(n_240),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g242 ( 
.A(n_147),
.B(n_243),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_149),
.Y(n_267)
);

INVx6_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_152),
.A2(n_153),
.B1(n_202),
.B2(n_206),
.Y(n_201)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_153),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_153),
.B(n_200),
.C(n_202),
.Y(n_244)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g240 ( 
.A1(n_156),
.A2(n_157),
.B1(n_161),
.B2(n_162),
.Y(n_240)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_161),
.A2(n_162),
.B1(n_209),
.B2(n_211),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_162),
.B(n_211),
.C(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_163),
.B(n_168),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_167),
.Y(n_163)
);

FAx1_ASAP7_75t_SL g488 ( 
.A(n_164),
.B(n_166),
.CI(n_167),
.CON(n_488),
.SN(n_488)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_169),
.Y(n_171)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_175),
.A2(n_478),
.B(n_495),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_296),
.B(n_477),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_177),
.B(n_247),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_177),
.B(n_247),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_231),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_178),
.B(n_232),
.C(n_235),
.Y(n_494)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_207),
.C(n_213),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_179),
.B(n_250),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_189),
.C(n_199),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g461 ( 
.A(n_180),
.B(n_462),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g180 ( 
.A(n_181),
.B(n_184),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_181),
.B(n_185),
.C(n_188),
.Y(n_212)
);

INVx5_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_189),
.A2(n_190),
.B1(n_199),
.B2(n_463),
.Y(n_462)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_193),
.C(n_197),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_191),
.B(n_197),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_193),
.B(n_452),
.Y(n_451)
);

BUFx3_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx5_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_199),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g206 ( 
.A(n_202),
.Y(n_206)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_204),
.Y(n_322)
);

INVx8_ASAP7_75t_L g341 ( 
.A(n_204),
.Y(n_341)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_205),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_213),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_209),
.Y(n_211)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_212),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_227),
.C(n_229),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_214),
.B(n_277),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_218),
.C(n_224),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_SL g258 ( 
.A(n_215),
.B(n_259),
.Y(n_258)
);

INVx6_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_219),
.B(n_224),
.Y(n_259)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx3_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g308 ( 
.A(n_222),
.Y(n_308)
);

INVx5_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

HB1xp67_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_227),
.B(n_229),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_241),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_237),
.B(n_239),
.C(n_241),
.Y(n_489)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_244),
.C(n_245),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_245),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_251),
.C(n_254),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_249),
.B(n_252),
.Y(n_472)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_254),
.B(n_472),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_275),
.C(n_278),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_256),
.B(n_465),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_260),
.C(n_264),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_257),
.A2(n_258),
.B1(n_443),
.B2(n_444),
.Y(n_442)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_260),
.A2(n_261),
.B(n_263),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_260),
.B(n_264),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_263),
.Y(n_260)
);

MAJx2_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_268),
.C(n_272),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_265),
.A2(n_266),
.B1(n_268),
.B2(n_269),
.Y(n_420)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

BUFx8_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_272),
.B(n_420),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_273),
.B(n_360),
.Y(n_359)
);

INVx6_ASAP7_75t_L g399 ( 
.A(n_274),
.Y(n_399)
);

AOI22xp33_ASAP7_75t_L g465 ( 
.A1(n_275),
.A2(n_276),
.B1(n_278),
.B2(n_466),
.Y(n_465)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_278),
.Y(n_466)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_291),
.C(n_295),
.Y(n_278)
);

INVx1_ASAP7_75t_SL g279 ( 
.A(n_280),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_280),
.B(n_454),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_284),
.C(n_288),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_281),
.B(n_432),
.Y(n_431)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_284),
.A2(n_288),
.B1(n_289),
.B2(n_433),
.Y(n_432)
);

INVx1_ASAP7_75t_SL g433 ( 
.A(n_284),
.Y(n_433)
);

INVx8_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

INVx3_ASAP7_75t_L g311 ( 
.A(n_286),
.Y(n_311)
);

BUFx5_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_287),
.Y(n_360)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g454 ( 
.A(n_291),
.B(n_295),
.Y(n_454)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

AOI21x1_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_470),
.B(n_476),
.Y(n_296)
);

OAI21x1_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_457),
.B(n_469),
.Y(n_297)
);

AOI21x1_ASAP7_75t_L g298 ( 
.A1(n_299),
.A2(n_439),
.B(n_456),
.Y(n_298)
);

OAI21x1_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_413),
.B(n_438),
.Y(n_299)
);

AOI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_301),
.A2(n_383),
.B(n_412),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g301 ( 
.A1(n_302),
.A2(n_352),
.B(n_382),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g302 ( 
.A1(n_303),
.A2(n_336),
.B(n_351),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g303 ( 
.A1(n_304),
.A2(n_316),
.B(n_335),
.Y(n_303)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_305),
.A2(n_312),
.B(n_315),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_306),
.B(n_310),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_310),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_309),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_307),
.B(n_313),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_307),
.B(n_309),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_318),
.Y(n_335)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_319),
.A2(n_320),
.B1(n_326),
.B2(n_327),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_319),
.B(n_329),
.C(n_331),
.Y(n_350)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_323),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_321),
.B(n_323),
.Y(n_344)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_328),
.A2(n_329),
.B1(n_331),
.B2(n_332),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_332),
.Y(n_331)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g336 ( 
.A(n_337),
.B(n_350),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_337),
.B(n_350),
.Y(n_351)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_338),
.B(n_345),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_344),
.Y(n_338)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_339),
.B(n_344),
.C(n_354),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_340),
.B(n_342),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g357 ( 
.A(n_340),
.B(n_342),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_345),
.Y(n_354)
);

BUFx24_ASAP7_75t_SL g504 ( 
.A(n_345),
.Y(n_504)
);

FAx1_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_348),
.CI(n_349),
.CON(n_345),
.SN(n_345)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_346),
.B(n_370),
.C(n_371),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_348),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_353),
.B(n_355),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_368),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_356),
.B(n_369),
.C(n_372),
.Y(n_411)
);

XOR2xp5_ASAP7_75t_L g356 ( 
.A(n_357),
.B(n_358),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_357),
.B(n_359),
.C(n_361),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_359),
.B(n_361),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_362),
.A2(n_363),
.B1(n_364),
.B2(n_367),
.Y(n_361)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_362),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g394 ( 
.A(n_363),
.B(n_367),
.Y(n_394)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XNOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_372),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_373),
.B(n_376),
.Y(n_372)
);

MAJx2_ASAP7_75t_L g410 ( 
.A(n_373),
.B(n_378),
.C(n_380),
.Y(n_410)
);

INVx3_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_377),
.A2(n_378),
.B1(n_380),
.B2(n_381),
.Y(n_376)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_377),
.Y(n_380)
);

INVx1_ASAP7_75t_SL g381 ( 
.A(n_378),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_384),
.B(n_411),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g412 ( 
.A(n_384),
.B(n_411),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_396),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_395),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_386),
.B(n_395),
.C(n_437),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_L g386 ( 
.A(n_387),
.B(n_394),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_392),
.Y(n_387)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_388),
.Y(n_427)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

INVx4_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

CKINVDCx14_ASAP7_75t_R g428 ( 
.A(n_392),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_394),
.B(n_427),
.C(n_428),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g437 ( 
.A(n_396),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_397),
.B(n_403),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_397),
.B(n_405),
.C(n_409),
.Y(n_416)
);

BUFx24_ASAP7_75t_SL g507 ( 
.A(n_397),
.Y(n_507)
);

FAx1_ASAP7_75t_SL g397 ( 
.A(n_398),
.B(n_400),
.CI(n_402),
.CON(n_397),
.SN(n_397)
);

MAJx2_ASAP7_75t_L g424 ( 
.A(n_398),
.B(n_400),
.C(n_402),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g403 ( 
.A1(n_404),
.A2(n_405),
.B1(n_409),
.B2(n_410),
.Y(n_403)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_408),
.Y(n_405)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_406),
.B(n_408),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g409 ( 
.A(n_410),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_436),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_414),
.B(n_436),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_425),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_416),
.B(n_417),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_416),
.B(n_417),
.C(n_425),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_421),
.B2(n_422),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_418),
.B(n_448),
.C(n_449),
.Y(n_447)
);

INVx1_ASAP7_75t_SL g418 ( 
.A(n_419),
.Y(n_418)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_423),
.B(n_424),
.Y(n_422)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_424),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_SL g425 ( 
.A(n_426),
.B(n_429),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_426),
.B(n_430),
.C(n_435),
.Y(n_445)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_430),
.A2(n_431),
.B1(n_434),
.B2(n_435),
.Y(n_429)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_430),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_431),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_455),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_SL g456 ( 
.A(n_440),
.B(n_455),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_446),
.Y(n_440)
);

XOR2xp5_ASAP7_75t_L g441 ( 
.A(n_442),
.B(n_445),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_442),
.B(n_445),
.C(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_443),
.Y(n_444)
);

INVxp67_ASAP7_75t_L g468 ( 
.A(n_446),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_447),
.B(n_450),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g459 ( 
.A(n_447),
.B(n_451),
.C(n_453),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_453),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_458),
.B(n_467),
.Y(n_457)
);

NAND2xp5_ASAP7_75t_L g469 ( 
.A(n_458),
.B(n_467),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_459),
.B(n_460),
.Y(n_458)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_459),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_464),
.Y(n_460)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_461),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_464),
.B(n_474),
.C(n_475),
.Y(n_473)
);

NAND2xp5_ASAP7_75t_SL g470 ( 
.A(n_471),
.B(n_473),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_471),
.B(n_473),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_490),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g495 ( 
.A1(n_479),
.A2(n_496),
.B(n_497),
.Y(n_495)
);

NOR2xp33_ASAP7_75t_SL g479 ( 
.A(n_480),
.B(n_483),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_483),
.Y(n_497)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_481),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_488),
.C(n_489),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g492 ( 
.A1(n_484),
.A2(n_485),
.B1(n_488),
.B2(n_493),
.Y(n_492)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_488),
.Y(n_493)
);

BUFx24_ASAP7_75t_SL g506 ( 
.A(n_488),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_492),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_491),
.B(n_494),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_491),
.B(n_494),
.Y(n_496)
);

BUFx4f_ASAP7_75t_SL g498 ( 
.A(n_499),
.Y(n_498)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_499),
.Y(n_502)
);

INVx13_ASAP7_75t_L g499 ( 
.A(n_500),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_503),
.Y(n_501)
);


endmodule