module real_jpeg_2225_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_288;
wire n_286;
wire n_215;
wire n_83;
wire n_249;
wire n_292;
wire n_221;
wire n_166;
wire n_176;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_291;
wire n_236;
wire n_47;
wire n_131;
wire n_281;
wire n_271;
wire n_276;
wire n_163;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_293;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_290;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_285;
wire n_160;
wire n_45;
wire n_211;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_294;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_198;
wire n_192;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_205;
wire n_258;
wire n_195;
wire n_289;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_278;
wire n_130;
wire n_144;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_226;
wire n_277;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_167;
wire n_202;
wire n_128;
wire n_179;
wire n_244;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_283;
wire n_85;
wire n_102;
wire n_181;
wire n_274;
wire n_101;
wire n_256;
wire n_182;
wire n_273;
wire n_96;
wire n_253;
wire n_269;
wire n_89;
wire n_16;

INVx2_ASAP7_75t_L g59 ( 
.A(n_0),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_1),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_2),
.Y(n_89)
);

OAI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_3),
.A2(n_32),
.B1(n_33),
.B2(n_40),
.Y(n_39)
);

CKINVDCx14_ASAP7_75t_R g40 ( 
.A(n_3),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_3),
.A2(n_23),
.B1(n_24),
.B2(n_40),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_3),
.A2(n_40),
.B1(n_58),
.B2(n_60),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_3),
.A2(n_40),
.B1(n_47),
.B2(n_48),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g36 ( 
.A1(n_4),
.A2(n_23),
.B1(n_24),
.B2(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_4),
.A2(n_37),
.B1(n_47),
.B2(n_48),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_4),
.A2(n_32),
.B1(n_33),
.B2(n_37),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_4),
.A2(n_37),
.B1(n_58),
.B2(n_60),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_4),
.B(n_29),
.C(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_4),
.B(n_31),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_4),
.B(n_44),
.C(n_48),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_4),
.B(n_89),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_4),
.B(n_56),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_4),
.B(n_57),
.C(n_60),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_4),
.B(n_50),
.Y(n_229)
);

BUFx4f_ASAP7_75t_L g44 ( 
.A(n_5),
.Y(n_44)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_L g22 ( 
.A1(n_7),
.A2(n_23),
.B1(n_24),
.B2(n_27),
.Y(n_22)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_7),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_7),
.A2(n_27),
.B1(n_32),
.B2(n_33),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_7),
.A2(n_27),
.B1(n_58),
.B2(n_60),
.Y(n_154)
);

BUFx16f_ASAP7_75t_L g57 ( 
.A(n_8),
.Y(n_57)
);

INVx2_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_11),
.A2(n_32),
.B1(n_33),
.B2(n_52),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_47),
.B1(n_48),
.B2(n_52),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_11),
.A2(n_23),
.B1(n_24),
.B2(n_52),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_11),
.A2(n_52),
.B1(n_58),
.B2(n_60),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_12),
.A2(n_15),
.B(n_292),
.Y(n_14)
);

BUFx10_ASAP7_75t_L g293 ( 
.A(n_12),
.Y(n_293)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_13),
.Y(n_49)
);

AOI21xp33_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_287),
.B(n_290),
.Y(n_15)
);

AO21x1_ASAP7_75t_L g16 ( 
.A1(n_17),
.A2(n_74),
.B(n_286),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_71),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_18),
.B(n_71),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_65),
.C(n_67),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_19),
.B(n_283),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_38),
.C(n_53),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_20),
.A2(n_95),
.B1(n_99),
.B2(n_100),
.Y(n_94)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_20),
.A2(n_100),
.B1(n_138),
.B2(n_156),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_20),
.B(n_138),
.C(n_148),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_20),
.A2(n_100),
.B1(n_273),
.B2(n_274),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_28),
.B1(n_31),
.B2(n_36),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g122 ( 
.A1(n_22),
.A2(n_68),
.B(n_70),
.Y(n_122)
);

O2A1O1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_23),
.A2(n_29),
.B(n_30),
.C(n_31),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_29),
.Y(n_30)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_24),
.B(n_151),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_28),
.B(n_36),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

AO22x1_ASAP7_75t_SL g31 ( 
.A1(n_29),
.A2(n_32),
.B1(n_33),
.B2(n_35),
.Y(n_31)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_31),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_32),
.A2(n_33),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_33),
.B(n_205),
.Y(n_204)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_36),
.B(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_38),
.A2(n_53),
.B1(n_260),
.B2(n_275),
.Y(n_274)
);

CKINVDCx16_ASAP7_75t_R g275 ( 
.A(n_38),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_41),
.B1(n_50),
.B2(n_51),
.Y(n_38)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_39),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_41),
.A2(n_50),
.B1(n_96),
.B2(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_42),
.B(n_46),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_42),
.B(n_98),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_42),
.A2(n_46),
.B(n_98),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

AOI22x1_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_46),
.A2(n_262),
.B(n_263),
.Y(n_261)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_47),
.A2(n_48),
.B1(n_57),
.B2(n_61),
.Y(n_63)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_48),
.B(n_222),
.Y(n_221)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

AO21x1_ASAP7_75t_L g95 ( 
.A1(n_50),
.A2(n_96),
.B(n_97),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_51),
.B(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_53),
.A2(n_260),
.B1(n_261),
.B2(n_264),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_53),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_53),
.B(n_122),
.C(n_261),
.Y(n_276)
);

AND2x2_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_64),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_62),
.Y(n_54)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_62),
.B1(n_84),
.B2(n_85),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_55),
.A2(n_107),
.B(n_108),
.Y(n_106)
);

OA22x2_ASAP7_75t_L g119 ( 
.A1(n_55),
.A2(n_62),
.B1(n_84),
.B2(n_85),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_55),
.A2(n_62),
.B(n_85),
.Y(n_164)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_56),
.B(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_56),
.A2(n_64),
.B1(n_110),
.B2(n_137),
.Y(n_136)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_57),
.Y(n_61)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_58),
.B(n_89),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_60),
.B(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_62),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_65),
.B(n_67),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_69),
.B(n_70),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_68),
.A2(n_69),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_68),
.B(n_72),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g287 ( 
.A(n_71),
.B(n_288),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_71),
.B(n_288),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_73),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g74 ( 
.A1(n_75),
.A2(n_281),
.B(n_285),
.Y(n_74)
);

AOI21xp33_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_252),
.B(n_278),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_142),
.B(n_251),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_123),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_78),
.B(n_123),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_101),
.C(n_112),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_79),
.B(n_101),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_93),
.B2(n_94),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_80),
.B(n_95),
.C(n_100),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_86),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_82),
.A2(n_83),
.B1(n_86),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_82),
.A2(n_83),
.B1(n_229),
.B2(n_230),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_82),
.A2(n_83),
.B1(n_202),
.B2(n_242),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_83),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_83),
.B(n_197),
.C(n_202),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_83),
.B(n_153),
.C(n_229),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_86),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_87),
.B(n_91),
.Y(n_104)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_88),
.A2(n_89),
.B1(n_117),
.B2(n_154),
.Y(n_153)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_90),
.A2(n_91),
.B(n_116),
.Y(n_115)
);

OA21x2_ASAP7_75t_L g173 ( 
.A1(n_91),
.A2(n_116),
.B(n_174),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_95),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_95),
.B(n_121),
.C(n_164),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_95),
.A2(n_99),
.B1(n_164),
.B2(n_169),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_95),
.A2(n_99),
.B1(n_118),
.B2(n_119),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_95),
.B(n_118),
.C(n_237),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_97),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_98),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_105),
.B1(n_106),
.B2(n_111),
.Y(n_101)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_102),
.B(n_106),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_102),
.A2(n_111),
.B1(n_131),
.B2(n_133),
.Y(n_130)
);

INVxp33_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_104),
.B(n_117),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g137 ( 
.A(n_107),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_110),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_111),
.A2(n_127),
.B(n_133),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_112),
.B(n_249),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_120),
.C(n_121),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_113),
.A2(n_114),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_118),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_115),
.A2(n_118),
.B1(n_119),
.B2(n_161),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_118),
.A2(n_119),
.B1(n_221),
.B2(n_223),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_118),
.B(n_223),
.Y(n_231)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_120),
.A2(n_121),
.B1(n_122),
.B2(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_120),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_121),
.A2(n_122),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_121),
.A2(n_122),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_121),
.A2(n_122),
.B1(n_271),
.B2(n_272),
.Y(n_270)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_122),
.B(n_272),
.C(n_276),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_141),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_134),
.B2(n_135),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_126),
.B(n_134),
.C(n_141),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_128),
.B1(n_129),
.B2(n_130),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_131),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_132),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_138),
.B(n_140),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_138),
.Y(n_140)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_138),
.B(n_172),
.C(n_173),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_138),
.A2(n_156),
.B1(n_198),
.B2(n_201),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_140),
.A2(n_256),
.B1(n_257),
.B2(n_265),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_140),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_143),
.A2(n_246),
.B(n_250),
.Y(n_142)
);

OAI211xp5_ASAP7_75t_L g143 ( 
.A1(n_144),
.A2(n_175),
.B(n_189),
.C(n_190),
.Y(n_143)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_165),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_145),
.B(n_165),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_157),
.B2(n_158),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_160),
.C(n_162),
.Y(n_177)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_149),
.B(n_152),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g170 ( 
.A1(n_149),
.A2(n_150),
.B1(n_152),
.B2(n_153),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_152),
.A2(n_153),
.B1(n_227),
.B2(n_228),
.Y(n_226)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_153),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_153),
.B(n_217),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_154),
.Y(n_174)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_164),
.Y(n_169)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_170),
.C(n_171),
.Y(n_165)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_166),
.B(n_195),
.Y(n_194)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g195 ( 
.A(n_170),
.B(n_171),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_172),
.A2(n_173),
.B1(n_199),
.B2(n_200),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_172),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_173),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_SL g190 ( 
.A(n_176),
.B(n_191),
.C(n_192),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_177),
.B(n_178),
.Y(n_176)
);

OR2x2_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_178),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_180),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_179),
.B(n_181),
.C(n_187),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_186),
.B2(n_187),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_208),
.B(n_245),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_194),
.B(n_196),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_197),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_198),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_200),
.B(n_220),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_206),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_203),
.A2(n_204),
.B1(n_206),
.B2(n_207),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_239),
.B(n_244),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_210),
.A2(n_233),
.B(n_238),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_225),
.B(n_232),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_219),
.B(n_224),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_216),
.B(n_218),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_221),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_231),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_231),
.Y(n_232)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_235),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_235),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_237),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_243),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_240),
.B(n_243),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_247),
.B(n_248),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_268),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_254),
.B(n_267),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_254),
.B(n_267),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_266),
.Y(n_254)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_257),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_257),
.B(n_265),
.C(n_266),
.Y(n_277)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g264 ( 
.A(n_261),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_268),
.A2(n_279),
.B(n_280),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_269),
.B(n_277),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_269),
.B(n_277),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_276),
.Y(n_269)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_284),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_282),
.B(n_284),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_291),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_294),
.Y(n_292)
);


endmodule