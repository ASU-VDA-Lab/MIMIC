module fake_jpeg_13411_n_599 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_599);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_599;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_349;
wire n_21;
wire n_393;
wire n_288;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_535;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx8_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_11),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx24_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_0),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_9),
.B(n_10),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_3),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

BUFx10_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_2),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_1),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_39),
.Y(n_58)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g148 ( 
.A(n_59),
.Y(n_148)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_39),
.Y(n_60)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_60),
.Y(n_145)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_45),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_61),
.Y(n_173)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_20),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_62),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_63),
.Y(n_134)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_30),
.Y(n_64)
);

CKINVDCx6p67_ASAP7_75t_R g195 ( 
.A(n_64),
.Y(n_195)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx3_ASAP7_75t_L g138 ( 
.A(n_65),
.Y(n_138)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_18),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_66),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_SL g136 ( 
.A(n_67),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_68),
.Y(n_157)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_69),
.Y(n_146)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_70),
.Y(n_161)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_45),
.Y(n_71)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_71),
.Y(n_152)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_72),
.Y(n_155)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_33),
.Y(n_74)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_74),
.Y(n_127)
);

BUFx24_ASAP7_75t_L g75 ( 
.A(n_30),
.Y(n_75)
);

BUFx24_ASAP7_75t_L g191 ( 
.A(n_75),
.Y(n_191)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_17),
.Y(n_76)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_76),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_41),
.B(n_16),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_77),
.B(n_93),
.Y(n_141)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_17),
.Y(n_78)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_78),
.Y(n_142)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx5_ASAP7_75t_L g188 ( 
.A(n_79),
.Y(n_188)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_18),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_80),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_35),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_81),
.Y(n_178)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_82),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_52),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g194 ( 
.A(n_83),
.Y(n_194)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_84),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_52),
.Y(n_85)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_86),
.Y(n_154)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_18),
.Y(n_87)
);

INVx6_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_88),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx6_ASAP7_75t_L g183 ( 
.A(n_89),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_90),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_54),
.Y(n_91)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_91),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_55),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_92),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_41),
.B(n_16),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_51),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_115),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_95),
.Y(n_190)
);

INVx11_ASAP7_75t_L g96 ( 
.A(n_30),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g135 ( 
.A(n_96),
.Y(n_135)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx8_ASAP7_75t_L g98 ( 
.A(n_21),
.Y(n_98)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_98),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_55),
.Y(n_99)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_19),
.B(n_15),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_100),
.B(n_13),
.Y(n_180)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_21),
.Y(n_101)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_101),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_56),
.Y(n_102)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_102),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_56),
.Y(n_103)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_104),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_56),
.Y(n_105)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_105),
.Y(n_174)
);

INVx8_ASAP7_75t_L g106 ( 
.A(n_21),
.Y(n_106)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_106),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_19),
.B(n_15),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_107),
.B(n_110),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_46),
.Y(n_108)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_108),
.Y(n_189)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_46),
.Y(n_109)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_109),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_32),
.B(n_14),
.Y(n_110)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_50),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_111),
.B(n_114),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_37),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g133 ( 
.A(n_112),
.B(n_113),
.Y(n_133)
);

INVx4_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_25),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_22),
.B(n_14),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_17),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_116),
.B(n_120),
.Y(n_139)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_46),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_117),
.B(n_118),
.Y(n_170)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_25),
.Y(n_118)
);

INVx8_ASAP7_75t_L g119 ( 
.A(n_51),
.Y(n_119)
);

INVx6_ASAP7_75t_SL g128 ( 
.A(n_119),
.Y(n_128)
);

INVx11_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_17),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_44),
.Y(n_153)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_25),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_44),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_115),
.A2(n_40),
.B1(n_32),
.B2(n_34),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_123),
.A2(n_124),
.B1(n_159),
.B2(n_162),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_66),
.A2(n_40),
.B1(n_34),
.B2(n_24),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g126 ( 
.A1(n_80),
.A2(n_26),
.B1(n_40),
.B2(n_57),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_126),
.A2(n_140),
.B1(n_147),
.B2(n_149),
.Y(n_263)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_31),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_129),
.B(n_132),
.Y(n_208)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_75),
.B(n_79),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_87),
.A2(n_101),
.B1(n_117),
.B2(n_108),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_76),
.A2(n_26),
.B1(n_24),
.B2(n_34),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_76),
.A2(n_26),
.B1(n_24),
.B2(n_51),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_59),
.A2(n_62),
.B1(n_51),
.B2(n_119),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_151),
.A2(n_181),
.B1(n_192),
.B2(n_99),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_153),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_109),
.A2(n_57),
.B1(n_53),
.B2(n_42),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_63),
.A2(n_53),
.B1(n_42),
.B2(n_38),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_62),
.A2(n_37),
.B1(n_44),
.B2(n_22),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_L g227 ( 
.A1(n_167),
.A2(n_196),
.B(n_29),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_175),
.B(n_27),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_73),
.B(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_179),
.B(n_182),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_180),
.B(n_186),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_98),
.A2(n_44),
.B1(n_37),
.B2(n_49),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_97),
.B(n_36),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_112),
.B(n_27),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g192 ( 
.A1(n_106),
.A2(n_44),
.B1(n_31),
.B2(n_49),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_68),
.B(n_28),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_193),
.B(n_1),
.Y(n_239)
);

A2O1A1Ixp33_ASAP7_75t_L g196 ( 
.A1(n_64),
.A2(n_43),
.B(n_47),
.C(n_38),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_81),
.B(n_29),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_85),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g202 ( 
.A1(n_126),
.A2(n_105),
.B1(n_103),
.B2(n_102),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g312 ( 
.A1(n_202),
.A2(n_242),
.B1(n_249),
.B2(n_253),
.Y(n_312)
);

INVx2_ASAP7_75t_SL g203 ( 
.A(n_191),
.Y(n_203)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_203),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_173),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_204),
.B(n_225),
.Y(n_281)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_127),
.Y(n_205)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

INVx4_ASAP7_75t_SL g206 ( 
.A(n_191),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g277 ( 
.A(n_206),
.B(n_213),
.Y(n_277)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_191),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_207),
.B(n_226),
.Y(n_280)
);

BUFx3_ASAP7_75t_L g209 ( 
.A(n_177),
.Y(n_209)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_209),
.Y(n_290)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_160),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g275 ( 
.A(n_210),
.Y(n_275)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_166),
.Y(n_211)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_211),
.Y(n_287)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_170),
.Y(n_212)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_212),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_214),
.A2(n_218),
.B(n_261),
.Y(n_326)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_165),
.Y(n_215)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

OAI22xp33_ASAP7_75t_SL g216 ( 
.A1(n_129),
.A2(n_95),
.B1(n_92),
.B2(n_91),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_216),
.A2(n_227),
.B1(n_258),
.B2(n_260),
.Y(n_301)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_160),
.Y(n_217)
);

INVx3_ASAP7_75t_L g289 ( 
.A(n_217),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_187),
.A2(n_90),
.B1(n_89),
.B2(n_86),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_169),
.Y(n_219)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_219),
.Y(n_274)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_220),
.Y(n_308)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_174),
.Y(n_222)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_168),
.B(n_47),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_223),
.B(n_246),
.Y(n_286)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

INVx2_ASAP7_75t_L g294 ( 
.A(n_224),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_187),
.Y(n_225)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_198),
.Y(n_228)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_228),
.Y(n_299)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_130),
.Y(n_229)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_229),
.Y(n_315)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_145),
.Y(n_230)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_230),
.Y(n_324)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_132),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_231),
.Y(n_279)
);

OAI22xp33_ASAP7_75t_L g232 ( 
.A1(n_181),
.A2(n_83),
.B1(n_28),
.B2(n_43),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_232),
.A2(n_188),
.B1(n_133),
.B2(n_199),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_177),
.Y(n_234)
);

INVx3_ASAP7_75t_L g298 ( 
.A(n_234),
.Y(n_298)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_146),
.Y(n_235)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_235),
.Y(n_322)
);

INVx11_ASAP7_75t_L g236 ( 
.A(n_135),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g325 ( 
.A(n_236),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_0),
.Y(n_237)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_237),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_134),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_238),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_239),
.B(n_243),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_196),
.B(n_1),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_240),
.B(n_256),
.Y(n_295)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_171),
.Y(n_241)
);

INVx3_ASAP7_75t_L g323 ( 
.A(n_241),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g242 ( 
.A1(n_161),
.A2(n_47),
.B1(n_14),
.B2(n_13),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_131),
.B(n_13),
.Y(n_243)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_137),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g273 ( 
.A(n_244),
.Y(n_273)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_171),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_245),
.B(n_247),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g246 ( 
.A(n_156),
.B(n_1),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_163),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_199),
.A2(n_12),
.B1(n_10),
.B2(n_3),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_184),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_250),
.Y(n_292)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_163),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_251),
.B(n_252),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_134),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_SL g253 ( 
.A1(n_161),
.A2(n_136),
.B1(n_142),
.B2(n_148),
.Y(n_253)
);

INVx5_ASAP7_75t_L g254 ( 
.A(n_144),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_254),
.B(n_255),
.Y(n_320)
);

INVx1_ASAP7_75t_SL g255 ( 
.A(n_195),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_164),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_139),
.B(n_1),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_257),
.B(n_264),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_SL g258 ( 
.A1(n_136),
.A2(n_12),
.B1(n_4),
.B2(n_5),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_197),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_259),
.B(n_265),
.Y(n_328)
);

OAI22xp33_ASAP7_75t_SL g260 ( 
.A1(n_151),
.A2(n_192),
.B1(n_147),
.B2(n_149),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g261 ( 
.A1(n_142),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_141),
.B(n_4),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_262),
.B(n_271),
.Y(n_302)
);

AND2x2_ASAP7_75t_SL g264 ( 
.A(n_144),
.B(n_5),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_197),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_143),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_266),
.A2(n_269),
.B1(n_195),
.B2(n_188),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_128),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_267),
.Y(n_296)
);

BUFx6f_ASAP7_75t_L g268 ( 
.A(n_157),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g305 ( 
.A(n_268),
.Y(n_305)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_148),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_269)
);

INVx6_ASAP7_75t_L g270 ( 
.A(n_157),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g307 ( 
.A(n_270),
.Y(n_307)
);

CKINVDCx14_ASAP7_75t_R g271 ( 
.A(n_195),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_282),
.B(n_247),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_231),
.A2(n_158),
.B1(n_143),
.B2(n_185),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_283),
.A2(n_285),
.B1(n_313),
.B2(n_317),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_284),
.A2(n_293),
.B1(n_310),
.B2(n_316),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_263),
.A2(n_154),
.B1(n_185),
.B2(n_183),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_201),
.A2(n_176),
.B1(n_150),
.B2(n_183),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_239),
.B(n_240),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_303),
.B(n_304),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_212),
.B(n_154),
.Y(n_304)
);

A2O1A1Ixp33_ASAP7_75t_L g309 ( 
.A1(n_208),
.A2(n_135),
.B(n_152),
.C(n_138),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_311),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_201),
.A2(n_150),
.B1(n_176),
.B2(n_194),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_213),
.B(n_158),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_232),
.A2(n_194),
.B1(n_178),
.B2(n_190),
.Y(n_313)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_218),
.A2(n_178),
.B1(n_190),
.B2(n_137),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_213),
.A2(n_125),
.B1(n_135),
.B2(n_8),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_223),
.B(n_125),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_318),
.B(n_251),
.Y(n_367)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_257),
.A2(n_8),
.B1(n_9),
.B2(n_233),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_321),
.A2(n_203),
.B1(n_266),
.B2(n_254),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_286),
.B(n_233),
.C(n_205),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_332),
.C(n_343),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_SL g331 ( 
.A(n_297),
.B(n_262),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_331),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_286),
.B(n_248),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_303),
.B(n_221),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_333),
.B(n_335),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_296),
.B(n_211),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_334),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_295),
.B(n_257),
.Y(n_335)
);

AOI22xp33_ASAP7_75t_SL g336 ( 
.A1(n_284),
.A2(n_203),
.B1(n_255),
.B2(n_217),
.Y(n_336)
);

AOI22xp33_ASAP7_75t_SL g381 ( 
.A1(n_336),
.A2(n_339),
.B1(n_359),
.B2(n_369),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_295),
.B(n_237),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_338),
.B(n_349),
.Y(n_377)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_278),
.Y(n_340)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_340),
.Y(n_375)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_278),
.Y(n_342)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_342),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_318),
.B(n_220),
.C(n_256),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_296),
.B(n_230),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_344),
.Y(n_398)
);

INVxp67_ASAP7_75t_L g345 ( 
.A(n_320),
.Y(n_345)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_345),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_326),
.A2(n_264),
.B(n_206),
.Y(n_347)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_347),
.A2(n_277),
.B(n_309),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g348 ( 
.A(n_327),
.B(n_264),
.C(n_246),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_355),
.C(n_365),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g349 ( 
.A(n_328),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_287),
.Y(n_350)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_350),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_280),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_351),
.B(n_358),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_310),
.A2(n_237),
.B1(n_246),
.B2(n_245),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_352),
.A2(n_357),
.B1(n_370),
.B2(n_276),
.Y(n_372)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

INVx1_ASAP7_75t_SL g383 ( 
.A(n_353),
.Y(n_383)
);

INVx3_ASAP7_75t_L g354 ( 
.A(n_291),
.Y(n_354)
);

INVx1_ASAP7_75t_SL g391 ( 
.A(n_354),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_306),
.B(n_235),
.C(n_229),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_301),
.A2(n_241),
.B1(n_215),
.B2(n_219),
.Y(n_356)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_356),
.A2(n_316),
.B1(n_312),
.B2(n_304),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g357 ( 
.A1(n_293),
.A2(n_222),
.B1(n_250),
.B2(n_210),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_308),
.Y(n_358)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_291),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_360),
.A2(n_317),
.B(n_277),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_314),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_361),
.B(n_362),
.Y(n_392)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_308),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_281),
.B(n_224),
.Y(n_363)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_363),
.Y(n_409)
);

INVx2_ASAP7_75t_L g364 ( 
.A(n_322),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g395 ( 
.A(n_364),
.B(n_366),
.Y(n_395)
);

AND2x2_ASAP7_75t_SL g365 ( 
.A(n_311),
.B(n_228),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_315),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_367),
.B(n_368),
.Y(n_397)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g369 ( 
.A(n_276),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_306),
.A2(n_270),
.B1(n_265),
.B2(n_259),
.Y(n_370)
);

INVx8_ASAP7_75t_L g371 ( 
.A(n_305),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_371),
.A2(n_305),
.B1(n_290),
.B2(n_298),
.Y(n_386)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_372),
.A2(n_376),
.B1(n_378),
.B2(n_390),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_374),
.A2(n_333),
.B1(n_338),
.B2(n_335),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_346),
.A2(n_301),
.B1(n_285),
.B2(n_326),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_346),
.A2(n_313),
.B1(n_282),
.B2(n_302),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_394),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g428 ( 
.A1(n_386),
.A2(n_396),
.B(n_399),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g390 ( 
.A1(n_347),
.A2(n_337),
.B1(n_341),
.B2(n_352),
.Y(n_390)
);

AOI22xp5_ASAP7_75t_L g393 ( 
.A1(n_329),
.A2(n_300),
.B1(n_277),
.B2(n_302),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_393),
.A2(n_407),
.B1(n_408),
.B2(n_355),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_337),
.A2(n_297),
.B1(n_307),
.B2(n_327),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_341),
.A2(n_367),
.B(n_360),
.Y(n_399)
);

AOI21xp5_ASAP7_75t_L g400 ( 
.A1(n_360),
.A2(n_273),
.B(n_279),
.Y(n_400)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_400),
.A2(n_405),
.B(n_406),
.Y(n_429)
);

MAJIxp5_ASAP7_75t_L g401 ( 
.A(n_330),
.B(n_324),
.C(n_315),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_401),
.B(n_299),
.C(n_294),
.Y(n_432)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_357),
.A2(n_307),
.B1(n_319),
.B2(n_324),
.Y(n_402)
);

AOI22x1_ASAP7_75t_L g415 ( 
.A1(n_402),
.A2(n_350),
.B1(n_353),
.B2(n_366),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_361),
.A2(n_238),
.B1(n_252),
.B2(n_268),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_404),
.B(n_371),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g405 ( 
.A1(n_343),
.A2(n_273),
.B(n_290),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_365),
.A2(n_292),
.B(n_298),
.Y(n_406)
);

AOI22xp5_ASAP7_75t_L g407 ( 
.A1(n_329),
.A2(n_356),
.B1(n_365),
.B2(n_339),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_365),
.A2(n_349),
.B1(n_340),
.B2(n_342),
.Y(n_408)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_395),
.Y(n_410)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_410),
.Y(n_452)
);

AOI22xp5_ASAP7_75t_L g451 ( 
.A1(n_411),
.A2(n_417),
.B1(n_394),
.B2(n_399),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_382),
.B(n_332),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_412),
.B(n_416),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g413 ( 
.A(n_380),
.Y(n_413)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_413),
.Y(n_457)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_395),
.Y(n_414)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_414),
.Y(n_458)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_415),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_382),
.B(n_348),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g418 ( 
.A1(n_376),
.A2(n_371),
.B1(n_358),
.B2(n_362),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_418),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_385),
.B(n_331),
.Y(n_419)
);

NOR2xp33_ASAP7_75t_SL g466 ( 
.A(n_419),
.B(n_426),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g420 ( 
.A(n_392),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_420),
.B(n_430),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g422 ( 
.A(n_383),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_422),
.B(n_438),
.Y(n_470)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_423),
.Y(n_460)
);

AO21x1_ASAP7_75t_L g424 ( 
.A1(n_399),
.A2(n_370),
.B(n_348),
.Y(n_424)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_424),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_392),
.B(n_368),
.Y(n_425)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_380),
.B(n_364),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_388),
.B(n_292),
.Y(n_427)
);

AO21x1_ASAP7_75t_L g447 ( 
.A1(n_427),
.A2(n_440),
.B(n_442),
.Y(n_447)
);

CKINVDCx14_ASAP7_75t_R g430 ( 
.A(n_388),
.Y(n_430)
);

XNOR2x1_ASAP7_75t_L g431 ( 
.A(n_389),
.B(n_236),
.Y(n_431)
);

XNOR2x1_ASAP7_75t_L g462 ( 
.A(n_431),
.B(n_389),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_432),
.B(n_433),
.Y(n_453)
);

MAJIxp5_ASAP7_75t_L g433 ( 
.A(n_382),
.B(n_289),
.C(n_325),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_375),
.Y(n_434)
);

INVxp67_ASAP7_75t_L g455 ( 
.A(n_434),
.Y(n_455)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g446 ( 
.A(n_435),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g436 ( 
.A(n_377),
.B(n_289),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g471 ( 
.A(n_436),
.B(n_405),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_408),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_437),
.Y(n_464)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_375),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_396),
.A2(n_275),
.B(n_299),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_398),
.B(n_275),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_441),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_397),
.B(n_354),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_397),
.B(n_323),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g468 ( 
.A(n_443),
.B(n_383),
.Y(n_468)
);

AOI32xp33_ASAP7_75t_SL g444 ( 
.A1(n_390),
.A2(n_359),
.A3(n_323),
.B1(n_234),
.B2(n_209),
.Y(n_444)
);

OAI21xp5_ASAP7_75t_SL g459 ( 
.A1(n_444),
.A2(n_400),
.B(n_408),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_SL g448 ( 
.A(n_416),
.B(n_412),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g479 ( 
.A(n_448),
.B(n_450),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_SL g450 ( 
.A(n_421),
.B(n_389),
.Y(n_450)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_451),
.A2(n_374),
.B1(n_381),
.B2(n_423),
.Y(n_497)
);

HB1xp67_ASAP7_75t_L g490 ( 
.A(n_459),
.Y(n_490)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_417),
.A2(n_378),
.B1(n_372),
.B2(n_402),
.Y(n_461)
);

OAI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_461),
.A2(n_463),
.B1(n_474),
.B2(n_476),
.Y(n_482)
);

XOR2xp5_ASAP7_75t_L g481 ( 
.A(n_462),
.B(n_469),
.Y(n_481)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_437),
.A2(n_402),
.B1(n_377),
.B2(n_409),
.Y(n_463)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_468),
.Y(n_478)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_401),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_473),
.Y(n_493)
);

OAI21xp5_ASAP7_75t_SL g472 ( 
.A1(n_428),
.A2(n_393),
.B(n_407),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_L g477 ( 
.A1(n_472),
.A2(n_428),
.B(n_429),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g473 ( 
.A(n_433),
.B(n_401),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g474 ( 
.A1(n_420),
.A2(n_409),
.B1(n_406),
.B2(n_407),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_410),
.A2(n_406),
.B1(n_398),
.B2(n_387),
.Y(n_476)
);

FAx1_ASAP7_75t_L g523 ( 
.A(n_477),
.B(n_491),
.CI(n_444),
.CON(n_523),
.SN(n_523)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_457),
.Y(n_480)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_480),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_475),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_483),
.B(n_484),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g484 ( 
.A1(n_454),
.A2(n_421),
.B(n_439),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_449),
.B(n_448),
.C(n_473),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_485),
.B(n_487),
.C(n_489),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_460),
.A2(n_429),
.B1(n_414),
.B2(n_439),
.Y(n_486)
);

OAI22xp5_ASAP7_75t_L g505 ( 
.A1(n_486),
.A2(n_502),
.B1(n_474),
.B2(n_476),
.Y(n_505)
);

MAJIxp5_ASAP7_75t_L g487 ( 
.A(n_449),
.B(n_432),
.C(n_436),
.Y(n_487)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_453),
.B(n_424),
.Y(n_488)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_488),
.B(n_500),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_453),
.B(n_373),
.C(n_393),
.Y(n_489)
);

OAI21xp5_ASAP7_75t_L g491 ( 
.A1(n_454),
.A2(n_440),
.B(n_427),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_470),
.Y(n_492)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_492),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_455),
.B(n_425),
.Y(n_494)
);

HB1xp67_ASAP7_75t_L g525 ( 
.A(n_494),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g495 ( 
.A(n_462),
.B(n_373),
.C(n_415),
.Y(n_495)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_495),
.B(n_496),
.C(n_498),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_450),
.B(n_415),
.C(n_422),
.Y(n_496)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_497),
.A2(n_499),
.B1(n_445),
.B2(n_456),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g498 ( 
.A(n_469),
.B(n_413),
.C(n_443),
.Y(n_498)
);

OAI22xp5_ASAP7_75t_L g499 ( 
.A1(n_461),
.A2(n_381),
.B1(n_374),
.B2(n_426),
.Y(n_499)
);

XOR2x1_ASAP7_75t_SL g500 ( 
.A(n_463),
.B(n_442),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_470),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_501),
.B(n_383),
.Y(n_526)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_470),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_471),
.B(n_438),
.C(n_434),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_503),
.B(n_498),
.C(n_500),
.Y(n_514)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_505),
.Y(n_530)
);

AOI22xp5_ASAP7_75t_SL g506 ( 
.A1(n_482),
.A2(n_445),
.B1(n_467),
.B2(n_466),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g536 ( 
.A(n_506),
.B(n_514),
.Y(n_536)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_487),
.B(n_493),
.Y(n_508)
);

XOR2xp5_ASAP7_75t_L g531 ( 
.A(n_508),
.B(n_510),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g527 ( 
.A(n_509),
.Y(n_527)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_493),
.B(n_451),
.Y(n_510)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_486),
.A2(n_456),
.B1(n_447),
.B2(n_464),
.Y(n_513)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_513),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_468),
.C(n_472),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_515),
.B(n_516),
.C(n_522),
.Y(n_535)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_503),
.B(n_458),
.C(n_452),
.Y(n_516)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_488),
.B(n_465),
.Y(n_517)
);

XNOR2xp5_ASAP7_75t_L g539 ( 
.A(n_517),
.B(n_519),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_489),
.B(n_457),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_SL g540 ( 
.A(n_518),
.B(n_521),
.Y(n_540)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_481),
.B(n_447),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g521 ( 
.A(n_495),
.B(n_459),
.Y(n_521)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_481),
.B(n_455),
.C(n_446),
.Y(n_522)
);

NAND2x1_ASAP7_75t_L g544 ( 
.A(n_523),
.B(n_478),
.Y(n_544)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_526),
.Y(n_534)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_516),
.Y(n_528)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_528),
.Y(n_546)
);

OR2x2_ASAP7_75t_L g529 ( 
.A(n_504),
.B(n_490),
.Y(n_529)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_529),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_482),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_537),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g537 ( 
.A(n_508),
.B(n_479),
.C(n_496),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_507),
.B(n_479),
.C(n_492),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_538),
.B(n_543),
.Y(n_553)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_524),
.A2(n_502),
.B1(n_491),
.B2(n_477),
.Y(n_541)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_541),
.A2(n_523),
.B1(n_525),
.B2(n_515),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_522),
.B(n_478),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g550 ( 
.A(n_542),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_512),
.B(n_484),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_544),
.B(n_511),
.Y(n_552)
);

BUFx24_ASAP7_75t_SL g545 ( 
.A(n_529),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_545),
.B(n_559),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_SL g547 ( 
.A(n_535),
.B(n_507),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_547),
.B(n_548),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_512),
.C(n_510),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_554),
.Y(n_569)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_552),
.B(n_539),
.Y(n_571)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_531),
.B(n_519),
.C(n_517),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_531),
.B(n_494),
.C(n_520),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_555),
.B(n_556),
.Y(n_572)
);

XNOR2xp5_ASAP7_75t_L g556 ( 
.A(n_536),
.B(n_523),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_534),
.B(n_480),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g564 ( 
.A(n_557),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_SL g558 ( 
.A1(n_527),
.A2(n_386),
.B1(n_403),
.B2(n_379),
.Y(n_558)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_558),
.B(n_541),
.Y(n_561)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_530),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_561),
.B(n_563),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g563 ( 
.A1(n_560),
.A2(n_533),
.B1(n_559),
.B2(n_550),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_549),
.B(n_540),
.Y(n_565)
);

NOR2xp33_ASAP7_75t_SL g575 ( 
.A(n_565),
.B(n_555),
.Y(n_575)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_551),
.B(n_538),
.C(n_536),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_568),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g568 ( 
.A(n_556),
.B(n_539),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g570 ( 
.A1(n_553),
.A2(n_537),
.B(n_542),
.Y(n_570)
);

XOR2xp5_ASAP7_75t_L g576 ( 
.A(n_570),
.B(n_571),
.Y(n_576)
);

OAI211xp5_ASAP7_75t_L g574 ( 
.A1(n_566),
.A2(n_546),
.B(n_544),
.C(n_548),
.Y(n_574)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

AOI22xp33_ASAP7_75t_SL g586 ( 
.A1(n_575),
.A2(n_576),
.B1(n_571),
.B2(n_581),
.Y(n_586)
);

AND2x2_ASAP7_75t_L g577 ( 
.A(n_569),
.B(n_554),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g588 ( 
.A(n_577),
.B(n_578),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_564),
.B(n_558),
.Y(n_578)
);

OAI21xp5_ASAP7_75t_SL g579 ( 
.A1(n_567),
.A2(n_552),
.B(n_391),
.Y(n_579)
);

XOR2xp5_ASAP7_75t_L g587 ( 
.A(n_579),
.B(n_568),
.Y(n_587)
);

AOI22xp33_ASAP7_75t_SL g580 ( 
.A1(n_563),
.A2(n_391),
.B1(n_403),
.B2(n_379),
.Y(n_580)
);

INVxp67_ASAP7_75t_L g583 ( 
.A(n_580),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_SL g582 ( 
.A(n_562),
.B(n_359),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_582),
.B(n_391),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_584),
.B(n_586),
.Y(n_591)
);

OAI21xp5_ASAP7_75t_SL g585 ( 
.A1(n_573),
.A2(n_572),
.B(n_571),
.Y(n_585)
);

A2O1A1Ixp33_ASAP7_75t_L g590 ( 
.A1(n_585),
.A2(n_578),
.B(n_581),
.C(n_561),
.Y(n_590)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_587),
.B(n_404),
.C(n_384),
.Y(n_592)
);

OAI21xp5_ASAP7_75t_SL g594 ( 
.A1(n_590),
.A2(n_593),
.B(n_588),
.Y(n_594)
);

INVxp67_ASAP7_75t_L g595 ( 
.A(n_592),
.Y(n_595)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_588),
.B(n_272),
.C(n_274),
.Y(n_593)
);

OAI22xp5_ASAP7_75t_L g596 ( 
.A1(n_594),
.A2(n_589),
.B1(n_591),
.B2(n_583),
.Y(n_596)
);

OAI22xp5_ASAP7_75t_L g597 ( 
.A1(n_596),
.A2(n_595),
.B1(n_272),
.B2(n_274),
.Y(n_597)
);

NOR3xp33_ASAP7_75t_L g598 ( 
.A(n_597),
.B(n_294),
.C(n_288),
.Y(n_598)
);

AOI21xp5_ASAP7_75t_L g599 ( 
.A1(n_598),
.A2(n_288),
.B(n_9),
.Y(n_599)
);


endmodule