module fake_jpeg_24608_n_203 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_203);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_203;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_14),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_SL g31 ( 
.A(n_3),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_7),
.Y(n_33)
);

INVx6_ASAP7_75t_SL g34 ( 
.A(n_23),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_29),
.Y(n_35)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_39),
.Y(n_53)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_37),
.A2(n_20),
.B1(n_23),
.B2(n_21),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.Y(n_38)
);

AND2x2_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_40),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_27),
.B(n_1),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g40 ( 
.A(n_24),
.B(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_24),
.Y(n_43)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_30),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_45),
.B(n_2),
.Y(n_74)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_22),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_38),
.B(n_30),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_47),
.B(n_52),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_40),
.B(n_27),
.Y(n_48)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_48),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_20),
.B1(n_23),
.B2(n_31),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_51),
.A2(n_57),
.B1(n_21),
.B2(n_32),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_30),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_R g82 ( 
.A(n_54),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_31),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_20),
.B1(n_21),
.B2(n_28),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_35),
.B(n_31),
.Y(n_59)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_34),
.B(n_19),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_19),
.Y(n_73)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_61),
.B(n_80),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_41),
.C(n_43),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_62),
.B(n_32),
.C(n_18),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_59),
.B(n_41),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_63),
.B(n_79),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_65),
.A2(n_66),
.B1(n_18),
.B2(n_28),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_44),
.A2(n_16),
.B1(n_33),
.B2(n_17),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_68),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_53),
.B(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_69),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g71 ( 
.A(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_73),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_72),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_81),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_L g75 ( 
.A1(n_51),
.A2(n_55),
.B1(n_44),
.B2(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_75),
.A2(n_47),
.B1(n_52),
.B2(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_53),
.B(n_55),
.Y(n_76)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_76),
.Y(n_90)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_49),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_77),
.B(n_78),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_56),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_29),
.Y(n_79)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_58),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_4),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_46),
.B(n_22),
.Y(n_83)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_83),
.Y(n_99)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_87),
.A2(n_98),
.B1(n_64),
.B2(n_67),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_48),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_91),
.B(n_61),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_78),
.B(n_46),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_92),
.B(n_106),
.C(n_84),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_74),
.B(n_29),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_102),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_73),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_103),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_72),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_97),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_58),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_65),
.Y(n_103)
);

FAx1_ASAP7_75t_SL g104 ( 
.A(n_62),
.B(n_19),
.CI(n_22),
.CON(n_104),
.SN(n_104)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_104),
.B(n_63),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_58),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_105),
.B(n_22),
.Y(n_127)
);

NOR3xp33_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_84),
.C(n_64),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_109),
.B(n_120),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_112),
.A2(n_115),
.B1(n_121),
.B2(n_99),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_89),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_113),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_107),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_114),
.B(n_119),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_103),
.A2(n_82),
.B1(n_75),
.B2(n_67),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_116),
.B(n_117),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_81),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_118),
.B(n_124),
.C(n_127),
.Y(n_131)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_108),
.Y(n_119)
);

NOR3xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_70),
.C(n_63),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_87),
.A2(n_70),
.B1(n_80),
.B2(n_77),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_86),
.Y(n_122)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_101),
.Y(n_125)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_125),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_90),
.B(n_33),
.Y(n_126)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_126),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_128),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_92),
.Y(n_129)
);

BUFx3_ASAP7_75t_L g146 ( 
.A(n_129),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_130),
.B(n_139),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_93),
.C(n_106),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_132),
.B(n_112),
.C(n_124),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_115),
.A2(n_105),
.B1(n_102),
.B2(n_96),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_137),
.B1(n_141),
.B2(n_4),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_129),
.A2(n_94),
.B(n_90),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_148),
.B(n_127),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_121),
.A2(n_95),
.B1(n_104),
.B2(n_88),
.Y(n_137)
);

AOI322xp5_ASAP7_75t_L g139 ( 
.A1(n_123),
.A2(n_104),
.A3(n_88),
.B1(n_93),
.B2(n_91),
.C1(n_99),
.C2(n_94),
.Y(n_139)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_111),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_147),
.B(n_25),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_125),
.A2(n_85),
.B1(n_26),
.B2(n_25),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_133),
.B(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_149),
.B(n_150),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_119),
.Y(n_150)
);

XOR2x2_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_118),
.Y(n_152)
);

OA21x2_ASAP7_75t_SL g167 ( 
.A1(n_152),
.A2(n_155),
.B(n_134),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_143),
.B(n_123),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_153),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_161),
.B1(n_162),
.B2(n_163),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_116),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_155),
.B(n_156),
.C(n_131),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_138),
.B(n_26),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_157),
.B(n_160),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_145),
.Y(n_158)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_138),
.B(n_17),
.Y(n_160)
);

A2O1A1Ixp33_ASAP7_75t_SL g161 ( 
.A1(n_146),
.A2(n_16),
.B(n_5),
.C(n_6),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_142),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_167),
.B(n_148),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_169),
.B(n_173),
.C(n_174),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_163),
.A2(n_140),
.B1(n_144),
.B2(n_136),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_171),
.B(n_137),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_156),
.B(n_132),
.C(n_135),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_151),
.C(n_134),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_175),
.B(n_177),
.Y(n_185)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_170),
.B(n_161),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_161),
.Y(n_178)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_164),
.B(n_161),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_179),
.B(n_180),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_165),
.B(n_9),
.Y(n_180)
);

AOI322xp5_ASAP7_75t_L g181 ( 
.A1(n_166),
.A2(n_15),
.A3(n_9),
.B1(n_10),
.B2(n_11),
.C1(n_13),
.C2(n_7),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_181),
.B(n_183),
.C(n_172),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_169),
.B(n_10),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_170),
.B1(n_171),
.B2(n_173),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_186),
.A2(n_172),
.B1(n_181),
.B2(n_164),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_189),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_182),
.B(n_174),
.C(n_165),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_191),
.B(n_193),
.C(n_187),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_186),
.B(n_15),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_188),
.B(n_13),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g196 ( 
.A(n_194),
.B(n_195),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_185),
.B(n_190),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_197),
.B(n_198),
.Y(n_200)
);

OAI321xp33_ASAP7_75t_L g198 ( 
.A1(n_193),
.A2(n_184),
.A3(n_192),
.B1(n_189),
.B2(n_5),
.C(n_8),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_6),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_199),
.B(n_8),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_201),
.B(n_196),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_202),
.B(n_200),
.Y(n_203)
);


endmodule