module fake_netlist_5_711_n_2183 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_220, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_219, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_221, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2183);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_220;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_219;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_221;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2183;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2031;
wire n_2076;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_798;
wire n_350;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_344;
wire n_1218;
wire n_1931;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_857;
wire n_832;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1891;
wire n_1662;
wire n_1711;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_604;
wire n_314;
wire n_368;
wire n_433;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_448;
wire n_259;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2131;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1363;
wire n_1301;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1439;
wire n_1312;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_356;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2008;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_1),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_16),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_51),
.Y(n_224)
);

INVx2_ASAP7_75t_SL g225 ( 
.A(n_125),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_135),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_44),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_113),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_87),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_30),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_141),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_152),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_107),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_150),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_55),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_153),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_45),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_168),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_108),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_27),
.Y(n_242)
);

INVx1_ASAP7_75t_SL g243 ( 
.A(n_29),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_49),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_140),
.Y(n_245)
);

BUFx2_ASAP7_75t_L g246 ( 
.A(n_73),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_20),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_26),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_155),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_144),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_170),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g252 ( 
.A(n_72),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_93),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_191),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_147),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_65),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_64),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_68),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_42),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_2),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_201),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_149),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_80),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_53),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_98),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_169),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_47),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_158),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_128),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_212),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_82),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_181),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_23),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g274 ( 
.A(n_20),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_56),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g276 ( 
.A(n_54),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_67),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_177),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_3),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_104),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_189),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_66),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_95),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g284 ( 
.A(n_57),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_18),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_16),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_30),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_79),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_100),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_2),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_182),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_142),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_37),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_87),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_220),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_33),
.Y(n_296)
);

BUFx2_ASAP7_75t_SL g297 ( 
.A(n_198),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_15),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_160),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_42),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_4),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_28),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_102),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_86),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_216),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_29),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_124),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_18),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_28),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_37),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_133),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_156),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g313 ( 
.A(n_185),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_64),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_32),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_31),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_85),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_203),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_75),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_47),
.Y(n_320)
);

INVx2_ASAP7_75t_SL g321 ( 
.A(n_213),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_199),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_165),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_209),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_69),
.Y(n_325)
);

BUFx6f_ASAP7_75t_L g326 ( 
.A(n_122),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_206),
.Y(n_327)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_23),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_74),
.Y(n_329)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_25),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_119),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_14),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_101),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_96),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_175),
.Y(n_335)
);

BUFx2_ASAP7_75t_L g336 ( 
.A(n_103),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_77),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_27),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_163),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_110),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_15),
.Y(n_341)
);

BUFx10_ASAP7_75t_L g342 ( 
.A(n_134),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_186),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_24),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_6),
.Y(n_345)
);

INVx1_ASAP7_75t_SL g346 ( 
.A(n_132),
.Y(n_346)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_136),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_106),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_172),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_6),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_13),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_33),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_112),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_79),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_162),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_131),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_97),
.Y(n_357)
);

CKINVDCx5p33_ASAP7_75t_R g358 ( 
.A(n_92),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_214),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_205),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_76),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_176),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_1),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_46),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_105),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_91),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_66),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g368 ( 
.A(n_46),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_48),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_217),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_59),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_120),
.Y(n_372)
);

BUFx10_ASAP7_75t_L g373 ( 
.A(n_114),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_58),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_3),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_215),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_195),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_9),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_196),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_10),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_171),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_9),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_70),
.Y(n_383)
);

CKINVDCx5p33_ASAP7_75t_R g384 ( 
.A(n_211),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_84),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_78),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_89),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_84),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_197),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_26),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_11),
.Y(n_391)
);

HB1xp67_ASAP7_75t_L g392 ( 
.A(n_115),
.Y(n_392)
);

INVx1_ASAP7_75t_SL g393 ( 
.A(n_89),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_130),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_154),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_194),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_146),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_208),
.Y(n_398)
);

CKINVDCx11_ASAP7_75t_R g399 ( 
.A(n_72),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g400 ( 
.A(n_139),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_56),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_41),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_178),
.Y(n_403)
);

BUFx5_ASAP7_75t_L g404 ( 
.A(n_14),
.Y(n_404)
);

INVx2_ASAP7_75t_SL g405 ( 
.A(n_48),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_121),
.Y(n_406)
);

INVx1_ASAP7_75t_SL g407 ( 
.A(n_174),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_80),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_166),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g410 ( 
.A(n_38),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_12),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_145),
.Y(n_412)
);

BUFx5_ASAP7_75t_L g413 ( 
.A(n_45),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_38),
.Y(n_414)
);

INVx2_ASAP7_75t_SL g415 ( 
.A(n_143),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_67),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_78),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_90),
.Y(n_418)
);

CKINVDCx5p33_ASAP7_75t_R g419 ( 
.A(n_71),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_77),
.Y(n_420)
);

BUFx2_ASAP7_75t_SL g421 ( 
.A(n_159),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_69),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_34),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_184),
.Y(n_424)
);

BUFx10_ASAP7_75t_L g425 ( 
.A(n_180),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_13),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_61),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_88),
.Y(n_428)
);

CKINVDCx16_ASAP7_75t_R g429 ( 
.A(n_74),
.Y(n_429)
);

INVx1_ASAP7_75t_SL g430 ( 
.A(n_94),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_39),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_204),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_22),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_76),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_34),
.Y(n_435)
);

CKINVDCx5p33_ASAP7_75t_R g436 ( 
.A(n_62),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_11),
.Y(n_437)
);

INVxp67_ASAP7_75t_SL g438 ( 
.A(n_392),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_276),
.Y(n_439)
);

INVxp67_ASAP7_75t_L g440 ( 
.A(n_246),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g441 ( 
.A(n_246),
.B(n_0),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_399),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_226),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_235),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_229),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_276),
.B(n_0),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_237),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_276),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_276),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_239),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_L g451 ( 
.A(n_336),
.B(n_4),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_276),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_227),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_252),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_245),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_250),
.Y(n_456)
);

CKINVDCx5p33_ASAP7_75t_R g457 ( 
.A(n_251),
.Y(n_457)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_232),
.Y(n_458)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_227),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_276),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_276),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_336),
.B(n_225),
.Y(n_462)
);

HB1xp67_ASAP7_75t_L g463 ( 
.A(n_429),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_255),
.Y(n_464)
);

INVxp67_ASAP7_75t_SL g465 ( 
.A(n_320),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_240),
.Y(n_466)
);

BUFx10_ASAP7_75t_L g467 ( 
.A(n_225),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_261),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_276),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_276),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_321),
.B(n_5),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_266),
.Y(n_472)
);

INVx2_ASAP7_75t_L g473 ( 
.A(n_404),
.Y(n_473)
);

CKINVDCx5p33_ASAP7_75t_R g474 ( 
.A(n_268),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_404),
.B(n_5),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_404),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_404),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_404),
.Y(n_478)
);

CKINVDCx5p33_ASAP7_75t_R g479 ( 
.A(n_270),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_281),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_404),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_404),
.Y(n_482)
);

BUFx6f_ASAP7_75t_SL g483 ( 
.A(n_241),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_404),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_404),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_321),
.B(n_7),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_291),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_241),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_289),
.Y(n_489)
);

CKINVDCx20_ASAP7_75t_R g490 ( 
.A(n_292),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_R g491 ( 
.A(n_312),
.B(n_347),
.Y(n_491)
);

INVxp33_ASAP7_75t_L g492 ( 
.A(n_236),
.Y(n_492)
);

CKINVDCx16_ASAP7_75t_R g493 ( 
.A(n_241),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_295),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_413),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_303),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_413),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_413),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_313),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_236),
.Y(n_500)
);

INVxp33_ASAP7_75t_SL g501 ( 
.A(n_222),
.Y(n_501)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_413),
.Y(n_502)
);

INVxp33_ASAP7_75t_L g503 ( 
.A(n_242),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_318),
.Y(n_504)
);

CKINVDCx5p33_ASAP7_75t_R g505 ( 
.A(n_322),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_413),
.Y(n_506)
);

CKINVDCx16_ASAP7_75t_R g507 ( 
.A(n_342),
.Y(n_507)
);

CKINVDCx16_ASAP7_75t_R g508 ( 
.A(n_342),
.Y(n_508)
);

INVxp33_ASAP7_75t_L g509 ( 
.A(n_242),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_413),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_413),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_362),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_323),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_413),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_327),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_413),
.Y(n_516)
);

CKINVDCx20_ASAP7_75t_R g517 ( 
.A(n_331),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_328),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_328),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_328),
.Y(n_520)
);

INVxp67_ASAP7_75t_L g521 ( 
.A(n_263),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_334),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g523 ( 
.A(n_263),
.Y(n_523)
);

INVx1_ASAP7_75t_L g524 ( 
.A(n_328),
.Y(n_524)
);

NOR2xp67_ASAP7_75t_L g525 ( 
.A(n_320),
.B(n_7),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_328),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_320),
.Y(n_527)
);

HB1xp67_ASAP7_75t_L g528 ( 
.A(n_224),
.Y(n_528)
);

BUFx2_ASAP7_75t_L g529 ( 
.A(n_284),
.Y(n_529)
);

CKINVDCx5p33_ASAP7_75t_R g530 ( 
.A(n_335),
.Y(n_530)
);

CKINVDCx5p33_ASAP7_75t_R g531 ( 
.A(n_340),
.Y(n_531)
);

CKINVDCx5p33_ASAP7_75t_R g532 ( 
.A(n_355),
.Y(n_532)
);

INVxp67_ASAP7_75t_L g533 ( 
.A(n_264),
.Y(n_533)
);

CKINVDCx5p33_ASAP7_75t_R g534 ( 
.A(n_356),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_223),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_L g536 ( 
.A(n_415),
.B(n_8),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_223),
.Y(n_537)
);

INVxp33_ASAP7_75t_SL g538 ( 
.A(n_230),
.Y(n_538)
);

CKINVDCx20_ASAP7_75t_R g539 ( 
.A(n_358),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_275),
.Y(n_540)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_275),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_359),
.Y(n_542)
);

INVxp67_ASAP7_75t_L g543 ( 
.A(n_264),
.Y(n_543)
);

INVxp67_ASAP7_75t_SL g544 ( 
.A(n_284),
.Y(n_544)
);

CKINVDCx5p33_ASAP7_75t_R g545 ( 
.A(n_360),
.Y(n_545)
);

CKINVDCx5p33_ASAP7_75t_R g546 ( 
.A(n_365),
.Y(n_546)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_415),
.B(n_8),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_330),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_366),
.Y(n_549)
);

INVxp33_ASAP7_75t_L g550 ( 
.A(n_271),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_330),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_271),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_285),
.Y(n_553)
);

CKINVDCx20_ASAP7_75t_R g554 ( 
.A(n_370),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g555 ( 
.A(n_228),
.B(n_10),
.Y(n_555)
);

CKINVDCx20_ASAP7_75t_R g556 ( 
.A(n_372),
.Y(n_556)
);

INVxp67_ASAP7_75t_L g557 ( 
.A(n_285),
.Y(n_557)
);

INVxp33_ASAP7_75t_L g558 ( 
.A(n_287),
.Y(n_558)
);

CKINVDCx5p33_ASAP7_75t_R g559 ( 
.A(n_376),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_518),
.Y(n_560)
);

INVxp67_ASAP7_75t_L g561 ( 
.A(n_454),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_518),
.Y(n_562)
);

NAND2x1_ASAP7_75t_L g563 ( 
.A(n_527),
.B(n_326),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_491),
.Y(n_564)
);

CKINVDCx5p33_ASAP7_75t_R g565 ( 
.A(n_517),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_539),
.Y(n_566)
);

BUFx8_ASAP7_75t_L g567 ( 
.A(n_483),
.Y(n_567)
);

CKINVDCx5p33_ASAP7_75t_R g568 ( 
.A(n_554),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_519),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_519),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_445),
.Y(n_571)
);

NOR2xp67_ASAP7_75t_L g572 ( 
.A(n_559),
.B(n_357),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g573 ( 
.A(n_443),
.B(n_269),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_444),
.B(n_447),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_463),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_520),
.Y(n_576)
);

BUFx2_ASAP7_75t_L g577 ( 
.A(n_529),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_SL g578 ( 
.A(n_488),
.B(n_342),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_520),
.Y(n_579)
);

OAI21x1_ASAP7_75t_L g580 ( 
.A1(n_452),
.A2(n_280),
.B(n_269),
.Y(n_580)
);

CKINVDCx5p33_ASAP7_75t_R g581 ( 
.A(n_556),
.Y(n_581)
);

AND2x4_ASAP7_75t_L g582 ( 
.A(n_465),
.B(n_525),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_450),
.Y(n_583)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_488),
.Y(n_584)
);

INVxp67_ASAP7_75t_L g585 ( 
.A(n_528),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_L g586 ( 
.A(n_455),
.B(n_280),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_456),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_524),
.Y(n_588)
);

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_457),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_464),
.Y(n_590)
);

INVxp67_ASAP7_75t_L g591 ( 
.A(n_529),
.Y(n_591)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_458),
.Y(n_592)
);

BUFx6f_ASAP7_75t_L g593 ( 
.A(n_526),
.Y(n_593)
);

INVxp67_ASAP7_75t_L g594 ( 
.A(n_544),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_468),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_472),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_474),
.Y(n_597)
);

OR2x2_ASAP7_75t_L g598 ( 
.A(n_440),
.B(n_405),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_479),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_452),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_527),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_473),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_446),
.Y(n_603)
);

INVx1_ASAP7_75t_SL g604 ( 
.A(n_466),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_489),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_475),
.Y(n_606)
);

CKINVDCx5p33_ASAP7_75t_R g607 ( 
.A(n_480),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_487),
.B(n_494),
.Y(n_608)
);

NAND2xp33_ASAP7_75t_L g609 ( 
.A(n_441),
.B(n_231),
.Y(n_609)
);

OAI21x1_ASAP7_75t_L g610 ( 
.A1(n_473),
.A2(n_395),
.B(n_394),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_439),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_496),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_439),
.Y(n_613)
);

INVx2_ASAP7_75t_L g614 ( 
.A(n_448),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_490),
.Y(n_615)
);

BUFx3_ASAP7_75t_L g616 ( 
.A(n_499),
.Y(n_616)
);

AND2x4_ASAP7_75t_L g617 ( 
.A(n_441),
.B(n_394),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_449),
.Y(n_618)
);

NAND2xp33_ASAP7_75t_R g619 ( 
.A(n_501),
.B(n_238),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_504),
.Y(n_620)
);

CKINVDCx5p33_ASAP7_75t_R g621 ( 
.A(n_505),
.Y(n_621)
);

AND2x2_ASAP7_75t_L g622 ( 
.A(n_462),
.B(n_492),
.Y(n_622)
);

BUFx6f_ASAP7_75t_L g623 ( 
.A(n_449),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_460),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_513),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_515),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_461),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_461),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_522),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_469),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_530),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_531),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_469),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_532),
.B(n_534),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_470),
.Y(n_635)
);

CKINVDCx5p33_ASAP7_75t_R g636 ( 
.A(n_542),
.Y(n_636)
);

INVxp33_ASAP7_75t_SL g637 ( 
.A(n_442),
.Y(n_637)
);

AND2x4_ASAP7_75t_L g638 ( 
.A(n_470),
.B(n_395),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_552),
.Y(n_639)
);

INVx6_ASAP7_75t_L g640 ( 
.A(n_467),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_538),
.B(n_234),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_545),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_R g643 ( 
.A(n_546),
.B(n_377),
.Y(n_643)
);

CKINVDCx5p33_ASAP7_75t_R g644 ( 
.A(n_549),
.Y(n_644)
);

BUFx8_ASAP7_75t_L g645 ( 
.A(n_483),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_476),
.Y(n_646)
);

INVx2_ASAP7_75t_L g647 ( 
.A(n_476),
.Y(n_647)
);

CKINVDCx5p33_ASAP7_75t_R g648 ( 
.A(n_512),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

INVx3_ASAP7_75t_L g650 ( 
.A(n_477),
.Y(n_650)
);

INVx1_ASAP7_75t_SL g651 ( 
.A(n_577),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_600),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_622),
.B(n_493),
.Y(n_653)
);

NAND2xp33_ASAP7_75t_L g654 ( 
.A(n_603),
.B(n_326),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_611),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_571),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_582),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_L g658 ( 
.A(n_582),
.B(n_438),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_600),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_594),
.B(n_493),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_602),
.Y(n_661)
);

AND2x4_ASAP7_75t_L g662 ( 
.A(n_582),
.B(n_552),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g663 ( 
.A(n_622),
.B(n_507),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_573),
.B(n_507),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_606),
.B(n_478),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_586),
.B(n_478),
.Y(n_666)
);

INVx4_ASAP7_75t_L g667 ( 
.A(n_611),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_577),
.B(n_508),
.Y(n_668)
);

INVx1_ASAP7_75t_SL g669 ( 
.A(n_604),
.Y(n_669)
);

INVx2_ASAP7_75t_SL g670 ( 
.A(n_598),
.Y(n_670)
);

AND2x6_ASAP7_75t_L g671 ( 
.A(n_617),
.B(n_233),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_628),
.Y(n_672)
);

AND2x4_ASAP7_75t_L g673 ( 
.A(n_617),
.B(n_553),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_633),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_591),
.B(n_508),
.Y(n_675)
);

OR2x6_ASAP7_75t_L g676 ( 
.A(n_616),
.B(n_451),
.Y(n_676)
);

INVx4_ASAP7_75t_L g677 ( 
.A(n_611),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_617),
.B(n_481),
.Y(n_678)
);

OAI21xp33_ASAP7_75t_SL g679 ( 
.A1(n_580),
.A2(n_486),
.B(n_471),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_646),
.B(n_481),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_L g681 ( 
.A(n_649),
.B(n_482),
.Y(n_681)
);

OR2x6_ASAP7_75t_L g682 ( 
.A(n_616),
.B(n_405),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_627),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_641),
.B(n_503),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_601),
.B(n_233),
.Y(n_685)
);

AOI22xp33_ASAP7_75t_L g686 ( 
.A1(n_638),
.A2(n_555),
.B1(n_536),
.B2(n_547),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_627),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_650),
.Y(n_688)
);

INVx5_ASAP7_75t_L g689 ( 
.A(n_611),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_611),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_627),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_650),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_585),
.B(n_467),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_650),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_602),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_598),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_613),
.Y(n_697)
);

BUFx6f_ASAP7_75t_L g698 ( 
.A(n_623),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_L g699 ( 
.A(n_572),
.B(n_484),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_R g700 ( 
.A(n_564),
.B(n_244),
.Y(n_700)
);

INVx2_ASAP7_75t_SL g701 ( 
.A(n_643),
.Y(n_701)
);

AOI22xp33_ASAP7_75t_L g702 ( 
.A1(n_638),
.A2(n_288),
.B1(n_293),
.B2(n_287),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_574),
.B(n_485),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_579),
.Y(n_704)
);

AND2x6_ASAP7_75t_L g705 ( 
.A(n_638),
.B(n_249),
.Y(n_705)
);

NAND2xp33_ASAP7_75t_SL g706 ( 
.A(n_619),
.B(n_315),
.Y(n_706)
);

CKINVDCx20_ASAP7_75t_R g707 ( 
.A(n_592),
.Y(n_707)
);

INVx3_ASAP7_75t_L g708 ( 
.A(n_623),
.Y(n_708)
);

OR2x2_ASAP7_75t_L g709 ( 
.A(n_561),
.B(n_509),
.Y(n_709)
);

INVx4_ASAP7_75t_SL g710 ( 
.A(n_640),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_608),
.B(n_495),
.Y(n_711)
);

INVx3_ASAP7_75t_L g712 ( 
.A(n_623),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_634),
.B(n_495),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_640),
.B(n_497),
.Y(n_714)
);

AND2x4_ASAP7_75t_L g715 ( 
.A(n_580),
.B(n_249),
.Y(n_715)
);

INVx5_ASAP7_75t_L g716 ( 
.A(n_635),
.Y(n_716)
);

AOI22xp5_ASAP7_75t_L g717 ( 
.A1(n_578),
.A2(n_609),
.B1(n_575),
.B2(n_620),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_583),
.B(n_406),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_613),
.Y(n_719)
);

INVx1_ASAP7_75t_SL g720 ( 
.A(n_565),
.Y(n_720)
);

AND3x2_ASAP7_75t_L g721 ( 
.A(n_626),
.B(n_293),
.C(n_288),
.Y(n_721)
);

AND2x4_ASAP7_75t_L g722 ( 
.A(n_610),
.B(n_253),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_639),
.B(n_553),
.Y(n_723)
);

AOI22xp5_ASAP7_75t_L g724 ( 
.A1(n_583),
.A2(n_483),
.B1(n_346),
.B2(n_400),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_640),
.B(n_497),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_L g726 ( 
.A(n_640),
.B(n_635),
.Y(n_726)
);

INVx6_ASAP7_75t_L g727 ( 
.A(n_567),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_639),
.A2(n_304),
.B1(n_306),
.B2(n_296),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_610),
.A2(n_304),
.B1(n_306),
.B2(n_296),
.Y(n_729)
);

NOR2xp33_ASAP7_75t_L g730 ( 
.A(n_562),
.B(n_467),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_579),
.Y(n_731)
);

NOR2xp33_ASAP7_75t_L g732 ( 
.A(n_569),
.B(n_467),
.Y(n_732)
);

INVx2_ASAP7_75t_L g733 ( 
.A(n_614),
.Y(n_733)
);

BUFx3_ASAP7_75t_L g734 ( 
.A(n_635),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_614),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_618),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_618),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_624),
.Y(n_738)
);

NOR2xp33_ASAP7_75t_L g739 ( 
.A(n_570),
.B(n_550),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_SL g740 ( 
.A(n_587),
.B(n_406),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_624),
.Y(n_741)
);

INVx4_ASAP7_75t_L g742 ( 
.A(n_635),
.Y(n_742)
);

NOR2xp33_ASAP7_75t_L g743 ( 
.A(n_576),
.B(n_558),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_630),
.Y(n_744)
);

INVx3_ASAP7_75t_L g745 ( 
.A(n_635),
.Y(n_745)
);

INVx4_ASAP7_75t_L g746 ( 
.A(n_593),
.Y(n_746)
);

INVx1_ASAP7_75t_L g747 ( 
.A(n_630),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_647),
.B(n_498),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_SL g749 ( 
.A(n_587),
.B(n_326),
.Y(n_749)
);

AOI22xp33_ASAP7_75t_L g750 ( 
.A1(n_647),
.A2(n_337),
.B1(n_344),
.B2(n_308),
.Y(n_750)
);

BUFx2_ASAP7_75t_L g751 ( 
.A(n_564),
.Y(n_751)
);

INVx1_ASAP7_75t_SL g752 ( 
.A(n_565),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_593),
.Y(n_753)
);

OR2x2_ASAP7_75t_L g754 ( 
.A(n_584),
.B(n_453),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_589),
.B(n_326),
.Y(n_755)
);

AO22x2_ASAP7_75t_L g756 ( 
.A1(n_563),
.A2(n_337),
.B1(n_344),
.B2(n_308),
.Y(n_756)
);

INVx2_ASAP7_75t_L g757 ( 
.A(n_560),
.Y(n_757)
);

AND2x4_ASAP7_75t_L g758 ( 
.A(n_588),
.B(n_314),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_SL g759 ( 
.A(n_589),
.B(n_326),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_560),
.Y(n_760)
);

BUFx2_ASAP7_75t_L g761 ( 
.A(n_648),
.Y(n_761)
);

OR2x6_ASAP7_75t_L g762 ( 
.A(n_563),
.B(n_297),
.Y(n_762)
);

NAND2xp5_ASAP7_75t_L g763 ( 
.A(n_593),
.B(n_498),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_593),
.Y(n_764)
);

BUFx2_ASAP7_75t_L g765 ( 
.A(n_648),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_590),
.B(n_253),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_593),
.Y(n_767)
);

INVx4_ASAP7_75t_L g768 ( 
.A(n_590),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_595),
.Y(n_769)
);

INVx5_ASAP7_75t_L g770 ( 
.A(n_567),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_595),
.B(n_596),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_596),
.B(n_502),
.Y(n_772)
);

INVx2_ASAP7_75t_L g773 ( 
.A(n_597),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_SL g774 ( 
.A(n_597),
.B(n_599),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_599),
.B(n_502),
.Y(n_775)
);

INVx2_ASAP7_75t_SL g776 ( 
.A(n_607),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_607),
.Y(n_777)
);

BUFx6f_ASAP7_75t_L g778 ( 
.A(n_612),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_612),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_621),
.Y(n_780)
);

INVx5_ASAP7_75t_L g781 ( 
.A(n_567),
.Y(n_781)
);

INVx3_ASAP7_75t_L g782 ( 
.A(n_621),
.Y(n_782)
);

OR2x2_ASAP7_75t_L g783 ( 
.A(n_625),
.B(n_459),
.Y(n_783)
);

INVx4_ASAP7_75t_SL g784 ( 
.A(n_645),
.Y(n_784)
);

BUFx6f_ASAP7_75t_L g785 ( 
.A(n_625),
.Y(n_785)
);

AOI22xp5_ASAP7_75t_L g786 ( 
.A1(n_629),
.A2(n_407),
.B1(n_430),
.B2(n_278),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_L g787 ( 
.A(n_629),
.B(n_506),
.Y(n_787)
);

INVx1_ASAP7_75t_L g788 ( 
.A(n_631),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_631),
.B(n_314),
.Y(n_789)
);

INVx4_ASAP7_75t_L g790 ( 
.A(n_632),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_632),
.Y(n_791)
);

INVx4_ASAP7_75t_L g792 ( 
.A(n_636),
.Y(n_792)
);

INVx1_ASAP7_75t_L g793 ( 
.A(n_636),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_642),
.B(n_506),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_642),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_644),
.Y(n_796)
);

BUFx3_ASAP7_75t_L g797 ( 
.A(n_644),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_L g798 ( 
.A(n_637),
.B(n_500),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_645),
.Y(n_799)
);

OR2x6_ASAP7_75t_L g800 ( 
.A(n_645),
.B(n_297),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_566),
.B(n_510),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_566),
.B(n_510),
.Y(n_802)
);

AND2x6_ASAP7_75t_L g803 ( 
.A(n_568),
.B(n_254),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_581),
.B(n_511),
.Y(n_804)
);

BUFx6f_ASAP7_75t_SL g805 ( 
.A(n_778),
.Y(n_805)
);

INVx2_ASAP7_75t_SL g806 ( 
.A(n_709),
.Y(n_806)
);

AOI22xp33_ASAP7_75t_L g807 ( 
.A1(n_715),
.A2(n_363),
.B1(n_364),
.B2(n_354),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_SL g808 ( 
.A(n_703),
.B(n_379),
.Y(n_808)
);

NOR2xp33_ASAP7_75t_L g809 ( 
.A(n_684),
.B(n_243),
.Y(n_809)
);

INVx3_ASAP7_75t_L g810 ( 
.A(n_657),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_657),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_723),
.Y(n_812)
);

AOI22xp5_ASAP7_75t_L g813 ( 
.A1(n_664),
.A2(n_389),
.B1(n_396),
.B2(n_384),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_772),
.B(n_274),
.Y(n_814)
);

AND2x6_ASAP7_75t_L g815 ( 
.A(n_715),
.B(n_262),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_723),
.Y(n_816)
);

OR2x2_ASAP7_75t_L g817 ( 
.A(n_670),
.B(n_581),
.Y(n_817)
);

OR2x2_ASAP7_75t_L g818 ( 
.A(n_696),
.B(n_368),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_775),
.B(n_397),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_SL g820 ( 
.A(n_787),
.B(n_398),
.Y(n_820)
);

NOR2xp67_ASAP7_75t_L g821 ( 
.A(n_701),
.B(n_521),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_L g822 ( 
.A(n_794),
.B(n_393),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_673),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_711),
.B(n_262),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_713),
.B(n_265),
.Y(n_825)
);

O2A1O1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_665),
.A2(n_533),
.B(n_543),
.C(n_523),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_801),
.B(n_247),
.Y(n_827)
);

AND2x2_ASAP7_75t_L g828 ( 
.A(n_653),
.B(n_557),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_673),
.Y(n_829)
);

OAI22xp5_ASAP7_75t_L g830 ( 
.A1(n_686),
.A2(n_311),
.B1(n_307),
.B2(n_305),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_SL g831 ( 
.A(n_662),
.B(n_409),
.Y(n_831)
);

NOR2xp33_ASAP7_75t_L g832 ( 
.A(n_802),
.B(n_248),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_662),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_652),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_678),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_804),
.B(n_658),
.Y(n_836)
);

BUFx5_ASAP7_75t_L g837 ( 
.A(n_705),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_666),
.B(n_265),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_SL g839 ( 
.A(n_664),
.B(n_412),
.Y(n_839)
);

AND2x2_ASAP7_75t_L g840 ( 
.A(n_663),
.B(n_605),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_672),
.B(n_272),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_660),
.B(n_418),
.Y(n_842)
);

INVx1_ASAP7_75t_L g843 ( 
.A(n_757),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_660),
.B(n_256),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_659),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_783),
.B(n_424),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_671),
.A2(n_421),
.B1(n_403),
.B2(n_324),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_679),
.A2(n_511),
.B(n_514),
.C(n_516),
.Y(n_848)
);

AOI22xp33_ASAP7_75t_L g849 ( 
.A1(n_715),
.A2(n_354),
.B1(n_386),
.B2(n_382),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_674),
.B(n_283),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_757),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_766),
.B(n_257),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_686),
.A2(n_717),
.B1(n_729),
.B2(n_786),
.Y(n_853)
);

AND2x4_ASAP7_75t_L g854 ( 
.A(n_758),
.B(n_338),
.Y(n_854)
);

AOI21xp33_ASAP7_75t_L g855 ( 
.A1(n_766),
.A2(n_305),
.B(n_299),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_722),
.Y(n_856)
);

INVx3_ASAP7_75t_L g857 ( 
.A(n_722),
.Y(n_857)
);

AOI22xp33_ASAP7_75t_L g858 ( 
.A1(n_722),
.A2(n_390),
.B1(n_386),
.B2(n_382),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_760),
.Y(n_859)
);

NOR2xp33_ASAP7_75t_L g860 ( 
.A(n_718),
.B(n_258),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_699),
.B(n_299),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_683),
.B(n_307),
.Y(n_862)
);

BUFx12f_ASAP7_75t_L g863 ( 
.A(n_778),
.Y(n_863)
);

O2A1O1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_718),
.A2(n_740),
.B(n_755),
.C(n_749),
.Y(n_864)
);

BUFx6f_ASAP7_75t_SL g865 ( 
.A(n_778),
.Y(n_865)
);

O2A1O1Ixp5_ASAP7_75t_L g866 ( 
.A1(n_687),
.A2(n_381),
.B(n_311),
.C(n_324),
.Y(n_866)
);

AND2x4_ASAP7_75t_L g867 ( 
.A(n_758),
.B(n_338),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_659),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_661),
.Y(n_869)
);

INVx2_ASAP7_75t_SL g870 ( 
.A(n_789),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_740),
.B(n_259),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_L g872 ( 
.A1(n_702),
.A2(n_364),
.B1(n_390),
.B2(n_422),
.Y(n_872)
);

BUFx6f_ASAP7_75t_L g873 ( 
.A(n_690),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_661),
.Y(n_874)
);

A2O1A1Ixp33_ASAP7_75t_L g875 ( 
.A1(n_739),
.A2(n_514),
.B(n_516),
.C(n_349),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_714),
.B(n_333),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_725),
.B(n_333),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_SL g878 ( 
.A(n_688),
.B(n_339),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_760),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_SL g880 ( 
.A(n_693),
.B(n_373),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_749),
.B(n_260),
.Y(n_881)
);

NOR2xp33_ASAP7_75t_L g882 ( 
.A(n_755),
.B(n_267),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_691),
.B(n_339),
.Y(n_883)
);

AND2x2_ASAP7_75t_L g884 ( 
.A(n_739),
.B(n_615),
.Y(n_884)
);

A2O1A1Ixp33_ASAP7_75t_L g885 ( 
.A1(n_743),
.A2(n_403),
.B(n_348),
.C(n_349),
.Y(n_885)
);

NOR2xp33_ASAP7_75t_L g886 ( 
.A(n_759),
.B(n_798),
.Y(n_886)
);

AND2x2_ASAP7_75t_L g887 ( 
.A(n_743),
.B(n_551),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_692),
.B(n_343),
.Y(n_888)
);

BUFx3_ASAP7_75t_L g889 ( 
.A(n_656),
.Y(n_889)
);

CKINVDCx5p33_ASAP7_75t_R g890 ( 
.A(n_707),
.Y(n_890)
);

NAND2xp5_ASAP7_75t_SL g891 ( 
.A(n_694),
.B(n_343),
.Y(n_891)
);

AND2x2_ASAP7_75t_L g892 ( 
.A(n_651),
.B(n_535),
.Y(n_892)
);

O2A1O1Ixp33_ASAP7_75t_L g893 ( 
.A1(n_759),
.A2(n_378),
.B(n_422),
.C(n_416),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_767),
.B(n_353),
.Y(n_894)
);

AOI22xp33_ASAP7_75t_L g895 ( 
.A1(n_702),
.A2(n_378),
.B1(n_380),
.B2(n_367),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_767),
.B(n_353),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_693),
.B(n_373),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_671),
.B(n_381),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_671),
.B(n_432),
.Y(n_899)
);

OR2x2_ASAP7_75t_L g900 ( 
.A(n_754),
.B(n_435),
.Y(n_900)
);

NOR2xp33_ASAP7_75t_L g901 ( 
.A(n_798),
.B(n_675),
.Y(n_901)
);

NOR3xp33_ASAP7_75t_L g902 ( 
.A(n_706),
.B(n_277),
.C(n_273),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_704),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_675),
.B(n_279),
.Y(n_904)
);

BUFx3_ASAP7_75t_L g905 ( 
.A(n_707),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_668),
.B(n_535),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_671),
.B(n_432),
.Y(n_907)
);

BUFx3_ASAP7_75t_L g908 ( 
.A(n_778),
.Y(n_908)
);

AND2x4_ASAP7_75t_L g909 ( 
.A(n_685),
.B(n_435),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_SL g910 ( 
.A(n_785),
.B(n_425),
.Y(n_910)
);

INVx2_ASAP7_75t_L g911 ( 
.A(n_695),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_671),
.B(n_421),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_SL g913 ( 
.A(n_785),
.B(n_425),
.Y(n_913)
);

BUFx5_ASAP7_75t_L g914 ( 
.A(n_705),
.Y(n_914)
);

INVx8_ASAP7_75t_L g915 ( 
.A(n_770),
.Y(n_915)
);

AND2x2_ASAP7_75t_L g916 ( 
.A(n_782),
.B(n_551),
.Y(n_916)
);

NOR2xp33_ASAP7_75t_L g917 ( 
.A(n_724),
.B(n_282),
.Y(n_917)
);

BUFx6f_ASAP7_75t_L g918 ( 
.A(n_690),
.Y(n_918)
);

A2O1A1Ixp33_ASAP7_75t_L g919 ( 
.A1(n_729),
.A2(n_363),
.B(n_380),
.C(n_367),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_704),
.Y(n_920)
);

INVx4_ASAP7_75t_L g921 ( 
.A(n_690),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_697),
.B(n_286),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_SL g923 ( 
.A(n_719),
.B(n_290),
.Y(n_923)
);

INVx2_ASAP7_75t_SL g924 ( 
.A(n_685),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_700),
.Y(n_925)
);

AOI22xp33_ASAP7_75t_L g926 ( 
.A1(n_728),
.A2(n_361),
.B1(n_387),
.B2(n_410),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_735),
.B(n_736),
.Y(n_927)
);

NAND2xp5_ASAP7_75t_SL g928 ( 
.A(n_738),
.B(n_294),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_695),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_782),
.B(n_537),
.Y(n_930)
);

BUFx3_ASAP7_75t_L g931 ( 
.A(n_761),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_741),
.B(n_298),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_733),
.Y(n_933)
);

AOI22xp33_ASAP7_75t_L g934 ( 
.A1(n_728),
.A2(n_423),
.B1(n_437),
.B2(n_300),
.Y(n_934)
);

NAND2xp5_ASAP7_75t_L g935 ( 
.A(n_747),
.B(n_301),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_731),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_731),
.Y(n_937)
);

INVx5_ASAP7_75t_L g938 ( 
.A(n_705),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_682),
.B(n_730),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_SL g940 ( 
.A(n_773),
.B(n_302),
.Y(n_940)
);

OR2x2_ASAP7_75t_L g941 ( 
.A(n_669),
.B(n_309),
.Y(n_941)
);

OR2x6_ASAP7_75t_L g942 ( 
.A(n_727),
.B(n_537),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_SL g943 ( 
.A(n_773),
.B(n_310),
.Y(n_943)
);

AOI22xp33_ASAP7_75t_L g944 ( 
.A1(n_750),
.A2(n_388),
.B1(n_317),
.B2(n_319),
.Y(n_944)
);

INVx4_ASAP7_75t_L g945 ( 
.A(n_690),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_726),
.A2(n_548),
.B(n_541),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_698),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_730),
.B(n_316),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_SL g949 ( 
.A(n_791),
.B(n_325),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_765),
.Y(n_950)
);

AOI22xp5_ASAP7_75t_L g951 ( 
.A1(n_803),
.A2(n_402),
.B1(n_332),
.B2(n_341),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_732),
.B(n_655),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_682),
.B(n_329),
.Y(n_953)
);

INVx8_ASAP7_75t_L g954 ( 
.A(n_770),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_732),
.B(n_345),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_SL g956 ( 
.A(n_791),
.B(n_350),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_655),
.B(n_351),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_685),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_733),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_708),
.B(n_352),
.Y(n_960)
);

NOR2xp33_ASAP7_75t_L g961 ( 
.A(n_682),
.B(n_369),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_737),
.B(n_371),
.Y(n_962)
);

NAND2xp5_ASAP7_75t_L g963 ( 
.A(n_708),
.B(n_374),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_737),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_857),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_857),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_836),
.B(n_803),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_856),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_856),
.B(n_795),
.Y(n_969)
);

NAND2xp5_ASAP7_75t_L g970 ( 
.A(n_836),
.B(n_803),
.Y(n_970)
);

HB1xp67_ASAP7_75t_L g971 ( 
.A(n_908),
.Y(n_971)
);

NOR2xp33_ASAP7_75t_L g972 ( 
.A(n_901),
.B(n_795),
.Y(n_972)
);

OAI321xp33_ASAP7_75t_L g973 ( 
.A1(n_830),
.A2(n_676),
.A3(n_750),
.B1(n_769),
.B2(n_793),
.C(n_788),
.Y(n_973)
);

A2O1A1Ixp33_ASAP7_75t_L g974 ( 
.A1(n_886),
.A2(n_706),
.B(n_796),
.C(n_771),
.Y(n_974)
);

OAI21xp5_ASAP7_75t_L g975 ( 
.A1(n_848),
.A2(n_681),
.B(n_680),
.Y(n_975)
);

OAI21xp5_ASAP7_75t_L g976 ( 
.A1(n_835),
.A2(n_748),
.B(n_763),
.Y(n_976)
);

O2A1O1Ixp5_ASAP7_75t_L g977 ( 
.A1(n_886),
.A2(n_796),
.B(n_745),
.C(n_712),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_901),
.B(n_768),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_L g979 ( 
.A1(n_853),
.A2(n_654),
.B(n_774),
.C(n_676),
.Y(n_979)
);

NAND2xp5_ASAP7_75t_L g980 ( 
.A(n_814),
.B(n_822),
.Y(n_980)
);

AND2x2_ASAP7_75t_L g981 ( 
.A(n_809),
.B(n_797),
.Y(n_981)
);

A2O1A1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_864),
.A2(n_771),
.B(n_780),
.C(n_777),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_856),
.A2(n_677),
.B(n_667),
.Y(n_983)
);

INVx2_ASAP7_75t_L g984 ( 
.A(n_843),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_851),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_856),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_806),
.Y(n_987)
);

NAND2xp5_ASAP7_75t_L g988 ( 
.A(n_814),
.B(n_803),
.Y(n_988)
);

AOI21xp5_ASAP7_75t_L g989 ( 
.A1(n_938),
.A2(n_742),
.B(n_734),
.Y(n_989)
);

INVx2_ASAP7_75t_SL g990 ( 
.A(n_892),
.Y(n_990)
);

AOI22xp5_ASAP7_75t_L g991 ( 
.A1(n_822),
.A2(n_803),
.B1(n_700),
.B2(n_705),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_827),
.B(n_832),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_L g993 ( 
.A(n_827),
.B(n_705),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_810),
.Y(n_994)
);

BUFx12f_ASAP7_75t_L g995 ( 
.A(n_863),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_921),
.A2(n_742),
.B(n_734),
.Y(n_996)
);

NOR2xp33_ASAP7_75t_L g997 ( 
.A(n_809),
.B(n_768),
.Y(n_997)
);

AOI21xp5_ASAP7_75t_L g998 ( 
.A1(n_921),
.A2(n_945),
.B(n_912),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_873),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_828),
.B(n_790),
.Y(n_1000)
);

NAND3xp33_ASAP7_75t_SL g1001 ( 
.A(n_934),
.B(n_720),
.C(n_752),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_837),
.B(n_790),
.Y(n_1002)
);

AND2x2_ASAP7_75t_L g1003 ( 
.A(n_906),
.B(n_797),
.Y(n_1003)
);

NOR2x1_ASAP7_75t_L g1004 ( 
.A(n_821),
.B(n_792),
.Y(n_1004)
);

OAI321xp33_ASAP7_75t_L g1005 ( 
.A1(n_852),
.A2(n_779),
.A3(n_800),
.B1(n_774),
.B2(n_799),
.C(n_776),
.Y(n_1005)
);

HB1xp67_ASAP7_75t_L g1006 ( 
.A(n_854),
.Y(n_1006)
);

CKINVDCx10_ASAP7_75t_R g1007 ( 
.A(n_805),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_832),
.B(n_744),
.Y(n_1008)
);

AO21x1_ASAP7_75t_L g1009 ( 
.A1(n_881),
.A2(n_654),
.B(n_764),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_810),
.Y(n_1010)
);

AOI22xp5_ASAP7_75t_L g1011 ( 
.A1(n_844),
.A2(n_792),
.B1(n_751),
.B2(n_712),
.Y(n_1011)
);

AO22x1_ASAP7_75t_L g1012 ( 
.A1(n_917),
.A2(n_781),
.B1(n_375),
.B2(n_428),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_916),
.B(n_756),
.Y(n_1013)
);

NOR2x1_ASAP7_75t_L g1014 ( 
.A(n_884),
.B(n_800),
.Y(n_1014)
);

AO32x2_ASAP7_75t_L g1015 ( 
.A1(n_924),
.A2(n_756),
.A3(n_746),
.B1(n_762),
.B2(n_721),
.Y(n_1015)
);

AOI21xp5_ASAP7_75t_L g1016 ( 
.A1(n_952),
.A2(n_698),
.B(n_689),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_859),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_879),
.Y(n_1018)
);

NOR3xp33_ASAP7_75t_L g1019 ( 
.A(n_852),
.B(n_433),
.C(n_385),
.Y(n_1019)
);

OAI22xp5_ASAP7_75t_L g1020 ( 
.A1(n_958),
.A2(n_849),
.B1(n_858),
.B2(n_807),
.Y(n_1020)
);

NOR3xp33_ASAP7_75t_L g1021 ( 
.A(n_917),
.B(n_434),
.C(n_391),
.Y(n_1021)
);

AOI22xp33_ASAP7_75t_SL g1022 ( 
.A1(n_925),
.A2(n_727),
.B1(n_781),
.B2(n_800),
.Y(n_1022)
);

NOR2x1_ASAP7_75t_L g1023 ( 
.A(n_942),
.B(n_762),
.Y(n_1023)
);

A2O1A1Ixp33_ASAP7_75t_L g1024 ( 
.A1(n_855),
.A2(n_383),
.B(n_401),
.C(n_408),
.Y(n_1024)
);

AOI21x1_ASAP7_75t_L g1025 ( 
.A1(n_876),
.A2(n_877),
.B(n_838),
.Y(n_1025)
);

O2A1O1Ixp33_ASAP7_75t_L g1026 ( 
.A1(n_919),
.A2(n_762),
.B(n_548),
.C(n_541),
.Y(n_1026)
);

NAND2xp5_ASAP7_75t_SL g1027 ( 
.A(n_837),
.B(n_710),
.Y(n_1027)
);

OAI21x1_ASAP7_75t_L g1028 ( 
.A1(n_933),
.A2(n_540),
.B(n_710),
.Y(n_1028)
);

NAND2xp5_ASAP7_75t_L g1029 ( 
.A(n_930),
.B(n_756),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_887),
.B(n_844),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_873),
.A2(n_947),
.B(n_918),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_918),
.A2(n_716),
.B(n_753),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_904),
.B(n_710),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_904),
.B(n_753),
.Y(n_1034)
);

AOI21x1_ASAP7_75t_L g1035 ( 
.A1(n_876),
.A2(n_540),
.B(n_753),
.Y(n_1035)
);

AOI21x1_ASAP7_75t_L g1036 ( 
.A1(n_877),
.A2(n_753),
.B(n_716),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_818),
.B(n_721),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_918),
.A2(n_781),
.B(n_411),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_918),
.A2(n_781),
.B(n_414),
.Y(n_1039)
);

AOI22xp5_ASAP7_75t_L g1040 ( 
.A1(n_939),
.A2(n_727),
.B1(n_784),
.B2(n_436),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_824),
.B(n_417),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_825),
.B(n_419),
.Y(n_1042)
);

AOI22xp5_ASAP7_75t_L g1043 ( 
.A1(n_939),
.A2(n_784),
.B1(n_431),
.B2(n_427),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_948),
.B(n_420),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_955),
.B(n_881),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_947),
.A2(n_426),
.B(n_161),
.Y(n_1046)
);

AOI22x1_ASAP7_75t_L g1047 ( 
.A1(n_811),
.A2(n_784),
.B1(n_221),
.B2(n_219),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_882),
.B(n_12),
.Y(n_1048)
);

AND2x2_ASAP7_75t_L g1049 ( 
.A(n_926),
.B(n_17),
.Y(n_1049)
);

INVx3_ASAP7_75t_L g1050 ( 
.A(n_947),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_903),
.Y(n_1051)
);

NOR2xp33_ASAP7_75t_L g1052 ( 
.A(n_860),
.B(n_17),
.Y(n_1052)
);

AO21x1_ASAP7_75t_L g1053 ( 
.A1(n_882),
.A2(n_19),
.B(n_21),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_947),
.A2(n_210),
.B(n_207),
.Y(n_1054)
);

INVxp67_ASAP7_75t_SL g1055 ( 
.A(n_833),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_808),
.B(n_19),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_894),
.A2(n_200),
.B(n_193),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_808),
.B(n_22),
.Y(n_1058)
);

NAND3xp33_ASAP7_75t_SL g1059 ( 
.A(n_934),
.B(n_24),
.C(n_25),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_L g1060 ( 
.A(n_860),
.B(n_31),
.Y(n_1060)
);

AOI22xp33_ASAP7_75t_L g1061 ( 
.A1(n_872),
.A2(n_32),
.B1(n_35),
.B2(n_36),
.Y(n_1061)
);

A2O1A1Ixp33_ASAP7_75t_L g1062 ( 
.A1(n_872),
.A2(n_35),
.B(n_36),
.C(n_39),
.Y(n_1062)
);

OAI22xp5_ASAP7_75t_L g1063 ( 
.A1(n_807),
.A2(n_192),
.B1(n_190),
.B2(n_188),
.Y(n_1063)
);

NOR2xp33_ASAP7_75t_L g1064 ( 
.A(n_871),
.B(n_40),
.Y(n_1064)
);

INVx4_ASAP7_75t_L g1065 ( 
.A(n_805),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_L g1066 ( 
.A(n_871),
.B(n_40),
.C(n_41),
.Y(n_1066)
);

INVxp67_ASAP7_75t_SL g1067 ( 
.A(n_823),
.Y(n_1067)
);

AOI21xp5_ASAP7_75t_L g1068 ( 
.A1(n_896),
.A2(n_187),
.B(n_183),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_815),
.A2(n_812),
.B1(n_816),
.B2(n_829),
.Y(n_1069)
);

NOR2xp33_ASAP7_75t_L g1070 ( 
.A(n_900),
.B(n_43),
.Y(n_1070)
);

INVx4_ASAP7_75t_L g1071 ( 
.A(n_865),
.Y(n_1071)
);

AND2x4_ASAP7_75t_L g1072 ( 
.A(n_870),
.B(n_137),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_SL g1073 ( 
.A(n_837),
.B(n_179),
.Y(n_1073)
);

NOR2xp33_ASAP7_75t_L g1074 ( 
.A(n_941),
.B(n_50),
.Y(n_1074)
);

AOI21xp5_ASAP7_75t_L g1075 ( 
.A1(n_927),
.A2(n_173),
.B(n_167),
.Y(n_1075)
);

INVx2_ASAP7_75t_L g1076 ( 
.A(n_834),
.Y(n_1076)
);

BUFx6f_ASAP7_75t_L g1077 ( 
.A(n_915),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_861),
.B(n_50),
.Y(n_1078)
);

AOI22xp5_ASAP7_75t_L g1079 ( 
.A1(n_815),
.A2(n_164),
.B1(n_157),
.B2(n_151),
.Y(n_1079)
);

A2O1A1Ixp33_ASAP7_75t_L g1080 ( 
.A1(n_895),
.A2(n_893),
.B(n_826),
.C(n_885),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_L g1081 ( 
.A(n_817),
.B(n_51),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_920),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_957),
.A2(n_148),
.B(n_138),
.Y(n_1083)
);

AOI22xp33_ASAP7_75t_L g1084 ( 
.A1(n_895),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_931),
.Y(n_1085)
);

CKINVDCx10_ASAP7_75t_R g1086 ( 
.A(n_865),
.Y(n_1086)
);

AOI21x1_ASAP7_75t_L g1087 ( 
.A1(n_936),
.A2(n_129),
.B(n_127),
.Y(n_1087)
);

INVx2_ASAP7_75t_L g1088 ( 
.A(n_845),
.Y(n_1088)
);

OAI22xp5_ASAP7_75t_L g1089 ( 
.A1(n_926),
.A2(n_126),
.B1(n_123),
.B2(n_118),
.Y(n_1089)
);

AOI21xp5_ASAP7_75t_L g1090 ( 
.A1(n_960),
.A2(n_117),
.B(n_116),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_937),
.Y(n_1091)
);

AOI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_963),
.A2(n_111),
.B(n_109),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_950),
.Y(n_1093)
);

INVx2_ASAP7_75t_L g1094 ( 
.A(n_868),
.Y(n_1094)
);

AND2x2_ASAP7_75t_L g1095 ( 
.A(n_840),
.B(n_52),
.Y(n_1095)
);

AND2x2_ASAP7_75t_SL g1096 ( 
.A(n_898),
.B(n_99),
.Y(n_1096)
);

A2O1A1Ixp33_ASAP7_75t_L g1097 ( 
.A1(n_951),
.A2(n_55),
.B(n_58),
.C(n_59),
.Y(n_1097)
);

NAND2x1p5_ASAP7_75t_L g1098 ( 
.A(n_959),
.B(n_60),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_964),
.Y(n_1099)
);

NOR3xp33_ASAP7_75t_L g1100 ( 
.A(n_910),
.B(n_60),
.C(n_61),
.Y(n_1100)
);

O2A1O1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_875),
.A2(n_891),
.B(n_878),
.C(n_962),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_819),
.B(n_62),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_869),
.Y(n_1103)
);

NOR2xp33_ASAP7_75t_L g1104 ( 
.A(n_839),
.B(n_63),
.Y(n_1104)
);

AOI22xp5_ASAP7_75t_L g1105 ( 
.A1(n_815),
.A2(n_63),
.B1(n_65),
.B2(n_68),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_820),
.B(n_70),
.Y(n_1106)
);

HB1xp67_ASAP7_75t_L g1107 ( 
.A(n_854),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_899),
.A2(n_71),
.B(n_75),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_907),
.A2(n_81),
.B(n_82),
.Y(n_1109)
);

AOI21xp5_ASAP7_75t_L g1110 ( 
.A1(n_831),
.A2(n_81),
.B(n_83),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_874),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_911),
.A2(n_83),
.B(n_85),
.Y(n_1112)
);

A2O1A1Ixp33_ASAP7_75t_L g1113 ( 
.A1(n_953),
.A2(n_88),
.B(n_961),
.C(n_944),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_929),
.Y(n_1114)
);

NOR2x1_ASAP7_75t_L g1115 ( 
.A(n_942),
.B(n_913),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_909),
.B(n_841),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_867),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_889),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_831),
.A2(n_932),
.B(n_922),
.Y(n_1119)
);

NAND2xp5_ASAP7_75t_L g1120 ( 
.A(n_909),
.B(n_850),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_935),
.A2(n_883),
.B(n_888),
.Y(n_1121)
);

NOR2xp33_ASAP7_75t_L g1122 ( 
.A(n_880),
.B(n_897),
.Y(n_1122)
);

CKINVDCx5p33_ASAP7_75t_R g1123 ( 
.A(n_890),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_815),
.B(n_862),
.Y(n_1124)
);

OAI21x1_ASAP7_75t_L g1125 ( 
.A1(n_946),
.A2(n_866),
.B(n_928),
.Y(n_1125)
);

AOI22xp33_ASAP7_75t_L g1126 ( 
.A1(n_815),
.A2(n_944),
.B1(n_902),
.B2(n_914),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_842),
.A2(n_923),
.B(n_846),
.Y(n_1127)
);

A2O1A1Ixp33_ASAP7_75t_L g1128 ( 
.A1(n_961),
.A2(n_867),
.B(n_847),
.C(n_813),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_940),
.B(n_956),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_943),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_949),
.Y(n_1131)
);

BUFx3_ASAP7_75t_L g1132 ( 
.A(n_905),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_837),
.A2(n_914),
.B(n_915),
.Y(n_1133)
);

O2A1O1Ixp5_ASAP7_75t_L g1134 ( 
.A1(n_837),
.A2(n_914),
.B(n_915),
.C(n_954),
.Y(n_1134)
);

O2A1O1Ixp33_ASAP7_75t_L g1135 ( 
.A1(n_942),
.A2(n_914),
.B(n_954),
.C(n_853),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_914),
.Y(n_1136)
);

OAI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_886),
.A2(n_853),
.B1(n_836),
.B2(n_857),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_836),
.B(n_835),
.Y(n_1138)
);

A2O1A1Ixp33_ASAP7_75t_L g1139 ( 
.A1(n_992),
.A2(n_980),
.B(n_1064),
.C(n_1052),
.Y(n_1139)
);

OAI21x1_ASAP7_75t_L g1140 ( 
.A1(n_1028),
.A2(n_1035),
.B(n_998),
.Y(n_1140)
);

NAND2xp5_ASAP7_75t_L g1141 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1141)
);

OAI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1137),
.A2(n_1064),
.B(n_1052),
.Y(n_1142)
);

NAND3xp33_ASAP7_75t_SL g1143 ( 
.A(n_997),
.B(n_1021),
.C(n_1113),
.Y(n_1143)
);

BUFx6f_ASAP7_75t_L g1144 ( 
.A(n_1077),
.Y(n_1144)
);

INVx2_ASAP7_75t_L g1145 ( 
.A(n_984),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_972),
.B(n_1045),
.Y(n_1146)
);

OAI21x1_ASAP7_75t_L g1147 ( 
.A1(n_1134),
.A2(n_1016),
.B(n_1133),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_993),
.A2(n_1136),
.B(n_1121),
.Y(n_1148)
);

OAI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_977),
.A2(n_975),
.B(n_972),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_978),
.B(n_1008),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_979),
.A2(n_1104),
.B(n_1060),
.C(n_1048),
.Y(n_1151)
);

AND2x4_ASAP7_75t_L g1152 ( 
.A(n_1006),
.B(n_1107),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_1018),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1104),
.A2(n_997),
.B(n_982),
.C(n_1113),
.Y(n_1154)
);

A2O1A1Ixp33_ASAP7_75t_L g1155 ( 
.A1(n_982),
.A2(n_978),
.B(n_1122),
.C(n_974),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1136),
.A2(n_1124),
.B(n_976),
.Y(n_1156)
);

AOI21x1_ASAP7_75t_L g1157 ( 
.A1(n_969),
.A2(n_1025),
.B(n_1119),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_987),
.Y(n_1158)
);

OAI21x1_ASAP7_75t_L g1159 ( 
.A1(n_996),
.A2(n_1031),
.B(n_1125),
.Y(n_1159)
);

CKINVDCx20_ASAP7_75t_R g1160 ( 
.A(n_1123),
.Y(n_1160)
);

AOI22xp5_ASAP7_75t_L g1161 ( 
.A1(n_1000),
.A2(n_1122),
.B1(n_981),
.B2(n_1003),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_989),
.A2(n_1032),
.B(n_983),
.Y(n_1162)
);

HB1xp67_ASAP7_75t_L g1163 ( 
.A(n_987),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_990),
.B(n_1000),
.Y(n_1164)
);

INVx1_ASAP7_75t_L g1165 ( 
.A(n_1018),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_974),
.A2(n_970),
.B(n_967),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1095),
.B(n_1049),
.Y(n_1167)
);

AND2x4_ASAP7_75t_L g1168 ( 
.A(n_1006),
.B(n_1107),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1013),
.A2(n_1029),
.B(n_988),
.Y(n_1169)
);

A2O1A1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_1074),
.A2(n_973),
.B(n_1127),
.C(n_1101),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1020),
.B(n_1116),
.Y(n_1171)
);

AOI21xp5_ASAP7_75t_L g1172 ( 
.A1(n_1033),
.A2(n_1135),
.B(n_1120),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1085),
.Y(n_1173)
);

OAI21xp5_ASAP7_75t_L g1174 ( 
.A1(n_1080),
.A2(n_1126),
.B(n_991),
.Y(n_1174)
);

NAND2xp5_ASAP7_75t_L g1175 ( 
.A(n_965),
.B(n_966),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1044),
.B(n_994),
.Y(n_1176)
);

BUFx6f_ASAP7_75t_L g1177 ( 
.A(n_1077),
.Y(n_1177)
);

HB1xp67_ASAP7_75t_L g1178 ( 
.A(n_1085),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_994),
.B(n_1010),
.Y(n_1179)
);

AOI22xp33_ASAP7_75t_L g1180 ( 
.A1(n_1059),
.A2(n_1089),
.B1(n_1019),
.B2(n_1056),
.Y(n_1180)
);

AND2x4_ASAP7_75t_L g1181 ( 
.A(n_1117),
.B(n_1055),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1027),
.A2(n_969),
.B(n_1073),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1027),
.A2(n_1073),
.B(n_1002),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1118),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_1002),
.A2(n_1128),
.B(n_1129),
.Y(n_1185)
);

AOI21xp5_ASAP7_75t_L g1186 ( 
.A1(n_1128),
.A2(n_1010),
.B(n_968),
.Y(n_1186)
);

O2A1O1Ixp5_ASAP7_75t_L g1187 ( 
.A1(n_1009),
.A2(n_1078),
.B(n_1057),
.C(n_1058),
.Y(n_1187)
);

CKINVDCx6p67_ASAP7_75t_R g1188 ( 
.A(n_1007),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1088),
.A2(n_1094),
.B(n_1087),
.Y(n_1189)
);

CKINVDCx20_ASAP7_75t_R g1190 ( 
.A(n_1118),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_L g1191 ( 
.A(n_985),
.B(n_1017),
.Y(n_1191)
);

AND2x4_ASAP7_75t_L g1192 ( 
.A(n_1117),
.B(n_1067),
.Y(n_1192)
);

INVx2_ASAP7_75t_SL g1193 ( 
.A(n_1093),
.Y(n_1193)
);

OAI21x1_ASAP7_75t_L g1194 ( 
.A1(n_1050),
.A2(n_1112),
.B(n_1082),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_986),
.A2(n_1126),
.B(n_999),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_999),
.Y(n_1196)
);

NAND2xp5_ASAP7_75t_L g1197 ( 
.A(n_1051),
.B(n_1091),
.Y(n_1197)
);

OAI22x1_ASAP7_75t_L g1198 ( 
.A1(n_1081),
.A2(n_1037),
.B1(n_1070),
.B2(n_1065),
.Y(n_1198)
);

INVx3_ASAP7_75t_L g1199 ( 
.A(n_999),
.Y(n_1199)
);

NAND3xp33_ASAP7_75t_L g1200 ( 
.A(n_1100),
.B(n_1070),
.C(n_1037),
.Y(n_1200)
);

AOI21xp5_ASAP7_75t_SL g1201 ( 
.A1(n_1077),
.A2(n_1063),
.B(n_1080),
.Y(n_1201)
);

A2O1A1Ixp33_ASAP7_75t_L g1202 ( 
.A1(n_1081),
.A2(n_1131),
.B(n_1130),
.C(n_1110),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1099),
.B(n_1041),
.Y(n_1203)
);

OA21x2_ASAP7_75t_L g1204 ( 
.A1(n_1103),
.A2(n_1102),
.B(n_1106),
.Y(n_1204)
);

INVx2_ASAP7_75t_L g1205 ( 
.A(n_1076),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1111),
.Y(n_1206)
);

OR2x2_ASAP7_75t_L g1207 ( 
.A(n_1001),
.B(n_1132),
.Y(n_1207)
);

NAND2xp5_ASAP7_75t_L g1208 ( 
.A(n_1042),
.B(n_1114),
.Y(n_1208)
);

AO31x2_ASAP7_75t_L g1209 ( 
.A1(n_1053),
.A2(n_1097),
.A3(n_1024),
.B(n_1062),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_971),
.B(n_1004),
.Y(n_1210)
);

OAI22xp5_ASAP7_75t_L g1211 ( 
.A1(n_1061),
.A2(n_1084),
.B1(n_1096),
.B2(n_1097),
.Y(n_1211)
);

BUFx6f_ASAP7_75t_SL g1212 ( 
.A(n_1065),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_971),
.B(n_1132),
.Y(n_1213)
);

BUFx2_ASAP7_75t_L g1214 ( 
.A(n_995),
.Y(n_1214)
);

AND2x4_ASAP7_75t_L g1215 ( 
.A(n_1115),
.B(n_1072),
.Y(n_1215)
);

OAI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_1069),
.A2(n_1026),
.B(n_1096),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1072),
.A2(n_1023),
.B(n_1083),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1024),
.A2(n_1109),
.A3(n_1108),
.B(n_1092),
.Y(n_1218)
);

AOI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1066),
.A2(n_1005),
.B(n_1105),
.Y(n_1219)
);

HB1xp67_ASAP7_75t_L g1220 ( 
.A(n_1071),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1011),
.A2(n_1079),
.B1(n_1022),
.B2(n_1098),
.Y(n_1221)
);

OAI22xp5_ASAP7_75t_L g1222 ( 
.A1(n_1098),
.A2(n_1043),
.B1(n_1040),
.B2(n_1014),
.Y(n_1222)
);

OAI21xp33_ASAP7_75t_L g1223 ( 
.A1(n_1038),
.A2(n_1039),
.B(n_1046),
.Y(n_1223)
);

INVx8_ASAP7_75t_L g1224 ( 
.A(n_1077),
.Y(n_1224)
);

AOI21xp5_ASAP7_75t_L g1225 ( 
.A1(n_1090),
.A2(n_1075),
.B(n_1068),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1054),
.A2(n_1047),
.B(n_1012),
.Y(n_1226)
);

BUFx6f_ASAP7_75t_L g1227 ( 
.A(n_1071),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_SL g1228 ( 
.A1(n_1015),
.A2(n_1135),
.B(n_1119),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1015),
.A2(n_1028),
.B(n_1036),
.Y(n_1229)
);

NAND2x1p5_ASAP7_75t_L g1230 ( 
.A(n_1086),
.B(n_1015),
.Y(n_1230)
);

AOI21xp5_ASAP7_75t_L g1231 ( 
.A1(n_1034),
.A2(n_857),
.B(n_856),
.Y(n_1231)
);

AOI21xp33_ASAP7_75t_L g1232 ( 
.A1(n_980),
.A2(n_992),
.B(n_1052),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_1085),
.Y(n_1233)
);

OAI21x1_ASAP7_75t_L g1234 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_1035),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_984),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_984),
.Y(n_1236)
);

A2O1A1Ixp33_ASAP7_75t_L g1237 ( 
.A1(n_992),
.A2(n_980),
.B(n_1064),
.C(n_1052),
.Y(n_1237)
);

NAND2x1p5_ASAP7_75t_L g1238 ( 
.A(n_1077),
.B(n_856),
.Y(n_1238)
);

BUFx6f_ASAP7_75t_L g1239 ( 
.A(n_1077),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1137),
.A2(n_848),
.B(n_679),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_SL g1241 ( 
.A1(n_1135),
.A2(n_1137),
.B(n_856),
.Y(n_1241)
);

NAND2xp5_ASAP7_75t_SL g1242 ( 
.A(n_1000),
.B(n_778),
.Y(n_1242)
);

OAI21x1_ASAP7_75t_L g1243 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_1035),
.Y(n_1243)
);

OAI21xp5_ASAP7_75t_L g1244 ( 
.A1(n_1137),
.A2(n_848),
.B(n_679),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_984),
.Y(n_1245)
);

AOI21x1_ASAP7_75t_SL g1246 ( 
.A1(n_1060),
.A2(n_1048),
.B(n_988),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_992),
.A2(n_980),
.B(n_1064),
.C(n_1052),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_999),
.Y(n_1248)
);

AO31x2_ASAP7_75t_L g1249 ( 
.A1(n_1009),
.A2(n_848),
.A3(n_1137),
.B(n_1064),
.Y(n_1249)
);

AND2x4_ASAP7_75t_L g1250 ( 
.A(n_1006),
.B(n_908),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1251)
);

OAI22xp5_ASAP7_75t_L g1252 ( 
.A1(n_1138),
.A2(n_980),
.B1(n_992),
.B2(n_1061),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_984),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1137),
.A2(n_848),
.B(n_679),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1255)
);

OAI22x1_ASAP7_75t_L g1256 ( 
.A1(n_1049),
.A2(n_901),
.B1(n_886),
.B2(n_980),
.Y(n_1256)
);

NAND2xp5_ASAP7_75t_SL g1257 ( 
.A(n_1000),
.B(n_778),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1138),
.A2(n_980),
.B1(n_992),
.B2(n_1061),
.Y(n_1258)
);

AOI21xp5_ASAP7_75t_L g1259 ( 
.A1(n_1034),
.A2(n_857),
.B(n_856),
.Y(n_1259)
);

OAI21x1_ASAP7_75t_L g1260 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_1035),
.Y(n_1260)
);

INVx2_ASAP7_75t_L g1261 ( 
.A(n_984),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1262)
);

INVx5_ASAP7_75t_L g1263 ( 
.A(n_999),
.Y(n_1263)
);

INVx4_ASAP7_75t_L g1264 ( 
.A(n_1077),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1265)
);

INVx2_ASAP7_75t_L g1266 ( 
.A(n_984),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1009),
.A2(n_848),
.A3(n_1137),
.B(n_1064),
.Y(n_1269)
);

OAI21x1_ASAP7_75t_L g1270 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_1035),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_L g1271 ( 
.A1(n_1034),
.A2(n_857),
.B(n_856),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_L g1272 ( 
.A1(n_1137),
.A2(n_848),
.B(n_679),
.Y(n_1272)
);

NAND2xp5_ASAP7_75t_L g1273 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1273)
);

INVx4_ASAP7_75t_L g1274 ( 
.A(n_1077),
.Y(n_1274)
);

AOI221xp5_ASAP7_75t_SL g1275 ( 
.A1(n_980),
.A2(n_830),
.B1(n_853),
.B2(n_1064),
.C(n_1052),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_1035),
.Y(n_1276)
);

AOI21xp33_ASAP7_75t_L g1277 ( 
.A1(n_980),
.A2(n_992),
.B(n_1052),
.Y(n_1277)
);

OAI21x1_ASAP7_75t_L g1278 ( 
.A1(n_1028),
.A2(n_1036),
.B(n_1035),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_1077),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1009),
.A2(n_848),
.A3(n_1137),
.B(n_1064),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_992),
.A2(n_980),
.B(n_1064),
.C(n_1052),
.Y(n_1281)
);

AND2x4_ASAP7_75t_L g1282 ( 
.A(n_1006),
.B(n_908),
.Y(n_1282)
);

A2O1A1Ixp33_ASAP7_75t_L g1283 ( 
.A1(n_992),
.A2(n_980),
.B(n_1064),
.C(n_1052),
.Y(n_1283)
);

BUFx12f_ASAP7_75t_L g1284 ( 
.A(n_995),
.Y(n_1284)
);

NOR2xp33_ASAP7_75t_L g1285 ( 
.A(n_980),
.B(n_992),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_1138),
.B(n_1030),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1190),
.Y(n_1288)
);

OAI21xp33_ASAP7_75t_L g1289 ( 
.A1(n_1139),
.A2(n_1247),
.B(n_1237),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1224),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1145),
.Y(n_1291)
);

NAND2x1p5_ASAP7_75t_L g1292 ( 
.A(n_1263),
.B(n_1264),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1233),
.Y(n_1293)
);

AOI21xp5_ASAP7_75t_L g1294 ( 
.A1(n_1172),
.A2(n_1156),
.B(n_1174),
.Y(n_1294)
);

AOI22xp33_ASAP7_75t_L g1295 ( 
.A1(n_1211),
.A2(n_1142),
.B1(n_1277),
.B2(n_1232),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1263),
.Y(n_1296)
);

AOI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1174),
.A2(n_1185),
.B(n_1149),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_1160),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1141),
.B(n_1251),
.Y(n_1299)
);

INVxp67_ASAP7_75t_L g1300 ( 
.A(n_1163),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1251),
.B(n_1255),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1255),
.B(n_1262),
.Y(n_1302)
);

BUFx2_ASAP7_75t_L g1303 ( 
.A(n_1213),
.Y(n_1303)
);

OAI22xp5_ASAP7_75t_SL g1304 ( 
.A1(n_1200),
.A2(n_1184),
.B1(n_1180),
.B2(n_1142),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1149),
.A2(n_1225),
.B(n_1170),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1262),
.B(n_1265),
.Y(n_1306)
);

BUFx3_ASAP7_75t_L g1307 ( 
.A(n_1227),
.Y(n_1307)
);

AND2x2_ASAP7_75t_L g1308 ( 
.A(n_1167),
.B(n_1164),
.Y(n_1308)
);

AOI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1151),
.A2(n_1201),
.B(n_1281),
.Y(n_1309)
);

INVx3_ASAP7_75t_L g1310 ( 
.A(n_1224),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1265),
.B(n_1267),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1263),
.Y(n_1312)
);

INVx2_ASAP7_75t_SL g1313 ( 
.A(n_1178),
.Y(n_1313)
);

NAND2xp5_ASAP7_75t_L g1314 ( 
.A(n_1267),
.B(n_1268),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1268),
.B(n_1273),
.Y(n_1315)
);

BUFx3_ASAP7_75t_L g1316 ( 
.A(n_1227),
.Y(n_1316)
);

NAND2x1p5_ASAP7_75t_L g1317 ( 
.A(n_1263),
.B(n_1264),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1273),
.B(n_1286),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1283),
.A2(n_1146),
.B1(n_1286),
.B2(n_1161),
.Y(n_1319)
);

O2A1O1Ixp5_ASAP7_75t_L g1320 ( 
.A1(n_1232),
.A2(n_1277),
.B(n_1154),
.C(n_1211),
.Y(n_1320)
);

INVx1_ASAP7_75t_L g1321 ( 
.A(n_1197),
.Y(n_1321)
);

AND2x2_ASAP7_75t_L g1322 ( 
.A(n_1152),
.B(n_1168),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1152),
.B(n_1168),
.Y(n_1323)
);

AND2x4_ASAP7_75t_L g1324 ( 
.A(n_1250),
.B(n_1282),
.Y(n_1324)
);

AOI21xp5_ASAP7_75t_SL g1325 ( 
.A1(n_1155),
.A2(n_1171),
.B(n_1258),
.Y(n_1325)
);

INVx4_ASAP7_75t_L g1326 ( 
.A(n_1224),
.Y(n_1326)
);

BUFx12f_ASAP7_75t_L g1327 ( 
.A(n_1284),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1146),
.B(n_1150),
.Y(n_1328)
);

AND2x4_ASAP7_75t_L g1329 ( 
.A(n_1250),
.B(n_1282),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1153),
.Y(n_1330)
);

NOR2xp33_ASAP7_75t_SL g1331 ( 
.A(n_1188),
.B(n_1212),
.Y(n_1331)
);

INVx2_ASAP7_75t_L g1332 ( 
.A(n_1261),
.Y(n_1332)
);

INVx6_ASAP7_75t_L g1333 ( 
.A(n_1227),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1274),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1266),
.Y(n_1335)
);

INVx3_ASAP7_75t_L g1336 ( 
.A(n_1274),
.Y(n_1336)
);

AND2x2_ASAP7_75t_L g1337 ( 
.A(n_1181),
.B(n_1192),
.Y(n_1337)
);

INVx3_ASAP7_75t_SL g1338 ( 
.A(n_1173),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1181),
.B(n_1192),
.Y(n_1339)
);

BUFx2_ASAP7_75t_L g1340 ( 
.A(n_1158),
.Y(n_1340)
);

BUFx4f_ASAP7_75t_SL g1341 ( 
.A(n_1214),
.Y(n_1341)
);

NOR2xp33_ASAP7_75t_L g1342 ( 
.A(n_1252),
.B(n_1258),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1165),
.Y(n_1343)
);

CKINVDCx5p33_ASAP7_75t_R g1344 ( 
.A(n_1212),
.Y(n_1344)
);

BUFx3_ASAP7_75t_L g1345 ( 
.A(n_1193),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1256),
.B(n_1215),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1235),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1203),
.B(n_1275),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_1203),
.B(n_1143),
.Y(n_1349)
);

INVx4_ASAP7_75t_L g1350 ( 
.A(n_1144),
.Y(n_1350)
);

NOR2xp33_ASAP7_75t_L g1351 ( 
.A(n_1171),
.B(n_1208),
.Y(n_1351)
);

BUFx4_ASAP7_75t_SL g1352 ( 
.A(n_1207),
.Y(n_1352)
);

CKINVDCx8_ASAP7_75t_R g1353 ( 
.A(n_1144),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1236),
.Y(n_1354)
);

AOI22xp5_ASAP7_75t_L g1355 ( 
.A1(n_1222),
.A2(n_1215),
.B1(n_1221),
.B2(n_1198),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1238),
.Y(n_1356)
);

OR2x6_ASAP7_75t_L g1357 ( 
.A(n_1144),
.B(n_1177),
.Y(n_1357)
);

NOR2x1_ASAP7_75t_L g1358 ( 
.A(n_1242),
.B(n_1257),
.Y(n_1358)
);

INVx2_ASAP7_75t_SL g1359 ( 
.A(n_1220),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1238),
.Y(n_1360)
);

BUFx6f_ASAP7_75t_L g1361 ( 
.A(n_1177),
.Y(n_1361)
);

AOI21xp5_ASAP7_75t_L g1362 ( 
.A1(n_1166),
.A2(n_1244),
.B(n_1272),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1219),
.A2(n_1221),
.B1(n_1222),
.B2(n_1254),
.Y(n_1363)
);

OR2x2_ASAP7_75t_L g1364 ( 
.A(n_1205),
.B(n_1206),
.Y(n_1364)
);

BUFx6f_ASAP7_75t_L g1365 ( 
.A(n_1177),
.Y(n_1365)
);

OR2x6_ASAP7_75t_L g1366 ( 
.A(n_1239),
.B(n_1279),
.Y(n_1366)
);

AOI22xp5_ASAP7_75t_L g1367 ( 
.A1(n_1176),
.A2(n_1210),
.B1(n_1202),
.B2(n_1217),
.Y(n_1367)
);

OR2x6_ASAP7_75t_L g1368 ( 
.A(n_1239),
.B(n_1279),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1245),
.Y(n_1369)
);

AOI21xp5_ASAP7_75t_L g1370 ( 
.A1(n_1166),
.A2(n_1240),
.B(n_1254),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1230),
.B(n_1253),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1176),
.B(n_1169),
.Y(n_1372)
);

OAI21xp5_ASAP7_75t_L g1373 ( 
.A1(n_1187),
.A2(n_1186),
.B(n_1169),
.Y(n_1373)
);

OA22x2_ASAP7_75t_L g1374 ( 
.A1(n_1216),
.A2(n_1228),
.B1(n_1244),
.B2(n_1240),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1230),
.B(n_1204),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_1179),
.Y(n_1376)
);

INVx2_ASAP7_75t_L g1377 ( 
.A(n_1175),
.Y(n_1377)
);

BUFx6f_ASAP7_75t_L g1378 ( 
.A(n_1239),
.Y(n_1378)
);

AOI21xp5_ASAP7_75t_L g1379 ( 
.A1(n_1231),
.A2(n_1259),
.B(n_1271),
.Y(n_1379)
);

NAND2xp5_ASAP7_75t_SL g1380 ( 
.A(n_1216),
.B(n_1219),
.Y(n_1380)
);

AO32x2_ASAP7_75t_L g1381 ( 
.A1(n_1209),
.A2(n_1249),
.A3(n_1280),
.B1(n_1269),
.B2(n_1246),
.Y(n_1381)
);

AOI221x1_ASAP7_75t_L g1382 ( 
.A1(n_1226),
.A2(n_1195),
.B1(n_1223),
.B2(n_1182),
.C(n_1183),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1204),
.B(n_1209),
.Y(n_1383)
);

A2O1A1Ixp33_ASAP7_75t_L g1384 ( 
.A1(n_1175),
.A2(n_1194),
.B(n_1179),
.C(n_1189),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1209),
.B(n_1248),
.Y(n_1385)
);

OR2x6_ASAP7_75t_L g1386 ( 
.A(n_1196),
.B(n_1199),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1196),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_SL g1388 ( 
.A(n_1157),
.B(n_1199),
.Y(n_1388)
);

BUFx2_ASAP7_75t_SL g1389 ( 
.A(n_1218),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1249),
.B(n_1280),
.Y(n_1390)
);

CKINVDCx11_ASAP7_75t_R g1391 ( 
.A(n_1218),
.Y(n_1391)
);

A2O1A1Ixp33_ASAP7_75t_L g1392 ( 
.A1(n_1229),
.A2(n_1159),
.B(n_1147),
.C(n_1162),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1249),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1269),
.B(n_1280),
.Y(n_1394)
);

AOI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1140),
.A2(n_1260),
.B(n_1270),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1276),
.Y(n_1396)
);

O2A1O1Ixp33_ASAP7_75t_L g1397 ( 
.A1(n_1278),
.A2(n_1237),
.B(n_1247),
.C(n_1139),
.Y(n_1397)
);

AOI21xp5_ASAP7_75t_L g1398 ( 
.A1(n_1148),
.A2(n_992),
.B(n_1241),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1148),
.A2(n_992),
.B(n_1241),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1224),
.Y(n_1400)
);

HB1xp67_ASAP7_75t_L g1401 ( 
.A(n_1163),
.Y(n_1401)
);

AOI221x1_ASAP7_75t_L g1402 ( 
.A1(n_1142),
.A2(n_1283),
.B1(n_1281),
.B2(n_1237),
.C(n_1247),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1145),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_1160),
.Y(n_1404)
);

O2A1O1Ixp5_ASAP7_75t_L g1405 ( 
.A1(n_1142),
.A2(n_992),
.B(n_1237),
.C(n_1139),
.Y(n_1405)
);

OA21x2_ASAP7_75t_L g1406 ( 
.A1(n_1174),
.A2(n_1166),
.B(n_1149),
.Y(n_1406)
);

NAND2x1_ASAP7_75t_L g1407 ( 
.A(n_1264),
.B(n_999),
.Y(n_1407)
);

AND2x2_ASAP7_75t_L g1408 ( 
.A(n_1167),
.B(n_981),
.Y(n_1408)
);

NOR2xp33_ASAP7_75t_R g1409 ( 
.A(n_1160),
.B(n_656),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1145),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1191),
.Y(n_1411)
);

AOI21xp5_ASAP7_75t_L g1412 ( 
.A1(n_1148),
.A2(n_992),
.B(n_1241),
.Y(n_1412)
);

OAI21xp33_ASAP7_75t_L g1413 ( 
.A1(n_1285),
.A2(n_980),
.B(n_926),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1191),
.Y(n_1414)
);

NAND2xp5_ASAP7_75t_L g1415 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1415)
);

AOI21xp5_ASAP7_75t_L g1416 ( 
.A1(n_1148),
.A2(n_992),
.B(n_1241),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1145),
.Y(n_1417)
);

AOI22xp5_ASAP7_75t_L g1418 ( 
.A1(n_1143),
.A2(n_992),
.B1(n_980),
.B2(n_925),
.Y(n_1418)
);

HB1xp67_ASAP7_75t_L g1419 ( 
.A(n_1163),
.Y(n_1419)
);

BUFx3_ASAP7_75t_L g1420 ( 
.A(n_1190),
.Y(n_1420)
);

NAND3xp33_ASAP7_75t_SL g1421 ( 
.A(n_1139),
.B(n_980),
.C(n_992),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1167),
.B(n_981),
.Y(n_1422)
);

INVx1_ASAP7_75t_L g1423 ( 
.A(n_1191),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1424)
);

INVx4_ASAP7_75t_R g1425 ( 
.A(n_1184),
.Y(n_1425)
);

AOI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1148),
.A2(n_992),
.B(n_1241),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1145),
.Y(n_1427)
);

AND2x4_ASAP7_75t_L g1428 ( 
.A(n_1152),
.B(n_1168),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1143),
.A2(n_992),
.B1(n_980),
.B2(n_925),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1191),
.Y(n_1430)
);

CKINVDCx20_ASAP7_75t_R g1431 ( 
.A(n_1160),
.Y(n_1431)
);

CKINVDCx20_ASAP7_75t_R g1432 ( 
.A(n_1160),
.Y(n_1432)
);

OR2x2_ASAP7_75t_L g1433 ( 
.A(n_1141),
.B(n_604),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1285),
.B(n_980),
.Y(n_1434)
);

NAND2xp5_ASAP7_75t_L g1435 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1435)
);

AND2x4_ASAP7_75t_L g1436 ( 
.A(n_1152),
.B(n_1168),
.Y(n_1436)
);

OA21x2_ASAP7_75t_L g1437 ( 
.A1(n_1174),
.A2(n_1166),
.B(n_1149),
.Y(n_1437)
);

AOI21xp5_ASAP7_75t_L g1438 ( 
.A1(n_1148),
.A2(n_992),
.B(n_1241),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1439)
);

NAND2xp5_ASAP7_75t_L g1440 ( 
.A(n_1285),
.B(n_1141),
.Y(n_1440)
);

INVx3_ASAP7_75t_SL g1441 ( 
.A(n_1188),
.Y(n_1441)
);

OAI21xp33_ASAP7_75t_L g1442 ( 
.A1(n_1285),
.A2(n_980),
.B(n_926),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1191),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1234),
.A2(n_1260),
.B(n_1243),
.Y(n_1444)
);

BUFx2_ASAP7_75t_L g1445 ( 
.A(n_1190),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1393),
.Y(n_1446)
);

INVx3_ASAP7_75t_L g1447 ( 
.A(n_1296),
.Y(n_1447)
);

OAI21x1_ASAP7_75t_L g1448 ( 
.A1(n_1395),
.A2(n_1444),
.B(n_1379),
.Y(n_1448)
);

AND2x2_ASAP7_75t_L g1449 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1449)
);

INVx2_ASAP7_75t_SL g1450 ( 
.A(n_1333),
.Y(n_1450)
);

CKINVDCx20_ASAP7_75t_R g1451 ( 
.A(n_1431),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1330),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_SL g1453 ( 
.A1(n_1434),
.A2(n_1304),
.B1(n_1342),
.B2(n_1349),
.Y(n_1453)
);

OAI22xp5_ASAP7_75t_L g1454 ( 
.A1(n_1434),
.A2(n_1287),
.B1(n_1435),
.B2(n_1415),
.Y(n_1454)
);

AOI21x1_ASAP7_75t_L g1455 ( 
.A1(n_1398),
.A2(n_1412),
.B(n_1399),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1343),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1351),
.B(n_1302),
.Y(n_1457)
);

AOI22xp33_ASAP7_75t_SL g1458 ( 
.A1(n_1342),
.A2(n_1374),
.B1(n_1309),
.B2(n_1409),
.Y(n_1458)
);

AOI22xp33_ASAP7_75t_SL g1459 ( 
.A1(n_1374),
.A2(n_1309),
.B1(n_1409),
.B2(n_1370),
.Y(n_1459)
);

BUFx3_ASAP7_75t_L g1460 ( 
.A(n_1307),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1385),
.Y(n_1461)
);

INVxp67_ASAP7_75t_L g1462 ( 
.A(n_1340),
.Y(n_1462)
);

OA21x2_ASAP7_75t_L g1463 ( 
.A1(n_1305),
.A2(n_1382),
.B(n_1294),
.Y(n_1463)
);

AOI22xp33_ASAP7_75t_L g1464 ( 
.A1(n_1413),
.A2(n_1442),
.B1(n_1363),
.B2(n_1289),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1337),
.B(n_1339),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1347),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1296),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1354),
.Y(n_1468)
);

INVx2_ASAP7_75t_L g1469 ( 
.A(n_1369),
.Y(n_1469)
);

INVx2_ASAP7_75t_SL g1470 ( 
.A(n_1333),
.Y(n_1470)
);

AOI22xp33_ASAP7_75t_L g1471 ( 
.A1(n_1363),
.A2(n_1421),
.B1(n_1380),
.B2(n_1295),
.Y(n_1471)
);

NAND2x1p5_ASAP7_75t_L g1472 ( 
.A(n_1367),
.B(n_1388),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_L g1473 ( 
.A1(n_1421),
.A2(n_1380),
.B1(n_1295),
.B2(n_1355),
.Y(n_1473)
);

INVx1_ASAP7_75t_L g1474 ( 
.A(n_1291),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1383),
.Y(n_1475)
);

AOI21x1_ASAP7_75t_L g1476 ( 
.A1(n_1398),
.A2(n_1412),
.B(n_1399),
.Y(n_1476)
);

AND2x2_ASAP7_75t_L g1477 ( 
.A(n_1299),
.B(n_1301),
.Y(n_1477)
);

AOI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1416),
.A2(n_1438),
.B(n_1426),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1316),
.Y(n_1479)
);

OAI21xp5_ASAP7_75t_L g1480 ( 
.A1(n_1405),
.A2(n_1429),
.B(n_1418),
.Y(n_1480)
);

HB1xp67_ASAP7_75t_SL g1481 ( 
.A(n_1298),
.Y(n_1481)
);

BUFx4f_ASAP7_75t_SL g1482 ( 
.A(n_1327),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1303),
.Y(n_1483)
);

NOR2xp33_ASAP7_75t_L g1484 ( 
.A(n_1433),
.B(n_1424),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1332),
.Y(n_1485)
);

CKINVDCx20_ASAP7_75t_R g1486 ( 
.A(n_1432),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1335),
.Y(n_1487)
);

OAI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1439),
.A2(n_1440),
.B1(n_1314),
.B2(n_1318),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1403),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1410),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1417),
.Y(n_1491)
);

HB1xp67_ASAP7_75t_L g1492 ( 
.A(n_1401),
.Y(n_1492)
);

HB1xp67_ASAP7_75t_L g1493 ( 
.A(n_1401),
.Y(n_1493)
);

AOI22xp33_ASAP7_75t_SL g1494 ( 
.A1(n_1362),
.A2(n_1370),
.B1(n_1319),
.B2(n_1408),
.Y(n_1494)
);

INVxp67_ASAP7_75t_SL g1495 ( 
.A(n_1419),
.Y(n_1495)
);

INVx3_ASAP7_75t_L g1496 ( 
.A(n_1296),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1427),
.Y(n_1497)
);

INVx2_ASAP7_75t_SL g1498 ( 
.A(n_1333),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1381),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1296),
.Y(n_1500)
);

OR2x6_ASAP7_75t_L g1501 ( 
.A(n_1325),
.B(n_1362),
.Y(n_1501)
);

CKINVDCx20_ASAP7_75t_R g1502 ( 
.A(n_1441),
.Y(n_1502)
);

INVx1_ASAP7_75t_SL g1503 ( 
.A(n_1288),
.Y(n_1503)
);

HB1xp67_ASAP7_75t_L g1504 ( 
.A(n_1419),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1321),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1364),
.Y(n_1506)
);

INVx3_ASAP7_75t_L g1507 ( 
.A(n_1312),
.Y(n_1507)
);

CKINVDCx11_ASAP7_75t_R g1508 ( 
.A(n_1441),
.Y(n_1508)
);

CKINVDCx6p67_ASAP7_75t_R g1509 ( 
.A(n_1338),
.Y(n_1509)
);

OR2x6_ASAP7_75t_L g1510 ( 
.A(n_1297),
.B(n_1389),
.Y(n_1510)
);

NOR2xp33_ASAP7_75t_L g1511 ( 
.A(n_1422),
.B(n_1322),
.Y(n_1511)
);

BUFx3_ASAP7_75t_L g1512 ( 
.A(n_1324),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1346),
.A2(n_1315),
.B1(n_1311),
.B2(n_1306),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1411),
.Y(n_1514)
);

OAI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1328),
.A2(n_1414),
.B1(n_1443),
.B2(n_1423),
.Y(n_1515)
);

AO21x2_ASAP7_75t_L g1516 ( 
.A1(n_1392),
.A2(n_1373),
.B(n_1297),
.Y(n_1516)
);

AOI22xp33_ASAP7_75t_L g1517 ( 
.A1(n_1391),
.A2(n_1308),
.B1(n_1348),
.B2(n_1371),
.Y(n_1517)
);

OA21x2_ASAP7_75t_L g1518 ( 
.A1(n_1402),
.A2(n_1392),
.B(n_1320),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1430),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1376),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1387),
.Y(n_1521)
);

CKINVDCx20_ASAP7_75t_R g1522 ( 
.A(n_1404),
.Y(n_1522)
);

AOI22xp33_ASAP7_75t_L g1523 ( 
.A1(n_1391),
.A2(n_1375),
.B1(n_1437),
.B2(n_1406),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1387),
.Y(n_1524)
);

OR2x2_ASAP7_75t_L g1525 ( 
.A(n_1372),
.B(n_1437),
.Y(n_1525)
);

NAND2x1_ASAP7_75t_L g1526 ( 
.A(n_1396),
.B(n_1358),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1320),
.Y(n_1527)
);

AOI22xp33_ASAP7_75t_L g1528 ( 
.A1(n_1428),
.A2(n_1436),
.B1(n_1323),
.B2(n_1329),
.Y(n_1528)
);

OAI21x1_ASAP7_75t_SL g1529 ( 
.A1(n_1397),
.A2(n_1350),
.B(n_1400),
.Y(n_1529)
);

AOI22xp33_ASAP7_75t_L g1530 ( 
.A1(n_1428),
.A2(n_1436),
.B1(n_1324),
.B2(n_1329),
.Y(n_1530)
);

OAI22xp5_ASAP7_75t_L g1531 ( 
.A1(n_1300),
.A2(n_1293),
.B1(n_1313),
.B2(n_1359),
.Y(n_1531)
);

OR2x2_ASAP7_75t_L g1532 ( 
.A(n_1390),
.B(n_1394),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1381),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1405),
.Y(n_1534)
);

AOI22xp33_ASAP7_75t_SL g1535 ( 
.A1(n_1331),
.A2(n_1445),
.B1(n_1420),
.B2(n_1341),
.Y(n_1535)
);

INVx3_ASAP7_75t_L g1536 ( 
.A(n_1312),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1386),
.Y(n_1537)
);

AOI22xp33_ASAP7_75t_L g1538 ( 
.A1(n_1341),
.A2(n_1345),
.B1(n_1360),
.B2(n_1356),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1386),
.Y(n_1539)
);

BUFx3_ASAP7_75t_L g1540 ( 
.A(n_1353),
.Y(n_1540)
);

NAND2x1_ASAP7_75t_L g1541 ( 
.A(n_1312),
.B(n_1360),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1386),
.Y(n_1542)
);

CKINVDCx11_ASAP7_75t_R g1543 ( 
.A(n_1338),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1361),
.Y(n_1544)
);

HB1xp67_ASAP7_75t_L g1545 ( 
.A(n_1357),
.Y(n_1545)
);

OAI22xp33_ASAP7_75t_L g1546 ( 
.A1(n_1344),
.A2(n_1352),
.B1(n_1400),
.B2(n_1326),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1356),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1384),
.B(n_1357),
.Y(n_1548)
);

OAI22xp5_ASAP7_75t_L g1549 ( 
.A1(n_1326),
.A2(n_1334),
.B1(n_1336),
.B2(n_1310),
.Y(n_1549)
);

OR2x2_ASAP7_75t_L g1550 ( 
.A(n_1357),
.B(n_1366),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1334),
.B(n_1336),
.Y(n_1551)
);

CKINVDCx6p67_ASAP7_75t_R g1552 ( 
.A(n_1366),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1361),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1292),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1290),
.A2(n_1310),
.B1(n_1292),
.B2(n_1317),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1290),
.A2(n_1350),
.B1(n_1361),
.B2(n_1365),
.Y(n_1556)
);

BUFx10_ASAP7_75t_L g1557 ( 
.A(n_1361),
.Y(n_1557)
);

CKINVDCx11_ASAP7_75t_R g1558 ( 
.A(n_1365),
.Y(n_1558)
);

BUFx2_ASAP7_75t_L g1559 ( 
.A(n_1366),
.Y(n_1559)
);

CKINVDCx5p33_ASAP7_75t_R g1560 ( 
.A(n_1352),
.Y(n_1560)
);

NAND2x1p5_ASAP7_75t_L g1561 ( 
.A(n_1407),
.B(n_1365),
.Y(n_1561)
);

AOI22xp33_ASAP7_75t_L g1562 ( 
.A1(n_1365),
.A2(n_1378),
.B1(n_1368),
.B2(n_1317),
.Y(n_1562)
);

OAI22xp5_ASAP7_75t_L g1563 ( 
.A1(n_1368),
.A2(n_1434),
.B1(n_980),
.B2(n_1415),
.Y(n_1563)
);

AO21x2_ASAP7_75t_L g1564 ( 
.A1(n_1368),
.A2(n_1378),
.B(n_1425),
.Y(n_1564)
);

INVx1_ASAP7_75t_L g1565 ( 
.A(n_1378),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1378),
.B(n_1349),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1434),
.B(n_925),
.Y(n_1567)
);

AOI22xp33_ASAP7_75t_SL g1568 ( 
.A1(n_1434),
.A2(n_578),
.B1(n_980),
.B2(n_992),
.Y(n_1568)
);

INVx3_ASAP7_75t_L g1569 ( 
.A(n_1296),
.Y(n_1569)
);

BUFx6f_ASAP7_75t_L g1570 ( 
.A(n_1296),
.Y(n_1570)
);

INVx3_ASAP7_75t_L g1571 ( 
.A(n_1296),
.Y(n_1571)
);

AO21x1_ASAP7_75t_L g1572 ( 
.A1(n_1309),
.A2(n_1142),
.B(n_1380),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1434),
.B(n_1285),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1330),
.Y(n_1574)
);

AOI21x1_ASAP7_75t_L g1575 ( 
.A1(n_1395),
.A2(n_1399),
.B(n_1398),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1434),
.B(n_1285),
.Y(n_1576)
);

BUFx2_ASAP7_75t_L g1577 ( 
.A(n_1303),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1303),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1434),
.B(n_1285),
.Y(n_1579)
);

AO21x2_ASAP7_75t_L g1580 ( 
.A1(n_1398),
.A2(n_1142),
.B(n_1399),
.Y(n_1580)
);

AOI22xp5_ASAP7_75t_L g1581 ( 
.A1(n_1413),
.A2(n_648),
.B1(n_980),
.B2(n_566),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1434),
.A2(n_980),
.B1(n_1415),
.B2(n_1287),
.Y(n_1582)
);

HB1xp67_ASAP7_75t_L g1583 ( 
.A(n_1401),
.Y(n_1583)
);

AND2x2_ASAP7_75t_L g1584 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1584)
);

BUFx6f_ASAP7_75t_L g1585 ( 
.A(n_1296),
.Y(n_1585)
);

AO21x1_ASAP7_75t_L g1586 ( 
.A1(n_1309),
.A2(n_1142),
.B(n_1380),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1413),
.A2(n_992),
.B1(n_1442),
.B2(n_1304),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1413),
.A2(n_992),
.B1(n_1442),
.B2(n_1304),
.Y(n_1588)
);

AOI21x1_ASAP7_75t_L g1589 ( 
.A1(n_1395),
.A2(n_1399),
.B(n_1398),
.Y(n_1589)
);

AO21x1_ASAP7_75t_L g1590 ( 
.A1(n_1309),
.A2(n_1142),
.B(n_1380),
.Y(n_1590)
);

AND2x4_ASAP7_75t_L g1591 ( 
.A(n_1337),
.B(n_1339),
.Y(n_1591)
);

AOI222xp33_ASAP7_75t_L g1592 ( 
.A1(n_1413),
.A2(n_1049),
.B1(n_1442),
.B2(n_980),
.C1(n_1211),
.C2(n_1059),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1377),
.Y(n_1593)
);

INVx2_ASAP7_75t_SL g1594 ( 
.A(n_1333),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1307),
.Y(n_1595)
);

INVx2_ASAP7_75t_SL g1596 ( 
.A(n_1333),
.Y(n_1596)
);

INVx1_ASAP7_75t_SL g1597 ( 
.A(n_1303),
.Y(n_1597)
);

BUFx3_ASAP7_75t_L g1598 ( 
.A(n_1307),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1330),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1434),
.B(n_1285),
.Y(n_1600)
);

BUFx6f_ASAP7_75t_L g1601 ( 
.A(n_1296),
.Y(n_1601)
);

OA21x2_ASAP7_75t_L g1602 ( 
.A1(n_1305),
.A2(n_1382),
.B(n_1294),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1434),
.B(n_1285),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1333),
.Y(n_1604)
);

BUFx3_ASAP7_75t_L g1605 ( 
.A(n_1307),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1413),
.A2(n_992),
.B1(n_1442),
.B2(n_1304),
.Y(n_1606)
);

INVx3_ASAP7_75t_L g1607 ( 
.A(n_1296),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1532),
.B(n_1461),
.Y(n_1608)
);

INVx1_ASAP7_75t_SL g1609 ( 
.A(n_1578),
.Y(n_1609)
);

HB1xp67_ASAP7_75t_L g1610 ( 
.A(n_1492),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1446),
.Y(n_1611)
);

OR2x6_ASAP7_75t_L g1612 ( 
.A(n_1501),
.B(n_1510),
.Y(n_1612)
);

INVx2_ASAP7_75t_SL g1613 ( 
.A(n_1493),
.Y(n_1613)
);

BUFx12f_ASAP7_75t_L g1614 ( 
.A(n_1508),
.Y(n_1614)
);

BUFx4f_ASAP7_75t_SL g1615 ( 
.A(n_1451),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1477),
.B(n_1484),
.Y(n_1616)
);

INVx2_ASAP7_75t_SL g1617 ( 
.A(n_1504),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1477),
.B(n_1454),
.Y(n_1618)
);

NAND2x1p5_ASAP7_75t_L g1619 ( 
.A(n_1548),
.B(n_1526),
.Y(n_1619)
);

AND2x2_ASAP7_75t_L g1620 ( 
.A(n_1532),
.B(n_1461),
.Y(n_1620)
);

AO21x2_ASAP7_75t_L g1621 ( 
.A1(n_1455),
.A2(n_1478),
.B(n_1476),
.Y(n_1621)
);

HB1xp67_ASAP7_75t_L g1622 ( 
.A(n_1583),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1483),
.Y(n_1623)
);

CKINVDCx20_ASAP7_75t_R g1624 ( 
.A(n_1451),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1525),
.Y(n_1625)
);

AND2x2_ASAP7_75t_L g1626 ( 
.A(n_1449),
.B(n_1584),
.Y(n_1626)
);

OR2x2_ASAP7_75t_L g1627 ( 
.A(n_1525),
.B(n_1475),
.Y(n_1627)
);

NOR2x1_ASAP7_75t_L g1628 ( 
.A(n_1515),
.B(n_1480),
.Y(n_1628)
);

OR2x6_ASAP7_75t_L g1629 ( 
.A(n_1501),
.B(n_1510),
.Y(n_1629)
);

BUFx2_ASAP7_75t_L g1630 ( 
.A(n_1548),
.Y(n_1630)
);

OAI21x1_ASAP7_75t_L g1631 ( 
.A1(n_1448),
.A2(n_1589),
.B(n_1575),
.Y(n_1631)
);

INVxp67_ASAP7_75t_L g1632 ( 
.A(n_1483),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1449),
.B(n_1584),
.Y(n_1633)
);

OAI21xp33_ASAP7_75t_SL g1634 ( 
.A1(n_1501),
.A2(n_1471),
.B(n_1464),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_L g1635 ( 
.A(n_1457),
.B(n_1582),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1577),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1523),
.B(n_1527),
.Y(n_1637)
);

HB1xp67_ASAP7_75t_L g1638 ( 
.A(n_1577),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1566),
.B(n_1459),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1566),
.B(n_1457),
.Y(n_1640)
);

BUFx4f_ASAP7_75t_SL g1641 ( 
.A(n_1486),
.Y(n_1641)
);

BUFx6f_ASAP7_75t_L g1642 ( 
.A(n_1570),
.Y(n_1642)
);

HB1xp67_ASAP7_75t_L g1643 ( 
.A(n_1495),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1499),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1458),
.B(n_1494),
.Y(n_1645)
);

AND2x6_ASAP7_75t_L g1646 ( 
.A(n_1527),
.B(n_1505),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1537),
.B(n_1542),
.Y(n_1647)
);

BUFx3_ASAP7_75t_L g1648 ( 
.A(n_1564),
.Y(n_1648)
);

BUFx2_ASAP7_75t_L g1649 ( 
.A(n_1472),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1473),
.B(n_1501),
.Y(n_1650)
);

AND2x2_ASAP7_75t_L g1651 ( 
.A(n_1453),
.B(n_1469),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1533),
.Y(n_1652)
);

INVx2_ASAP7_75t_L g1653 ( 
.A(n_1463),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1533),
.Y(n_1654)
);

AND2x2_ASAP7_75t_L g1655 ( 
.A(n_1469),
.B(n_1518),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1472),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1472),
.Y(n_1657)
);

INVx1_ASAP7_75t_L g1658 ( 
.A(n_1510),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1510),
.Y(n_1659)
);

AND2x2_ASAP7_75t_L g1660 ( 
.A(n_1518),
.B(n_1534),
.Y(n_1660)
);

OAI21x1_ASAP7_75t_L g1661 ( 
.A1(n_1526),
.A2(n_1529),
.B(n_1463),
.Y(n_1661)
);

INVx3_ASAP7_75t_L g1662 ( 
.A(n_1516),
.Y(n_1662)
);

AND2x4_ASAP7_75t_L g1663 ( 
.A(n_1542),
.B(n_1539),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1514),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1519),
.Y(n_1665)
);

AO21x2_ASAP7_75t_L g1666 ( 
.A1(n_1580),
.A2(n_1572),
.B(n_1590),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1452),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1520),
.Y(n_1668)
);

OA21x2_ASAP7_75t_L g1669 ( 
.A1(n_1572),
.A2(n_1590),
.B(n_1586),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1456),
.Y(n_1670)
);

HB1xp67_ASAP7_75t_L g1671 ( 
.A(n_1597),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1466),
.Y(n_1672)
);

INVxp67_ASAP7_75t_L g1673 ( 
.A(n_1511),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1488),
.B(n_1573),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1468),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1518),
.B(n_1586),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1518),
.B(n_1593),
.Y(n_1677)
);

OR2x6_ASAP7_75t_L g1678 ( 
.A(n_1529),
.B(n_1463),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1574),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1576),
.B(n_1579),
.Y(n_1680)
);

INVx2_ASAP7_75t_SL g1681 ( 
.A(n_1521),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1580),
.A2(n_1516),
.B(n_1599),
.Y(n_1682)
);

HB1xp67_ASAP7_75t_L g1683 ( 
.A(n_1559),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1559),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1587),
.A2(n_1588),
.B(n_1606),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1602),
.Y(n_1686)
);

BUFx2_ASAP7_75t_L g1687 ( 
.A(n_1524),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1513),
.B(n_1602),
.Y(n_1688)
);

BUFx2_ASAP7_75t_L g1689 ( 
.A(n_1545),
.Y(n_1689)
);

NAND2xp5_ASAP7_75t_L g1690 ( 
.A(n_1600),
.B(n_1603),
.Y(n_1690)
);

BUFx2_ASAP7_75t_L g1691 ( 
.A(n_1580),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1563),
.B(n_1506),
.Y(n_1692)
);

INVxp67_ASAP7_75t_L g1693 ( 
.A(n_1462),
.Y(n_1693)
);

OR2x6_ASAP7_75t_L g1694 ( 
.A(n_1554),
.B(n_1541),
.Y(n_1694)
);

AND2x4_ASAP7_75t_L g1695 ( 
.A(n_1547),
.B(n_1485),
.Y(n_1695)
);

HB1xp67_ASAP7_75t_L g1696 ( 
.A(n_1550),
.Y(n_1696)
);

OA21x2_ASAP7_75t_L g1697 ( 
.A1(n_1517),
.A2(n_1491),
.B(n_1487),
.Y(n_1697)
);

INVx2_ASAP7_75t_SL g1698 ( 
.A(n_1557),
.Y(n_1698)
);

OAI21x1_ASAP7_75t_L g1699 ( 
.A1(n_1541),
.A2(n_1549),
.B(n_1497),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1497),
.B(n_1474),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1568),
.B(n_1567),
.Y(n_1701)
);

INVx2_ASAP7_75t_L g1702 ( 
.A(n_1489),
.Y(n_1702)
);

INVx1_ASAP7_75t_L g1703 ( 
.A(n_1490),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1557),
.Y(n_1704)
);

OR2x6_ASAP7_75t_L g1705 ( 
.A(n_1555),
.B(n_1601),
.Y(n_1705)
);

INVx6_ASAP7_75t_L g1706 ( 
.A(n_1557),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1592),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1531),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1465),
.B(n_1591),
.Y(n_1709)
);

OR2x2_ASAP7_75t_L g1710 ( 
.A(n_1503),
.B(n_1581),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1544),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1553),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1565),
.Y(n_1713)
);

INVx1_ASAP7_75t_SL g1714 ( 
.A(n_1486),
.Y(n_1714)
);

AO21x1_ASAP7_75t_SL g1715 ( 
.A1(n_1562),
.A2(n_1551),
.B(n_1538),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1570),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1608),
.B(n_1591),
.Y(n_1717)
);

AOI22xp33_ASAP7_75t_L g1718 ( 
.A1(n_1707),
.A2(n_1591),
.B1(n_1465),
.B2(n_1535),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1608),
.B(n_1465),
.Y(n_1719)
);

HB1xp67_ASAP7_75t_L g1720 ( 
.A(n_1625),
.Y(n_1720)
);

AND2x2_ASAP7_75t_L g1721 ( 
.A(n_1620),
.B(n_1447),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1620),
.B(n_1607),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1688),
.B(n_1607),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1688),
.B(n_1640),
.Y(n_1724)
);

AND2x4_ASAP7_75t_L g1725 ( 
.A(n_1612),
.B(n_1607),
.Y(n_1725)
);

BUFx4f_ASAP7_75t_L g1726 ( 
.A(n_1685),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1653),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1640),
.B(n_1536),
.Y(n_1728)
);

BUFx3_ASAP7_75t_L g1729 ( 
.A(n_1648),
.Y(n_1729)
);

AOI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1707),
.A2(n_1546),
.B1(n_1560),
.B2(n_1502),
.Y(n_1730)
);

INVx2_ASAP7_75t_SL g1731 ( 
.A(n_1648),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1674),
.B(n_1536),
.Y(n_1732)
);

OAI22xp5_ASAP7_75t_L g1733 ( 
.A1(n_1701),
.A2(n_1560),
.B1(n_1552),
.B2(n_1509),
.Y(n_1733)
);

INVx2_ASAP7_75t_L g1734 ( 
.A(n_1611),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1630),
.B(n_1496),
.Y(n_1735)
);

BUFx3_ASAP7_75t_L g1736 ( 
.A(n_1619),
.Y(n_1736)
);

HB1xp67_ASAP7_75t_L g1737 ( 
.A(n_1682),
.Y(n_1737)
);

OR2x6_ASAP7_75t_L g1738 ( 
.A(n_1612),
.B(n_1561),
.Y(n_1738)
);

OAI31xp33_ASAP7_75t_L g1739 ( 
.A1(n_1645),
.A2(n_1710),
.A3(n_1680),
.B(n_1690),
.Y(n_1739)
);

AND2x2_ASAP7_75t_L g1740 ( 
.A(n_1630),
.B(n_1496),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1655),
.B(n_1496),
.Y(n_1741)
);

AOI32xp33_ASAP7_75t_L g1742 ( 
.A1(n_1645),
.A2(n_1540),
.A3(n_1528),
.B1(n_1512),
.B2(n_1530),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1660),
.B(n_1676),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1660),
.B(n_1507),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1626),
.B(n_1633),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1626),
.B(n_1569),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1618),
.B(n_1569),
.Y(n_1747)
);

AOI22xp33_ASAP7_75t_L g1748 ( 
.A1(n_1685),
.A2(n_1512),
.B1(n_1508),
.B2(n_1543),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1639),
.B(n_1500),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1639),
.B(n_1507),
.Y(n_1750)
);

INVxp67_ASAP7_75t_L g1751 ( 
.A(n_1643),
.Y(n_1751)
);

OR2x2_ASAP7_75t_L g1752 ( 
.A(n_1627),
.B(n_1509),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1627),
.B(n_1450),
.Y(n_1753)
);

BUFx4f_ASAP7_75t_L g1754 ( 
.A(n_1685),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1677),
.B(n_1571),
.Y(n_1755)
);

OR2x2_ASAP7_75t_L g1756 ( 
.A(n_1682),
.B(n_1604),
.Y(n_1756)
);

AND2x2_ASAP7_75t_L g1757 ( 
.A(n_1696),
.B(n_1467),
.Y(n_1757)
);

BUFx2_ASAP7_75t_L g1758 ( 
.A(n_1646),
.Y(n_1758)
);

BUFx6f_ASAP7_75t_L g1759 ( 
.A(n_1629),
.Y(n_1759)
);

AOI22xp33_ASAP7_75t_L g1760 ( 
.A1(n_1685),
.A2(n_1628),
.B1(n_1634),
.B2(n_1650),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1621),
.A2(n_1601),
.B(n_1570),
.Y(n_1761)
);

HB1xp67_ASAP7_75t_L g1762 ( 
.A(n_1682),
.Y(n_1762)
);

OR2x2_ASAP7_75t_L g1763 ( 
.A(n_1637),
.B(n_1596),
.Y(n_1763)
);

AND2x4_ASAP7_75t_L g1764 ( 
.A(n_1629),
.B(n_1658),
.Y(n_1764)
);

OR2x2_ASAP7_75t_L g1765 ( 
.A(n_1637),
.B(n_1596),
.Y(n_1765)
);

AOI222xp33_ASAP7_75t_L g1766 ( 
.A1(n_1634),
.A2(n_1482),
.B1(n_1543),
.B2(n_1502),
.C1(n_1540),
.C2(n_1522),
.Y(n_1766)
);

NOR2x1_ASAP7_75t_L g1767 ( 
.A(n_1628),
.B(n_1571),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1650),
.A2(n_1522),
.B1(n_1605),
.B2(n_1479),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1686),
.Y(n_1769)
);

BUFx3_ASAP7_75t_L g1770 ( 
.A(n_1619),
.Y(n_1770)
);

AND2x2_ASAP7_75t_L g1771 ( 
.A(n_1676),
.B(n_1570),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1658),
.B(n_1594),
.Y(n_1772)
);

BUFx2_ASAP7_75t_L g1773 ( 
.A(n_1646),
.Y(n_1773)
);

AND2x4_ASAP7_75t_L g1774 ( 
.A(n_1629),
.B(n_1601),
.Y(n_1774)
);

AND2x4_ASAP7_75t_SL g1775 ( 
.A(n_1705),
.B(n_1552),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1747),
.B(n_1616),
.Y(n_1776)
);

OAI221xp5_ASAP7_75t_L g1777 ( 
.A1(n_1739),
.A2(n_1710),
.B1(n_1635),
.B2(n_1692),
.C(n_1708),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1739),
.B(n_1692),
.C(n_1657),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1747),
.B(n_1610),
.Y(n_1779)
);

NAND3xp33_ASAP7_75t_L g1780 ( 
.A(n_1766),
.B(n_1657),
.C(n_1656),
.Y(n_1780)
);

AND2x2_ASAP7_75t_SL g1781 ( 
.A(n_1726),
.B(n_1669),
.Y(n_1781)
);

NOR3xp33_ASAP7_75t_L g1782 ( 
.A(n_1733),
.B(n_1651),
.C(n_1693),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1751),
.B(n_1622),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1724),
.B(n_1659),
.Y(n_1784)
);

NAND3xp33_ASAP7_75t_L g1785 ( 
.A(n_1766),
.B(n_1656),
.C(n_1697),
.Y(n_1785)
);

NAND4xp25_ASAP7_75t_L g1786 ( 
.A(n_1732),
.B(n_1651),
.C(n_1632),
.D(n_1673),
.Y(n_1786)
);

NAND3xp33_ASAP7_75t_L g1787 ( 
.A(n_1748),
.B(n_1697),
.C(n_1663),
.Y(n_1787)
);

NAND3xp33_ASAP7_75t_L g1788 ( 
.A(n_1748),
.B(n_1697),
.C(n_1663),
.Y(n_1788)
);

AND2x2_ASAP7_75t_L g1789 ( 
.A(n_1724),
.B(n_1678),
.Y(n_1789)
);

NAND3xp33_ASAP7_75t_L g1790 ( 
.A(n_1760),
.B(n_1697),
.C(n_1663),
.Y(n_1790)
);

AND2x2_ASAP7_75t_L g1791 ( 
.A(n_1743),
.B(n_1678),
.Y(n_1791)
);

NAND2xp5_ASAP7_75t_SL g1792 ( 
.A(n_1726),
.B(n_1647),
.Y(n_1792)
);

NAND3xp33_ASAP7_75t_L g1793 ( 
.A(n_1760),
.B(n_1663),
.C(n_1647),
.Y(n_1793)
);

NOR3xp33_ASAP7_75t_L g1794 ( 
.A(n_1733),
.B(n_1689),
.C(n_1714),
.Y(n_1794)
);

BUFx2_ASAP7_75t_SL g1795 ( 
.A(n_1757),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1751),
.B(n_1623),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1732),
.B(n_1636),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1743),
.B(n_1678),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1767),
.B(n_1742),
.C(n_1768),
.Y(n_1799)
);

OAI221xp5_ASAP7_75t_SL g1800 ( 
.A1(n_1742),
.A2(n_1609),
.B1(n_1705),
.B2(n_1678),
.C(n_1691),
.Y(n_1800)
);

NAND3xp33_ASAP7_75t_L g1801 ( 
.A(n_1767),
.B(n_1768),
.C(n_1730),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1753),
.B(n_1638),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_SL g1803 ( 
.A(n_1726),
.B(n_1647),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1743),
.B(n_1678),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1753),
.B(n_1668),
.Y(n_1805)
);

NAND3xp33_ASAP7_75t_L g1806 ( 
.A(n_1730),
.B(n_1647),
.C(n_1649),
.Y(n_1806)
);

NAND2xp5_ASAP7_75t_L g1807 ( 
.A(n_1721),
.B(n_1613),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1752),
.B(n_1615),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1723),
.B(n_1689),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1721),
.B(n_1613),
.Y(n_1810)
);

AOI221xp5_ASAP7_75t_L g1811 ( 
.A1(n_1726),
.A2(n_1671),
.B1(n_1617),
.B2(n_1684),
.C(n_1683),
.Y(n_1811)
);

NAND2xp5_ASAP7_75t_L g1812 ( 
.A(n_1722),
.B(n_1617),
.Y(n_1812)
);

NAND3xp33_ASAP7_75t_L g1813 ( 
.A(n_1718),
.B(n_1649),
.C(n_1669),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_SL g1814 ( 
.A(n_1754),
.B(n_1695),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1745),
.B(n_1687),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1754),
.B(n_1695),
.Y(n_1816)
);

OAI22xp5_ASAP7_75t_L g1817 ( 
.A1(n_1718),
.A2(n_1705),
.B1(n_1624),
.B2(n_1641),
.Y(n_1817)
);

NAND3xp33_ASAP7_75t_L g1818 ( 
.A(n_1752),
.B(n_1765),
.C(n_1763),
.Y(n_1818)
);

AND2x2_ASAP7_75t_L g1819 ( 
.A(n_1771),
.B(n_1644),
.Y(n_1819)
);

OAI22xp5_ASAP7_75t_L g1820 ( 
.A1(n_1754),
.A2(n_1705),
.B1(n_1556),
.B2(n_1614),
.Y(n_1820)
);

NAND3xp33_ASAP7_75t_L g1821 ( 
.A(n_1763),
.B(n_1669),
.C(n_1679),
.Y(n_1821)
);

NOR2xp33_ASAP7_75t_L g1822 ( 
.A(n_1717),
.B(n_1614),
.Y(n_1822)
);

NAND2xp5_ASAP7_75t_L g1823 ( 
.A(n_1765),
.B(n_1681),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1717),
.B(n_1681),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_L g1825 ( 
.A(n_1719),
.B(n_1667),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1744),
.B(n_1652),
.Y(n_1826)
);

OA21x2_ASAP7_75t_L g1827 ( 
.A1(n_1737),
.A2(n_1631),
.B(n_1661),
.Y(n_1827)
);

AND2x2_ASAP7_75t_L g1828 ( 
.A(n_1744),
.B(n_1652),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1744),
.B(n_1654),
.Y(n_1829)
);

AOI22xp33_ASAP7_75t_L g1830 ( 
.A1(n_1754),
.A2(n_1715),
.B1(n_1705),
.B2(n_1709),
.Y(n_1830)
);

OAI22xp33_ASAP7_75t_SL g1831 ( 
.A1(n_1738),
.A2(n_1700),
.B1(n_1672),
.B2(n_1675),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_SL g1832 ( 
.A(n_1759),
.B(n_1736),
.Y(n_1832)
);

NOR2xp33_ASAP7_75t_L g1833 ( 
.A(n_1719),
.B(n_1481),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_L g1834 ( 
.A(n_1772),
.B(n_1669),
.C(n_1675),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1749),
.B(n_1667),
.Y(n_1835)
);

NOR2xp33_ASAP7_75t_L g1836 ( 
.A(n_1746),
.B(n_1460),
.Y(n_1836)
);

NAND3xp33_ASAP7_75t_L g1837 ( 
.A(n_1772),
.B(n_1679),
.C(n_1672),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_SL g1838 ( 
.A(n_1759),
.B(n_1695),
.Y(n_1838)
);

OAI21xp5_ASAP7_75t_L g1839 ( 
.A1(n_1761),
.A2(n_1699),
.B(n_1694),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1750),
.B(n_1670),
.Y(n_1840)
);

OAI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1775),
.A2(n_1694),
.B1(n_1664),
.B2(n_1665),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_L g1842 ( 
.A(n_1756),
.B(n_1670),
.C(n_1665),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_SL g1843 ( 
.A(n_1759),
.B(n_1695),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1741),
.B(n_1654),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1741),
.B(n_1662),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1750),
.B(n_1664),
.Y(n_1846)
);

NAND3xp33_ASAP7_75t_L g1847 ( 
.A(n_1756),
.B(n_1703),
.C(n_1700),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1728),
.B(n_1703),
.Y(n_1848)
);

NAND2xp33_ASAP7_75t_SL g1849 ( 
.A(n_1759),
.B(n_1642),
.Y(n_1849)
);

NAND2xp5_ASAP7_75t_L g1850 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1761),
.A2(n_1699),
.B(n_1694),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1727),
.Y(n_1852)
);

AND2x4_ASAP7_75t_L g1853 ( 
.A(n_1791),
.B(n_1759),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1852),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1791),
.B(n_1758),
.Y(n_1855)
);

INVx2_ASAP7_75t_L g1856 ( 
.A(n_1852),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1776),
.B(n_1819),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1826),
.Y(n_1858)
);

AND2x4_ASAP7_75t_L g1859 ( 
.A(n_1798),
.B(n_1759),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1784),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1798),
.B(n_1758),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1804),
.B(n_1731),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1804),
.B(n_1773),
.Y(n_1863)
);

AND2x4_ASAP7_75t_L g1864 ( 
.A(n_1832),
.B(n_1731),
.Y(n_1864)
);

AND2x4_ASAP7_75t_L g1865 ( 
.A(n_1832),
.B(n_1731),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1826),
.Y(n_1866)
);

AND2x2_ASAP7_75t_L g1867 ( 
.A(n_1789),
.B(n_1795),
.Y(n_1867)
);

BUFx3_ASAP7_75t_L g1868 ( 
.A(n_1796),
.Y(n_1868)
);

OR2x2_ASAP7_75t_L g1869 ( 
.A(n_1797),
.B(n_1720),
.Y(n_1869)
);

INVx2_ASAP7_75t_L g1870 ( 
.A(n_1828),
.Y(n_1870)
);

BUFx2_ASAP7_75t_L g1871 ( 
.A(n_1849),
.Y(n_1871)
);

AND2x2_ASAP7_75t_SL g1872 ( 
.A(n_1781),
.B(n_1773),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1828),
.Y(n_1873)
);

INVxp67_ASAP7_75t_L g1874 ( 
.A(n_1783),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1829),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1789),
.B(n_1764),
.Y(n_1876)
);

AND2x4_ASAP7_75t_L g1877 ( 
.A(n_1792),
.B(n_1729),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1829),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1844),
.B(n_1734),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1844),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1845),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1779),
.B(n_1805),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1802),
.Y(n_1883)
);

INVx3_ASAP7_75t_L g1884 ( 
.A(n_1827),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1835),
.B(n_1734),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1840),
.B(n_1846),
.Y(n_1886)
);

INVx2_ASAP7_75t_SL g1887 ( 
.A(n_1809),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1842),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1818),
.Y(n_1889)
);

INVx1_ASAP7_75t_L g1890 ( 
.A(n_1837),
.Y(n_1890)
);

AND2x2_ASAP7_75t_L g1891 ( 
.A(n_1781),
.B(n_1729),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1823),
.B(n_1735),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1847),
.Y(n_1893)
);

AND2x4_ASAP7_75t_L g1894 ( 
.A(n_1792),
.B(n_1729),
.Y(n_1894)
);

INVx2_ASAP7_75t_SL g1895 ( 
.A(n_1807),
.Y(n_1895)
);

OR2x2_ASAP7_75t_L g1896 ( 
.A(n_1815),
.B(n_1769),
.Y(n_1896)
);

INVx1_ASAP7_75t_L g1897 ( 
.A(n_1848),
.Y(n_1897)
);

AND2x2_ASAP7_75t_L g1898 ( 
.A(n_1803),
.B(n_1755),
.Y(n_1898)
);

INVx3_ASAP7_75t_L g1899 ( 
.A(n_1827),
.Y(n_1899)
);

INVx1_ASAP7_75t_L g1900 ( 
.A(n_1850),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1825),
.Y(n_1901)
);

AND2x4_ASAP7_75t_SL g1902 ( 
.A(n_1794),
.B(n_1738),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1803),
.B(n_1814),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1814),
.B(n_1755),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1834),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1849),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1827),
.Y(n_1907)
);

AND2x4_ASAP7_75t_L g1908 ( 
.A(n_1816),
.B(n_1736),
.Y(n_1908)
);

NAND2xp5_ASAP7_75t_L g1909 ( 
.A(n_1821),
.B(n_1734),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1890),
.B(n_1810),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1890),
.B(n_1812),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1872),
.B(n_1816),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1856),
.Y(n_1913)
);

OR2x2_ASAP7_75t_L g1914 ( 
.A(n_1905),
.B(n_1893),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1870),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1870),
.Y(n_1916)
);

NAND2xp67_ASAP7_75t_SL g1917 ( 
.A(n_1891),
.B(n_1811),
.Y(n_1917)
);

INVx2_ASAP7_75t_L g1918 ( 
.A(n_1856),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1870),
.Y(n_1919)
);

AND2x2_ASAP7_75t_L g1920 ( 
.A(n_1872),
.B(n_1839),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1872),
.B(n_1851),
.Y(n_1921)
);

INVx1_ASAP7_75t_L g1922 ( 
.A(n_1854),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1867),
.B(n_1838),
.Y(n_1923)
);

NOR2x1_ASAP7_75t_SL g1924 ( 
.A(n_1903),
.B(n_1790),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1868),
.B(n_1778),
.Y(n_1925)
);

AND2x2_ASAP7_75t_L g1926 ( 
.A(n_1867),
.B(n_1838),
.Y(n_1926)
);

NAND2xp5_ASAP7_75t_L g1927 ( 
.A(n_1868),
.B(n_1824),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1880),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1880),
.Y(n_1929)
);

INVx1_ASAP7_75t_L g1930 ( 
.A(n_1858),
.Y(n_1930)
);

AND2x2_ASAP7_75t_L g1931 ( 
.A(n_1853),
.B(n_1859),
.Y(n_1931)
);

INVx1_ASAP7_75t_L g1932 ( 
.A(n_1858),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_L g1933 ( 
.A(n_1868),
.B(n_1782),
.Y(n_1933)
);

OA211x2_ASAP7_75t_L g1934 ( 
.A1(n_1909),
.A2(n_1801),
.B(n_1799),
.C(n_1813),
.Y(n_1934)
);

AND2x2_ASAP7_75t_SL g1935 ( 
.A(n_1871),
.B(n_1775),
.Y(n_1935)
);

OAI31xp33_ASAP7_75t_L g1936 ( 
.A1(n_1889),
.A2(n_1777),
.A3(n_1800),
.B(n_1788),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1866),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1856),
.Y(n_1938)
);

NAND4xp25_ASAP7_75t_L g1939 ( 
.A(n_1905),
.B(n_1785),
.C(n_1780),
.D(n_1786),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1866),
.Y(n_1940)
);

NAND3xp33_ASAP7_75t_L g1941 ( 
.A(n_1893),
.B(n_1787),
.C(n_1806),
.Y(n_1941)
);

OR2x2_ASAP7_75t_L g1942 ( 
.A(n_1888),
.B(n_1843),
.Y(n_1942)
);

INVx2_ASAP7_75t_L g1943 ( 
.A(n_1881),
.Y(n_1943)
);

NAND4xp25_ASAP7_75t_L g1944 ( 
.A(n_1888),
.B(n_1793),
.C(n_1830),
.D(n_1808),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_L g1945 ( 
.A(n_1883),
.B(n_1836),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_L g1946 ( 
.A(n_1874),
.B(n_1831),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1873),
.Y(n_1947)
);

INVx1_ASAP7_75t_L g1948 ( 
.A(n_1873),
.Y(n_1948)
);

BUFx2_ASAP7_75t_L g1949 ( 
.A(n_1871),
.Y(n_1949)
);

INVx1_ASAP7_75t_SL g1950 ( 
.A(n_1882),
.Y(n_1950)
);

AND2x4_ASAP7_75t_L g1951 ( 
.A(n_1891),
.B(n_1853),
.Y(n_1951)
);

OR2x2_ASAP7_75t_L g1952 ( 
.A(n_1909),
.B(n_1843),
.Y(n_1952)
);

AND2x2_ASAP7_75t_L g1953 ( 
.A(n_1853),
.B(n_1738),
.Y(n_1953)
);

OR2x2_ASAP7_75t_L g1954 ( 
.A(n_1869),
.B(n_1737),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1875),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1875),
.Y(n_1956)
);

INVx1_ASAP7_75t_L g1957 ( 
.A(n_1854),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1878),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1901),
.B(n_1735),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1881),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_L g1961 ( 
.A(n_1901),
.B(n_1740),
.Y(n_1961)
);

NOR2xp67_ASAP7_75t_SL g1962 ( 
.A(n_1903),
.B(n_1736),
.Y(n_1962)
);

OR2x2_ASAP7_75t_L g1963 ( 
.A(n_1869),
.B(n_1762),
.Y(n_1963)
);

INVx1_ASAP7_75t_L g1964 ( 
.A(n_1878),
.Y(n_1964)
);

INVx1_ASAP7_75t_L g1965 ( 
.A(n_1879),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1895),
.B(n_1740),
.Y(n_1966)
);

OR2x2_ASAP7_75t_L g1967 ( 
.A(n_1896),
.B(n_1762),
.Y(n_1967)
);

OR2x2_ASAP7_75t_L g1968 ( 
.A(n_1914),
.B(n_1879),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1922),
.Y(n_1969)
);

NOR2xp67_ASAP7_75t_L g1970 ( 
.A(n_1912),
.B(n_1853),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1922),
.Y(n_1971)
);

AND2x2_ASAP7_75t_L g1972 ( 
.A(n_1935),
.B(n_1906),
.Y(n_1972)
);

BUFx2_ASAP7_75t_L g1973 ( 
.A(n_1949),
.Y(n_1973)
);

OR2x2_ASAP7_75t_L g1974 ( 
.A(n_1914),
.B(n_1857),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_L g1975 ( 
.A(n_1950),
.B(n_1897),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1957),
.Y(n_1976)
);

AND2x2_ASAP7_75t_L g1977 ( 
.A(n_1935),
.B(n_1906),
.Y(n_1977)
);

AND2x2_ASAP7_75t_L g1978 ( 
.A(n_1912),
.B(n_1859),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1917),
.B(n_1822),
.Y(n_1979)
);

NAND2xp5_ASAP7_75t_L g1980 ( 
.A(n_1910),
.B(n_1897),
.Y(n_1980)
);

NOR2xp67_ASAP7_75t_L g1981 ( 
.A(n_1941),
.B(n_1859),
.Y(n_1981)
);

NOR2xp33_ASAP7_75t_SL g1982 ( 
.A(n_1936),
.B(n_1820),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1911),
.B(n_1925),
.Y(n_1983)
);

INVxp67_ASAP7_75t_SL g1984 ( 
.A(n_1924),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1957),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1928),
.Y(n_1986)
);

AOI22xp5_ASAP7_75t_L g1987 ( 
.A1(n_1934),
.A2(n_1902),
.B1(n_1817),
.B2(n_1908),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1929),
.Y(n_1988)
);

OAI21xp33_ASAP7_75t_L g1989 ( 
.A1(n_1939),
.A2(n_1921),
.B(n_1920),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1930),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_L g1991 ( 
.A(n_1944),
.B(n_1859),
.Y(n_1991)
);

INVx1_ASAP7_75t_L g1992 ( 
.A(n_1932),
.Y(n_1992)
);

OR2x2_ASAP7_75t_L g1993 ( 
.A(n_1946),
.B(n_1857),
.Y(n_1993)
);

INVx1_ASAP7_75t_L g1994 ( 
.A(n_1937),
.Y(n_1994)
);

INVx1_ASAP7_75t_SL g1995 ( 
.A(n_1949),
.Y(n_1995)
);

INVx1_ASAP7_75t_L g1996 ( 
.A(n_1940),
.Y(n_1996)
);

NAND4xp25_ASAP7_75t_SL g1997 ( 
.A(n_1920),
.B(n_1861),
.C(n_1863),
.D(n_1855),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1921),
.A2(n_1902),
.B1(n_1908),
.B2(n_1877),
.Y(n_1998)
);

OR2x2_ASAP7_75t_L g1999 ( 
.A(n_1952),
.B(n_1896),
.Y(n_1999)
);

INVx2_ASAP7_75t_L g2000 ( 
.A(n_1913),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1947),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1931),
.B(n_1876),
.Y(n_2002)
);

NOR2xp33_ASAP7_75t_L g2003 ( 
.A(n_1933),
.B(n_1833),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1948),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1931),
.B(n_1876),
.Y(n_2005)
);

INVx1_ASAP7_75t_L g2006 ( 
.A(n_1955),
.Y(n_2006)
);

INVx2_ASAP7_75t_L g2007 ( 
.A(n_1913),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_L g2008 ( 
.A(n_1942),
.B(n_1895),
.Y(n_2008)
);

INVx1_ASAP7_75t_L g2009 ( 
.A(n_1956),
.Y(n_2009)
);

INVxp67_ASAP7_75t_L g2010 ( 
.A(n_1942),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1927),
.B(n_1900),
.Y(n_2011)
);

AND2x2_ASAP7_75t_L g2012 ( 
.A(n_1924),
.B(n_1855),
.Y(n_2012)
);

AND2x4_ASAP7_75t_SL g2013 ( 
.A(n_1951),
.B(n_1908),
.Y(n_2013)
);

AND2x2_ASAP7_75t_L g2014 ( 
.A(n_1951),
.B(n_1861),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1952),
.B(n_1900),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1958),
.Y(n_2016)
);

INVx1_ASAP7_75t_L g2017 ( 
.A(n_1964),
.Y(n_2017)
);

AOI22xp33_ASAP7_75t_L g2018 ( 
.A1(n_1945),
.A2(n_1902),
.B1(n_1715),
.B2(n_1666),
.Y(n_2018)
);

AND2x4_ASAP7_75t_L g2019 ( 
.A(n_1951),
.B(n_1908),
.Y(n_2019)
);

BUFx2_ASAP7_75t_L g2020 ( 
.A(n_1917),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1966),
.A2(n_1775),
.B1(n_1894),
.B2(n_1877),
.Y(n_2021)
);

INVx1_ASAP7_75t_L g2022 ( 
.A(n_1969),
.Y(n_2022)
);

AND2x2_ASAP7_75t_L g2023 ( 
.A(n_2012),
.B(n_1953),
.Y(n_2023)
);

OAI22xp5_ASAP7_75t_L g2024 ( 
.A1(n_2020),
.A2(n_1926),
.B1(n_1923),
.B2(n_1894),
.Y(n_2024)
);

NOR2x1_ASAP7_75t_L g2025 ( 
.A(n_1979),
.B(n_1981),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_2012),
.B(n_1953),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1971),
.Y(n_2027)
);

INVx2_ASAP7_75t_L g2028 ( 
.A(n_1973),
.Y(n_2028)
);

BUFx8_ASAP7_75t_SL g2029 ( 
.A(n_1972),
.Y(n_2029)
);

OAI22xp5_ASAP7_75t_L g2030 ( 
.A1(n_1984),
.A2(n_1926),
.B1(n_1923),
.B2(n_1894),
.Y(n_2030)
);

AOI22xp33_ASAP7_75t_L g2031 ( 
.A1(n_1982),
.A2(n_1989),
.B1(n_1991),
.B2(n_1997),
.Y(n_2031)
);

INVx1_ASAP7_75t_SL g2032 ( 
.A(n_1972),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_2013),
.B(n_1962),
.Y(n_2033)
);

INVx2_ASAP7_75t_L g2034 ( 
.A(n_2000),
.Y(n_2034)
);

OAI21xp33_ASAP7_75t_SL g2035 ( 
.A1(n_1970),
.A2(n_1965),
.B(n_1916),
.Y(n_2035)
);

INVx1_ASAP7_75t_SL g2036 ( 
.A(n_1977),
.Y(n_2036)
);

NAND2xp5_ASAP7_75t_L g2037 ( 
.A(n_1983),
.B(n_1959),
.Y(n_2037)
);

INVx1_ASAP7_75t_L g2038 ( 
.A(n_1976),
.Y(n_2038)
);

OAI21xp33_ASAP7_75t_SL g2039 ( 
.A1(n_1991),
.A2(n_1919),
.B(n_1915),
.Y(n_2039)
);

HB1xp67_ASAP7_75t_L g2040 ( 
.A(n_1995),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_L g2041 ( 
.A(n_2010),
.B(n_1961),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1985),
.Y(n_2042)
);

INVx2_ASAP7_75t_L g2043 ( 
.A(n_2000),
.Y(n_2043)
);

INVx4_ASAP7_75t_L g2044 ( 
.A(n_2013),
.Y(n_2044)
);

NOR2xp33_ASAP7_75t_L g2045 ( 
.A(n_2003),
.B(n_1993),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1986),
.Y(n_2046)
);

BUFx6f_ASAP7_75t_L g2047 ( 
.A(n_2007),
.Y(n_2047)
);

INVx1_ASAP7_75t_L g2048 ( 
.A(n_1988),
.Y(n_2048)
);

OR2x2_ASAP7_75t_L g2049 ( 
.A(n_1974),
.B(n_1954),
.Y(n_2049)
);

AND2x2_ASAP7_75t_L g2050 ( 
.A(n_1977),
.B(n_1962),
.Y(n_2050)
);

INVx1_ASAP7_75t_SL g2051 ( 
.A(n_2019),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_L g2052 ( 
.A(n_2003),
.B(n_1898),
.Y(n_2052)
);

AOI22xp33_ASAP7_75t_L g2053 ( 
.A1(n_2019),
.A2(n_1738),
.B1(n_1894),
.B2(n_1877),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1990),
.Y(n_2054)
);

OR2x2_ASAP7_75t_L g2055 ( 
.A(n_1974),
.B(n_1954),
.Y(n_2055)
);

NAND2xp33_ASAP7_75t_L g2056 ( 
.A(n_1987),
.B(n_1841),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1978),
.B(n_1943),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1992),
.Y(n_2058)
);

INVx1_ASAP7_75t_L g2059 ( 
.A(n_1994),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1996),
.Y(n_2060)
);

INVx3_ASAP7_75t_SL g2061 ( 
.A(n_2019),
.Y(n_2061)
);

INVx1_ASAP7_75t_L g2062 ( 
.A(n_2001),
.Y(n_2062)
);

AOI21xp33_ASAP7_75t_SL g2063 ( 
.A1(n_2031),
.A2(n_2021),
.B(n_1998),
.Y(n_2063)
);

OAI31xp33_ASAP7_75t_L g2064 ( 
.A1(n_2045),
.A2(n_2018),
.A3(n_1978),
.B(n_2014),
.Y(n_2064)
);

AOI211xp5_ASAP7_75t_L g2065 ( 
.A1(n_2056),
.A2(n_2008),
.B(n_2015),
.C(n_1975),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_2032),
.B(n_2014),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_2036),
.B(n_1980),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_2040),
.B(n_2002),
.Y(n_2068)
);

HB1xp67_ASAP7_75t_L g2069 ( 
.A(n_2028),
.Y(n_2069)
);

INVx1_ASAP7_75t_L g2070 ( 
.A(n_2022),
.Y(n_2070)
);

AND2x2_ASAP7_75t_L g2071 ( 
.A(n_2025),
.B(n_2002),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_2022),
.Y(n_2072)
);

NAND4xp25_ASAP7_75t_L g2073 ( 
.A(n_2051),
.B(n_2028),
.C(n_2050),
.D(n_2044),
.Y(n_2073)
);

OAI32xp33_ASAP7_75t_L g2074 ( 
.A1(n_2035),
.A2(n_1968),
.A3(n_1999),
.B1(n_2018),
.B2(n_2009),
.Y(n_2074)
);

NAND4xp75_ASAP7_75t_L g2075 ( 
.A(n_2039),
.B(n_2005),
.C(n_2006),
.D(n_2004),
.Y(n_2075)
);

INVx1_ASAP7_75t_L g2076 ( 
.A(n_2027),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_2027),
.Y(n_2077)
);

INVx1_ASAP7_75t_L g2078 ( 
.A(n_2038),
.Y(n_2078)
);

OAI322xp33_ASAP7_75t_L g2079 ( 
.A1(n_2046),
.A2(n_1968),
.A3(n_1999),
.B1(n_2016),
.B2(n_2017),
.C1(n_2011),
.C2(n_2007),
.Y(n_2079)
);

NOR2xp33_ASAP7_75t_R g2080 ( 
.A(n_2056),
.B(n_1460),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_2029),
.B(n_2005),
.Y(n_2081)
);

A2O1A1Ixp33_ASAP7_75t_L g2082 ( 
.A1(n_2050),
.A2(n_1865),
.B(n_1864),
.C(n_1877),
.Y(n_2082)
);

INVx2_ASAP7_75t_SL g2083 ( 
.A(n_2061),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_2044),
.B(n_1864),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2038),
.Y(n_2085)
);

AOI22xp33_ASAP7_75t_L g2086 ( 
.A1(n_2044),
.A2(n_1738),
.B1(n_1774),
.B2(n_1725),
.Y(n_2086)
);

A2O1A1Ixp33_ASAP7_75t_L g2087 ( 
.A1(n_2052),
.A2(n_1865),
.B(n_1864),
.C(n_1770),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_2042),
.Y(n_2088)
);

INVx1_ASAP7_75t_L g2089 ( 
.A(n_2042),
.Y(n_2089)
);

NOR2xp33_ASAP7_75t_L g2090 ( 
.A(n_2037),
.B(n_1886),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2048),
.Y(n_2091)
);

INVx1_ASAP7_75t_L g2092 ( 
.A(n_2048),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_2061),
.B(n_1943),
.Y(n_2093)
);

AOI22xp33_ASAP7_75t_L g2094 ( 
.A1(n_2064),
.A2(n_2062),
.B1(n_2061),
.B2(n_2024),
.Y(n_2094)
);

INVx1_ASAP7_75t_L g2095 ( 
.A(n_2069),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2083),
.B(n_2023),
.Y(n_2096)
);

INVx1_ASAP7_75t_SL g2097 ( 
.A(n_2071),
.Y(n_2097)
);

NAND2x1_ASAP7_75t_L g2098 ( 
.A(n_2071),
.B(n_2033),
.Y(n_2098)
);

AND2x2_ASAP7_75t_L g2099 ( 
.A(n_2081),
.B(n_2023),
.Y(n_2099)
);

INVx1_ASAP7_75t_L g2100 ( 
.A(n_2070),
.Y(n_2100)
);

AOI22xp5_ASAP7_75t_L g2101 ( 
.A1(n_2073),
.A2(n_2083),
.B1(n_2075),
.B2(n_2084),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2093),
.B(n_2026),
.Y(n_2102)
);

INVx1_ASAP7_75t_SL g2103 ( 
.A(n_2080),
.Y(n_2103)
);

NAND2xp5_ASAP7_75t_L g2104 ( 
.A(n_2068),
.B(n_2026),
.Y(n_2104)
);

OR2x2_ASAP7_75t_L g2105 ( 
.A(n_2066),
.B(n_2041),
.Y(n_2105)
);

OR2x2_ASAP7_75t_L g2106 ( 
.A(n_2067),
.B(n_2049),
.Y(n_2106)
);

AND2x2_ASAP7_75t_L g2107 ( 
.A(n_2093),
.B(n_2033),
.Y(n_2107)
);

NAND2x1_ASAP7_75t_SL g2108 ( 
.A(n_2091),
.B(n_2057),
.Y(n_2108)
);

INVx1_ASAP7_75t_L g2109 ( 
.A(n_2072),
.Y(n_2109)
);

OR2x2_ASAP7_75t_L g2110 ( 
.A(n_2090),
.B(n_2049),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2084),
.B(n_2057),
.Y(n_2111)
);

NAND2xp33_ASAP7_75t_SL g2112 ( 
.A(n_2080),
.B(n_2030),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_L g2113 ( 
.A(n_2065),
.B(n_2054),
.Y(n_2113)
);

OR2x6_ASAP7_75t_L g2114 ( 
.A(n_2075),
.B(n_1479),
.Y(n_2114)
);

AND2x2_ASAP7_75t_SL g2115 ( 
.A(n_2092),
.B(n_2047),
.Y(n_2115)
);

AND2x2_ASAP7_75t_L g2116 ( 
.A(n_2082),
.B(n_2053),
.Y(n_2116)
);

OAI21xp5_ASAP7_75t_L g2117 ( 
.A1(n_2094),
.A2(n_2063),
.B(n_2074),
.Y(n_2117)
);

AOI221x1_ASAP7_75t_L g2118 ( 
.A1(n_2095),
.A2(n_2089),
.B1(n_2088),
.B2(n_2076),
.C(n_2077),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_L g2119 ( 
.A(n_2097),
.B(n_2078),
.Y(n_2119)
);

OAI211xp5_ASAP7_75t_SL g2120 ( 
.A1(n_2094),
.A2(n_2082),
.B(n_2085),
.C(n_2087),
.Y(n_2120)
);

OAI21xp5_ASAP7_75t_SL g2121 ( 
.A1(n_2101),
.A2(n_2086),
.B(n_2087),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_2115),
.Y(n_2122)
);

OAI22xp33_ASAP7_75t_L g2123 ( 
.A1(n_2114),
.A2(n_2055),
.B1(n_2047),
.B2(n_2054),
.Y(n_2123)
);

NOR3xp33_ASAP7_75t_L g2124 ( 
.A(n_2113),
.B(n_2079),
.C(n_2059),
.Y(n_2124)
);

AOI322xp5_ASAP7_75t_L g2125 ( 
.A1(n_2112),
.A2(n_2060),
.A3(n_2059),
.B1(n_2058),
.B2(n_2034),
.C1(n_2043),
.C2(n_2047),
.Y(n_2125)
);

OAI211xp5_ASAP7_75t_L g2126 ( 
.A1(n_2108),
.A2(n_2060),
.B(n_2058),
.C(n_2043),
.Y(n_2126)
);

AOI31xp33_ASAP7_75t_L g2127 ( 
.A1(n_2103),
.A2(n_2055),
.A3(n_2034),
.B(n_1865),
.Y(n_2127)
);

AOI221xp5_ASAP7_75t_L g2128 ( 
.A1(n_2112),
.A2(n_2047),
.B1(n_1884),
.B2(n_1899),
.C(n_1907),
.Y(n_2128)
);

AOI22xp33_ASAP7_75t_L g2129 ( 
.A1(n_2114),
.A2(n_2099),
.B1(n_2116),
.B2(n_2107),
.Y(n_2129)
);

NAND5xp2_ASAP7_75t_L g2130 ( 
.A(n_2099),
.B(n_1863),
.C(n_1904),
.D(n_1898),
.E(n_1711),
.Y(n_2130)
);

OAI221xp5_ASAP7_75t_SL g2131 ( 
.A1(n_2114),
.A2(n_1963),
.B1(n_1884),
.B2(n_1899),
.C(n_1907),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_SL g2132 ( 
.A1(n_2115),
.A2(n_2047),
.B1(n_1598),
.B2(n_1605),
.Y(n_2132)
);

NAND4xp25_ASAP7_75t_L g2133 ( 
.A(n_2117),
.B(n_2096),
.C(n_2104),
.D(n_2105),
.Y(n_2133)
);

NOR2x1_ASAP7_75t_L g2134 ( 
.A(n_2122),
.B(n_2098),
.Y(n_2134)
);

OAI322xp33_ASAP7_75t_L g2135 ( 
.A1(n_2123),
.A2(n_2109),
.A3(n_2100),
.B1(n_2106),
.B2(n_2110),
.C1(n_2116),
.C2(n_2111),
.Y(n_2135)
);

NAND2xp5_ASAP7_75t_L g2136 ( 
.A(n_2129),
.B(n_2107),
.Y(n_2136)
);

AND2x2_ASAP7_75t_L g2137 ( 
.A(n_2125),
.B(n_2102),
.Y(n_2137)
);

NOR3xp33_ASAP7_75t_L g2138 ( 
.A(n_2120),
.B(n_2111),
.C(n_2102),
.Y(n_2138)
);

NOR2x1_ASAP7_75t_SL g2139 ( 
.A(n_2126),
.B(n_1963),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2119),
.Y(n_2140)
);

NOR2x1p5_ASAP7_75t_L g2141 ( 
.A(n_2127),
.B(n_1595),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_2118),
.Y(n_2142)
);

OAI211xp5_ASAP7_75t_SL g2143 ( 
.A1(n_2124),
.A2(n_1558),
.B(n_1967),
.C(n_1884),
.Y(n_2143)
);

OA22x2_ASAP7_75t_L g2144 ( 
.A1(n_2121),
.A2(n_1864),
.B1(n_1865),
.B2(n_1960),
.Y(n_2144)
);

NOR3xp33_ASAP7_75t_SL g2145 ( 
.A(n_2132),
.B(n_2131),
.C(n_2128),
.Y(n_2145)
);

AOI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2124),
.A2(n_1598),
.B1(n_1595),
.B2(n_1558),
.Y(n_2146)
);

NOR2xp67_ASAP7_75t_L g2147 ( 
.A(n_2130),
.B(n_1918),
.Y(n_2147)
);

AOI211xp5_ASAP7_75t_L g2148 ( 
.A1(n_2135),
.A2(n_1967),
.B(n_1899),
.C(n_1884),
.Y(n_2148)
);

NAND2xp5_ASAP7_75t_L g2149 ( 
.A(n_2138),
.B(n_1960),
.Y(n_2149)
);

OAI211xp5_ASAP7_75t_L g2150 ( 
.A1(n_2146),
.A2(n_1899),
.B(n_1498),
.C(n_1470),
.Y(n_2150)
);

NOR2x1_ASAP7_75t_L g2151 ( 
.A(n_2142),
.B(n_2134),
.Y(n_2151)
);

NAND2xp5_ASAP7_75t_L g2152 ( 
.A(n_2137),
.B(n_1918),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_L g2153 ( 
.A(n_2146),
.B(n_1470),
.C(n_1498),
.Y(n_2153)
);

OR3x1_ASAP7_75t_L g2154 ( 
.A(n_2143),
.B(n_1716),
.C(n_1712),
.Y(n_2154)
);

AOI22xp5_ASAP7_75t_L g2155 ( 
.A1(n_2151),
.A2(n_2136),
.B1(n_2133),
.B2(n_2144),
.Y(n_2155)
);

AOI22xp5_ASAP7_75t_L g2156 ( 
.A1(n_2154),
.A2(n_2141),
.B1(n_2140),
.B2(n_2147),
.Y(n_2156)
);

HB1xp67_ASAP7_75t_L g2157 ( 
.A(n_2149),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_2152),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2153),
.Y(n_2159)
);

INVx1_ASAP7_75t_L g2160 ( 
.A(n_2148),
.Y(n_2160)
);

AOI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_2150),
.A2(n_2145),
.B1(n_2139),
.B2(n_1938),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2151),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2162),
.Y(n_2163)
);

NAND3xp33_ASAP7_75t_L g2164 ( 
.A(n_2155),
.B(n_1594),
.C(n_1907),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_2158),
.B(n_1938),
.Y(n_2165)
);

NOR2x1p5_ASAP7_75t_L g2166 ( 
.A(n_2159),
.B(n_1585),
.Y(n_2166)
);

HB1xp67_ASAP7_75t_L g2167 ( 
.A(n_2157),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2160),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2163),
.B(n_2167),
.Y(n_2169)
);

INVx1_ASAP7_75t_L g2170 ( 
.A(n_2166),
.Y(n_2170)
);

INVxp67_ASAP7_75t_L g2171 ( 
.A(n_2164),
.Y(n_2171)
);

XOR2xp5_ASAP7_75t_L g2172 ( 
.A(n_2169),
.B(n_2168),
.Y(n_2172)
);

NAND4xp25_ASAP7_75t_L g2173 ( 
.A(n_2172),
.B(n_2169),
.C(n_2171),
.D(n_2170),
.Y(n_2173)
);

HB1xp67_ASAP7_75t_L g2174 ( 
.A(n_2173),
.Y(n_2174)
);

AOI22xp5_ASAP7_75t_L g2175 ( 
.A1(n_2173),
.A2(n_2161),
.B1(n_2156),
.B2(n_2165),
.Y(n_2175)
);

AO22x1_ASAP7_75t_L g2176 ( 
.A1(n_2174),
.A2(n_1585),
.B1(n_1698),
.B2(n_1704),
.Y(n_2176)
);

OAI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_2175),
.A2(n_1886),
.B(n_1892),
.Y(n_2177)
);

AOI21xp5_ASAP7_75t_L g2178 ( 
.A1(n_2176),
.A2(n_1887),
.B(n_1885),
.Y(n_2178)
);

NOR2x1_ASAP7_75t_L g2179 ( 
.A(n_2177),
.B(n_1585),
.Y(n_2179)
);

AOI221xp5_ASAP7_75t_L g2180 ( 
.A1(n_2178),
.A2(n_1887),
.B1(n_1862),
.B2(n_1713),
.C(n_1711),
.Y(n_2180)
);

AOI22xp5_ASAP7_75t_L g2181 ( 
.A1(n_2180),
.A2(n_2179),
.B1(n_1860),
.B2(n_1862),
.Y(n_2181)
);

OAI221xp5_ASAP7_75t_R g2182 ( 
.A1(n_2181),
.A2(n_1860),
.B1(n_1706),
.B2(n_1862),
.C(n_1704),
.Y(n_2182)
);

AOI211xp5_ASAP7_75t_L g2183 ( 
.A1(n_2182),
.A2(n_1585),
.B(n_1698),
.C(n_1642),
.Y(n_2183)
);


endmodule