module fake_netlist_6_281_n_195 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_195);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_195;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_193;
wire n_147;
wire n_154;
wire n_191;
wire n_88;
wire n_98;
wire n_113;
wire n_63;
wire n_39;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_153;
wire n_168;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_160;
wire n_90;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_32;
wire n_130;
wire n_99;
wire n_66;
wire n_78;
wire n_84;
wire n_85;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_67;
wire n_37;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_97;
wire n_94;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_194;
wire n_171;
wire n_192;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_30),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_7),
.Y(n_36)
);

NOR2xp67_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_14),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

INVxp67_ASAP7_75t_SL g46 ( 
.A(n_15),
.Y(n_46)
);

INVxp67_ASAP7_75t_SL g47 ( 
.A(n_10),
.Y(n_47)
);

INVxp67_ASAP7_75t_SL g48 ( 
.A(n_2),
.Y(n_48)
);

BUFx2_ASAP7_75t_L g49 ( 
.A(n_10),
.Y(n_49)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx16_ASAP7_75t_R g51 ( 
.A(n_25),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_5),
.Y(n_52)
);

INVx4_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_51),
.B(n_1),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_38),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_42),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_45),
.Y(n_72)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_53),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g77 ( 
.A(n_74),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

AO22x2_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_48),
.B1(n_46),
.B2(n_50),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_57),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

AO22x2_ASAP7_75t_L g89 ( 
.A1(n_73),
.A2(n_50),
.B1(n_53),
.B2(n_51),
.Y(n_89)
);

CKINVDCx5p33_ASAP7_75t_R g90 ( 
.A(n_74),
.Y(n_90)
);

AO22x2_ASAP7_75t_L g91 ( 
.A1(n_72),
.A2(n_37),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_81),
.B(n_60),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_74),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_88),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_77),
.B(n_68),
.Y(n_96)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_78),
.A2(n_55),
.B(n_72),
.C(n_63),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_79),
.B(n_55),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_36),
.B1(n_32),
.B2(n_71),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_75),
.B(n_63),
.Y(n_102)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_82),
.B(n_68),
.Y(n_103)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_71),
.B(n_60),
.C(n_63),
.Y(n_104)
);

INVxp67_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_75),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_89),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_89),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_99),
.A2(n_68),
.B(n_87),
.C(n_86),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_101),
.A2(n_102),
.B(n_75),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_98),
.Y(n_111)
);

A2O1A1Ixp33_ASAP7_75t_L g112 ( 
.A1(n_105),
.A2(n_92),
.B(n_100),
.C(n_103),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

AND2x4_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

NAND2xp33_ASAP7_75t_L g115 ( 
.A(n_106),
.B(n_75),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g116 ( 
.A(n_111),
.B(n_100),
.Y(n_116)
);

AND2x4_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_103),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_106),
.B(n_80),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_114),
.B(n_111),
.Y(n_119)
);

A2O1A1Ixp33_ASAP7_75t_L g120 ( 
.A1(n_112),
.A2(n_104),
.B(n_108),
.C(n_37),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_113),
.Y(n_121)
);

BUFx12f_ASAP7_75t_L g122 ( 
.A(n_116),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_117),
.Y(n_123)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_121),
.Y(n_124)
);

NAND3xp33_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_74),
.C(n_118),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_121),
.Y(n_126)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_119),
.Y(n_127)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_123),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

INVxp67_ASAP7_75t_SL g130 ( 
.A(n_123),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_123),
.Y(n_131)
);

NOR3xp33_ASAP7_75t_L g132 ( 
.A(n_122),
.B(n_118),
.C(n_117),
.Y(n_132)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_122),
.A2(n_115),
.B(n_110),
.Y(n_133)
);

INVx2_ASAP7_75t_SL g134 ( 
.A(n_119),
.Y(n_134)
);

OR2x6_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_114),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_134),
.B(n_89),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_132),
.A2(n_80),
.B1(n_91),
.B2(n_33),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_129),
.B(n_80),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_129),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_124),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_127),
.A2(n_91),
.B1(n_52),
.B2(n_39),
.Y(n_141)
);

HB1xp67_ASAP7_75t_L g142 ( 
.A(n_134),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_140),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_142),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g146 ( 
.A(n_139),
.B(n_135),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_138),
.B(n_127),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_127),
.Y(n_148)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_125),
.Y(n_149)
);

BUFx2_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_127),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_144),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_146),
.B(n_126),
.Y(n_154)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_146),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_143),
.Y(n_156)
);

INVx1_ASAP7_75t_SL g157 ( 
.A(n_145),
.Y(n_157)
);

OAI221xp5_ASAP7_75t_L g158 ( 
.A1(n_152),
.A2(n_62),
.B1(n_70),
.B2(n_69),
.C(n_65),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_148),
.B(n_124),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_147),
.B(n_151),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_126),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_156),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_149),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_149),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_154),
.B(n_130),
.Y(n_165)
);

HB1xp67_ASAP7_75t_L g166 ( 
.A(n_153),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_58),
.Y(n_167)
);

NAND4xp75_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_58),
.C(n_70),
.D(n_69),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_159),
.B(n_131),
.Y(n_170)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_166),
.Y(n_171)
);

OAI21x1_ASAP7_75t_SL g172 ( 
.A1(n_163),
.A2(n_61),
.B(n_65),
.Y(n_172)
);

AOI221xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_160),
.B1(n_158),
.B2(n_61),
.C(n_62),
.Y(n_173)
);

NOR3xp33_ASAP7_75t_L g174 ( 
.A(n_167),
.B(n_56),
.C(n_161),
.Y(n_174)
);

NAND3x1_ASAP7_75t_L g175 ( 
.A(n_164),
.B(n_161),
.C(n_56),
.Y(n_175)
);

NOR2x1_ASAP7_75t_L g176 ( 
.A(n_162),
.B(n_169),
.Y(n_176)
);

OAI322xp33_ASAP7_75t_L g177 ( 
.A1(n_170),
.A2(n_64),
.A3(n_66),
.B1(n_6),
.B2(n_8),
.C1(n_9),
.C2(n_1),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_165),
.A2(n_131),
.B(n_128),
.Y(n_178)
);

AND3x4_ASAP7_75t_L g179 ( 
.A(n_174),
.B(n_168),
.C(n_128),
.Y(n_179)
);

NOR2x1_ASAP7_75t_L g180 ( 
.A(n_176),
.B(n_166),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_171),
.Y(n_181)
);

AOI221xp5_ASAP7_75t_L g182 ( 
.A1(n_177),
.A2(n_64),
.B1(n_66),
.B2(n_83),
.C(n_84),
.Y(n_182)
);

NAND5xp2_ASAP7_75t_L g183 ( 
.A(n_173),
.B(n_85),
.C(n_8),
.D(n_9),
.E(n_11),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_175),
.A2(n_66),
.B1(n_64),
.B2(n_5),
.Y(n_184)
);

NOR2xp67_ASAP7_75t_L g185 ( 
.A(n_178),
.B(n_11),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_172),
.Y(n_186)
);

NAND5xp2_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_16),
.C(n_19),
.D(n_21),
.E(n_23),
.Y(n_187)
);

AOI221xp5_ASAP7_75t_L g188 ( 
.A1(n_184),
.A2(n_66),
.B1(n_93),
.B2(n_95),
.C(n_29),
.Y(n_188)
);

AOI322xp5_ASAP7_75t_L g189 ( 
.A1(n_180),
.A2(n_66),
.A3(n_27),
.B1(n_28),
.B2(n_31),
.C1(n_26),
.C2(n_93),
.Y(n_189)
);

AOI322xp5_ASAP7_75t_L g190 ( 
.A1(n_183),
.A2(n_93),
.A3(n_95),
.B1(n_101),
.B2(n_110),
.C1(n_186),
.C2(n_181),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_188),
.B(n_179),
.Y(n_191)
);

OR2x2_ASAP7_75t_L g192 ( 
.A(n_187),
.B(n_185),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_191),
.Y(n_193)
);

OAI222xp33_ASAP7_75t_L g194 ( 
.A1(n_192),
.A2(n_190),
.B1(n_189),
.B2(n_93),
.C1(n_101),
.C2(n_95),
.Y(n_194)
);

AOI221xp5_ASAP7_75t_L g195 ( 
.A1(n_193),
.A2(n_95),
.B1(n_101),
.B2(n_194),
.C(n_191),
.Y(n_195)
);


endmodule