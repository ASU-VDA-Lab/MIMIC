module fake_jpeg_9644_n_269 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_269);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_269;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_175;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_192;
wire n_156;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

INVx5_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx11_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_11),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_37),
.Y(n_43)
);

INVxp67_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_19),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_40),
.B(n_28),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_26),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_42),
.B(n_48),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_40),
.B(n_26),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_50),
.B(n_53),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_26),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_59),
.Y(n_74)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_33),
.Y(n_54)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_34),
.A2(n_16),
.B1(n_22),
.B2(n_21),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_56),
.A2(n_16),
.B1(n_22),
.B2(n_18),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_57),
.B(n_28),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_27),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g60 ( 
.A1(n_34),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_23),
.B1(n_30),
.B2(n_24),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_61),
.A2(n_69),
.B(n_87),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_42),
.B(n_39),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_62),
.B(n_76),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_51),
.A2(n_19),
.B1(n_23),
.B2(n_31),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_63),
.A2(n_82),
.B1(n_27),
.B2(n_25),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_57),
.B(n_32),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g95 ( 
.A(n_66),
.B(n_67),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_0),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_47),
.A2(n_23),
.B1(n_31),
.B2(n_29),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_72),
.B1(n_84),
.B2(n_58),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_45),
.A2(n_29),
.B1(n_31),
.B2(n_18),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_47),
.A2(n_30),
.B1(n_29),
.B2(n_18),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_73),
.A2(n_53),
.B1(n_49),
.B2(n_54),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_75),
.A2(n_46),
.B1(n_38),
.B2(n_8),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_27),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_77),
.B(n_46),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_86),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_44),
.B(n_17),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_79),
.B(n_81),
.Y(n_100)
);

AOI32xp33_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_24),
.A3(n_38),
.B1(n_25),
.B2(n_27),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_1),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_44),
.B(n_17),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_44),
.A2(n_24),
.B1(n_27),
.B2(n_25),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_50),
.B(n_17),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_83),
.B(n_88),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_45),
.A2(n_27),
.B1(n_25),
.B2(n_17),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_55),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_45),
.A2(n_10),
.B1(n_15),
.B2(n_14),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_55),
.B(n_9),
.Y(n_88)
);

AO21x1_ASAP7_75t_SL g132 ( 
.A1(n_90),
.A2(n_94),
.B(n_71),
.Y(n_132)
);

O2A1O1Ixp33_ASAP7_75t_L g91 ( 
.A1(n_75),
.A2(n_53),
.B(n_49),
.C(n_54),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_91),
.A2(n_114),
.B(n_88),
.Y(n_122)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_71),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_92),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g93 ( 
.A(n_62),
.B(n_0),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_93),
.A2(n_81),
.B(n_79),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_74),
.A2(n_58),
.B1(n_52),
.B2(n_46),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_96),
.A2(n_107),
.B1(n_64),
.B2(n_71),
.Y(n_133)
);

AND2x6_ASAP7_75t_L g99 ( 
.A(n_74),
.B(n_12),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_99),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_68),
.B(n_52),
.C(n_58),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_111),
.C(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_17),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_103),
.B(n_106),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_85),
.Y(n_138)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_105),
.B(n_82),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_38),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_108),
.B(n_76),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_78),
.A2(n_38),
.B1(n_6),
.B2(n_9),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_109),
.A2(n_110),
.B1(n_72),
.B2(n_73),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_63),
.A2(n_5),
.B1(n_13),
.B2(n_12),
.Y(n_110)
);

MAJx2_ASAP7_75t_L g111 ( 
.A(n_68),
.B(n_0),
.C(n_1),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_70),
.B(n_0),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_113),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_69),
.B(n_1),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_116),
.A2(n_139),
.B1(n_109),
.B2(n_100),
.Y(n_152)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_117),
.B(n_121),
.Y(n_146)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_96),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_118),
.B(n_124),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_98),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_122),
.B(n_137),
.Y(n_151)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_90),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_129),
.Y(n_153)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_92),
.Y(n_125)
);

INVx3_ASAP7_75t_SL g160 ( 
.A(n_125),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_145)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_99),
.Y(n_127)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_127),
.Y(n_156)
);

OAI22x1_ASAP7_75t_L g130 ( 
.A1(n_89),
.A2(n_80),
.B1(n_69),
.B2(n_65),
.Y(n_130)
);

MAJx2_ASAP7_75t_L g131 ( 
.A(n_101),
.B(n_69),
.C(n_66),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_134),
.B(n_135),
.Y(n_150)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_141),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_138),
.A2(n_112),
.B1(n_93),
.B2(n_111),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_105),
.A2(n_64),
.B1(n_86),
.B2(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_94),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_141),
.A2(n_104),
.B1(n_114),
.B2(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_142),
.A2(n_143),
.B1(n_119),
.B2(n_121),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_132),
.A2(n_89),
.B1(n_102),
.B2(n_64),
.Y(n_143)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_130),
.A2(n_102),
.B(n_111),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_144),
.A2(n_3),
.B(n_5),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_136),
.B(n_95),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_147),
.B(n_148),
.Y(n_172)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_149),
.B(n_157),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_152),
.A2(n_127),
.B1(n_119),
.B2(n_122),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_123),
.A2(n_118),
.B1(n_134),
.B2(n_138),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_133),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_93),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_140),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_159),
.A2(n_131),
.B(n_137),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_128),
.B(n_100),
.Y(n_161)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_161),
.Y(n_185)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_120),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_162),
.B(n_164),
.Y(n_173)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_115),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_163),
.B(n_166),
.Y(n_175)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_116),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_167),
.B(n_125),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_128),
.B(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_169),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_146),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_170),
.B(n_174),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_171),
.A2(n_188),
.B1(n_142),
.B2(n_148),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_150),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_190),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_162),
.B(n_95),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_179),
.B(n_153),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g181 ( 
.A(n_160),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_166),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_182),
.B(n_165),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_183),
.A2(n_191),
.B1(n_192),
.B2(n_152),
.Y(n_198)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_151),
.B(n_1),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_187),
.A2(n_169),
.B(n_161),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_167),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_164),
.B(n_9),
.Y(n_189)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_143),
.A2(n_2),
.B1(n_5),
.B2(n_6),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_157),
.A2(n_2),
.B1(n_12),
.B2(n_13),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g193 ( 
.A(n_168),
.B(n_151),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_193),
.B(n_156),
.C(n_154),
.Y(n_199)
);

OA21x2_ASAP7_75t_SL g194 ( 
.A1(n_172),
.A2(n_159),
.B(n_168),
.Y(n_194)
);

OAI21xp33_ASAP7_75t_L g215 ( 
.A1(n_194),
.A2(n_170),
.B(n_176),
.Y(n_215)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_181),
.Y(n_195)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_195),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_198),
.A2(n_212),
.B1(n_188),
.B2(n_180),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_199),
.B(n_205),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_200),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_193),
.B(n_159),
.C(n_154),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_207),
.C(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_203),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_191),
.Y(n_223)
);

XNOR2x1_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_150),
.Y(n_205)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_206),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_145),
.Y(n_207)
);

CKINVDCx14_ASAP7_75t_R g209 ( 
.A(n_173),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_210),
.Y(n_219)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_192),
.Y(n_211)
);

INVx13_ASAP7_75t_L g214 ( 
.A(n_211),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_180),
.A2(n_158),
.B1(n_2),
.B2(n_14),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_171),
.B(n_183),
.Y(n_213)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_215),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_223),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g221 ( 
.A1(n_202),
.A2(n_174),
.B(n_186),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_221),
.A2(n_178),
.B(n_197),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_186),
.B1(n_178),
.B2(n_185),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_197),
.B1(n_187),
.B2(n_190),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_223),
.B(n_204),
.Y(n_230)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_195),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_196),
.B(n_185),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_230),
.B(n_233),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_225),
.B(n_201),
.C(n_199),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_231),
.B(n_232),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_217),
.C(n_216),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_217),
.B(n_213),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_207),
.C(n_205),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_236),
.Y(n_248)
);

A2O1A1Ixp33_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_206),
.B(n_212),
.C(n_173),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_235),
.B(n_218),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_175),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_238),
.B(n_226),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_239),
.B(n_221),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g245 ( 
.A1(n_240),
.A2(n_220),
.B1(n_214),
.B2(n_224),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g253 ( 
.A1(n_241),
.A2(n_249),
.B1(n_235),
.B2(n_219),
.Y(n_253)
);

OAI21x1_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_237),
.B(n_234),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_245),
.B(n_219),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g246 ( 
.A(n_229),
.Y(n_246)
);

OR2x2_ASAP7_75t_L g255 ( 
.A(n_246),
.B(n_247),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_243),
.B(n_232),
.C(n_231),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_250),
.B(n_254),
.Y(n_260)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_252),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_253),
.B(n_256),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_248),
.B(n_208),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_227),
.B(n_220),
.Y(n_256)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_251),
.A2(n_246),
.B(n_244),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_258),
.B(n_252),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_255),
.B(n_233),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_255),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_262),
.A2(n_263),
.B1(n_257),
.B2(n_214),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_260),
.B(n_250),
.C(n_259),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_244),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

OAI21xp33_ASAP7_75t_R g268 ( 
.A1(n_267),
.A2(n_182),
.B(n_255),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_268),
.B(n_182),
.Y(n_269)
);


endmodule