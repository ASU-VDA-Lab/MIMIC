module fake_jpeg_18875_n_39 (n_3, n_2, n_1, n_0, n_4, n_5, n_39);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_39;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx3_ASAP7_75t_L g6 ( 
.A(n_3),
.Y(n_6)
);

CKINVDCx20_ASAP7_75t_R g7 ( 
.A(n_0),
.Y(n_7)
);

BUFx6f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

NOR2xp33_ASAP7_75t_L g9 ( 
.A(n_0),
.B(n_4),
.Y(n_9)
);

NOR2xp33_ASAP7_75t_L g10 ( 
.A(n_2),
.B(n_3),
.Y(n_10)
);

INVx2_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_11),
.Y(n_12)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_13),
.B(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_9),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_14),
.B(n_7),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_SL g15 ( 
.A(n_7),
.B(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_15),
.B(n_10),
.Y(n_18)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g23 ( 
.A(n_17),
.B(n_18),
.Y(n_23)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_19),
.Y(n_21)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_21),
.Y(n_28)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_20),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_24),
.Y(n_26)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_21),
.A2(n_12),
.B1(n_11),
.B2(n_15),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_25),
.B(n_27),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_14),
.C(n_12),
.Y(n_27)
);

NOR4xp25_ASAP7_75t_L g30 ( 
.A(n_28),
.B(n_27),
.C(n_26),
.D(n_14),
.Y(n_30)
);

XNOR2xp5_ASAP7_75t_L g33 ( 
.A(n_30),
.B(n_13),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_31),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_33),
.B(n_13),
.Y(n_35)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_32),
.A2(n_29),
.B(n_4),
.Y(n_34)
);

MAJx2_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_35),
.C(n_33),
.Y(n_36)
);

A2O1A1Ixp33_ASAP7_75t_L g37 ( 
.A1(n_36),
.A2(n_8),
.B(n_5),
.C(n_0),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_5),
.B(n_8),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_38),
.B(n_16),
.Y(n_39)
);


endmodule