module fake_jpeg_5362_n_327 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_327);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_327;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx11_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx8_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_28),
.B(n_30),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_29),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_25),
.Y(n_32)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_32),
.Y(n_45)
);

HB1xp67_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_34),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_35),
.Y(n_43)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_37),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_19),
.B(n_6),
.Y(n_38)
);

NAND2xp33_ASAP7_75t_SL g53 ( 
.A(n_38),
.B(n_19),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_42),
.Y(n_65)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_49),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_51),
.Y(n_77)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_29),
.Y(n_52)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

AND2x4_ASAP7_75t_L g70 ( 
.A(n_53),
.B(n_38),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_39),
.A2(n_18),
.B1(n_13),
.B2(n_53),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_58),
.A2(n_67),
.B1(n_70),
.B2(n_71),
.Y(n_89)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_54),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_59),
.B(n_64),
.Y(n_84)
);

BUFx4f_ASAP7_75t_SL g62 ( 
.A(n_52),
.Y(n_62)
);

BUFx5_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_38),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_63),
.B(n_27),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_56),
.A2(n_36),
.B1(n_18),
.B2(n_20),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_69),
.Y(n_98)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_56),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_13),
.B1(n_45),
.B2(n_44),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_42),
.Y(n_72)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_44),
.A2(n_13),
.B1(n_22),
.B2(n_15),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_73),
.A2(n_75),
.B1(n_22),
.B2(n_15),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_74),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_13),
.B1(n_16),
.B2(n_17),
.Y(n_75)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_63),
.B(n_50),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_79),
.B(n_100),
.Y(n_103)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx11_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_65),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_81),
.B(n_87),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_82),
.A2(n_66),
.B1(n_76),
.B2(n_72),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_74),
.Y(n_85)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

O2A1O1Ixp33_ASAP7_75t_SL g86 ( 
.A1(n_70),
.A2(n_20),
.B(n_19),
.C(n_24),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_86),
.A2(n_17),
.B(n_16),
.Y(n_117)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_62),
.Y(n_87)
);

A2O1A1Ixp33_ASAP7_75t_L g88 ( 
.A1(n_70),
.A2(n_24),
.B(n_49),
.C(n_27),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_88),
.B(n_96),
.Y(n_121)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_57),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_75),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_70),
.A2(n_45),
.B1(n_55),
.B2(n_43),
.Y(n_94)
);

AOI21xp5_ASAP7_75t_L g104 ( 
.A1(n_94),
.A2(n_99),
.B(n_68),
.Y(n_104)
);

INVx3_ASAP7_75t_L g95 ( 
.A(n_64),
.Y(n_95)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_69),
.A2(n_24),
.B1(n_22),
.B2(n_15),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_74),
.B(n_46),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g101 ( 
.A(n_57),
.Y(n_101)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_66),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_104),
.A2(n_116),
.B(n_117),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_113),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_96),
.B(n_48),
.C(n_61),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_114),
.C(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_93),
.B(n_78),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_118),
.Y(n_135)
);

AO21x2_ASAP7_75t_SL g109 ( 
.A1(n_88),
.A2(n_35),
.B(n_21),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_109),
.A2(n_119),
.B1(n_84),
.B2(n_95),
.Y(n_138)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_110),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_27),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_79),
.B(n_60),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_97),
.Y(n_115)
);

INVxp67_ASAP7_75t_SL g132 ( 
.A(n_115),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_89),
.A2(n_16),
.B(n_17),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_86),
.B(n_59),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_81),
.A2(n_60),
.B1(n_77),
.B2(n_26),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_86),
.A2(n_77),
.B1(n_26),
.B2(n_21),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_120),
.A2(n_84),
.B1(n_92),
.B2(n_101),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_100),
.A2(n_27),
.B(n_14),
.Y(n_122)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_122),
.A2(n_14),
.B(n_26),
.Y(n_150)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_124),
.B(n_91),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_121),
.A2(n_82),
.B(n_98),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_125),
.A2(n_128),
.B(n_14),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_90),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_127),
.B(n_131),
.Y(n_177)
);

AOI32xp33_ASAP7_75t_SL g128 ( 
.A1(n_109),
.A2(n_27),
.A3(n_90),
.B1(n_87),
.B2(n_80),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_129),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_130),
.B(n_144),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_105),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_105),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_134),
.Y(n_163)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_111),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_137),
.Y(n_167)
);

OAI21xp33_ASAP7_75t_SL g162 ( 
.A1(n_138),
.A2(n_120),
.B(n_119),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_123),
.B(n_83),
.Y(n_139)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_123),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_140),
.B(n_141),
.Y(n_171)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_109),
.A2(n_118),
.B1(n_121),
.B2(n_117),
.Y(n_142)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g143 ( 
.A(n_103),
.B(n_27),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_107),
.C(n_14),
.Y(n_164)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_103),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_106),
.B(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_145),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_83),
.Y(n_146)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_146),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_147),
.A2(n_107),
.B1(n_115),
.B2(n_112),
.Y(n_165)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_106),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_108),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g160 ( 
.A1(n_150),
.A2(n_122),
.B(n_124),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_109),
.B1(n_104),
.B2(n_113),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_152),
.A2(n_158),
.B1(n_165),
.B2(n_178),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_144),
.B(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_156),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_127),
.A2(n_109),
.B1(n_113),
.B2(n_116),
.Y(n_158)
);

OA21x2_ASAP7_75t_L g203 ( 
.A1(n_160),
.A2(n_162),
.B(n_174),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_164),
.B(n_85),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_126),
.A2(n_136),
.B(n_148),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_143),
.Y(n_191)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_139),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_168),
.B(n_167),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_169),
.A2(n_173),
.B1(n_131),
.B2(n_134),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_135),
.B(n_14),
.Y(n_170)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_170),
.Y(n_183)
);

A2O1A1Ixp33_ASAP7_75t_L g172 ( 
.A1(n_126),
.A2(n_112),
.B(n_102),
.C(n_14),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_172),
.B(n_140),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_136),
.A2(n_91),
.B(n_111),
.Y(n_173)
);

OA22x2_ASAP7_75t_L g174 ( 
.A1(n_128),
.A2(n_26),
.B1(n_21),
.B2(n_14),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_0),
.Y(n_175)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_175),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_130),
.B(n_112),
.C(n_102),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_164),
.C(n_153),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_102),
.B1(n_21),
.B2(n_91),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_179),
.B(n_190),
.C(n_191),
.Y(n_220)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_155),
.Y(n_180)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_180),
.Y(n_207)
);

INVxp33_ASAP7_75t_L g184 ( 
.A(n_155),
.Y(n_184)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_184),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_154),
.A2(n_142),
.B1(n_138),
.B2(n_125),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_186),
.A2(n_200),
.B1(n_174),
.B2(n_157),
.Y(n_212)
);

INVx5_ASAP7_75t_L g187 ( 
.A(n_174),
.Y(n_187)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_187),
.Y(n_228)
);

OAI22x1_ASAP7_75t_L g188 ( 
.A1(n_174),
.A2(n_146),
.B1(n_145),
.B2(n_132),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_188),
.A2(n_174),
.B1(n_172),
.B2(n_157),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_189),
.B(n_161),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_143),
.C(n_150),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_193),
.A2(n_196),
.B1(n_199),
.B2(n_158),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_176),
.B(n_141),
.C(n_133),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_194),
.B(n_198),
.Y(n_222)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_171),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_195),
.B(n_197),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_133),
.B1(n_149),
.B2(n_129),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_132),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_154),
.A2(n_137),
.B1(n_2),
.B2(n_3),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_158),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_201),
.B(n_202),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_167),
.Y(n_202)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_177),
.Y(n_204)
);

INVx13_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_205),
.B(n_164),
.Y(n_221)
);

XNOR2x1_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_166),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_206),
.B(n_227),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_208),
.A2(n_212),
.B1(n_227),
.B2(n_163),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_211),
.A2(n_213),
.B1(n_226),
.B2(n_172),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g213 ( 
.A1(n_188),
.A2(n_159),
.B1(n_161),
.B2(n_174),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g214 ( 
.A(n_194),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g229 ( 
.A1(n_214),
.A2(n_218),
.B(n_169),
.Y(n_229)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_215),
.Y(n_232)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_187),
.Y(n_217)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_217),
.Y(n_237)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_181),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_189),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_219),
.B(n_170),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_221),
.B(n_205),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_185),
.B(n_175),
.Y(n_223)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_223),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_199),
.A2(n_152),
.B1(n_165),
.B2(n_178),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_181),
.A2(n_163),
.B1(n_160),
.B2(n_152),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_210),
.B(n_224),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_230),
.A2(n_239),
.B1(n_162),
.B2(n_209),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_220),
.B(n_179),
.C(n_198),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_231),
.B(n_235),
.C(n_236),
.Y(n_259)
);

OR2x2_ASAP7_75t_L g233 ( 
.A(n_215),
.B(n_180),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_233),
.B(n_243),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_222),
.B(n_190),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_234),
.B(n_245),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_220),
.B(n_156),
.C(n_182),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_207),
.B(n_183),
.C(n_186),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_225),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_246),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_218),
.A2(n_168),
.B1(n_151),
.B2(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_240),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_207),
.B(n_184),
.C(n_159),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_247),
.C(n_248),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_242),
.A2(n_228),
.B1(n_212),
.B2(n_203),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_222),
.B(n_200),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_217),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_216),
.B(n_214),
.C(n_206),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_216),
.B(n_151),
.C(n_203),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_223),
.Y(n_257)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_250),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_241),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_253),
.A2(n_256),
.B(n_261),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_248),
.A2(n_228),
.B1(n_211),
.B2(n_226),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_254),
.A2(n_247),
.B1(n_244),
.B2(n_237),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_262),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_8),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_209),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_234),
.B(n_85),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_231),
.B(n_85),
.C(n_2),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_235),
.C(n_2),
.Y(n_270)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_265),
.A2(n_266),
.B(n_267),
.Y(n_284)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_236),
.Y(n_266)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_249),
.B(n_7),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_268),
.Y(n_277)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_269),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_270),
.A2(n_272),
.B(n_276),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_259),
.B(n_1),
.C(n_2),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_271),
.B(n_273),
.C(n_274),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_251),
.B(n_7),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_1),
.C(n_3),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_260),
.B(n_1),
.C(n_4),
.Y(n_274)
);

INVxp67_ASAP7_75t_SL g276 ( 
.A(n_267),
.Y(n_276)
);

OAI321xp33_ASAP7_75t_L g278 ( 
.A1(n_250),
.A2(n_12),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_8),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_278),
.A2(n_12),
.B1(n_4),
.B2(n_6),
.Y(n_289)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_255),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_280),
.B(n_263),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_281),
.B(n_6),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_253),
.A2(n_9),
.B1(n_4),
.B2(n_5),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_282),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_297)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_286),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_291),
.Y(n_305)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_283),
.B(n_252),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_288),
.B(n_296),
.C(n_10),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_289),
.B(n_294),
.Y(n_302)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_275),
.A2(n_260),
.B(n_284),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_290),
.B(n_293),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_277),
.A2(n_257),
.B1(n_264),
.B2(n_262),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_279),
.B(n_252),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g296 ( 
.A(n_283),
.B(n_9),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_297),
.B(n_273),
.Y(n_306)
);

INVx11_ASAP7_75t_L g298 ( 
.A(n_296),
.Y(n_298)
);

INVx11_ASAP7_75t_L g312 ( 
.A(n_298),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_288),
.B(n_295),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_307),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_292),
.B(n_274),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_303),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_281),
.B1(n_270),
.B2(n_271),
.Y(n_304)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_304),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_306),
.B(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_285),
.B(n_10),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_285),
.C(n_1),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_314),
.B(n_302),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_307),
.B(n_11),
.C(n_12),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_311),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_316),
.A2(n_317),
.B(n_318),
.Y(n_321)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_315),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_L g319 ( 
.A1(n_313),
.A2(n_299),
.B(n_301),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_SL g320 ( 
.A1(n_319),
.A2(n_310),
.B(n_313),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_320),
.B(n_315),
.Y(n_322)
);

AOI21xp5_ASAP7_75t_L g323 ( 
.A1(n_322),
.A2(n_309),
.B(n_321),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_323),
.A2(n_304),
.B(n_312),
.Y(n_324)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_324),
.A2(n_312),
.B(n_298),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_325),
.B(n_314),
.C(n_11),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_326),
.B(n_12),
.Y(n_327)
);


endmodule