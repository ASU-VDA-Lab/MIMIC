module fake_jpeg_13537_n_525 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_525);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_293;
wire n_38;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_11),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_2),
.Y(n_17)
);

BUFx5_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_6),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_8),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_11),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_12),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_9),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_10),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_2),
.Y(n_43)
);

INVx13_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_29),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g103 ( 
.A(n_46),
.B(n_48),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_21),
.B(n_6),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_47),
.B(n_54),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_20),
.Y(n_49)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_49),
.Y(n_105)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_20),
.Y(n_50)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_50),
.Y(n_108)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_51),
.Y(n_120)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_21),
.B(n_6),
.Y(n_54)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_18),
.Y(n_55)
);

INVx5_ASAP7_75t_L g133 ( 
.A(n_55),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_15),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_56),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_57),
.B(n_64),
.Y(n_112)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_58),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_36),
.B(n_5),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_59),
.B(n_75),
.Y(n_126)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_60),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_15),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_29),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_65),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_15),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_66),
.Y(n_110)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_67),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_25),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_68),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_42),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_70),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_71),
.Y(n_149)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_16),
.Y(n_72)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx3_ASAP7_75t_SL g73 ( 
.A(n_25),
.Y(n_73)
);

CKINVDCx6p67_ASAP7_75t_R g114 ( 
.A(n_73),
.Y(n_114)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_25),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_74),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_29),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_42),
.Y(n_76)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_39),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_24),
.B(n_5),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_78),
.B(n_82),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_43),
.Y(n_79)
);

INVx8_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx3_ASAP7_75t_L g144 ( 
.A(n_81),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_24),
.B(n_5),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_41),
.Y(n_83)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_83),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_17),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_84),
.B(n_85),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_27),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_26),
.B(n_7),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_86),
.B(n_90),
.Y(n_140)
);

INVx2_ASAP7_75t_SL g87 ( 
.A(n_39),
.Y(n_87)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_87),
.Y(n_148)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_88),
.Y(n_116)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_31),
.Y(n_89)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_26),
.B(n_7),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_17),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_91),
.B(n_32),
.Y(n_134)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_20),
.B(n_7),
.Y(n_92)
);

A2O1A1Ixp33_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_27),
.B(n_33),
.C(n_32),
.Y(n_102)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_93),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_43),
.Y(n_94)
);

BUFx12f_ASAP7_75t_L g118 ( 
.A(n_94),
.Y(n_118)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_102),
.B(n_124),
.Y(n_200)
);

INVx6_ASAP7_75t_SL g107 ( 
.A(n_46),
.Y(n_107)
);

INVx13_ASAP7_75t_L g185 ( 
.A(n_107),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_87),
.A2(n_28),
.B1(n_37),
.B2(n_31),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_111),
.A2(n_73),
.B1(n_55),
.B2(n_58),
.Y(n_169)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g193 ( 
.A(n_117),
.Y(n_193)
);

BUFx10_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_119),
.Y(n_159)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_69),
.Y(n_121)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_121),
.Y(n_168)
);

INVx6_ASAP7_75t_SL g123 ( 
.A(n_48),
.Y(n_123)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_123),
.Y(n_157)
);

HAxp5_ASAP7_75t_SL g124 ( 
.A(n_92),
.B(n_91),
.CON(n_124),
.SN(n_124)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_70),
.Y(n_127)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_57),
.Y(n_131)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_131),
.Y(n_184)
);

INVx13_ASAP7_75t_L g132 ( 
.A(n_64),
.Y(n_132)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_134),
.B(n_147),
.Y(n_161)
);

INVx11_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_84),
.B(n_23),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_138),
.B(n_33),
.Y(n_181)
);

BUFx4f_ASAP7_75t_SL g139 ( 
.A(n_53),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g160 ( 
.A(n_139),
.Y(n_160)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_72),
.Y(n_141)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_88),
.Y(n_143)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_143),
.Y(n_172)
);

OR2x2_ASAP7_75t_L g147 ( 
.A(n_52),
.B(n_28),
.Y(n_147)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_136),
.Y(n_158)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_158),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_103),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_162),
.B(n_166),
.Y(n_213)
);

INVx3_ASAP7_75t_L g163 ( 
.A(n_131),
.Y(n_163)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_163),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_152),
.B(n_67),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g167 ( 
.A(n_112),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_167),
.B(n_178),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_169),
.B(n_198),
.Y(n_226)
);

INVx3_ASAP7_75t_L g170 ( 
.A(n_118),
.Y(n_170)
);

INVx3_ASAP7_75t_L g235 ( 
.A(n_170),
.Y(n_235)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

BUFx3_ASAP7_75t_L g214 ( 
.A(n_171),
.Y(n_214)
);

INVx11_ASAP7_75t_L g173 ( 
.A(n_119),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_173),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_119),
.Y(n_174)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_174),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_142),
.A2(n_94),
.B1(n_81),
.B2(n_79),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_175),
.A2(n_180),
.B1(n_182),
.B2(n_191),
.Y(n_206)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_95),
.Y(n_176)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_176),
.Y(n_211)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_177),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_152),
.B(n_75),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_101),
.Y(n_179)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_179),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_106),
.A2(n_49),
.B1(n_50),
.B2(n_63),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_181),
.B(n_189),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_126),
.A2(n_93),
.B1(n_56),
.B2(n_45),
.Y(n_182)
);

INVx2_ASAP7_75t_SL g183 ( 
.A(n_120),
.Y(n_183)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_183),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_126),
.B(n_60),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_188),
.Y(n_202)
);

CKINVDCx12_ASAP7_75t_R g187 ( 
.A(n_132),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_187),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_147),
.B(n_65),
.Y(n_188)
);

OAI32xp33_ASAP7_75t_L g189 ( 
.A1(n_150),
.A2(n_83),
.A3(n_76),
.B1(n_68),
.B2(n_74),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_140),
.B(n_89),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_190),
.B(n_192),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_97),
.A2(n_61),
.B1(n_71),
.B2(n_66),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_148),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_115),
.A2(n_62),
.B1(n_51),
.B2(n_80),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_194),
.A2(n_196),
.B1(n_130),
.B2(n_133),
.Y(n_232)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_195),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_129),
.A2(n_37),
.B1(n_31),
.B2(n_35),
.Y(n_196)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_104),
.Y(n_197)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_125),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_122),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_199),
.B(n_201),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_114),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_186),
.B(n_150),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_209),
.B(n_223),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_111),
.B1(n_124),
.B2(n_114),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_212),
.A2(n_227),
.B1(n_233),
.B2(n_174),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_193),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_215),
.B(n_220),
.Y(n_240)
);

A2O1A1Ixp33_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_113),
.B(n_114),
.C(n_139),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_225),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_200),
.B(n_145),
.C(n_137),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_218),
.C(n_219),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_177),
.B(n_105),
.C(n_108),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_181),
.B(n_113),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_173),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_161),
.B(n_136),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_179),
.B(n_144),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_189),
.A2(n_110),
.B1(n_151),
.B2(n_149),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_109),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_175),
.A2(n_110),
.B1(n_151),
.B2(n_149),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_155),
.B(n_128),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_174),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_225),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_243),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g241 ( 
.A(n_204),
.Y(n_241)
);

INVx1_ASAP7_75t_SL g298 ( 
.A(n_241),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_234),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_221),
.A2(n_191),
.B1(n_194),
.B2(n_99),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_244),
.A2(n_247),
.B1(n_253),
.B2(n_232),
.Y(n_286)
);

INVx13_ASAP7_75t_L g245 ( 
.A(n_205),
.Y(n_245)
);

CKINVDCx14_ASAP7_75t_R g288 ( 
.A(n_245),
.Y(n_288)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_208),
.Y(n_246)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_246),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_221),
.A2(n_98),
.B1(n_99),
.B2(n_100),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_255),
.Y(n_276)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_214),
.Y(n_249)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_249),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_202),
.B(n_156),
.C(n_199),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_250),
.B(n_203),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_184),
.B(n_163),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g297 ( 
.A1(n_251),
.A2(n_228),
.B(n_204),
.Y(n_297)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_208),
.Y(n_252)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_252),
.Y(n_279)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_236),
.Y(n_254)
);

INVx2_ASAP7_75t_L g272 ( 
.A(n_254),
.Y(n_272)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_224),
.Y(n_256)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_202),
.B(n_155),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_258),
.B(n_261),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_209),
.A2(n_185),
.B(n_157),
.Y(n_259)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_259),
.Y(n_299)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_224),
.Y(n_260)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_260),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_219),
.B(n_165),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_210),
.B(n_155),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_262),
.B(n_264),
.Y(n_300)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_229),
.Y(n_264)
);

INVx13_ASAP7_75t_L g265 ( 
.A(n_205),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_265),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_210),
.B(n_195),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_266),
.B(n_267),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_213),
.B(n_157),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_L g268 ( 
.A(n_223),
.B(n_185),
.C(n_171),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_268),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_227),
.A2(n_172),
.B1(n_165),
.B2(n_154),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_206),
.Y(n_277)
);

XNOR2x1_ASAP7_75t_L g271 ( 
.A(n_238),
.B(n_217),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_271),
.B(n_273),
.Y(n_326)
);

XNOR2x1_ASAP7_75t_L g273 ( 
.A(n_238),
.B(n_212),
.Y(n_273)
);

XOR2x2_ASAP7_75t_L g275 ( 
.A(n_257),
.B(n_230),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_293),
.Y(n_324)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_277),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_239),
.B(n_230),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_243),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_241),
.A2(n_184),
.B1(n_220),
.B2(n_222),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_284),
.A2(n_286),
.B1(n_291),
.B2(n_295),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_261),
.B(n_234),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_290),
.C(n_296),
.Y(n_308)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_254),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_289),
.Y(n_312)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_257),
.B(n_218),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_244),
.A2(n_226),
.B1(n_206),
.B2(n_233),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_247),
.A2(n_226),
.B1(n_237),
.B2(n_203),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_250),
.B(n_229),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g334 ( 
.A1(n_297),
.A2(n_159),
.B(n_222),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_242),
.A2(n_226),
.B(n_231),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_302),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_303),
.B(n_311),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_276),
.A2(n_242),
.B1(n_253),
.B2(n_258),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_304),
.A2(n_330),
.B1(n_295),
.B2(n_302),
.Y(n_348)
);

BUFx5_ASAP7_75t_L g305 ( 
.A(n_289),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g340 ( 
.A(n_305),
.Y(n_340)
);

INVx6_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g363 ( 
.A(n_306),
.Y(n_363)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_292),
.B(n_267),
.Y(n_309)
);

NAND3xp33_ASAP7_75t_L g341 ( 
.A(n_309),
.B(n_310),
.C(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_275),
.B(n_266),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_280),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_276),
.A2(n_255),
.B1(n_269),
.B2(n_251),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_313),
.B(n_316),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_271),
.B(n_262),
.C(n_248),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_314),
.B(n_323),
.C(n_328),
.Y(n_352)
);

NOR2xp33_ASAP7_75t_SL g315 ( 
.A(n_282),
.B(n_265),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_240),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_291),
.A2(n_240),
.B1(n_253),
.B2(n_241),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_317),
.Y(n_347)
);

AND2x6_ASAP7_75t_L g318 ( 
.A(n_273),
.B(n_265),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_318),
.B(n_320),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_299),
.A2(n_252),
.B1(n_246),
.B2(n_260),
.Y(n_319)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_319),
.A2(n_334),
.B(n_160),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_215),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_321),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_286),
.A2(n_256),
.B1(n_263),
.B2(n_236),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_322),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_172),
.C(n_154),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_298),
.B(n_207),
.Y(n_325)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_325),
.Y(n_339)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_297),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_327),
.B(n_294),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_296),
.B(n_231),
.C(n_235),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_277),
.A2(n_236),
.B1(n_207),
.B2(n_197),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_331),
.Y(n_342)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_279),
.Y(n_333)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_333),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_293),
.B(n_235),
.C(n_245),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_335),
.B(n_183),
.C(n_211),
.Y(n_368)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_283),
.Y(n_336)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_336),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g337 ( 
.A(n_308),
.B(n_326),
.Y(n_337)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_337),
.B(n_351),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_307),
.A2(n_299),
.B(n_287),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_L g379 ( 
.A1(n_343),
.A2(n_357),
.B(n_360),
.Y(n_379)
);

NOR4xp25_ASAP7_75t_L g344 ( 
.A(n_316),
.B(n_245),
.C(n_285),
.D(n_288),
.Y(n_344)
);

FAx1_ASAP7_75t_SL g394 ( 
.A(n_344),
.B(n_44),
.CI(n_96),
.CON(n_394),
.SN(n_394)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_348),
.A2(n_359),
.B1(n_367),
.B2(n_313),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_308),
.B(n_298),
.Y(n_351)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_321),
.Y(n_355)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_355),
.Y(n_372)
);

CKINVDCx16_ASAP7_75t_R g356 ( 
.A(n_325),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_356),
.B(n_361),
.Y(n_385)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_303),
.Y(n_358)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g359 ( 
.A1(n_329),
.A2(n_281),
.B1(n_283),
.B2(n_272),
.Y(n_359)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_307),
.A2(n_278),
.B(n_272),
.Y(n_360)
);

INVxp67_ASAP7_75t_L g361 ( 
.A(n_334),
.Y(n_361)
);

A2O1A1O1Ixp25_ASAP7_75t_L g362 ( 
.A1(n_314),
.A2(n_183),
.B(n_164),
.C(n_159),
.D(n_160),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_362),
.B(n_366),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g371 ( 
.A(n_364),
.Y(n_371)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_365),
.Y(n_380)
);

INVxp67_ASAP7_75t_L g366 ( 
.A(n_335),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g367 ( 
.A1(n_304),
.A2(n_249),
.B1(n_158),
.B2(n_214),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_368),
.B(n_323),
.C(n_326),
.Y(n_370)
);

NOR2xp33_ASAP7_75t_L g369 ( 
.A(n_349),
.B(n_328),
.Y(n_369)
);

NAND3xp33_ASAP7_75t_L g409 ( 
.A(n_369),
.B(n_363),
.C(n_14),
.Y(n_409)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_370),
.B(n_375),
.C(n_376),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g374 ( 
.A(n_351),
.B(n_324),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g416 ( 
.A(n_374),
.B(n_388),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_352),
.B(n_324),
.C(n_317),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_352),
.B(n_332),
.C(n_318),
.Y(n_376)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_378),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g381 ( 
.A1(n_347),
.A2(n_322),
.B1(n_306),
.B2(n_330),
.Y(n_381)
);

HB1xp67_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_350),
.A2(n_319),
.B1(n_312),
.B2(n_305),
.Y(n_382)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_382),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_337),
.B(n_211),
.C(n_170),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_383),
.B(n_384),
.C(n_393),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_366),
.B(n_198),
.C(n_176),
.Y(n_384)
);

OAI21xp33_ASAP7_75t_L g386 ( 
.A1(n_353),
.A2(n_249),
.B(n_164),
.Y(n_386)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_386),
.Y(n_418)
);

AOI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_361),
.A2(n_312),
.B1(n_109),
.B2(n_96),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_387),
.A2(n_340),
.B1(n_363),
.B2(n_362),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_168),
.Y(n_388)
);

INVxp67_ASAP7_75t_SL g389 ( 
.A(n_342),
.Y(n_389)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_389),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_339),
.B(n_168),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_392),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_348),
.B(n_347),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_368),
.B(n_104),
.C(n_153),
.Y(n_393)
);

OR2x2_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_37),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_338),
.B(n_153),
.C(n_128),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_395),
.B(n_396),
.C(n_397),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_360),
.B(n_100),
.C(n_98),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_346),
.B(n_22),
.C(n_40),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_354),
.Y(n_398)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_398),
.Y(n_419)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_379),
.A2(n_364),
.B(n_350),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g430 ( 
.A1(n_399),
.A2(n_387),
.B(n_371),
.Y(n_430)
);

XNOR2xp5_ASAP7_75t_L g400 ( 
.A(n_375),
.B(n_367),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_400),
.B(n_411),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_359),
.Y(n_401)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_401),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_SL g402 ( 
.A(n_373),
.B(n_341),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_423),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_377),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_403),
.B(n_406),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_345),
.Y(n_404)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_404),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_405),
.A2(n_396),
.B1(n_394),
.B2(n_40),
.Y(n_438)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_390),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_380),
.B(n_340),
.Y(n_408)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_408),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_409),
.B(n_424),
.Y(n_432)
);

OAI21xp33_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_14),
.B(n_13),
.Y(n_411)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_413),
.A2(n_35),
.B1(n_34),
.B2(n_40),
.Y(n_442)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_386),
.Y(n_421)
);

INVx2_ASAP7_75t_L g434 ( 
.A(n_421),
.Y(n_434)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_373),
.B(n_44),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_392),
.B(n_14),
.Y(n_424)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_370),
.B(n_44),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g431 ( 
.A(n_425),
.B(n_384),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_400),
.B(n_383),
.C(n_376),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_427),
.B(n_435),
.Y(n_466)
);

BUFx2_ASAP7_75t_L g428 ( 
.A(n_407),
.Y(n_428)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_428),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g453 ( 
.A(n_430),
.B(n_437),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g460 ( 
.A(n_431),
.B(n_423),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_420),
.B(n_393),
.C(n_395),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_410),
.B(n_397),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_438),
.A2(n_413),
.B1(n_415),
.B2(n_418),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_SL g440 ( 
.A(n_417),
.B(n_13),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_440),
.B(n_9),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_420),
.B(n_412),
.C(n_410),
.Y(n_441)
);

MAJIxp5_ASAP7_75t_L g463 ( 
.A(n_441),
.B(n_446),
.C(n_422),
.Y(n_463)
);

OR2x2_ASAP7_75t_L g458 ( 
.A(n_442),
.B(n_405),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_419),
.B(n_22),
.Y(n_443)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_443),
.Y(n_451)
);

AO21x1_ASAP7_75t_L g445 ( 
.A1(n_418),
.A2(n_13),
.B(n_14),
.Y(n_445)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_445),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_412),
.B(n_38),
.C(n_22),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_414),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_447)
);

HB1xp67_ASAP7_75t_L g455 ( 
.A(n_447),
.Y(n_455)
);

OAI22xp5_ASAP7_75t_SL g448 ( 
.A1(n_414),
.A2(n_38),
.B1(n_35),
.B2(n_34),
.Y(n_448)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_448),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_35),
.Y(n_449)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_449),
.Y(n_462)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_428),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_454),
.B(n_456),
.Y(n_470)
);

XNOR2xp5_ASAP7_75t_SL g457 ( 
.A(n_429),
.B(n_402),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g473 ( 
.A(n_457),
.B(n_460),
.Y(n_473)
);

HB1xp67_ASAP7_75t_L g474 ( 
.A(n_458),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_435),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_459),
.B(n_464),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g483 ( 
.A1(n_461),
.A2(n_462),
.B1(n_455),
.B2(n_468),
.Y(n_483)
);

XNOR2xp5_ASAP7_75t_L g476 ( 
.A(n_463),
.B(n_431),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_SL g464 ( 
.A1(n_427),
.A2(n_399),
.B(n_416),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g465 ( 
.A(n_437),
.B(n_425),
.C(n_422),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_465),
.B(n_467),
.Y(n_480)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_433),
.Y(n_467)
);

OAI21xp5_ASAP7_75t_L g469 ( 
.A1(n_466),
.A2(n_463),
.B(n_434),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_469),
.A2(n_481),
.B(n_465),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g471 ( 
.A(n_459),
.B(n_432),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_471),
.B(n_472),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_454),
.B(n_436),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_476),
.B(n_478),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_453),
.B(n_439),
.Y(n_477)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_477),
.B(n_4),
.Y(n_493)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_458),
.Y(n_478)
);

O2A1O1Ixp33_ASAP7_75t_SL g479 ( 
.A1(n_452),
.A2(n_401),
.B(n_404),
.C(n_426),
.Y(n_479)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_479),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_453),
.B(n_446),
.C(n_439),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_450),
.B(n_444),
.Y(n_482)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_482),
.Y(n_486)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_483),
.Y(n_489)
);

FAx1_ASAP7_75t_SL g484 ( 
.A(n_457),
.B(n_424),
.CI(n_429),
.CON(n_484),
.SN(n_484)
);

OAI22xp5_ASAP7_75t_L g491 ( 
.A1(n_484),
.A2(n_445),
.B1(n_448),
.B2(n_447),
.Y(n_491)
);

NOR3xp33_ASAP7_75t_L g485 ( 
.A(n_475),
.B(n_430),
.C(n_451),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g500 ( 
.A(n_485),
.B(n_488),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g499 ( 
.A(n_487),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_476),
.B(n_460),
.C(n_438),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_491),
.B(n_0),
.Y(n_508)
);

OR2x6_ASAP7_75t_SL g503 ( 
.A(n_493),
.B(n_477),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_474),
.A2(n_4),
.B(n_10),
.Y(n_494)
);

AOI21xp5_ASAP7_75t_L g507 ( 
.A1(n_494),
.A2(n_496),
.B(n_9),
.Y(n_507)
);

OAI21xp5_ASAP7_75t_SL g496 ( 
.A1(n_480),
.A2(n_9),
.B(n_1),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_470),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_497),
.B(n_498),
.Y(n_501)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_483),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_492),
.B(n_481),
.Y(n_502)
);

OR2x2_ASAP7_75t_L g509 ( 
.A(n_502),
.B(n_505),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g515 ( 
.A1(n_503),
.A2(n_504),
.B(n_506),
.Y(n_515)
);

NOR2xp67_ASAP7_75t_L g504 ( 
.A(n_486),
.B(n_473),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_495),
.B(n_479),
.C(n_484),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_488),
.B(n_489),
.Y(n_506)
);

OAI211xp5_ASAP7_75t_L g511 ( 
.A1(n_507),
.A2(n_490),
.B(n_494),
.C(n_2),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_508),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_501),
.B(n_490),
.Y(n_510)
);

AOI31xp33_ASAP7_75t_L g519 ( 
.A1(n_510),
.A2(n_511),
.A3(n_514),
.B(n_0),
.Y(n_519)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_500),
.Y(n_513)
);

AOI322xp5_ASAP7_75t_L g516 ( 
.A1(n_513),
.A2(n_507),
.A3(n_493),
.B1(n_34),
.B2(n_39),
.C1(n_3),
.C2(n_1),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g514 ( 
.A(n_499),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g521 ( 
.A(n_516),
.B(n_517),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_509),
.A2(n_34),
.B(n_1),
.Y(n_517)
);

OAI21xp5_ASAP7_75t_L g518 ( 
.A1(n_515),
.A2(n_512),
.B(n_1),
.Y(n_518)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_519),
.Y(n_520)
);

OAI21xp5_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_0),
.B(n_3),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_L g523 ( 
.A(n_522),
.B(n_0),
.Y(n_523)
);

OAI21xp5_ASAP7_75t_L g524 ( 
.A1(n_523),
.A2(n_520),
.B(n_3),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_3),
.Y(n_525)
);


endmodule