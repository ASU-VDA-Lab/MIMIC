module fake_jpeg_24452_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_1),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

AND2x2_ASAP7_75t_SL g23 ( 
.A(n_3),
.B(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_12),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_7),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVxp67_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

AOI21xp33_ASAP7_75t_L g37 ( 
.A1(n_23),
.A2(n_14),
.B(n_13),
.Y(n_37)
);

HAxp5_ASAP7_75t_SL g68 ( 
.A(n_37),
.B(n_40),
.CON(n_68),
.SN(n_68)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_38),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_26),
.B(n_0),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx2_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_28),
.Y(n_45)
);

BUFx24_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_46),
.Y(n_100)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_48),
.B(n_49),
.Y(n_73)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_50),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_23),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_23),
.Y(n_83)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_53),
.B(n_62),
.Y(n_97)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_55),
.Y(n_87)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_44),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_18),
.B1(n_30),
.B2(n_28),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_58),
.Y(n_90)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_60),
.Y(n_109)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

INVx2_ASAP7_75t_SL g93 ( 
.A(n_61),
.Y(n_93)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_38),
.Y(n_62)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_64),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_42),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_65),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_60),
.A2(n_18),
.B1(n_27),
.B2(n_30),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_70),
.Y(n_117)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_52),
.Y(n_71)
);

INVx8_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_72),
.A2(n_86),
.B1(n_98),
.B2(n_99),
.Y(n_123)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_76),
.Y(n_113)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_77),
.B(n_80),
.Y(n_132)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_68),
.A2(n_23),
.B(n_20),
.Y(n_78)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_78),
.B(n_10),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_27),
.B1(n_16),
.B2(n_33),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_79),
.Y(n_126)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

A2O1A1Ixp33_ASAP7_75t_L g82 ( 
.A1(n_68),
.A2(n_23),
.B(n_32),
.C(n_36),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_82),
.B(n_83),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_36),
.B1(n_16),
.B2(n_42),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_84),
.A2(n_85),
.B1(n_107),
.B2(n_26),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_55),
.A2(n_16),
.B1(n_42),
.B2(n_33),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_47),
.A2(n_20),
.B1(n_34),
.B2(n_33),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_54),
.A2(n_19),
.B1(n_25),
.B2(n_34),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_88),
.A2(n_26),
.B1(n_35),
.B2(n_13),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_69),
.B(n_31),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_89),
.Y(n_119)
);

OA22x2_ASAP7_75t_L g92 ( 
.A1(n_58),
.A2(n_43),
.B1(n_41),
.B2(n_39),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_92),
.A2(n_66),
.B1(n_43),
.B2(n_41),
.Y(n_116)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_56),
.Y(n_94)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_48),
.A2(n_19),
.B1(n_25),
.B2(n_17),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_95),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_138)
);

OR2x2_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_17),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_106),
.Y(n_137)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_67),
.A2(n_17),
.B1(n_24),
.B2(n_19),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_59),
.A2(n_29),
.B1(n_25),
.B2(n_35),
.Y(n_99)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_67),
.A2(n_29),
.B(n_41),
.C(n_39),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_62),
.A2(n_29),
.B1(n_35),
.B2(n_24),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_104),
.A2(n_108),
.B1(n_12),
.B2(n_11),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_63),
.B(n_43),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_66),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_L g108 ( 
.A1(n_63),
.A2(n_24),
.B1(n_31),
.B2(n_22),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g110 ( 
.A(n_66),
.B(n_0),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_110),
.B(n_26),
.C(n_14),
.Y(n_125)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_71),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_112),
.B(n_120),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g146 ( 
.A1(n_116),
.A2(n_121),
.B1(n_133),
.B2(n_134),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_83),
.B(n_43),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_118),
.B(n_125),
.C(n_130),
.Y(n_162)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_90),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_110),
.A2(n_29),
.B1(n_22),
.B2(n_35),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_71),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_122),
.B(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_124),
.B(n_129),
.Y(n_156)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_83),
.B(n_41),
.C(n_39),
.Y(n_130)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_131),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_82),
.A2(n_39),
.B1(n_1),
.B2(n_2),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_81),
.A2(n_13),
.B1(n_12),
.B2(n_11),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_97),
.B1(n_93),
.B2(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_136),
.B(n_139),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_138),
.A2(n_99),
.B1(n_104),
.B2(n_110),
.Y(n_152)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_97),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_140),
.B(n_109),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_132),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_142),
.B(n_150),
.Y(n_179)
);

OA22x2_ASAP7_75t_L g143 ( 
.A1(n_116),
.A2(n_103),
.B1(n_92),
.B2(n_95),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_143),
.A2(n_117),
.B1(n_126),
.B2(n_125),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g144 ( 
.A(n_119),
.B(n_89),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_144),
.B(n_147),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_158),
.B1(n_170),
.B2(n_172),
.Y(n_184)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_105),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_149),
.B(n_160),
.Y(n_173)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_113),
.Y(n_150)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_115),
.A2(n_105),
.B(n_72),
.C(n_96),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_151),
.A2(n_157),
.B(n_163),
.Y(n_177)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_153),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_119),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_164),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_128),
.A2(n_93),
.B1(n_102),
.B2(n_75),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_101),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_136),
.B(n_96),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_101),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_161),
.B(n_165),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_128),
.A2(n_91),
.B(n_102),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_140),
.B(n_107),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_166),
.B(n_167),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_139),
.B(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_127),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_168),
.Y(n_191)
);

BUFx8_ASAP7_75t_L g169 ( 
.A(n_112),
.Y(n_169)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_169),
.Y(n_192)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_127),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_123),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_171),
.B(n_0),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g172 ( 
.A1(n_123),
.A2(n_93),
.B1(n_75),
.B2(n_91),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_174),
.A2(n_183),
.B1(n_143),
.B2(n_168),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_117),
.B1(n_126),
.B2(n_138),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_175),
.A2(n_176),
.B1(n_185),
.B2(n_199),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_165),
.A2(n_129),
.B1(n_87),
.B2(n_92),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_114),
.C(n_100),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_178),
.B(n_196),
.C(n_203),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g181 ( 
.A(n_167),
.B(n_92),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_181),
.B(n_200),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_164),
.A2(n_114),
.B1(n_87),
.B2(n_94),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_147),
.A2(n_111),
.B1(n_80),
.B2(n_100),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g216 ( 
.A1(n_188),
.A2(n_151),
.B(n_156),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_149),
.B(n_0),
.Y(n_190)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_190),
.Y(n_206)
);

OR2x2_ASAP7_75t_L g193 ( 
.A(n_154),
.B(n_71),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_194),
.Y(n_226)
);

OR2x2_ASAP7_75t_L g194 ( 
.A(n_160),
.B(n_90),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_162),
.B(n_111),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_161),
.B(n_141),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

AND2x6_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_163),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g230 ( 
.A1(n_198),
.A2(n_201),
.B(n_169),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_145),
.A2(n_77),
.B1(n_74),
.B2(n_127),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_166),
.B(n_10),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g201 ( 
.A(n_142),
.B(n_1),
.Y(n_201)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_152),
.B(n_122),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_191),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_204),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_191),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_205),
.B(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_209),
.B(n_216),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_179),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_196),
.B(n_157),
.C(n_158),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_211),
.B(n_221),
.Y(n_241)
);

NAND3xp33_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_144),
.C(n_150),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_212),
.B(n_214),
.Y(n_237)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_195),
.A2(n_172),
.B1(n_155),
.B2(n_143),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_217),
.A2(n_218),
.B1(n_174),
.B2(n_177),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_176),
.A2(n_143),
.B1(n_155),
.B2(n_146),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g219 ( 
.A(n_183),
.Y(n_219)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_219),
.Y(n_234)
);

CKINVDCx14_ASAP7_75t_R g220 ( 
.A(n_185),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_223),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_178),
.B(n_148),
.C(n_146),
.Y(n_221)
);

AO21x1_ASAP7_75t_L g233 ( 
.A1(n_222),
.A2(n_230),
.B(n_228),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g223 ( 
.A(n_188),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_173),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_224),
.B(n_228),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_170),
.C(n_169),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_225),
.B(n_227),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_197),
.B(n_169),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_193),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_173),
.Y(n_229)
);

NOR4xp25_ASAP7_75t_L g231 ( 
.A(n_229),
.B(n_190),
.C(n_182),
.D(n_186),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_233),
.Y(n_265)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_235),
.B(n_238),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_236),
.A2(n_242),
.B(n_243),
.Y(n_252)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_227),
.Y(n_238)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_226),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_240),
.B(n_246),
.Y(n_259)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_226),
.A2(n_177),
.B(n_198),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_230),
.A2(n_229),
.B(n_224),
.Y(n_243)
);

XNOR2x1_ASAP7_75t_L g244 ( 
.A(n_207),
.B(n_203),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_244),
.B(n_215),
.Y(n_261)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_205),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_216),
.A2(n_175),
.B(n_194),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_247),
.A2(n_182),
.B(n_213),
.Y(n_258)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_204),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_204),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_192),
.Y(n_253)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_253),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g254 ( 
.A(n_232),
.Y(n_254)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_254),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_241),
.B(n_207),
.Y(n_255)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_255),
.B(n_260),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_243),
.B(n_202),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g273 ( 
.A(n_256),
.B(n_239),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_258),
.A2(n_245),
.B(n_234),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_244),
.B(n_215),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_261),
.B(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_214),
.B1(n_213),
.B2(n_209),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_262),
.A2(n_234),
.B1(n_245),
.B2(n_235),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_221),
.C(n_211),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_264),
.B(n_266),
.C(n_269),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_251),
.B(n_208),
.C(n_206),
.Y(n_266)
);

HB1xp67_ASAP7_75t_L g267 ( 
.A(n_246),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_267),
.B(n_192),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_248),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_181),
.Y(n_269)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_270),
.Y(n_294)
);

MAJx2_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_280),
.C(n_247),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_283),
.C(n_271),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_252),
.A2(n_240),
.B(n_249),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_276),
.B(n_279),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_249),
.Y(n_276)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_277),
.A2(n_258),
.B(n_265),
.Y(n_285)
);

XNOR2x1_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_238),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_L g290 ( 
.A1(n_282),
.A2(n_201),
.B(n_200),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_269),
.Y(n_283)
);

OAI322xp33_ASAP7_75t_L g284 ( 
.A1(n_280),
.A2(n_263),
.A3(n_187),
.B1(n_257),
.B2(n_259),
.C1(n_261),
.C2(n_260),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_284),
.A2(n_289),
.B(n_276),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_285),
.A2(n_287),
.B(n_2),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_292),
.Y(n_300)
);

AO21x1_ASAP7_75t_L g287 ( 
.A1(n_277),
.A2(n_233),
.B(n_236),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_288),
.B(n_290),
.Y(n_296)
);

OAI322xp33_ASAP7_75t_L g289 ( 
.A1(n_272),
.A2(n_266),
.A3(n_255),
.B1(n_237),
.B2(n_208),
.C1(n_206),
.C2(n_268),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g292 ( 
.A(n_275),
.B(n_217),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_271),
.B(n_281),
.C(n_274),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_293),
.B(n_4),
.Y(n_302)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_295),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_294),
.A2(n_270),
.B1(n_278),
.B2(n_199),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_297),
.B(n_299),
.C(n_302),
.Y(n_303)
);

NOR3xp33_ASAP7_75t_L g298 ( 
.A(n_291),
.B(n_283),
.C(n_281),
.Y(n_298)
);

NOR4xp25_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_4),
.C(n_5),
.D(n_6),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g301 ( 
.A1(n_287),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_301),
.A2(n_285),
.B1(n_5),
.B2(n_6),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_292),
.C(n_286),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_304),
.B(n_306),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g309 ( 
.A1(n_305),
.A2(n_299),
.B1(n_297),
.B2(n_300),
.Y(n_309)
);

NOR3xp33_ASAP7_75t_L g311 ( 
.A(n_309),
.B(n_310),
.C(n_307),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_303),
.Y(n_310)
);

OAI21x1_ASAP7_75t_L g313 ( 
.A1(n_311),
.A2(n_312),
.B(n_6),
.Y(n_313)
);

NOR3xp33_ASAP7_75t_L g312 ( 
.A(n_308),
.B(n_300),
.C(n_7),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_313),
.B(n_8),
.C(n_9),
.Y(n_314)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_314),
.B(n_8),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_8),
.Y(n_316)
);


endmodule