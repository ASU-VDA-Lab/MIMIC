module fake_jpeg_13337_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g11 ( 
.A(n_0),
.Y(n_11)
);

INVx2_ASAP7_75t_SL g12 ( 
.A(n_9),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_23),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_25),
.Y(n_43)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_13),
.B(n_1),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_32),
.Y(n_38)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

BUFx4f_ASAP7_75t_SL g33 ( 
.A(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_33),
.B(n_25),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_35),
.B(n_36),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_20),
.C(n_14),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_20),
.C(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_42),
.Y(n_51)
);

AO22x2_ASAP7_75t_SL g41 ( 
.A1(n_26),
.A2(n_17),
.B1(n_2),
.B2(n_1),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_41),
.A2(n_27),
.B1(n_28),
.B2(n_44),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_33),
.B(n_18),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_18),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_33),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_52),
.Y(n_68)
);

A2O1A1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_38),
.A2(n_29),
.B(n_16),
.C(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_49),
.B(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_50),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_34),
.B(n_22),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_17),
.Y(n_54)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_54),
.B(n_57),
.C(n_58),
.Y(n_61)
);

INVxp67_ASAP7_75t_SL g55 ( 
.A(n_43),
.Y(n_55)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_55),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_21),
.Y(n_56)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_15),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_27),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_39),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_31),
.B(n_2),
.Y(n_67)
);

XNOR2x1_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_45),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_60),
.B(n_65),
.C(n_69),
.Y(n_77)
);

AND2x6_ASAP7_75t_L g63 ( 
.A(n_51),
.B(n_8),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_3),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g65 ( 
.A(n_59),
.B(n_37),
.C(n_16),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_67),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_58),
.B(n_24),
.C(n_2),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_57),
.A2(n_24),
.B1(n_4),
.B2(n_5),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g73 ( 
.A1(n_71),
.A2(n_47),
.B1(n_54),
.B2(n_58),
.Y(n_73)
);

OR2x2_ASAP7_75t_L g72 ( 
.A(n_66),
.B(n_49),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_73),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_50),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_75),
.B(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_5),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_68),
.A2(n_24),
.B1(n_6),
.B2(n_9),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_70),
.Y(n_79)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_73),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_78),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_77),
.Y(n_89)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_89),
.B(n_90),
.Y(n_96)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_74),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_82),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_91),
.B(n_92),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_88),
.Y(n_93)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_93),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_84),
.B1(n_81),
.B2(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_95),
.B(n_83),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_98),
.B(n_99),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_77),
.B1(n_82),
.B2(n_63),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_96),
.B(n_90),
.C(n_97),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_96),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_102),
.B(n_65),
.C(n_69),
.Y(n_103)
);

AO21x1_ASAP7_75t_L g105 ( 
.A1(n_103),
.A2(n_104),
.B(n_67),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_62),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_62),
.Y(n_106)
);


endmodule