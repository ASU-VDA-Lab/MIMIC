module fake_jpeg_982_n_198 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_198);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_198;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

INVx8_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

INVx3_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_1),
.B(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx11_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_6),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_13),
.B(n_0),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx10_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_11),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_37),
.B(n_38),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_14),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_39),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_25),
.Y(n_42)
);

INVx5_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_29),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_43),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_44),
.Y(n_71)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_26),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_28),
.B(n_14),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_46),
.B(n_21),
.Y(n_73)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_47),
.Y(n_63)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_48),
.Y(n_69)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_50),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_23),
.B(n_2),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_20),
.C(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_52),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_54),
.B(n_55),
.Y(n_74)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_56),
.A2(n_33),
.B(n_32),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_62),
.B(n_2),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_16),
.C(n_32),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_64),
.B(n_80),
.C(n_84),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_42),
.Y(n_66)
);

CKINVDCx5p33_ASAP7_75t_R g103 ( 
.A(n_66),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_52),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_68),
.B(n_73),
.Y(n_107)
);

OR2x4_ASAP7_75t_L g108 ( 
.A(n_70),
.B(n_31),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g89 ( 
.A(n_72),
.Y(n_89)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_21),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_77),
.B(n_79),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_41),
.B(n_16),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_47),
.A2(n_27),
.B(n_22),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_SL g82 ( 
.A1(n_48),
.A2(n_33),
.B(n_31),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_82),
.A2(n_22),
.B(n_30),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_19),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_83),
.B(n_27),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_31),
.C(n_30),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_84),
.A2(n_40),
.B1(n_53),
.B2(n_36),
.Y(n_87)
);

AO21x2_ASAP7_75t_L g126 ( 
.A1(n_87),
.A2(n_71),
.B(n_67),
.Y(n_126)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_88),
.B(n_109),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_65),
.A2(n_44),
.B1(n_43),
.B2(n_26),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_90),
.A2(n_98),
.B1(n_101),
.B2(n_59),
.Y(n_130)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g118 ( 
.A(n_93),
.Y(n_118)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_95),
.B(n_96),
.Y(n_123)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_69),
.B(n_54),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_97),
.B(n_100),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_76),
.A2(n_50),
.B1(n_39),
.B2(n_15),
.Y(n_98)
);

O2A1O1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_82),
.A2(n_31),
.B(n_26),
.C(n_34),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_99),
.B(n_66),
.Y(n_116)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_76),
.A2(n_15),
.B1(n_31),
.B2(n_25),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_60),
.B(n_12),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_102),
.B(n_105),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_4),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_85),
.B(n_11),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_74),
.A2(n_85),
.B(n_57),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_106),
.A2(n_61),
.B(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_108),
.B(n_3),
.Y(n_120)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_74),
.Y(n_109)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_57),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_112),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

OAI21xp33_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_120),
.B(n_125),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_88),
.A2(n_78),
.B1(n_71),
.B2(n_67),
.Y(n_115)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_115),
.A2(n_116),
.B1(n_89),
.B2(n_58),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_110),
.B(n_78),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_100),
.C(n_96),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_110),
.B(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_121),
.B(n_128),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_103),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_126),
.A2(n_130),
.B1(n_133),
.B2(n_101),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_127),
.B(n_129),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_97),
.B(n_59),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_91),
.B(n_4),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_107),
.B(n_15),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_132),
.B(n_92),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_109),
.A2(n_58),
.B1(n_66),
.B2(n_34),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_129),
.B(n_104),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_142),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_122),
.A2(n_99),
.B(n_106),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_137),
.A2(n_148),
.B(n_126),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_121),
.B(n_97),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_138),
.B(n_139),
.C(n_140),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_119),
.B(n_94),
.C(n_93),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_112),
.C(n_111),
.Y(n_141)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_141),
.B(n_117),
.C(n_118),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_131),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_143),
.Y(n_153)
);

FAx1_ASAP7_75t_SL g144 ( 
.A(n_122),
.B(n_103),
.CI(n_98),
.CON(n_144),
.SN(n_144)
);

AOI322xp5_ASAP7_75t_L g154 ( 
.A1(n_144),
.A2(n_124),
.A3(n_120),
.B1(n_128),
.B2(n_113),
.C1(n_123),
.C2(n_126),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_145),
.A2(n_151),
.B1(n_126),
.B2(n_124),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_92),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_146),
.B(n_147),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_117),
.Y(n_149)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_125),
.B(n_116),
.Y(n_152)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_152),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_154),
.A2(n_157),
.B1(n_151),
.B2(n_142),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_141),
.Y(n_173)
);

AO21x1_ASAP7_75t_L g160 ( 
.A1(n_136),
.A2(n_123),
.B(n_126),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_160),
.B(n_163),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_150),
.A2(n_133),
.B(n_118),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_161),
.B(n_144),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_136),
.B(n_89),
.C(n_130),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_164),
.B(n_139),
.C(n_140),
.Y(n_168)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_149),
.Y(n_165)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_165),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_166),
.A2(n_162),
.B(n_152),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_167),
.B(n_170),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_168),
.B(n_173),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_159),
.B(n_134),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_143),
.C(n_138),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_172),
.B(n_174),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_156),
.B(n_148),
.C(n_145),
.Y(n_174)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_171),
.A2(n_162),
.A3(n_159),
.B1(n_160),
.B2(n_175),
.C1(n_153),
.C2(n_163),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_169),
.B(n_153),
.Y(n_181)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_181),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_175),
.A2(n_164),
.B1(n_161),
.B2(n_158),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g186 ( 
.A(n_182),
.Y(n_186)
);

AOI31xp67_ASAP7_75t_L g184 ( 
.A1(n_180),
.A2(n_174),
.A3(n_168),
.B(n_165),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_SL g190 ( 
.A(n_184),
.B(n_182),
.Y(n_190)
);

FAx1_ASAP7_75t_R g185 ( 
.A(n_178),
.B(n_173),
.CI(n_144),
.CON(n_185),
.SN(n_185)
);

NAND3xp33_ASAP7_75t_L g191 ( 
.A(n_185),
.B(n_155),
.C(n_126),
.Y(n_191)
);

NOR2xp67_ASAP7_75t_SL g188 ( 
.A(n_187),
.B(n_176),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_188),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_186),
.B(n_176),
.C(n_179),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_189),
.B(n_190),
.C(n_191),
.Y(n_194)
);

AOI322xp5_ASAP7_75t_L g193 ( 
.A1(n_190),
.A2(n_185),
.A3(n_183),
.B1(n_155),
.B2(n_9),
.C1(n_5),
.C2(n_8),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_193),
.B(n_6),
.C(n_8),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_195),
.B(n_196),
.C(n_192),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g196 ( 
.A1(n_194),
.A2(n_6),
.B(n_8),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g198 ( 
.A(n_197),
.B(n_9),
.Y(n_198)
);


endmodule