module fake_jpeg_8581_n_118 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_118);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_118;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_116;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx8_ASAP7_75t_L g42 ( 
.A(n_38),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_39),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_27),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_10),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_8),
.Y(n_48)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_0),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_9),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx6f_ASAP7_75t_SL g55 ( 
.A(n_14),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_19),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_55),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_61),
.B(n_2),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_56),
.Y(n_62)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_52),
.Y(n_63)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_45),
.B(n_0),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_66),
.B(n_2),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_44),
.B(n_1),
.Y(n_67)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_67),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_68),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_69),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_58),
.Y(n_70)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_70),
.Y(n_73)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_66),
.A2(n_49),
.B1(n_54),
.B2(n_42),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_75),
.A2(n_84),
.B1(n_85),
.B2(n_88),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_76),
.B(n_81),
.Y(n_91)
);

AND2x2_ASAP7_75t_L g77 ( 
.A(n_66),
.B(n_1),
.Y(n_77)
);

NOR2x1_ASAP7_75t_R g100 ( 
.A(n_77),
.B(n_20),
.Y(n_100)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_79),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_57),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_SL g92 ( 
.A(n_83),
.B(n_87),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g84 ( 
.A1(n_63),
.A2(n_48),
.B1(n_46),
.B2(n_43),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_63),
.A2(n_60),
.B1(n_53),
.B2(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_65),
.A2(n_42),
.B1(n_3),
.B2(n_5),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_89),
.B(n_21),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_73),
.A2(n_3),
.B1(n_4),
.B2(n_7),
.Y(n_94)
);

NOR2x1_ASAP7_75t_R g103 ( 
.A(n_94),
.B(n_97),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_85),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_82),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g98 ( 
.A1(n_90),
.A2(n_11),
.B1(n_12),
.B2(n_15),
.Y(n_98)
);

OA22x2_ASAP7_75t_L g99 ( 
.A1(n_80),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_72),
.B(n_22),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_92),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_74),
.C(n_91),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_106),
.B(n_96),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_107),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_108),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_109),
.B(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_102),
.B1(n_103),
.B2(n_100),
.Y(n_111)
);

OAI321xp33_ASAP7_75t_L g112 ( 
.A1(n_111),
.A2(n_99),
.A3(n_93),
.B1(n_98),
.B2(n_101),
.C(n_71),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_112),
.B(n_99),
.C(n_86),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_113),
.B(n_25),
.Y(n_114)
);

MAJx2_ASAP7_75t_L g115 ( 
.A(n_114),
.B(n_26),
.C(n_28),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_31),
.C(n_32),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_116),
.B(n_33),
.C(n_34),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g118 ( 
.A(n_117),
.B(n_35),
.Y(n_118)
);


endmodule