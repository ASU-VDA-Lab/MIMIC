module real_aes_2224_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_792;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_571;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_537;
wire n_320;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_578;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_774;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_781;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_505;
wire n_502;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_785;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_637;
wire n_526;
wire n_155;
wire n_243;
wire n_692;
wire n_789;
wire n_268;
wire n_544;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_546;
wire n_151;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_0), .B(n_147), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g155 ( .A1(n_1), .A2(n_156), .B(n_161), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_2), .B(n_107), .Y(n_106) );
CKINVDCx20_ASAP7_75t_R g793 ( .A(n_3), .Y(n_793) );
NAND2xp5_ASAP7_75t_SL g201 ( .A(n_4), .B(n_163), .Y(n_201) );
INVx1_ASAP7_75t_L g154 ( .A(n_5), .Y(n_154) );
NAND2xp5_ASAP7_75t_L g229 ( .A(n_6), .B(n_163), .Y(n_229) );
NAND2xp5_ASAP7_75t_SL g556 ( .A(n_7), .B(n_173), .Y(n_556) );
INVx1_ASAP7_75t_L g536 ( .A(n_8), .Y(n_536) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_9), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g125 ( .A(n_10), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g502 ( .A(n_11), .Y(n_502) );
NAND2xp33_ASAP7_75t_L g190 ( .A(n_12), .B(n_165), .Y(n_190) );
INVx2_ASAP7_75t_L g144 ( .A(n_13), .Y(n_144) );
AOI221x1_ASAP7_75t_L g236 ( .A1(n_14), .A2(n_26), .B1(n_147), .B2(n_156), .C(n_237), .Y(n_236) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_15), .Y(n_108) );
NAND2xp5_ASAP7_75t_SL g186 ( .A(n_16), .B(n_147), .Y(n_186) );
AO21x2_ASAP7_75t_L g183 ( .A1(n_17), .A2(n_184), .B(n_185), .Y(n_183) );
INVx1_ASAP7_75t_L g564 ( .A(n_18), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_19), .B(n_167), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g177 ( .A(n_20), .B(n_163), .Y(n_177) );
AO21x1_ASAP7_75t_L g196 ( .A1(n_21), .A2(n_147), .B(n_197), .Y(n_196) );
NOR2xp33_ASAP7_75t_SL g103 ( .A(n_22), .B(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g124 ( .A(n_22), .Y(n_124) );
INVx1_ASAP7_75t_L g562 ( .A(n_23), .Y(n_562) );
INVx1_ASAP7_75t_SL g484 ( .A(n_24), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g552 ( .A(n_25), .B(n_148), .Y(n_552) );
NAND2x1_ASAP7_75t_L g209 ( .A(n_27), .B(n_163), .Y(n_209) );
AOI33xp33_ASAP7_75t_L g522 ( .A1(n_28), .A2(n_54), .A3(n_467), .B1(n_472), .B2(n_523), .B3(n_524), .Y(n_522) );
NAND2x1_ASAP7_75t_L g228 ( .A(n_29), .B(n_165), .Y(n_228) );
INVx1_ASAP7_75t_L g495 ( .A(n_30), .Y(n_495) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_31), .A2(n_88), .B(n_144), .Y(n_143) );
OR2x2_ASAP7_75t_L g169 ( .A(n_31), .B(n_88), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_32), .B(n_475), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_33), .B(n_165), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_34), .B(n_163), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_35), .B(n_165), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_36), .A2(n_156), .B(n_217), .Y(n_216) );
AND2x2_ASAP7_75t_L g153 ( .A(n_37), .B(n_154), .Y(n_153) );
AND2x2_ASAP7_75t_L g157 ( .A(n_37), .B(n_158), .Y(n_157) );
INVx1_ASAP7_75t_L g466 ( .A(n_37), .Y(n_466) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_38), .B(n_106), .C(n_108), .Y(n_105) );
OR2x6_ASAP7_75t_L g122 ( .A(n_38), .B(n_123), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g498 ( .A(n_39), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g220 ( .A(n_40), .B(n_147), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_41), .B(n_475), .Y(n_509) );
AOI22xp5_ASAP7_75t_L g545 ( .A1(n_42), .A2(n_142), .B1(n_173), .B2(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_43), .B(n_554), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_44), .B(n_148), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_45), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g218 ( .A(n_46), .B(n_165), .Y(n_218) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_47), .B(n_184), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_48), .B(n_148), .Y(n_537) );
AOI21xp5_ASAP7_75t_L g226 ( .A1(n_49), .A2(n_156), .B(n_227), .Y(n_226) );
CKINVDCx5p33_ASAP7_75t_R g549 ( .A(n_50), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g800 ( .A1(n_51), .A2(n_84), .B1(n_801), .B2(n_802), .Y(n_800) );
CKINVDCx20_ASAP7_75t_R g802 ( .A(n_51), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_52), .A2(n_79), .B1(n_784), .B2(n_785), .Y(n_783) );
CKINVDCx20_ASAP7_75t_R g785 ( .A(n_52), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_53), .B(n_165), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_55), .B(n_148), .Y(n_513) );
INVx1_ASAP7_75t_L g150 ( .A(n_56), .Y(n_150) );
INVx1_ASAP7_75t_L g160 ( .A(n_56), .Y(n_160) );
AND2x2_ASAP7_75t_L g514 ( .A(n_57), .B(n_167), .Y(n_514) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_58), .A2(n_74), .B1(n_464), .B2(n_475), .C(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_59), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g239 ( .A(n_60), .B(n_163), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_61), .B(n_142), .Y(n_504) );
AOI21xp5_ASAP7_75t_SL g463 ( .A1(n_62), .A2(n_464), .B(n_469), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g207 ( .A1(n_63), .A2(n_156), .B(n_208), .Y(n_207) );
INVx1_ASAP7_75t_L g559 ( .A(n_64), .Y(n_559) );
AO21x1_ASAP7_75t_L g198 ( .A1(n_65), .A2(n_156), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_SL g146 ( .A(n_66), .B(n_147), .Y(n_146) );
INVx1_ASAP7_75t_L g512 ( .A(n_67), .Y(n_512) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_68), .B(n_147), .Y(n_230) );
AOI21xp5_ASAP7_75t_L g510 ( .A1(n_69), .A2(n_464), .B(n_511), .Y(n_510) );
AND2x2_ASAP7_75t_L g221 ( .A(n_70), .B(n_168), .Y(n_221) );
INVx1_ASAP7_75t_L g152 ( .A(n_71), .Y(n_152) );
INVx1_ASAP7_75t_L g158 ( .A(n_71), .Y(n_158) );
AND2x2_ASAP7_75t_L g232 ( .A(n_72), .B(n_141), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_73), .B(n_475), .Y(n_525) );
AND2x2_ASAP7_75t_L g486 ( .A(n_75), .B(n_141), .Y(n_486) );
INVx1_ASAP7_75t_L g560 ( .A(n_76), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_77), .A2(n_464), .B(n_483), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g550 ( .A1(n_78), .A2(n_464), .B(n_517), .C(n_551), .Y(n_550) );
CKINVDCx20_ASAP7_75t_R g784 ( .A(n_79), .Y(n_784) );
INVx1_ASAP7_75t_L g104 ( .A(n_80), .Y(n_104) );
AND2x2_ASAP7_75t_L g140 ( .A(n_81), .B(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_82), .B(n_147), .Y(n_179) );
AND2x2_ASAP7_75t_SL g461 ( .A(n_83), .B(n_141), .Y(n_461) );
INVx1_ASAP7_75t_L g801 ( .A(n_84), .Y(n_801) );
AOI22xp5_ASAP7_75t_L g519 ( .A1(n_85), .A2(n_464), .B1(n_520), .B2(n_521), .Y(n_519) );
AND2x2_ASAP7_75t_L g197 ( .A(n_86), .B(n_173), .Y(n_197) );
INVxp33_ASAP7_75t_L g809 ( .A(n_87), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_89), .B(n_165), .Y(n_178) );
AND2x2_ASAP7_75t_L g213 ( .A(n_90), .B(n_141), .Y(n_213) );
INVx1_ASAP7_75t_L g470 ( .A(n_91), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_92), .B(n_163), .Y(n_219) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_93), .A2(n_156), .B(n_176), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_94), .B(n_165), .Y(n_238) );
AND2x2_ASAP7_75t_L g526 ( .A(n_95), .B(n_141), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_96), .B(n_163), .Y(n_162) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_97), .A2(n_493), .B(n_494), .C(n_497), .Y(n_492) );
BUFx2_ASAP7_75t_L g113 ( .A(n_98), .Y(n_113) );
BUFx2_ASAP7_75t_SL g796 ( .A(n_98), .Y(n_796) );
AOI21xp5_ASAP7_75t_L g187 ( .A1(n_99), .A2(n_156), .B(n_188), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_100), .B(n_148), .Y(n_473) );
AOI21xp33_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_109), .B(n_808), .Y(n_101) );
INVx2_ASAP7_75t_L g812 ( .A(n_102), .Y(n_812) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g123 ( .A(n_104), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_L g120 ( .A(n_108), .B(n_121), .Y(n_120) );
AND2x6_ASAP7_75t_SL g130 ( .A(n_108), .B(n_122), .Y(n_130) );
OR2x6_ASAP7_75t_SL g450 ( .A(n_108), .B(n_121), .Y(n_450) );
OR2x2_ASAP7_75t_L g792 ( .A(n_108), .B(n_122), .Y(n_792) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_126), .B(n_794), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g110 ( .A(n_111), .B(n_114), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g111 ( .A(n_112), .Y(n_111) );
CKINVDCx20_ASAP7_75t_R g112 ( .A(n_113), .Y(n_112) );
INVxp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g797 ( .A1(n_115), .A2(n_798), .B(n_805), .Y(n_797) );
NOR2xp33_ASAP7_75t_SL g115 ( .A(n_116), .B(n_125), .Y(n_115) );
INVx1_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_119), .Y(n_118) );
BUFx3_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
BUFx2_ASAP7_75t_R g807 ( .A(n_120), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g121 ( .A(n_122), .Y(n_121) );
OAI222xp33_ASAP7_75t_L g126 ( .A1(n_127), .A2(n_783), .B1(n_786), .B2(n_787), .C1(n_792), .C2(n_793), .Y(n_126) );
AOI22x1_ASAP7_75t_L g127 ( .A1(n_128), .A2(n_131), .B1(n_449), .B2(n_451), .Y(n_127) );
INVx3_ASAP7_75t_SL g128 ( .A(n_129), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
CKINVDCx11_ASAP7_75t_R g791 ( .A(n_130), .Y(n_791) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
INVx3_ASAP7_75t_L g790 ( .A(n_132), .Y(n_790) );
INVx1_ASAP7_75t_L g799 ( .A(n_132), .Y(n_799) );
AND2x4_ASAP7_75t_L g132 ( .A(n_133), .B(n_358), .Y(n_132) );
NOR4xp25_ASAP7_75t_L g133 ( .A(n_134), .B(n_276), .C(n_302), .D(n_342), .Y(n_133) );
OAI211xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_191), .B(n_222), .C(n_262), .Y(n_134) );
INVxp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_170), .Y(n_136) );
AND2x2_ASAP7_75t_L g429 ( .A(n_137), .B(n_430), .Y(n_429) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_138), .B(n_170), .Y(n_296) );
BUFx2_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x2_ASAP7_75t_L g223 ( .A(n_139), .B(n_224), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_139), .B(n_249), .Y(n_248) );
INVx5_ASAP7_75t_L g282 ( .A(n_139), .Y(n_282) );
NOR2x1_ASAP7_75t_SL g324 ( .A(n_139), .B(n_171), .Y(n_324) );
AND2x2_ASAP7_75t_L g380 ( .A(n_139), .B(n_183), .Y(n_380) );
OR2x6_ASAP7_75t_L g139 ( .A(n_140), .B(n_145), .Y(n_139) );
INVx3_ASAP7_75t_L g212 ( .A(n_141), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g491 ( .A1(n_141), .A2(n_212), .B1(n_492), .B2(n_498), .Y(n_491) );
INVx4_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_142), .B(n_501), .Y(n_500) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx4f_ASAP7_75t_L g184 ( .A(n_143), .Y(n_184) );
AND2x2_ASAP7_75t_SL g168 ( .A(n_144), .B(n_169), .Y(n_168) );
AND2x4_ASAP7_75t_L g173 ( .A(n_144), .B(n_169), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_155), .B(n_167), .Y(n_145) );
AND2x4_ASAP7_75t_L g147 ( .A(n_148), .B(n_153), .Y(n_147) );
INVx1_ASAP7_75t_L g496 ( .A(n_148), .Y(n_496) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_151), .Y(n_148) );
AND2x6_ASAP7_75t_L g165 ( .A(n_149), .B(n_158), .Y(n_165) );
INVx2_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g163 ( .A(n_151), .B(n_160), .Y(n_163) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx5_ASAP7_75t_L g166 ( .A(n_153), .Y(n_166) );
HB1xp67_ASAP7_75t_L g497 ( .A(n_153), .Y(n_497) );
AND2x2_ASAP7_75t_L g159 ( .A(n_154), .B(n_160), .Y(n_159) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_154), .Y(n_477) );
AND2x6_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
BUFx3_ASAP7_75t_L g478 ( .A(n_157), .Y(n_478) );
INVx2_ASAP7_75t_L g468 ( .A(n_158), .Y(n_468) );
AND2x4_ASAP7_75t_L g464 ( .A(n_159), .B(n_465), .Y(n_464) );
INVx2_ASAP7_75t_L g472 ( .A(n_160), .Y(n_472) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_162), .A2(n_164), .B(n_166), .Y(n_161) );
INVxp67_ASAP7_75t_L g565 ( .A(n_163), .Y(n_565) );
INVxp67_ASAP7_75t_L g563 ( .A(n_165), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g176 ( .A1(n_166), .A2(n_177), .B(n_178), .Y(n_176) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_166), .A2(n_189), .B(n_190), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_166), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_166), .A2(n_209), .B(n_210), .Y(n_208) );
AOI21xp5_ASAP7_75t_L g217 ( .A1(n_166), .A2(n_218), .B(n_219), .Y(n_217) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_166), .A2(n_228), .B(n_229), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_166), .A2(n_238), .B(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g469 ( .A1(n_166), .A2(n_470), .B(n_471), .C(n_473), .Y(n_469) );
O2A1O1Ixp33_ASAP7_75t_SL g483 ( .A1(n_166), .A2(n_471), .B(n_484), .C(n_485), .Y(n_483) );
O2A1O1Ixp33_ASAP7_75t_L g511 ( .A1(n_166), .A2(n_471), .B(n_512), .C(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g520 ( .A(n_166), .Y(n_520) );
O2A1O1Ixp33_ASAP7_75t_SL g535 ( .A1(n_166), .A2(n_471), .B(n_536), .C(n_537), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_166), .A2(n_552), .B(n_553), .Y(n_551) );
NOR2xp33_ASAP7_75t_L g566 ( .A(n_166), .B(n_173), .Y(n_566) );
CKINVDCx5p33_ASAP7_75t_R g231 ( .A(n_167), .Y(n_231) );
OA21x2_ASAP7_75t_L g235 ( .A1(n_167), .A2(n_236), .B(n_240), .Y(n_235) );
OA21x2_ASAP7_75t_L g275 ( .A1(n_167), .A2(n_236), .B(n_240), .Y(n_275) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_168), .Y(n_167) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_182), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_171), .B(n_183), .Y(n_252) );
AND2x2_ASAP7_75t_L g313 ( .A(n_171), .B(n_282), .Y(n_313) );
AO21x2_ASAP7_75t_L g171 ( .A1(n_172), .A2(n_174), .B(n_180), .Y(n_171) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_172), .B(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g266 ( .A1(n_172), .A2(n_174), .B(n_180), .Y(n_266) );
INVx1_ASAP7_75t_SL g172 ( .A(n_173), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g185 ( .A1(n_173), .A2(n_186), .B(n_187), .Y(n_185) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_173), .B(n_203), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g462 ( .A1(n_173), .A2(n_463), .B(n_474), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_175), .B(n_179), .Y(n_174) );
AND2x2_ASAP7_75t_L g325 ( .A(n_182), .B(n_249), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_182), .B(n_330), .Y(n_329) );
OR2x2_ASAP7_75t_L g369 ( .A(n_182), .B(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g402 ( .A(n_182), .B(n_223), .Y(n_402) );
INVx2_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
INVx1_ASAP7_75t_L g246 ( .A(n_183), .Y(n_246) );
AND2x2_ASAP7_75t_L g279 ( .A(n_183), .B(n_280), .Y(n_279) );
BUFx3_ASAP7_75t_L g314 ( .A(n_183), .Y(n_314) );
OR2x2_ASAP7_75t_L g390 ( .A(n_183), .B(n_249), .Y(n_390) );
INVx2_ASAP7_75t_SL g517 ( .A(n_184), .Y(n_517) );
OA21x2_ASAP7_75t_L g533 ( .A1(n_184), .A2(n_534), .B(n_538), .Y(n_533) );
INVx1_ASAP7_75t_SL g191 ( .A(n_192), .Y(n_191) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_204), .Y(n_192) );
AOI211x1_ASAP7_75t_SL g319 ( .A1(n_193), .A2(n_311), .B(n_320), .C(n_322), .Y(n_319) );
AND2x2_ASAP7_75t_SL g364 ( .A(n_193), .B(n_365), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_193), .B(n_362), .Y(n_409) );
BUFx2_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx2_ASAP7_75t_L g259 ( .A(n_194), .Y(n_259) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx2_ASAP7_75t_L g234 ( .A(n_195), .Y(n_234) );
OAI21x1_ASAP7_75t_SL g195 ( .A1(n_196), .A2(n_198), .B(n_202), .Y(n_195) );
INVx1_ASAP7_75t_L g203 ( .A(n_197), .Y(n_203) );
AOI322xp5_ASAP7_75t_L g222 ( .A1(n_204), .A2(n_223), .A3(n_233), .B1(n_241), .B2(n_244), .C1(n_250), .C2(n_253), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_204), .B(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_214), .Y(n_204) );
INVx2_ASAP7_75t_L g257 ( .A(n_205), .Y(n_257) );
INVxp67_ASAP7_75t_L g299 ( .A(n_205), .Y(n_299) );
BUFx3_ASAP7_75t_L g363 ( .A(n_205), .Y(n_363) );
AO21x2_ASAP7_75t_L g205 ( .A1(n_206), .A2(n_212), .B(n_213), .Y(n_205) );
AO21x2_ASAP7_75t_L g243 ( .A1(n_206), .A2(n_212), .B(n_213), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_211), .Y(n_206) );
AO21x2_ASAP7_75t_L g214 ( .A1(n_212), .A2(n_215), .B(n_221), .Y(n_214) );
AO21x2_ASAP7_75t_L g261 ( .A1(n_212), .A2(n_215), .B(n_221), .Y(n_261) );
AO21x2_ASAP7_75t_L g507 ( .A1(n_212), .A2(n_508), .B(n_514), .Y(n_507) );
AO21x2_ASAP7_75t_L g530 ( .A1(n_212), .A2(n_508), .B(n_514), .Y(n_530) );
INVx2_ASAP7_75t_L g272 ( .A(n_214), .Y(n_272) );
AND2x2_ASAP7_75t_L g321 ( .A(n_214), .B(n_235), .Y(n_321) );
AND2x2_ASAP7_75t_L g365 ( .A(n_214), .B(n_274), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_216), .B(n_220), .Y(n_215) );
AND2x2_ASAP7_75t_L g250 ( .A(n_223), .B(n_251), .Y(n_250) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_223), .B(n_435), .Y(n_434) );
AND2x2_ASAP7_75t_SL g444 ( .A(n_223), .B(n_279), .Y(n_444) );
INVx4_ASAP7_75t_L g249 ( .A(n_224), .Y(n_249) );
AND2x2_ASAP7_75t_L g281 ( .A(n_224), .B(n_282), .Y(n_281) );
HB1xp67_ASAP7_75t_L g334 ( .A(n_224), .Y(n_334) );
AO21x2_ASAP7_75t_L g224 ( .A1(n_225), .A2(n_231), .B(n_232), .Y(n_224) );
NAND2xp5_ASAP7_75t_L g225 ( .A(n_226), .B(n_230), .Y(n_225) );
AO21x2_ASAP7_75t_L g479 ( .A1(n_231), .A2(n_480), .B(n_486), .Y(n_479) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_233), .B(n_318), .Y(n_343) );
INVx1_ASAP7_75t_SL g382 ( .A(n_233), .Y(n_382) );
AND2x4_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
AND2x4_ASAP7_75t_L g273 ( .A(n_234), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_234), .B(n_272), .Y(n_341) );
AND2x2_ASAP7_75t_L g393 ( .A(n_234), .B(n_243), .Y(n_393) );
OR2x2_ASAP7_75t_L g417 ( .A(n_234), .B(n_235), .Y(n_417) );
AND2x2_ASAP7_75t_L g241 ( .A(n_235), .B(n_242), .Y(n_241) );
AND2x2_ASAP7_75t_L g291 ( .A(n_235), .B(n_272), .Y(n_291) );
AND2x2_ASAP7_75t_SL g347 ( .A(n_235), .B(n_259), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_241), .B(n_354), .Y(n_371) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
BUFx2_ASAP7_75t_L g306 ( .A(n_243), .Y(n_306) );
AND2x4_ASAP7_75t_SL g346 ( .A(n_243), .B(n_260), .Y(n_346) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_247), .Y(n_244) );
OR2x2_ASAP7_75t_L g294 ( .A(n_245), .B(n_248), .Y(n_294) );
INVx1_ASAP7_75t_L g245 ( .A(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g263 ( .A(n_246), .B(n_264), .Y(n_263) );
AND2x2_ASAP7_75t_L g411 ( .A(n_246), .B(n_324), .Y(n_411) );
AND2x2_ASAP7_75t_L g427 ( .A(n_246), .B(n_281), .Y(n_427) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
AOI311xp33_ASAP7_75t_L g397 ( .A1(n_248), .A2(n_336), .A3(n_398), .B(n_400), .C(n_407), .Y(n_397) );
AND2x4_ASAP7_75t_L g264 ( .A(n_249), .B(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g268 ( .A(n_249), .Y(n_268) );
NAND2x1p5_ASAP7_75t_L g338 ( .A(n_249), .B(n_282), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_249), .B(n_368), .Y(n_367) );
AND2x2_ASAP7_75t_L g381 ( .A(n_249), .B(n_368), .Y(n_381) );
AND2x2_ASAP7_75t_L g267 ( .A(n_251), .B(n_268), .Y(n_267) );
INVxp67_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
INVxp67_ASAP7_75t_SL g285 ( .A(n_252), .Y(n_285) );
OR2x2_ASAP7_75t_L g374 ( .A(n_252), .B(n_338), .Y(n_374) );
INVx1_ASAP7_75t_L g430 ( .A(n_252), .Y(n_430) );
INVx1_ASAP7_75t_SL g253 ( .A(n_254), .Y(n_253) );
OR2x2_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g339 ( .A(n_256), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g353 ( .A(n_256), .B(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g428 ( .A(n_256), .B(n_301), .Y(n_428) );
BUFx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
AND2x2_ASAP7_75t_L g271 ( .A(n_257), .B(n_272), .Y(n_271) );
AND2x2_ASAP7_75t_L g290 ( .A(n_257), .B(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g352 ( .A(n_258), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g407 ( .A1(n_258), .A2(n_408), .B1(n_409), .B2(n_410), .Y(n_407) );
OR2x2_ASAP7_75t_L g258 ( .A(n_259), .B(n_260), .Y(n_258) );
AND2x2_ASAP7_75t_L g301 ( .A(n_259), .B(n_272), .Y(n_301) );
AND2x4_ASAP7_75t_L g354 ( .A(n_259), .B(n_261), .Y(n_354) );
INVx2_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
OAI21xp33_ASAP7_75t_SL g262 ( .A1(n_263), .A2(n_267), .B(n_269), .Y(n_262) );
AOI22xp5_ASAP7_75t_L g348 ( .A1(n_263), .A2(n_349), .B1(n_353), .B2(n_355), .Y(n_348) );
AND2x2_ASAP7_75t_SL g308 ( .A(n_264), .B(n_282), .Y(n_308) );
INVx2_ASAP7_75t_L g370 ( .A(n_264), .Y(n_370) );
AND2x2_ASAP7_75t_L g384 ( .A(n_264), .B(n_380), .Y(n_384) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g280 ( .A(n_266), .Y(n_280) );
INVx1_ASAP7_75t_L g333 ( .A(n_266), .Y(n_333) );
INVx1_ASAP7_75t_L g284 ( .A(n_268), .Y(n_284) );
AND3x2_ASAP7_75t_L g312 ( .A(n_268), .B(n_313), .C(n_314), .Y(n_312) );
INVx1_ASAP7_75t_SL g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g376 ( .A(n_271), .Y(n_376) );
AND2x2_ASAP7_75t_L g304 ( .A(n_273), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g375 ( .A(n_273), .B(n_376), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g386 ( .A1(n_273), .A2(n_387), .B1(n_391), .B2(n_394), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g425 ( .A(n_273), .B(n_421), .Y(n_425) );
BUFx2_ASAP7_75t_L g316 ( .A(n_274), .Y(n_316) );
INVx2_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx2_ASAP7_75t_L g287 ( .A(n_275), .Y(n_287) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_275), .Y(n_406) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_277), .A2(n_286), .B1(n_288), .B2(n_289), .C(n_292), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_283), .Y(n_277) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx1_ASAP7_75t_L g368 ( .A(n_280), .Y(n_368) );
INVx2_ASAP7_75t_SL g357 ( .A(n_281), .Y(n_357) );
AND2x2_ASAP7_75t_L g439 ( .A(n_281), .B(n_306), .Y(n_439) );
INVx4_ASAP7_75t_L g330 ( .A(n_282), .Y(n_330) );
INVx1_ASAP7_75t_L g288 ( .A(n_283), .Y(n_288) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
AND2x4_ASAP7_75t_L g399 ( .A(n_287), .B(n_354), .Y(n_399) );
INVx1_ASAP7_75t_SL g438 ( .A(n_287), .Y(n_438) );
AND2x2_ASAP7_75t_L g443 ( .A(n_287), .B(n_346), .Y(n_443) );
INVx1_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
INVx1_ASAP7_75t_L g385 ( .A(n_291), .Y(n_385) );
OAI21xp5_ASAP7_75t_SL g292 ( .A1(n_293), .A2(n_295), .B(n_297), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OR2x2_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
INVx1_ASAP7_75t_L g318 ( .A(n_299), .Y(n_318) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x2_ASAP7_75t_L g315 ( .A(n_301), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g405 ( .A(n_301), .B(n_406), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g302 ( .A1(n_303), .A2(n_307), .B(n_309), .C(n_326), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g398 ( .A(n_305), .B(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g322 ( .A(n_306), .B(n_321), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_306), .B(n_416), .Y(n_415) );
AND2x2_ASAP7_75t_L g431 ( .A(n_306), .B(n_354), .Y(n_431) );
OAI221xp5_ASAP7_75t_SL g342 ( .A1(n_307), .A2(n_331), .B1(n_343), .B2(n_344), .C(n_348), .Y(n_342) );
INVx3_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
AND2x2_ASAP7_75t_L g413 ( .A(n_308), .B(n_314), .Y(n_413) );
OAI32xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_315), .A3(n_317), .B1(n_319), .B2(n_323), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
INVx2_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVxp67_ASAP7_75t_SL g403 ( .A(n_313), .Y(n_403) );
INVx2_ASAP7_75t_L g336 ( .A(n_314), .Y(n_336) );
O2A1O1Ixp33_ASAP7_75t_L g445 ( .A1(n_314), .A2(n_366), .B(n_446), .C(n_447), .Y(n_445) );
INVx1_ASAP7_75t_L g351 ( .A(n_316), .Y(n_351) );
OR2x2_ASAP7_75t_L g447 ( .A(n_316), .B(n_448), .Y(n_447) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_320), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx1_ASAP7_75t_L g408 ( .A(n_323), .Y(n_408) );
AND2x2_ASAP7_75t_L g323 ( .A(n_324), .B(n_325), .Y(n_323) );
INVx1_ASAP7_75t_L g389 ( .A(n_324), .Y(n_389) );
OAI21xp33_ASAP7_75t_SL g326 ( .A1(n_327), .A2(n_335), .B(n_339), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
OR2x2_ASAP7_75t_L g328 ( .A(n_329), .B(n_331), .Y(n_328) );
OR2x2_ASAP7_75t_L g366 ( .A(n_329), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_330), .B(n_333), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
AOI221xp5_ASAP7_75t_L g432 ( .A1(n_332), .A2(n_364), .B1(n_433), .B2(n_436), .C(n_440), .Y(n_432) );
INVx2_ASAP7_75t_L g435 ( .A(n_332), .Y(n_435) );
INVx2_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
OR2x2_ASAP7_75t_L g356 ( .A(n_336), .B(n_357), .Y(n_356) );
AND2x4_ASAP7_75t_L g423 ( .A(n_336), .B(n_381), .Y(n_423) );
INVx2_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
INVxp67_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_347), .Y(n_345) );
INVx1_ASAP7_75t_L g421 ( .A(n_346), .Y(n_421) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_351), .B(n_352), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_354), .B(n_384), .Y(n_441) );
INVx2_ASAP7_75t_L g448 ( .A(n_354), .Y(n_448) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g418 ( .A1(n_356), .A2(n_419), .B1(n_422), .B2(n_424), .C(n_426), .Y(n_418) );
AND5x1_ASAP7_75t_L g358 ( .A(n_359), .B(n_397), .C(n_412), .D(n_432), .E(n_442), .Y(n_358) );
NOR2xp33_ASAP7_75t_SL g359 ( .A(n_360), .B(n_377), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_361), .A2(n_366), .B1(n_369), .B2(n_371), .C(n_372), .Y(n_360) );
NAND2xp5_ASAP7_75t_SL g361 ( .A(n_362), .B(n_364), .Y(n_361) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_373), .B(n_375), .Y(n_372) );
INVx2_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
OAI221xp5_ASAP7_75t_SL g377 ( .A1(n_378), .A2(n_382), .B1(n_383), .B2(n_385), .C(n_386), .Y(n_377) );
INVx1_ASAP7_75t_SL g378 ( .A(n_379), .Y(n_378) );
AND2x4_ASAP7_75t_L g379 ( .A(n_380), .B(n_381), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g420 ( .A(n_382), .B(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_SL g387 ( .A(n_388), .Y(n_387) );
OR2x2_ASAP7_75t_L g388 ( .A(n_389), .B(n_390), .Y(n_388) );
OR2x2_ASAP7_75t_L g395 ( .A(n_390), .B(n_396), .Y(n_395) );
CKINVDCx16_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
INVx2_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
AOI21xp33_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_403), .B(n_404), .Y(n_400) );
INVx1_ASAP7_75t_SL g401 ( .A(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_413), .A2(n_414), .B(n_418), .Y(n_412) );
INVx1_ASAP7_75t_SL g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_SL g416 ( .A(n_417), .Y(n_416) );
INVxp67_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
INVxp67_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
AOI22xp5_ASAP7_75t_L g426 ( .A1(n_427), .A2(n_428), .B1(n_429), .B2(n_431), .Y(n_426) );
O2A1O1Ixp33_ASAP7_75t_L g442 ( .A1(n_428), .A2(n_443), .B(n_444), .C(n_445), .Y(n_442) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx1_ASAP7_75t_L g446 ( .A(n_439), .Y(n_446) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_SL g789 ( .A(n_449), .Y(n_789) );
CKINVDCx11_ASAP7_75t_R g449 ( .A(n_450), .Y(n_449) );
OAI22x1_ASAP7_75t_L g788 ( .A1(n_451), .A2(n_789), .B1(n_790), .B2(n_791), .Y(n_788) );
INVx1_ASAP7_75t_SL g451 ( .A(n_452), .Y(n_451) );
AND3x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_673), .C(n_736), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_637), .Y(n_454) );
NOR3xp33_ASAP7_75t_L g455 ( .A(n_456), .B(n_578), .C(n_607), .Y(n_455) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_457), .B(n_567), .Y(n_456) );
AOI22xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_487), .B1(n_527), .B2(n_539), .Y(n_457) );
NAND2x1_ASAP7_75t_L g722 ( .A(n_458), .B(n_568), .Y(n_722) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_479), .Y(n_459) );
INVx2_ASAP7_75t_L g541 ( .A(n_460), .Y(n_541) );
INVx4_ASAP7_75t_L g583 ( .A(n_460), .Y(n_583) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_460), .Y(n_603) );
AND2x4_ASAP7_75t_L g614 ( .A(n_460), .B(n_582), .Y(n_614) );
AND2x2_ASAP7_75t_L g620 ( .A(n_460), .B(n_544), .Y(n_620) );
NOR2x1_ASAP7_75t_SL g750 ( .A(n_460), .B(n_555), .Y(n_750) );
OR2x6_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_L g503 ( .A(n_464), .Y(n_503) );
NOR2x1p5_ASAP7_75t_L g465 ( .A(n_466), .B(n_467), .Y(n_465) );
INVx1_ASAP7_75t_L g524 ( .A(n_467), .Y(n_524) );
INVx3_ASAP7_75t_L g467 ( .A(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g471 ( .A(n_468), .B(n_472), .Y(n_471) );
INVxp67_ASAP7_75t_L g493 ( .A(n_471), .Y(n_493) );
INVx2_ASAP7_75t_L g554 ( .A(n_471), .Y(n_554) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_471), .A2(n_496), .B1(n_559), .B2(n_560), .Y(n_558) );
AND2x2_ASAP7_75t_L g476 ( .A(n_472), .B(n_477), .Y(n_476) );
INVxp33_ASAP7_75t_L g523 ( .A(n_472), .Y(n_523) );
INVx1_ASAP7_75t_L g505 ( .A(n_475), .Y(n_505) );
AND2x4_ASAP7_75t_L g475 ( .A(n_476), .B(n_478), .Y(n_475) );
INVx1_ASAP7_75t_L g547 ( .A(n_476), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_478), .Y(n_548) );
INVx2_ASAP7_75t_L g586 ( .A(n_479), .Y(n_586) );
HB1xp67_ASAP7_75t_L g600 ( .A(n_479), .Y(n_600) );
INVx1_ASAP7_75t_L g611 ( .A(n_479), .Y(n_611) );
HB1xp67_ASAP7_75t_L g623 ( .A(n_479), .Y(n_623) );
AND2x2_ASAP7_75t_L g655 ( .A(n_479), .B(n_555), .Y(n_655) );
AND2x2_ASAP7_75t_L g687 ( .A(n_479), .B(n_571), .Y(n_687) );
INVx1_ASAP7_75t_L g694 ( .A(n_479), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g480 ( .A(n_481), .B(n_482), .Y(n_480) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_506), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
AND2x2_ASAP7_75t_L g636 ( .A(n_489), .B(n_575), .Y(n_636) );
INVx2_ASAP7_75t_L g710 ( .A(n_489), .Y(n_710) );
AND2x2_ASAP7_75t_L g733 ( .A(n_489), .B(n_506), .Y(n_733) );
INVx1_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_490), .B(n_530), .Y(n_574) );
INVx2_ASAP7_75t_L g595 ( .A(n_490), .Y(n_595) );
AND2x4_ASAP7_75t_L g617 ( .A(n_490), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g652 ( .A(n_490), .Y(n_652) );
AND2x2_ASAP7_75t_L g729 ( .A(n_490), .B(n_533), .Y(n_729) );
OR2x2_ASAP7_75t_L g490 ( .A(n_491), .B(n_499), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_495), .B(n_496), .Y(n_494) );
OAI22xp5_ASAP7_75t_L g499 ( .A1(n_500), .A2(n_503), .B1(n_504), .B2(n_505), .Y(n_499) );
INVx1_ASAP7_75t_L g501 ( .A(n_502), .Y(n_501) );
INVx1_ASAP7_75t_L g700 ( .A(n_506), .Y(n_700) );
AND2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_515), .Y(n_506) );
NOR2xp67_ASAP7_75t_L g625 ( .A(n_507), .B(n_595), .Y(n_625) );
AND2x2_ASAP7_75t_L g630 ( .A(n_507), .B(n_595), .Y(n_630) );
INVx2_ASAP7_75t_L g643 ( .A(n_507), .Y(n_643) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_507), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_510), .Y(n_508) );
AND2x4_ASAP7_75t_L g616 ( .A(n_515), .B(n_529), .Y(n_616) );
AND2x2_ASAP7_75t_L g631 ( .A(n_515), .B(n_632), .Y(n_631) );
INVx1_ASAP7_75t_L g684 ( .A(n_515), .Y(n_684) );
INVx2_ASAP7_75t_L g515 ( .A(n_516), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_516), .B(n_533), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g688 ( .A(n_516), .B(n_530), .Y(n_688) );
AO21x2_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_518), .B(n_526), .Y(n_516) );
AO21x2_ASAP7_75t_L g577 ( .A1(n_517), .A2(n_518), .B(n_526), .Y(n_577) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_519), .B(n_525), .Y(n_518) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
INVxp33_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
NAND2x1p5_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx3_ASAP7_75t_L g592 ( .A(n_529), .Y(n_592) );
INVx3_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
HB1xp67_ASAP7_75t_L g590 ( .A(n_530), .Y(n_590) );
AND2x2_ASAP7_75t_L g759 ( .A(n_530), .B(n_760), .Y(n_759) );
INVx3_ASAP7_75t_L g647 ( .A(n_531), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g779 ( .A(n_531), .B(n_684), .Y(n_779) );
BUFx3_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g594 ( .A(n_532), .B(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
AND2x4_ASAP7_75t_L g575 ( .A(n_533), .B(n_576), .Y(n_575) );
INVx2_ASAP7_75t_L g618 ( .A(n_533), .Y(n_618) );
INVxp67_ASAP7_75t_L g632 ( .A(n_533), .Y(n_632) );
INVx1_ASAP7_75t_L g692 ( .A(n_533), .Y(n_692) );
HB1xp67_ASAP7_75t_L g760 ( .A(n_533), .Y(n_760) );
INVx1_ASAP7_75t_L g744 ( .A(n_539), .Y(n_744) );
NOR2x1_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
NOR2x1_ASAP7_75t_L g664 ( .A(n_540), .B(n_665), .Y(n_664) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g698 ( .A(n_541), .B(n_570), .Y(n_698) );
OR2x2_ASAP7_75t_L g734 ( .A(n_542), .B(n_735), .Y(n_734) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g716 ( .A(n_543), .B(n_694), .Y(n_716) );
AND2x2_ASAP7_75t_L g768 ( .A(n_543), .B(n_603), .Y(n_768) );
AND2x2_ASAP7_75t_L g543 ( .A(n_544), .B(n_555), .Y(n_543) );
AND2x4_ASAP7_75t_L g570 ( .A(n_544), .B(n_571), .Y(n_570) );
INVx1_ASAP7_75t_L g582 ( .A(n_544), .Y(n_582) );
INVx2_ASAP7_75t_L g599 ( .A(n_544), .Y(n_599) );
HB1xp67_ASAP7_75t_L g777 ( .A(n_544), .Y(n_777) );
AND2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_550), .Y(n_544) );
NOR3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_548), .C(n_549), .Y(n_546) );
INVx3_ASAP7_75t_L g571 ( .A(n_555), .Y(n_571) );
INVx2_ASAP7_75t_L g665 ( .A(n_555), .Y(n_665) );
AND2x4_ASAP7_75t_L g555 ( .A(n_556), .B(n_557), .Y(n_555) );
OAI21xp5_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B(n_566), .Y(n_557) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_563), .B1(n_564), .B2(n_565), .Y(n_561) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_572), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g662 ( .A(n_569), .B(n_645), .Y(n_662) );
NOR2x1_ASAP7_75t_L g704 ( .A(n_569), .B(n_583), .Y(n_704) );
INVx4_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_570), .B(n_645), .Y(n_782) );
AND2x2_ASAP7_75t_L g598 ( .A(n_571), .B(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g612 ( .A(n_571), .Y(n_612) );
AOI22xp5_ASAP7_75t_SL g660 ( .A1(n_572), .A2(n_661), .B1(n_662), .B2(n_663), .Y(n_660) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_575), .Y(n_572) );
NAND2x1p5_ASAP7_75t_L g657 ( .A(n_573), .B(n_631), .Y(n_657) );
INVx2_ASAP7_75t_SL g573 ( .A(n_574), .Y(n_573) );
OR2x2_ASAP7_75t_L g718 ( .A(n_574), .B(n_606), .Y(n_718) );
AND2x2_ASAP7_75t_L g588 ( .A(n_575), .B(n_589), .Y(n_588) );
AND2x4_ASAP7_75t_L g624 ( .A(n_575), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g720 ( .A(n_575), .B(n_710), .Y(n_720) );
INVx2_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
AND2x4_ASAP7_75t_L g642 ( .A(n_577), .B(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g668 ( .A(n_577), .Y(n_668) );
AND2x2_ASAP7_75t_L g758 ( .A(n_577), .B(n_595), .Y(n_758) );
OAI221xp5_ASAP7_75t_L g578 ( .A1(n_579), .A2(n_587), .B1(n_591), .B2(n_596), .C(n_601), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_581), .B(n_584), .Y(n_580) );
INVx1_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_581), .B(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g774 ( .A(n_581), .B(n_655), .Y(n_774) );
AND2x4_ASAP7_75t_L g581 ( .A(n_582), .B(n_583), .Y(n_581) );
NOR2xp67_ASAP7_75t_SL g627 ( .A(n_583), .B(n_628), .Y(n_627) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_583), .Y(n_640) );
OR2x2_ASAP7_75t_L g724 ( .A(n_583), .B(n_725), .Y(n_724) );
AND2x4_ASAP7_75t_SL g776 ( .A(n_583), .B(n_777), .Y(n_776) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx3_ASAP7_75t_L g645 ( .A(n_585), .Y(n_645) );
INVx2_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_586), .Y(n_735) );
INVx1_ASAP7_75t_L g587 ( .A(n_588), .Y(n_587) );
AOI221x1_ASAP7_75t_L g675 ( .A1(n_588), .A2(n_676), .B1(n_678), .B2(n_681), .C(n_685), .Y(n_675) );
AND2x2_ASAP7_75t_L g661 ( .A(n_589), .B(n_617), .Y(n_661) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OR2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_593), .Y(n_591) );
AND2x2_ASAP7_75t_L g604 ( .A(n_592), .B(n_605), .Y(n_604) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_592), .B(n_594), .Y(n_731) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_600), .Y(n_597) );
AND2x2_ASAP7_75t_SL g602 ( .A(n_598), .B(n_603), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_598), .B(n_611), .Y(n_628) );
INVx2_ASAP7_75t_L g635 ( .A(n_598), .Y(n_635) );
INVx1_ASAP7_75t_L g680 ( .A(n_599), .Y(n_680) );
BUFx2_ASAP7_75t_L g769 ( .A(n_600), .Y(n_769) );
NAND2xp33_ASAP7_75t_SL g601 ( .A(n_602), .B(n_604), .Y(n_601) );
OR2x6_ASAP7_75t_L g634 ( .A(n_603), .B(n_635), .Y(n_634) );
AND2x2_ASAP7_75t_L g715 ( .A(n_603), .B(n_655), .Y(n_715) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_608), .B(n_626), .Y(n_607) );
AOI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_615), .B1(n_619), .B2(n_624), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_610), .B(n_613), .Y(n_609) );
AND2x2_ASAP7_75t_SL g672 ( .A(n_610), .B(n_614), .Y(n_672) );
AND2x4_ASAP7_75t_L g678 ( .A(n_610), .B(n_679), .Y(n_678) );
AND2x4_ASAP7_75t_SL g610 ( .A(n_611), .B(n_612), .Y(n_610) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_611), .Y(n_703) );
INVx2_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_614), .B(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_614), .B(n_645), .Y(n_677) );
HB1xp67_ASAP7_75t_L g761 ( .A(n_614), .Y(n_761) );
AND2x2_ASAP7_75t_L g615 ( .A(n_616), .B(n_617), .Y(n_615) );
AND2x2_ASAP7_75t_L g708 ( .A(n_616), .B(n_709), .Y(n_708) );
INVx3_ASAP7_75t_L g669 ( .A(n_617), .Y(n_669) );
NAND2x1_ASAP7_75t_SL g713 ( .A(n_617), .B(n_668), .Y(n_713) );
AND2x2_ASAP7_75t_L g747 ( .A(n_617), .B(n_642), .Y(n_747) );
AND2x2_ASAP7_75t_L g619 ( .A(n_620), .B(n_621), .Y(n_619) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_627), .A2(n_629), .B1(n_633), .B2(n_636), .Y(n_626) );
BUFx2_ASAP7_75t_L g742 ( .A(n_628), .Y(n_742) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_629), .A2(n_698), .B1(n_772), .B2(n_781), .Y(n_780) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
NAND2x1p5_ASAP7_75t_L g683 ( .A(n_630), .B(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g650 ( .A(n_631), .B(n_651), .Y(n_650) );
INVx2_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
NAND3xp33_ASAP7_75t_L g766 ( .A(n_635), .B(n_767), .C(n_769), .Y(n_766) );
INVx1_ASAP7_75t_L g670 ( .A(n_636), .Y(n_670) );
AOI211x1_ASAP7_75t_L g637 ( .A1(n_638), .A2(n_646), .B(n_648), .C(n_666), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_640), .B(n_641), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g697 ( .A(n_641), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .Y(n_641) );
AND2x2_ASAP7_75t_L g728 ( .A(n_642), .B(n_729), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_642), .B(n_709), .Y(n_740) );
AND2x2_ASAP7_75t_L g772 ( .A(n_642), .B(n_710), .Y(n_772) );
INVx1_ASAP7_75t_L g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g753 ( .A(n_645), .Y(n_753) );
INVx1_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
OR2x2_ASAP7_75t_L g682 ( .A(n_647), .B(n_683), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_649), .B(n_660), .Y(n_648) );
AOI22xp5_ASAP7_75t_SL g649 ( .A1(n_650), .A2(n_653), .B1(n_656), .B2(n_658), .Y(n_649) );
BUFx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
AND2x2_ASAP7_75t_L g690 ( .A(n_652), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g705 ( .A(n_652), .Y(n_705) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
AND2x2_ASAP7_75t_SL g775 ( .A(n_655), .B(n_776), .Y(n_775) );
INVx3_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
INVxp67_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
HB1xp67_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
AND2x2_ASAP7_75t_L g711 ( .A(n_664), .B(n_694), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g666 ( .A1(n_667), .A2(n_670), .B(n_671), .Y(n_666) );
OR2x2_ASAP7_75t_L g667 ( .A(n_668), .B(n_669), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_668), .B(n_690), .Y(n_765) );
OR2x2_ASAP7_75t_L g743 ( .A(n_669), .B(n_688), .Y(n_743) );
INVx1_ASAP7_75t_SL g671 ( .A(n_672), .Y(n_671) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
NAND3x1_ASAP7_75t_L g674 ( .A(n_675), .B(n_695), .C(n_719), .Y(n_674) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_678), .A2(n_708), .B1(n_711), .B2(n_712), .Y(n_707) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_679), .B(n_694), .Y(n_693) );
INVx2_ASAP7_75t_SL g752 ( .A(n_679), .Y(n_752) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_679), .B(n_753), .Y(n_756) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
OAI222xp33_ASAP7_75t_L g739 ( .A1(n_683), .A2(n_740), .B1(n_741), .B2(n_742), .C1(n_743), .C2(n_744), .Y(n_739) );
OAI22xp5_ASAP7_75t_L g685 ( .A1(n_686), .A2(n_688), .B1(n_689), .B2(n_693), .Y(n_685) );
INVx1_ASAP7_75t_SL g725 ( .A(n_687), .Y(n_725) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
AND2x2_ASAP7_75t_L g762 ( .A(n_691), .B(n_758), .Y(n_762) );
NOR2x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_706), .Y(n_695) );
AOI21xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_699), .B(n_705), .Y(n_696) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_704), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_714), .Y(n_706) );
INVx1_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_713), .B(n_727), .Y(n_726) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_715), .A2(n_716), .B(n_717), .Y(n_714) );
INVx1_ASAP7_75t_L g741 ( .A(n_716), .Y(n_741) );
INVx1_ASAP7_75t_SL g717 ( .A(n_718), .Y(n_717) );
AOI221xp5_ASAP7_75t_L g719 ( .A1(n_720), .A2(n_721), .B1(n_723), .B2(n_726), .C(n_730), .Y(n_719) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
INVxp67_ASAP7_75t_L g723 ( .A(n_724), .Y(n_723) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g730 ( .A1(n_731), .A2(n_732), .B(n_734), .Y(n_730) );
INVx1_ASAP7_75t_L g732 ( .A(n_733), .Y(n_732) );
INVxp67_ASAP7_75t_SL g736 ( .A(n_737), .Y(n_736) );
NAND3x1_ASAP7_75t_L g737 ( .A(n_738), .B(n_763), .C(n_770), .Y(n_737) );
NOR2x1_ASAP7_75t_L g738 ( .A(n_739), .B(n_745), .Y(n_738) );
NAND2xp5_ASAP7_75t_L g745 ( .A(n_746), .B(n_754), .Y(n_745) );
NAND2xp5_ASAP7_75t_SL g746 ( .A(n_747), .B(n_748), .Y(n_746) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_751), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_749), .B(n_756), .Y(n_755) );
INVx1_ASAP7_75t_L g749 ( .A(n_750), .Y(n_749) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_753), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_757), .B1(n_761), .B2(n_762), .Y(n_754) );
AND2x4_ASAP7_75t_L g757 ( .A(n_758), .B(n_759), .Y(n_757) );
NAND2xp5_ASAP7_75t_SL g763 ( .A(n_764), .B(n_766), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g770 ( .A(n_771), .B(n_780), .Y(n_770) );
AOI22xp5_ASAP7_75t_SL g771 ( .A1(n_772), .A2(n_773), .B1(n_775), .B2(n_778), .Y(n_771) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
INVxp67_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g786 ( .A(n_783), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
INVx1_ASAP7_75t_L g803 ( .A(n_790), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_797), .Y(n_794) );
CKINVDCx5p33_ASAP7_75t_R g795 ( .A(n_796), .Y(n_795) );
OAI22xp5_ASAP7_75t_SL g798 ( .A1(n_799), .A2(n_800), .B1(n_803), .B2(n_804), .Y(n_798) );
INVx1_ASAP7_75t_L g804 ( .A(n_800), .Y(n_804) );
INVx1_ASAP7_75t_SL g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_SL g806 ( .A(n_807), .Y(n_806) );
NOR2xp33_ASAP7_75t_L g808 ( .A(n_809), .B(n_810), .Y(n_808) );
HB1xp67_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
endmodule