module real_jpeg_14735_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;

BUFx2_ASAP7_75t_L g87 ( 
.A(n_0),
.Y(n_87)
);

BUFx4f_ASAP7_75t_L g52 ( 
.A(n_1),
.Y(n_52)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_2),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_3),
.A2(n_63),
.B1(n_64),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_3),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_3),
.A2(n_28),
.B1(n_30),
.B2(n_130),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_36),
.B1(n_38),
.B2(n_130),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g226 ( 
.A1(n_3),
.A2(n_48),
.B1(n_53),
.B2(n_130),
.Y(n_226)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_4),
.Y(n_37)
);

INVx11_ASAP7_75t_L g50 ( 
.A(n_5),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_6),
.A2(n_28),
.B1(n_30),
.B2(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_6),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_6),
.A2(n_36),
.B1(n_38),
.B2(n_136),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_6),
.A2(n_48),
.B1(n_53),
.B2(n_136),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_6),
.A2(n_63),
.B1(n_64),
.B2(n_136),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_L g42 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_43),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_7),
.A2(n_43),
.B1(n_63),
.B2(n_64),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_7),
.A2(n_36),
.B1(n_38),
.B2(n_43),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_7),
.A2(n_43),
.B1(n_48),
.B2(n_53),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_9),
.A2(n_63),
.B1(n_64),
.B2(n_67),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_9),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_9),
.A2(n_28),
.B1(n_30),
.B2(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_9),
.A2(n_48),
.B1(n_53),
.B2(n_67),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g177 ( 
.A1(n_9),
.A2(n_36),
.B1(n_38),
.B2(n_67),
.Y(n_177)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_10),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_11),
.A2(n_63),
.B1(n_64),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_11),
.Y(n_128)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_11),
.A2(n_60),
.B(n_63),
.C(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_11),
.B(n_102),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_11),
.A2(n_36),
.B1(n_38),
.B2(n_128),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_11),
.A2(n_85),
.B1(n_88),
.B2(n_226),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_11),
.B(n_82),
.Y(n_239)
);

BUFx8_ASAP7_75t_L g60 ( 
.A(n_12),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_13),
.A2(n_28),
.B1(n_30),
.B2(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_13),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_13),
.A2(n_63),
.B1(n_64),
.B2(n_134),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_13),
.A2(n_36),
.B1(n_38),
.B2(n_134),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_L g218 ( 
.A1(n_13),
.A2(n_48),
.B1(n_53),
.B2(n_134),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_14),
.A2(n_36),
.B1(n_38),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_14),
.A2(n_48),
.B1(n_53),
.B2(n_57),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_14),
.A2(n_57),
.B1(n_63),
.B2(n_64),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_14),
.A2(n_28),
.B1(n_30),
.B2(n_57),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_15),
.A2(n_28),
.B1(n_29),
.B2(n_30),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_15),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_15),
.A2(n_29),
.B1(n_36),
.B2(n_38),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_15),
.A2(n_29),
.B1(n_63),
.B2(n_64),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_15),
.A2(n_29),
.B1(n_48),
.B2(n_53),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_119),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_118),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_103),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_20),
.B(n_103),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_73),
.C(n_83),
.Y(n_20)
);

FAx1_ASAP7_75t_SL g305 ( 
.A(n_21),
.B(n_73),
.CI(n_83),
.CON(n_305),
.SN(n_305)
);

OAI22xp5_ASAP7_75t_SL g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_72),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_24),
.B(n_45),
.C(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_31),
.B(n_40),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_27),
.A2(n_32),
.B1(n_80),
.B2(n_82),
.Y(n_79)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_28),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g39 ( 
.A1(n_28),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_28),
.A2(n_30),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g189 ( 
.A(n_28),
.B(n_128),
.CON(n_189),
.SN(n_189)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_30),
.A2(n_61),
.B(n_128),
.Y(n_144)
);

NOR3xp33_ASAP7_75t_L g190 ( 
.A(n_30),
.B(n_35),
.C(n_36),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_31),
.A2(n_33),
.B1(n_155),
.B2(n_157),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_31),
.A2(n_112),
.B(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_32),
.B(n_115),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_32),
.A2(n_82),
.B1(n_133),
.B2(n_135),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_32),
.A2(n_82),
.B1(n_156),
.B2(n_189),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g267 ( 
.A1(n_32),
.A2(n_41),
.B(n_113),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_39),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_33),
.B(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_33),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_33),
.A2(n_81),
.B(n_114),
.Y(n_283)
);

OA22x2_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_36),
.B2(n_38),
.Y(n_33)
);

O2A1O1Ixp33_ASAP7_75t_SL g187 ( 
.A1(n_34),
.A2(n_38),
.B(n_188),
.C(n_190),
.Y(n_187)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g38 ( 
.A(n_36),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_36),
.A2(n_38),
.B1(n_51),
.B2(n_52),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_38),
.B(n_210),
.Y(n_209)
);

INVxp33_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_42),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_44),
.A2(n_45),
.B1(n_111),
.B2(n_116),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_54),
.B(n_56),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_46),
.B(n_56),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_46),
.A2(n_54),
.B1(n_195),
.B2(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_46),
.A2(n_54),
.B1(n_212),
.B2(n_213),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_46),
.A2(n_54),
.B1(n_203),
.B2(n_213),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_46),
.A2(n_54),
.B1(n_94),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_47),
.B(n_55),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_47),
.B(n_78),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_47),
.A2(n_76),
.B(n_177),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_47),
.B(n_128),
.Y(n_229)
);

OA22x2_ASAP7_75t_L g47 ( 
.A1(n_48),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_47)
);

CKINVDCx6p67_ASAP7_75t_R g53 ( 
.A(n_48),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_51),
.B(n_53),
.C(n_128),
.Y(n_210)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_53),
.B(n_87),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_53),
.B(n_224),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_54),
.B(n_77),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_54),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_54),
.A2(n_56),
.B(n_95),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_54),
.Y(n_193)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_58),
.A2(n_72),
.B1(n_106),
.B2(n_117),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_62),
.B(n_68),
.Y(n_58)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_59),
.B(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_59),
.A2(n_98),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx11_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_61),
.B1(n_63),
.B2(n_64),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_62),
.Y(n_108)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_71),
.Y(n_68)
);

CKINVDCx14_ASAP7_75t_R g98 ( 
.A(n_69),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_69),
.A2(n_102),
.B1(n_108),
.B2(n_109),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_69),
.A2(n_102),
.B1(n_127),
.B2(n_129),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_69),
.A2(n_102),
.B1(n_166),
.B2(n_269),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_71),
.B(n_102),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_73),
.A2(n_74),
.B(n_79),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_76),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_75),
.A2(n_193),
.B(n_194),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_82),
.B(n_113),
.Y(n_112)
);

AOI21xp33_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_91),
.B(n_96),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_84),
.B(n_92),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g276 ( 
.A1(n_84),
.A2(n_92),
.B1(n_93),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_84),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_84),
.A2(n_96),
.B1(n_97),
.B2(n_277),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_88),
.B(n_89),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_85),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_85),
.A2(n_88),
.B1(n_218),
.B2(n_226),
.Y(n_228)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_85),
.A2(n_220),
.B(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_86),
.A2(n_87),
.B1(n_140),
.B2(n_142),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_86),
.B(n_150),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_86),
.A2(n_90),
.B(n_175),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_86),
.A2(n_87),
.B1(n_217),
.B2(n_219),
.Y(n_216)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_87),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_87),
.B(n_90),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_88),
.A2(n_141),
.B(n_149),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_88),
.B(n_151),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_88),
.B(n_128),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_91),
.B(n_298),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_101),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g284 ( 
.A1(n_98),
.A2(n_285),
.B(n_286),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_100),
.B(n_102),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_106),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_110),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_111),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_114),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_302),
.B(n_306),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_291),
.B(n_301),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g121 ( 
.A1(n_122),
.A2(n_272),
.B(n_290),
.Y(n_121)
);

O2A1O1Ixp33_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_179),
.B(n_254),
.C(n_271),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_158),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g180 ( 
.A(n_124),
.B(n_158),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_138),
.C(n_147),
.Y(n_124)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_125),
.B(n_251),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_126),
.B(n_132),
.C(n_137),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_129),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_137),
.Y(n_131)
);

CKINVDCx14_ASAP7_75t_R g157 ( 
.A(n_133),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_135),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_138),
.B(n_147),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_138)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_139),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_142),
.Y(n_173)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_143),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_145),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_152),
.C(n_154),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_148),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g260 ( 
.A(n_149),
.B(n_236),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_SL g196 ( 
.A(n_154),
.B(n_197),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_170),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_159),
.B(n_171),
.C(n_178),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g159 ( 
.A1(n_160),
.A2(n_161),
.B1(n_162),
.B2(n_169),
.Y(n_159)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_160),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_163),
.B(n_167),
.C(n_169),
.Y(n_256)
);

CKINVDCx14_ASAP7_75t_R g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_178),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_172),
.B(n_176),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_177),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_249),
.B(n_253),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_204),
.B(n_248),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_199),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_184),
.B(n_199),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_196),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_192),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_186),
.B(n_192),
.C(n_196),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_187),
.B(n_191),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_SL g200 ( 
.A(n_187),
.B(n_191),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_201),
.C(n_202),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g244 ( 
.A(n_200),
.B(n_245),
.Y(n_244)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_202),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_243),
.B(n_247),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_232),
.B(n_242),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_221),
.B(n_231),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_216),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_208),
.B(n_216),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_209),
.A2(n_211),
.B1(n_214),
.B2(n_215),
.Y(n_208)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_211),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_211),
.B(n_214),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_220),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_227),
.B(n_230),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_225),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_228),
.B(n_229),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_234),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_233),
.B(n_234),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_235),
.B(n_237),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_235),
.B(n_238),
.C(n_241),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_240),
.B2(n_241),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_240),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_244),
.B(n_246),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_246),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_250),
.B(n_252),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_255),
.B(n_270),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_255),
.B(n_270),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_257),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_256),
.B(n_258),
.C(n_264),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_264),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_259),
.A2(n_260),
.B1(n_261),
.B2(n_263),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_259),
.B(n_263),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_260),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_261),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_267),
.C(n_268),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g285 ( 
.A(n_269),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_274),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_273),
.B(n_274),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_289),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_278),
.B1(n_287),
.B2(n_288),
.Y(n_275)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_276),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_276),
.B(n_288),
.C(n_289),
.Y(n_300)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_278),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_279),
.B(n_283),
.C(n_284),
.Y(n_294)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_300),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_292),
.B(n_300),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_295),
.B2(n_299),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_293),
.B(n_296),
.C(n_297),
.Y(n_304)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_294),
.Y(n_293)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_295),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_304),
.B(n_305),
.Y(n_307)
);

BUFx24_ASAP7_75t_SL g309 ( 
.A(n_305),
.Y(n_309)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);


endmodule