module fake_jpeg_20850_n_277 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_277);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_277;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_96;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_13),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_5),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_25),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_36),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_L g41 ( 
.A1(n_37),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_41)
);

AO22x1_ASAP7_75t_SL g61 ( 
.A1(n_41),
.A2(n_51),
.B1(n_36),
.B2(n_40),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_36),
.A2(n_32),
.B1(n_18),
.B2(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_43),
.A2(n_52),
.B1(n_35),
.B2(n_16),
.Y(n_81)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_45),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_46),
.B(n_39),
.Y(n_70)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_35),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_35),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_37),
.A2(n_18),
.B1(n_32),
.B2(n_17),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_36),
.A2(n_32),
.B1(n_17),
.B2(n_16),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_16),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_54),
.B(n_57),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_31),
.B1(n_25),
.B2(n_29),
.Y(n_55)
);

AOI222xp33_ASAP7_75t_L g60 ( 
.A1(n_55),
.A2(n_56),
.B1(n_39),
.B2(n_33),
.C1(n_30),
.C2(n_19),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_38),
.A2(n_31),
.B1(n_30),
.B2(n_29),
.Y(n_56)
);

A2O1A1Ixp33_ASAP7_75t_L g57 ( 
.A1(n_38),
.A2(n_31),
.B(n_24),
.C(n_26),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_60),
.A2(n_69),
.B1(n_70),
.B2(n_80),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_61),
.A2(n_47),
.B1(n_48),
.B2(n_45),
.Y(n_98)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVxp67_ASAP7_75t_L g63 ( 
.A(n_44),
.Y(n_63)
);

INVx13_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx13_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_64),
.B(n_66),
.Y(n_93)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_65),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_54),
.Y(n_66)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_68),
.B(n_69),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_53),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_70),
.B(n_72),
.Y(n_95)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_58),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_71),
.B(n_74),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_34),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_44),
.B(n_36),
.Y(n_73)
);

OAI32xp33_ASAP7_75t_L g113 ( 
.A1(n_73),
.A2(n_77),
.A3(n_79),
.B1(n_40),
.B2(n_34),
.Y(n_113)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_42),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_24),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_75),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_40),
.Y(n_77)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_78),
.A2(n_82),
.B1(n_83),
.B2(n_40),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_57),
.B(n_40),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_57),
.B(n_38),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_80),
.A2(n_85),
.B(n_49),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_81),
.A2(n_35),
.B1(n_21),
.B2(n_27),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_43),
.A2(n_30),
.B1(n_29),
.B2(n_19),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_47),
.A2(n_27),
.B1(n_19),
.B2(n_21),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_41),
.B(n_24),
.Y(n_84)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_47),
.B(n_26),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_24),
.Y(n_87)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_88),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_73),
.B(n_26),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g137 ( 
.A1(n_89),
.A2(n_50),
.B(n_67),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_90),
.A2(n_107),
.B(n_50),
.Y(n_131)
);

MAJx2_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_52),
.C(n_35),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_85),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_98),
.A2(n_61),
.B1(n_86),
.B2(n_65),
.Y(n_121)
);

HB1xp67_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_100),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_102),
.A2(n_103),
.B1(n_99),
.B2(n_105),
.Y(n_135)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_27),
.B1(n_21),
.B2(n_34),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_104),
.A2(n_76),
.B1(n_77),
.B2(n_60),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_76),
.A2(n_24),
.B(n_26),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_59),
.Y(n_108)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_108),
.Y(n_117)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_59),
.Y(n_109)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_109),
.Y(n_128)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_72),
.Y(n_112)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_112),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_85),
.Y(n_125)
);

AND2x6_ASAP7_75t_L g114 ( 
.A(n_80),
.B(n_20),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_114),
.B(n_79),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_115),
.Y(n_116)
);

NOR3xp33_ASAP7_75t_SL g165 ( 
.A(n_118),
.B(n_23),
.C(n_22),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_119),
.A2(n_121),
.B1(n_122),
.B2(n_130),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_104),
.B(n_64),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_120),
.B(n_129),
.C(n_139),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_112),
.A2(n_61),
.B1(n_86),
.B2(n_71),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_105),
.B1(n_101),
.B2(n_113),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_123),
.A2(n_135),
.B1(n_28),
.B2(n_23),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_23),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_109),
.B1(n_108),
.B2(n_92),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_91),
.B(n_20),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_126),
.B(n_127),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g127 ( 
.A(n_97),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_95),
.B(n_26),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_114),
.A2(n_68),
.B1(n_78),
.B2(n_74),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_143),
.Y(n_161)
);

OR2x6_ASAP7_75t_L g132 ( 
.A(n_94),
.B(n_50),
.Y(n_132)
);

OA21x2_ASAP7_75t_L g172 ( 
.A1(n_132),
.A2(n_0),
.B(n_15),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_107),
.A2(n_0),
.B(n_28),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_133),
.A2(n_143),
.B(n_89),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_93),
.B(n_10),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_134),
.B(n_136),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_95),
.B(n_96),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_137),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g139 ( 
.A(n_90),
.B(n_23),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g140 ( 
.A(n_110),
.Y(n_140)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_140),
.Y(n_144)
);

CKINVDCx16_ASAP7_75t_R g141 ( 
.A(n_106),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_106),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_89),
.B(n_91),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_L g177 ( 
.A1(n_145),
.A2(n_161),
.B(n_170),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_146),
.B(n_147),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_117),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_149),
.B(n_153),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_125),
.A2(n_102),
.B1(n_92),
.B2(n_110),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_152),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_132),
.A2(n_111),
.B1(n_50),
.B2(n_28),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_128),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_142),
.Y(n_154)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_154),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_155),
.B(n_158),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_111),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_156),
.Y(n_190)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_142),
.Y(n_157)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_157),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_135),
.B(n_28),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_159),
.B(n_172),
.Y(n_191)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_122),
.Y(n_160)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_160),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_162),
.B(n_139),
.Y(n_183)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_140),
.Y(n_164)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_167),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_116),
.A2(n_8),
.B1(n_1),
.B2(n_2),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_0),
.B(n_1),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_116),
.A2(n_0),
.B(n_1),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_171),
.A2(n_137),
.B(n_127),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_160),
.A2(n_132),
.B1(n_131),
.B2(n_121),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_168),
.B(n_124),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_178),
.B(n_168),
.C(n_162),
.Y(n_200)
);

MAJx2_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_120),
.C(n_129),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_180),
.B(n_183),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_154),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_181),
.B(n_186),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_185),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_163),
.B(n_3),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g188 ( 
.A(n_161),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_188),
.B(n_172),
.Y(n_201)
);

AOI21xp33_ASAP7_75t_L g189 ( 
.A1(n_170),
.A2(n_3),
.B(n_4),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_189),
.A2(n_7),
.B(n_9),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_171),
.A2(n_4),
.B(n_5),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_192),
.A2(n_4),
.B(n_6),
.Y(n_209)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_144),
.Y(n_195)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_195),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_194),
.A2(n_166),
.B1(n_155),
.B2(n_172),
.Y(n_198)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_198),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_200),
.B(n_204),
.Y(n_221)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_201),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_178),
.B(n_147),
.C(n_150),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_203),
.C(n_207),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_166),
.C(n_167),
.Y(n_203)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_165),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_174),
.A2(n_152),
.B1(n_151),
.B2(n_157),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_206),
.A2(n_175),
.B1(n_174),
.B2(n_184),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_177),
.B(n_148),
.C(n_151),
.Y(n_207)
);

XOR2x2_ASAP7_75t_L g208 ( 
.A(n_180),
.B(n_164),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_208),
.B(n_213),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_211),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_190),
.B(n_144),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_210),
.B(n_186),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_177),
.B(n_15),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_176),
.Y(n_214)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_214),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_215),
.A2(n_194),
.B1(n_191),
.B2(n_192),
.Y(n_228)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_179),
.Y(n_216)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_216),
.Y(n_229)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_217),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_199),
.B(n_181),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_218),
.B(n_219),
.Y(n_233)
);

AO221x1_ASAP7_75t_L g219 ( 
.A1(n_204),
.A2(n_187),
.B1(n_193),
.B2(n_184),
.C(n_196),
.Y(n_219)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_205),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_232),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_225),
.A2(n_202),
.B1(n_197),
.B2(n_182),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_228),
.A2(n_213),
.B1(n_182),
.B2(n_185),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_200),
.B(n_173),
.C(n_179),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_231),
.B(n_222),
.C(n_227),
.Y(n_237)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_206),
.Y(n_232)
);

FAx1_ASAP7_75t_SL g234 ( 
.A(n_227),
.B(n_208),
.CI(n_212),
.CON(n_234),
.SN(n_234)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_234),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_226),
.B(n_211),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_235),
.B(n_236),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_237),
.B(n_242),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_187),
.Y(n_238)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_238),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_212),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_239),
.B(n_221),
.Y(n_247)
);

NAND2xp33_ASAP7_75t_L g240 ( 
.A(n_223),
.B(n_215),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_240),
.B(n_241),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_222),
.B(n_207),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_247),
.B(n_239),
.C(n_242),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g249 ( 
.A(n_233),
.Y(n_249)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_249),
.Y(n_255)
);

NAND2x1_ASAP7_75t_L g250 ( 
.A(n_234),
.B(n_231),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_250),
.B(n_237),
.Y(n_258)
);

NAND4xp25_ASAP7_75t_SL g251 ( 
.A(n_243),
.B(n_230),
.C(n_228),
.D(n_244),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_251),
.B(n_252),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_224),
.Y(n_252)
);

AOI21x1_ASAP7_75t_SL g256 ( 
.A1(n_245),
.A2(n_220),
.B(n_232),
.Y(n_256)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_256),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_258),
.B(n_262),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g259 ( 
.A1(n_254),
.A2(n_225),
.B1(n_203),
.B2(n_229),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_259),
.B(n_260),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_246),
.A2(n_196),
.B1(n_193),
.B2(n_209),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_SL g261 ( 
.A1(n_246),
.A2(n_252),
.B(n_248),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_234),
.Y(n_265)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_265),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_255),
.B(n_253),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g270 ( 
.A1(n_266),
.A2(n_268),
.A3(n_261),
.B1(n_262),
.B2(n_256),
.C1(n_14),
.C2(n_10),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_9),
.Y(n_268)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_263),
.A2(n_12),
.B(n_13),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_271),
.B(n_272),
.Y(n_274)
);

OAI21x1_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_14),
.B(n_15),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_273),
.B(n_269),
.C(n_267),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_275),
.A2(n_274),
.B(n_264),
.Y(n_276)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_276),
.B(n_14),
.Y(n_277)
);


endmodule