module fake_jpeg_5607_n_164 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_164);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_9),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_13),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g20 ( 
.A(n_4),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx1_ASAP7_75t_SL g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_5),
.Y(n_30)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_31),
.Y(n_70)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx5_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_36),
.B(n_37),
.Y(n_56)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_39),
.Y(n_64)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_14),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx6_ASAP7_75t_SL g42 ( 
.A(n_18),
.Y(n_42)
);

INVx1_ASAP7_75t_SL g61 ( 
.A(n_42),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_43),
.B(n_21),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_18),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_44),
.B(n_20),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_42),
.B(n_23),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_47),
.B(n_49),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_39),
.A2(n_20),
.B1(n_17),
.B2(n_22),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_50),
.A2(n_16),
.B1(n_12),
.B2(n_11),
.Y(n_89)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_41),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_57),
.Y(n_82)
);

OR2x2_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_30),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g93 ( 
.A(n_53),
.B(n_54),
.Y(n_93)
);

NOR2xp67_ASAP7_75t_L g54 ( 
.A(n_33),
.B(n_24),
.Y(n_54)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_36),
.B(n_22),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_33),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_58),
.B(n_72),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_31),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_60),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_38),
.B(n_28),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_34),
.B(n_28),
.C(n_27),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_62),
.B(n_30),
.C(n_17),
.Y(n_79)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_66),
.Y(n_87)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_0),
.Y(n_94)
);

OR2x4_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_24),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_69),
.A2(n_15),
.B(n_26),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_15),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_29),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_44),
.B(n_27),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_74),
.B(n_79),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_71),
.B1(n_69),
.B2(n_57),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_89),
.B1(n_93),
.B2(n_92),
.Y(n_108)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

OA22x2_ASAP7_75t_L g77 ( 
.A1(n_51),
.A2(n_50),
.B1(n_63),
.B2(n_68),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_81),
.B1(n_55),
.B2(n_66),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_29),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_61),
.Y(n_96)
);

OAI22x1_ASAP7_75t_SL g81 ( 
.A1(n_63),
.A2(n_20),
.B1(n_21),
.B2(n_24),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_3),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_62),
.B(n_26),
.Y(n_85)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g86 ( 
.A1(n_56),
.A2(n_16),
.B(n_1),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_86),
.A2(n_52),
.B(n_45),
.Y(n_97)
);

BUFx2_ASAP7_75t_L g88 ( 
.A(n_48),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_65),
.B(n_8),
.C(n_1),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_8),
.C(n_2),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_55),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_48),
.B1(n_70),
.B2(n_4),
.Y(n_100)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_94),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

INVx2_ASAP7_75t_SL g115 ( 
.A(n_95),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_109),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_97),
.A2(n_103),
.B(n_86),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_100),
.B1(n_89),
.B2(n_90),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_99),
.B(n_108),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_74),
.B(n_61),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_102),
.B(n_107),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_84),
.A2(n_70),
.B(n_46),
.Y(n_103)
);

AND2x6_ASAP7_75t_L g106 ( 
.A(n_77),
.B(n_45),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g121 ( 
.A(n_106),
.B(n_108),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_82),
.B(n_0),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_73),
.B(n_5),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_78),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_106),
.B(n_93),
.C(n_77),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_116),
.C(n_127),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_77),
.C(n_80),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_117),
.A2(n_109),
.B(n_101),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g119 ( 
.A(n_103),
.B(n_81),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_122),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_120),
.B(n_123),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g123 ( 
.A(n_110),
.B(n_80),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_112),
.B(n_79),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_125),
.B(n_126),
.Y(n_136)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_96),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_98),
.B(n_87),
.Y(n_127)
);

MAJx2_ASAP7_75t_L g128 ( 
.A(n_117),
.B(n_101),
.C(n_109),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_138),
.C(n_105),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_116),
.A2(n_113),
.B(n_121),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_129),
.A2(n_135),
.B(n_124),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_130),
.B(n_133),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_131),
.B(n_120),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_115),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_118),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_136),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_139),
.B(n_143),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_129),
.B(n_127),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_140),
.B(n_142),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_134),
.A2(n_119),
.B1(n_122),
.B2(n_114),
.Y(n_141)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_147),
.C(n_137),
.Y(n_148)
);

OAI31xp33_ASAP7_75t_L g146 ( 
.A1(n_128),
.A2(n_95),
.A3(n_83),
.B(n_105),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_146),
.A2(n_99),
.B1(n_111),
.B2(n_104),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_104),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_137),
.B1(n_131),
.B2(n_130),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_151),
.B(n_140),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_146),
.B(n_144),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_149),
.B(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_154),
.B(n_149),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_155),
.B(n_150),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_157),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_L g161 ( 
.A1(n_159),
.A2(n_160),
.B(n_148),
.Y(n_161)
);

AOI21xp33_ASAP7_75t_L g163 ( 
.A1(n_161),
.A2(n_162),
.B(n_158),
.Y(n_163)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_158),
.A2(n_153),
.A3(n_152),
.B1(n_157),
.B2(n_151),
.C1(n_150),
.C2(n_88),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_6),
.Y(n_164)
);


endmodule