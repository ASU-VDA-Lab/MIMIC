module fake_jpeg_12199_n_180 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_180);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_180;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_8),
.Y(n_12)
);

BUFx5_ASAP7_75t_L g13 ( 
.A(n_9),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_7),
.B(n_9),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_8),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_12),
.B(n_11),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_36),
.B(n_52),
.Y(n_76)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

CKINVDCx16_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_26),
.Y(n_38)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_39),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_47),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_13),
.Y(n_42)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

INVx4_ASAP7_75t_SL g44 ( 
.A(n_25),
.Y(n_44)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_18),
.B(n_7),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_45),
.B(n_50),
.Y(n_63)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_46),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_0),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_23),
.Y(n_48)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_27),
.Y(n_49)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_49),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_22),
.B(n_0),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_28),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_1),
.Y(n_53)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_53),
.Y(n_69)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVxp33_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_56),
.Y(n_85)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_14),
.Y(n_57)
);

OR2x2_ASAP7_75t_L g73 ( 
.A(n_57),
.B(n_58),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_15),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_31),
.B(n_1),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_60),
.Y(n_88)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_15),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_20),
.B(n_30),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_SL g91 ( 
.A1(n_61),
.A2(n_44),
.B(n_48),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_56),
.A2(n_20),
.B1(n_30),
.B2(n_29),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_65),
.A2(n_71),
.B1(n_75),
.B2(n_86),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_19),
.B1(n_29),
.B2(n_24),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_46),
.B1(n_58),
.B2(n_21),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_34),
.A2(n_19),
.B1(n_24),
.B2(n_21),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_83),
.B1(n_72),
.B2(n_70),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_31),
.B1(n_3),
.B2(n_4),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_42),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_42),
.A2(n_39),
.B1(n_41),
.B2(n_37),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_91),
.B(n_97),
.Y(n_135)
);

AND2x2_ASAP7_75t_SL g93 ( 
.A(n_74),
.B(n_48),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g130 ( 
.A(n_93),
.Y(n_130)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx2_ASAP7_75t_L g117 ( 
.A(n_94),
.Y(n_117)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_78),
.Y(n_95)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_85),
.B1(n_77),
.B2(n_90),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g120 ( 
.A1(n_96),
.A2(n_105),
.B1(n_110),
.B2(n_84),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_66),
.B(n_63),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_74),
.Y(n_98)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_98),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g99 ( 
.A(n_61),
.B(n_88),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_99),
.B(n_102),
.Y(n_116)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_100),
.Y(n_133)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_90),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_103),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_106),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_73),
.Y(n_106)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_89),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_107),
.B(n_109),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_69),
.B(n_76),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_112),
.B(n_113),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_88),
.B(n_73),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_75),
.A2(n_65),
.B1(n_64),
.B2(n_70),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_64),
.B(n_82),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_115),
.B(n_112),
.Y(n_124)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_70),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_78),
.B(n_80),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g115 ( 
.A(n_80),
.Y(n_115)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_91),
.B(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_105),
.A2(n_82),
.B1(n_89),
.B2(n_84),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_122),
.B(n_125),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_62),
.B1(n_106),
.B2(n_92),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_123),
.A2(n_126),
.B1(n_128),
.B2(n_130),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_124),
.A2(n_130),
.B(n_126),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_110),
.A2(n_92),
.B1(n_111),
.B2(n_101),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_93),
.A2(n_102),
.B1(n_98),
.B2(n_103),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_100),
.B1(n_94),
.B2(n_93),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_127),
.B(n_125),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_104),
.A2(n_115),
.B1(n_108),
.B2(n_107),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g137 ( 
.A(n_135),
.B(n_95),
.C(n_116),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_137),
.B(n_145),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_133),
.Y(n_138)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_138),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g141 ( 
.A(n_116),
.B(n_129),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_144),
.Y(n_153)
);

AOI21xp5_ASAP7_75t_SL g151 ( 
.A1(n_142),
.A2(n_143),
.B(n_121),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_119),
.A2(n_129),
.B(n_124),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_119),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_131),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_147),
.B(n_123),
.Y(n_152)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_131),
.Y(n_148)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_148),
.Y(n_159)
);

CKINVDCx14_ASAP7_75t_R g154 ( 
.A(n_149),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_136),
.B(n_128),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_150),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_151),
.B(n_147),
.C(n_149),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_155),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_SL g155 ( 
.A1(n_143),
.A2(n_120),
.B(n_134),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_160),
.B(n_137),
.C(n_142),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_162),
.B(n_165),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_153),
.B(n_141),
.Y(n_163)
);

HB1xp67_ASAP7_75t_L g170 ( 
.A(n_163),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_159),
.B(n_148),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_166),
.B1(n_158),
.B2(n_132),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_157),
.B(n_134),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_161),
.A2(n_154),
.B1(n_152),
.B2(n_146),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_169),
.B1(n_156),
.B2(n_118),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_162),
.A2(n_146),
.B1(n_158),
.B2(n_140),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_171),
.B(n_170),
.Y(n_173)
);

O2A1O1Ixp33_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_140),
.B(n_155),
.C(n_151),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_172),
.B(n_173),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_174),
.B(n_168),
.C(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_176),
.B(n_138),
.Y(n_178)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_175),
.A2(n_172),
.A3(n_168),
.B1(n_145),
.B2(n_138),
.C1(n_122),
.C2(n_117),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_177),
.B(n_178),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_179),
.B(n_117),
.Y(n_180)
);


endmodule