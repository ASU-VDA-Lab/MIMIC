module real_jpeg_23911_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_216;
wire n_128;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_0),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_1),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx8_ASAP7_75t_SL g58 ( 
.A(n_3),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_4),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_4),
.B(n_73),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_4),
.B(n_28),
.C(n_40),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_4),
.A2(n_37),
.B1(n_38),
.B2(n_164),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_4),
.B(n_86),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g236 ( 
.A1(n_4),
.A2(n_25),
.B1(n_234),
.B2(n_237),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_59),
.B1(n_60),
.B2(n_80),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_5),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_80),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_5),
.A2(n_64),
.B1(n_65),
.B2(n_80),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_80),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_6),
.A2(n_37),
.B1(n_38),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_49),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_49),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_6),
.A2(n_49),
.B1(n_59),
.B2(n_60),
.Y(n_115)
);

OAI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_7),
.A2(n_59),
.B1(n_60),
.B2(n_160),
.Y(n_159)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_7),
.Y(n_160)
);

OAI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_7),
.A2(n_64),
.B1(n_65),
.B2(n_160),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_160),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_160),
.Y(n_227)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_9),
.A2(n_27),
.B1(n_28),
.B2(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_9),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_9),
.A2(n_33),
.B1(n_63),
.B2(n_64),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_9),
.A2(n_33),
.B1(n_37),
.B2(n_38),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_9),
.A2(n_33),
.B1(n_59),
.B2(n_60),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_10),
.A2(n_37),
.B1(n_38),
.B2(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_10),
.A2(n_45),
.B1(n_59),
.B2(n_60),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_45),
.Y(n_150)
);

INVx13_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

NAND3xp33_ASAP7_75t_L g186 ( 
.A(n_11),
.B(n_58),
.C(n_59),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_12),
.A2(n_63),
.B1(n_64),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_12),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_12),
.A2(n_59),
.B1(n_60),
.B2(n_120),
.Y(n_161)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_120),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_120),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g167 ( 
.A1(n_13),
.A2(n_65),
.B1(n_70),
.B2(n_168),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_13),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_168),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_13),
.A2(n_37),
.B1(n_38),
.B2(n_168),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_168),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_14),
.Y(n_39)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx6_ASAP7_75t_L g103 ( 
.A(n_15),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_141),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_140),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_20),
.B(n_122),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_75),
.C(n_96),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_21),
.A2(n_75),
.B1(n_76),
.B2(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_21),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_50),
.B2(n_74),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_22),
.A2(n_51),
.B(n_53),
.Y(n_139)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_34),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_24),
.A2(n_51),
.B1(n_52),
.B2(n_53),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_24),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_24),
.A2(n_34),
.B1(n_51),
.B2(n_299),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_31),
.B(n_32),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_L g148 ( 
.A1(n_25),
.A2(n_149),
.B(n_151),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g215 ( 
.A1(n_25),
.A2(n_101),
.B(n_216),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_25),
.A2(n_153),
.B1(n_227),
.B2(n_234),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_25),
.A2(n_32),
.B(n_151),
.Y(n_253)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_26),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_26),
.A2(n_150),
.B1(n_152),
.B2(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_26),
.A2(n_152),
.B1(n_226),
.B2(n_228),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_29),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g42 ( 
.A1(n_27),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_27),
.B(n_240),
.Y(n_239)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx5_ASAP7_75t_L g238 ( 
.A(n_30),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_31),
.B(n_164),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_32),
.Y(n_104)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_34),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_SL g34 ( 
.A1(n_35),
.A2(n_43),
.B(n_46),
.Y(n_34)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_35),
.A2(n_42),
.B(n_133),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_35),
.A2(n_42),
.B1(n_213),
.B2(n_222),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_35),
.A2(n_89),
.B(n_272),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_42),
.Y(n_35)
);

OAI22xp33_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_38),
.B1(n_40),
.B2(n_41),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_37),
.A2(n_38),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

O2A1O1Ixp33_ASAP7_75t_L g248 ( 
.A1(n_37),
.A2(n_84),
.B(n_249),
.C(n_251),
.Y(n_248)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_38),
.B(n_209),
.Y(n_208)
);

NOR3xp33_ASAP7_75t_L g251 ( 
.A(n_38),
.B(n_59),
.C(n_83),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_SL g40 ( 
.A(n_41),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_42),
.B(n_48),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_42),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_42),
.A2(n_92),
.B(n_110),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_42),
.B(n_164),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_44),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_44),
.A2(n_91),
.B1(n_93),
.B2(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g157 ( 
.A1(n_47),
.A2(n_90),
.B(n_93),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_48),
.Y(n_94)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_66),
.B(n_68),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_54),
.A2(n_118),
.B(n_121),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_54),
.A2(n_56),
.B1(n_167),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_55),
.B(n_69),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_55),
.A2(n_73),
.B1(n_163),
.B2(n_166),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_55),
.A2(n_73),
.B1(n_119),
.B2(n_174),
.Y(n_290)
);

AND2x2_ASAP7_75t_SL g55 ( 
.A(n_56),
.B(n_62),
.Y(n_55)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_56),
.A2(n_127),
.B(n_128),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g62 ( 
.A1(n_57),
.A2(n_58),
.B1(n_63),
.B2(n_64),
.Y(n_62)
);

A2O1A1Ixp33_ASAP7_75t_L g185 ( 
.A1(n_57),
.A2(n_60),
.B(n_165),
.C(n_186),
.Y(n_185)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_59),
.A2(n_60),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

HAxp5_ASAP7_75t_SL g250 ( 
.A(n_60),
.B(n_164),
.CON(n_250),
.SN(n_250)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx11_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_65),
.Y(n_70)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_65),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_67),
.B(n_73),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_69),
.B(n_73),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_70),
.B(n_164),
.Y(n_165)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

OAI21xp33_ASAP7_75t_L g163 ( 
.A1(n_72),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_88),
.B(n_95),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_77),
.B(n_88),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_81),
.B1(n_86),
.B2(n_87),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g112 ( 
.A1(n_79),
.A2(n_85),
.B(n_113),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_114),
.Y(n_113)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_81),
.A2(n_87),
.B(n_136),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_81),
.A2(n_86),
.B1(n_159),
.B2(n_161),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_81),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_81),
.A2(n_86),
.B1(n_199),
.B2(n_250),
.Y(n_255)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_81),
.A2(n_136),
.B(n_179),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_85),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_115),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_85),
.A2(n_177),
.B1(n_198),
.B2(n_200),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_86),
.B(n_179),
.Y(n_178)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_92),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_90),
.B(n_91),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_90),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_91),
.A2(n_93),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_91),
.A2(n_93),
.B1(n_257),
.B2(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_95),
.A2(n_124),
.B1(n_137),
.B2(n_138),
.Y(n_123)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_95),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_96),
.A2(n_97),
.B1(n_309),
.B2(n_311),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_111),
.C(n_116),
.Y(n_97)
);

XNOR2xp5_ASAP7_75t_SL g300 ( 
.A(n_98),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_107),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_99),
.A2(n_100),
.B1(n_107),
.B2(n_108),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_101),
.B(n_105),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_104),
.Y(n_101)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g154 ( 
.A(n_103),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_103),
.A2(n_105),
.B(n_184),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_106),
.B(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_111),
.A2(n_112),
.B1(n_116),
.B2(n_117),
.Y(n_301)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_139),
.Y(n_122)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_124),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_129),
.B2(n_130),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_134),
.B2(n_135),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_142),
.A2(n_306),
.B(n_312),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_294),
.B(n_305),
.Y(n_142)
);

O2A1O1Ixp33_ASAP7_75t_SL g143 ( 
.A1(n_144),
.A2(n_201),
.B(n_282),
.C(n_293),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_188),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_145),
.B(n_188),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_169),
.Y(n_145)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_156),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_147),
.B(n_156),
.C(n_169),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_155),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_148),
.B(n_155),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_150),
.Y(n_149)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_158),
.C(n_162),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_158),
.Y(n_190)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_159),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_161),
.Y(n_176)
);

XOR2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_190),
.Y(n_189)
);

CKINVDCx14_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_170),
.A2(n_171),
.B1(n_180),
.B2(n_187),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_172),
.B(n_175),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_172),
.B(n_175),
.C(n_187),
.Y(n_292)
);

CKINVDCx14_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_177),
.B(n_178),
.Y(n_175)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_180),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_185),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_185),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_191),
.C(n_193),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_189),
.B(n_278),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_191),
.B(n_193),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.C(n_197),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_194),
.Y(n_267)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_197),
.B(n_266),
.Y(n_265)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_202),
.B(n_281),
.Y(n_201)
);

AOI21xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_276),
.B(n_280),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_261),
.B(n_275),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_205),
.A2(n_244),
.B(n_260),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_223),
.B(n_243),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_214),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_214),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_210),
.Y(n_207)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_208),
.B(n_210),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_217),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_215),
.B(n_218),
.C(n_221),
.Y(n_259)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_216),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_218),
.A2(n_219),
.B1(n_220),
.B2(n_221),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g257 ( 
.A(n_222),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_230),
.B(n_242),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_229),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_225),
.B(n_229),
.Y(n_242)
);

CKINVDCx14_ASAP7_75t_R g226 ( 
.A(n_227),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_231),
.A2(n_235),
.B(n_241),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_232),
.B(n_233),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_236),
.B(n_239),
.Y(n_235)
);

INVx5_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_245),
.B(n_259),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_245),
.B(n_259),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_246),
.B(n_255),
.C(n_256),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_252),
.B2(n_253),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_247),
.B(n_253),
.Y(n_270)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_263),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_268),
.B2(n_269),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_271),
.C(n_273),
.Y(n_279)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_269)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_270),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_277),
.B(n_279),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_277),
.B(n_279),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_284),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_283),
.B(n_284),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_292),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_287),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_287),
.C(n_292),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_288),
.B(n_290),
.C(n_291),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_296),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_295),
.B(n_296),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_304),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_298),
.A2(n_300),
.B1(n_302),
.B2(n_303),
.Y(n_297)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_298),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_298),
.B(n_303),
.C(n_304),
.Y(n_307)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_307),
.B(n_308),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_307),
.B(n_308),
.Y(n_312)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_309),
.Y(n_311)
);


endmodule