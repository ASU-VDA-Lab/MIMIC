module fake_aes_7083_n_11 (n_1, n_2, n_0, n_11);
input n_1;
input n_2;
input n_0;
output n_11;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_7;
wire n_10;
wire n_8;
INVx4_ASAP7_75t_L g3 ( .A(n_1), .Y(n_3) );
CKINVDCx5p33_ASAP7_75t_R g4 ( .A(n_1), .Y(n_4) );
OAI22xp5_ASAP7_75t_L g5 ( .A1(n_4), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_5) );
INVx2_ASAP7_75t_L g6 ( .A(n_3), .Y(n_6) );
OAI22xp33_ASAP7_75t_L g7 ( .A1(n_5), .A2(n_3), .B1(n_1), .B2(n_2), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
OAI211xp5_ASAP7_75t_L g9 ( .A1(n_8), .A2(n_3), .B(n_6), .C(n_2), .Y(n_9) );
OAI22xp5_ASAP7_75t_L g10 ( .A1(n_9), .A2(n_8), .B1(n_3), .B2(n_2), .Y(n_10) );
AOI222xp33_ASAP7_75t_L g11 ( .A1(n_10), .A2(n_0), .B1(n_3), .B2(n_8), .C1(n_7), .C2(n_5), .Y(n_11) );
endmodule