module fake_jpeg_8288_n_225 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_225);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_225;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx8_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_1),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_1),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

BUFx4f_ASAP7_75t_SL g36 ( 
.A(n_32),
.Y(n_36)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_40),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

BUFx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_25),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_25),
.Y(n_41)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

AND2x4_ASAP7_75t_L g43 ( 
.A(n_35),
.B(n_0),
.Y(n_43)
);

AO22x1_ASAP7_75t_L g60 ( 
.A1(n_43),
.A2(n_34),
.B1(n_24),
.B2(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_31),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_47),
.B(n_33),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_43),
.A2(n_34),
.B1(n_24),
.B2(n_35),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_56),
.B1(n_59),
.B2(n_27),
.Y(n_87)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_50),
.Y(n_73)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_52),
.Y(n_72)
);

CKINVDCx12_ASAP7_75t_R g52 ( 
.A(n_43),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_18),
.B1(n_17),
.B2(n_23),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_18),
.B1(n_17),
.B2(n_23),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_28),
.B1(n_21),
.B2(n_26),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_44),
.A2(n_18),
.B1(n_20),
.B2(n_22),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_60),
.B(n_61),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_22),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_37),
.Y(n_62)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_62),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_28),
.B1(n_30),
.B2(n_29),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_63),
.A2(n_0),
.B(n_2),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_67),
.B(n_68),
.Y(n_80)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_37),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_69),
.B(n_40),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_42),
.B(n_34),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_42),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_75),
.B(n_91),
.Y(n_103)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_76),
.B(n_77),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_53),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_66),
.B(n_31),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_79),
.B(n_82),
.Y(n_105)
);

AO21x1_ASAP7_75t_SL g121 ( 
.A1(n_81),
.A2(n_6),
.B(n_7),
.Y(n_121)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_59),
.Y(n_82)
);

A2O1A1Ixp33_ASAP7_75t_L g83 ( 
.A1(n_50),
.A2(n_26),
.B(n_21),
.C(n_29),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g119 ( 
.A(n_83),
.B(n_5),
.Y(n_119)
);

OAI21xp5_ASAP7_75t_SL g84 ( 
.A1(n_71),
.A2(n_60),
.B(n_48),
.Y(n_84)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_84),
.B(n_97),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_53),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_85),
.B(n_88),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_60),
.A2(n_33),
.B1(n_30),
.B2(n_24),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_86),
.A2(n_92),
.B1(n_93),
.B2(n_49),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_82),
.B1(n_98),
.B2(n_89),
.Y(n_106)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_70),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_89),
.B(n_99),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_61),
.B(n_41),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_55),
.A2(n_39),
.B1(n_41),
.B2(n_3),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_55),
.A2(n_39),
.B1(n_2),
.B2(n_3),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_7),
.B(n_8),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_67),
.B(n_3),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_56),
.B(n_4),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_98),
.B(n_6),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_64),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_54),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_100),
.B(n_54),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_90),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_109),
.Y(n_144)
);

A2O1A1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_74),
.A2(n_72),
.B(n_91),
.C(n_94),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_104),
.B(n_118),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_106),
.B(n_86),
.Y(n_133)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_112),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_87),
.A2(n_51),
.B1(n_65),
.B2(n_69),
.Y(n_114)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_114),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_80),
.B(n_65),
.Y(n_115)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_115),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_90),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_116),
.B(n_119),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_80),
.B(n_49),
.Y(n_117)
);

CKINVDCx16_ASAP7_75t_R g126 ( 
.A(n_117),
.Y(n_126)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_75),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_120),
.A2(n_121),
.B1(n_124),
.B2(n_85),
.Y(n_145)
);

FAx1_ASAP7_75t_SL g130 ( 
.A(n_122),
.B(n_93),
.CI(n_83),
.CON(n_130),
.SN(n_130)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_6),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_97),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_113),
.B(n_84),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_128),
.C(n_132),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_113),
.B(n_74),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_130),
.B(n_139),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_131),
.B(n_133),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_73),
.C(n_88),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_103),
.B(n_73),
.C(n_99),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g149 ( 
.A(n_134),
.B(n_136),
.Y(n_149)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_103),
.B(n_81),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_123),
.B(n_97),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_138),
.B(n_140),
.Y(n_167)
);

INVx13_ASAP7_75t_L g139 ( 
.A(n_102),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_106),
.B(n_76),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_116),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_143),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g143 ( 
.A(n_110),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_101),
.B1(n_119),
.B2(n_110),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g146 ( 
.A1(n_121),
.A2(n_100),
.B(n_77),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_146),
.A2(n_117),
.B1(n_101),
.B2(n_108),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_127),
.A2(n_111),
.B(n_124),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_128),
.Y(n_168)
);

AOI322xp5_ASAP7_75t_SL g154 ( 
.A1(n_135),
.A2(n_104),
.A3(n_105),
.B1(n_107),
.B2(n_111),
.C1(n_121),
.C2(n_115),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_154),
.B(n_156),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_140),
.A2(n_114),
.B1(n_104),
.B2(n_105),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_155),
.A2(n_159),
.B1(n_137),
.B2(n_147),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_144),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_142),
.B(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_157),
.B(n_164),
.Y(n_172)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_139),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_158),
.B(n_161),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_137),
.A2(n_109),
.B1(n_120),
.B2(n_122),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_160),
.A2(n_166),
.B1(n_145),
.B2(n_146),
.Y(n_183)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_132),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_162),
.B(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_134),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_146),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_153),
.Y(n_188)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_171),
.B(n_175),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_158),
.B(n_129),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_173),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_125),
.C(n_133),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_174),
.B(n_182),
.C(n_130),
.Y(n_195)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_160),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_136),
.C(n_138),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_151),
.C(n_149),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_164),
.B(n_126),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_179),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_178),
.A2(n_180),
.B1(n_167),
.B2(n_161),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g179 ( 
.A(n_150),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_167),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_149),
.B(n_131),
.C(n_95),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g186 ( 
.A(n_183),
.B(n_159),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_184),
.B(n_189),
.C(n_192),
.Y(n_197)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_186),
.B(n_195),
.Y(n_202)
);

XOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_168),
.B(n_151),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_188),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_174),
.B(n_163),
.C(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_191),
.B(n_193),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_176),
.B(n_155),
.Y(n_192)
);

NAND3xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_130),
.C(n_148),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_194),
.B(n_171),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_201),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g198 ( 
.A1(n_190),
.A2(n_175),
.B(n_169),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_198),
.A2(n_143),
.B(n_96),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_185),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_192),
.B(n_182),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_203),
.B(n_148),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g204 ( 
.A1(n_187),
.A2(n_172),
.B(n_181),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_204),
.B(n_169),
.Y(n_207)
);

AOI322xp5_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_178),
.A3(n_195),
.B1(n_189),
.B2(n_184),
.C1(n_181),
.C2(n_188),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_205),
.B(n_208),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_207),
.A2(n_197),
.B(n_202),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_198),
.B(n_95),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_210),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_197),
.A2(n_13),
.B1(n_16),
.B2(n_15),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_211),
.A2(n_202),
.B1(n_16),
.B2(n_15),
.Y(n_212)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_212),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_214),
.B(n_9),
.Y(n_219)
);

AOI322xp5_ASAP7_75t_L g216 ( 
.A1(n_208),
.A2(n_203),
.A3(n_200),
.B1(n_90),
.B2(n_12),
.C1(n_11),
.C2(n_10),
.Y(n_216)
);

O2A1O1Ixp33_ASAP7_75t_SL g217 ( 
.A1(n_216),
.A2(n_206),
.B(n_210),
.C(n_12),
.Y(n_217)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_217),
.B(n_216),
.C(n_11),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_213),
.A2(n_200),
.B(n_9),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_218),
.B(n_219),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_221),
.B(n_220),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_223),
.B(n_222),
.Y(n_224)
);

FAx1_ASAP7_75t_SL g225 ( 
.A(n_224),
.B(n_215),
.CI(n_219),
.CON(n_225),
.SN(n_225)
);


endmodule