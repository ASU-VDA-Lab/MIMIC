module real_jpeg_33296_n_18 (n_17, n_8, n_0, n_2, n_579, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_579;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_556;
wire n_507;
wire n_57;
wire n_157;
wire n_560;
wire n_84;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_487;
wire n_242;
wire n_493;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_546;
wire n_531;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_0),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g277 ( 
.A(n_0),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_0),
.Y(n_315)
);

BUFx3_ASAP7_75t_L g329 ( 
.A(n_0),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_1),
.Y(n_559)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_2),
.B(n_40),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_2),
.B(n_61),
.Y(n_60)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_2),
.B(n_150),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_2),
.B(n_172),
.Y(n_171)
);

AND2x2_ASAP7_75t_SL g207 ( 
.A(n_2),
.B(n_208),
.Y(n_207)
);

AND2x2_ASAP7_75t_L g358 ( 
.A(n_2),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_SL g408 ( 
.A(n_2),
.B(n_210),
.Y(n_408)
);

AND2x2_ASAP7_75t_L g470 ( 
.A(n_2),
.B(n_471),
.Y(n_470)
);

NOR2xp33_ASAP7_75t_L g558 ( 
.A(n_3),
.B(n_559),
.Y(n_558)
);

CKINVDCx11_ASAP7_75t_R g570 ( 
.A(n_3),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_4),
.B(n_30),
.Y(n_29)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_4),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g92 ( 
.A(n_4),
.B(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_4),
.B(n_155),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_4),
.B(n_222),
.Y(n_221)
);

AND2x2_ASAP7_75t_SL g272 ( 
.A(n_4),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_4),
.B(n_312),
.Y(n_311)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_5),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_5),
.Y(n_170)
);

BUFx3_ASAP7_75t_L g474 ( 
.A(n_5),
.Y(n_474)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_6),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_6),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_6),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_6),
.B(n_169),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_6),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_SL g295 ( 
.A(n_6),
.B(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_6),
.B(n_310),
.Y(n_309)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_7),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_7),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_8),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_9),
.B(n_34),
.Y(n_33)
);

AND2x4_ASAP7_75t_L g163 ( 
.A(n_9),
.B(n_164),
.Y(n_163)
);

NAND2x1_ASAP7_75t_L g191 ( 
.A(n_9),
.B(n_192),
.Y(n_191)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_9),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_9),
.B(n_416),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_9),
.B(n_465),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_9),
.B(n_507),
.Y(n_506)
);

INVxp67_ASAP7_75t_L g531 ( 
.A(n_9),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_10),
.B(n_102),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g115 ( 
.A(n_10),
.B(n_116),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_10),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_10),
.B(n_93),
.Y(n_205)
);

AND2x2_ASAP7_75t_L g374 ( 
.A(n_10),
.B(n_262),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_10),
.B(n_403),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_10),
.B(n_486),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g516 ( 
.A(n_10),
.B(n_169),
.Y(n_516)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_11),
.Y(n_85)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_11),
.Y(n_95)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_11),
.Y(n_373)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_12),
.Y(n_53)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_12),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_13),
.B(n_52),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_13),
.B(n_65),
.Y(n_64)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_13),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_13),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_13),
.B(n_300),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_13),
.B(n_322),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_13),
.B(n_328),
.Y(n_327)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_14),
.Y(n_194)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_14),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_15),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g360 ( 
.A(n_15),
.Y(n_360)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_34),
.Y(n_42)
);

AND2x4_ASAP7_75t_SL g56 ( 
.A(n_16),
.B(n_57),
.Y(n_56)
);

AND2x2_ASAP7_75t_L g79 ( 
.A(n_16),
.B(n_80),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_16),
.B(n_76),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_16),
.B(n_99),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g235 ( 
.A(n_16),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_16),
.B(n_380),
.Y(n_379)
);

AND2x2_ASAP7_75t_SL g391 ( 
.A(n_16),
.B(n_392),
.Y(n_391)
);

AND2x2_ASAP7_75t_SL g81 ( 
.A(n_17),
.B(n_82),
.Y(n_81)
);

AND2x2_ASAP7_75t_SL g109 ( 
.A(n_17),
.B(n_110),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_17),
.B(n_138),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_17),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_17),
.B(n_239),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_17),
.B(n_242),
.Y(n_241)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_17),
.B(n_276),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_17),
.B(n_222),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_571),
.Y(n_18)
);

AOI321xp33_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_447),
.A3(n_545),
.B1(n_560),
.B2(n_564),
.C(n_579),
.Y(n_19)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_20),
.Y(n_572)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

OA21x2_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_343),
.B(n_440),
.Y(n_22)
);

NAND3xp33_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_176),
.C(n_223),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_131),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_25),
.B(n_131),
.Y(n_442)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_70),
.C(n_106),
.Y(n_25)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_26),
.B(n_71),
.Y(n_227)
);

XOR2x2_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_54),
.Y(n_26)
);

XOR2xp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_36),
.Y(n_27)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_28),
.B(n_54),
.C(n_175),
.Y(n_174)
);

OA21x2_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_33),
.B(n_35),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_33),
.Y(n_35)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_31),
.Y(n_404)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g161 ( 
.A(n_35),
.B(n_162),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_35),
.B(n_160),
.C(n_162),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_36),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_43),
.C(n_50),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_37),
.A2(n_38),
.B1(n_231),
.B2(n_232),
.Y(n_230)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_38),
.A2(n_220),
.B(n_376),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_42),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_39),
.A2(n_101),
.B1(n_104),
.B2(n_105),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g104 ( 
.A(n_39),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_39),
.B(n_105),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_39),
.A2(n_104),
.B1(n_220),
.B2(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_39),
.B(n_42),
.Y(n_376)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_40),
.Y(n_310)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_41),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_41),
.Y(n_243)
);

INVx1_ASAP7_75t_SL g218 ( 
.A(n_42),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_42),
.A2(n_218),
.B1(n_241),
.B2(n_280),
.Y(n_279)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_42),
.A2(n_378),
.B(n_383),
.Y(n_377)
);

OAI221xp5_ASAP7_75t_L g383 ( 
.A1(n_42),
.A2(n_235),
.B1(n_379),
.B2(n_381),
.C(n_382),
.Y(n_383)
);

MAJx2_ASAP7_75t_L g388 ( 
.A(n_42),
.B(n_379),
.C(n_381),
.Y(n_388)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_43),
.A2(n_44),
.B1(n_50),
.B2(n_51),
.Y(n_231)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx3_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_49),
.Y(n_141)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_52),
.Y(n_507)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_53),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_53),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_55),
.B(n_64),
.C(n_68),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g487 ( 
.A1(n_55),
.A2(n_56),
.B1(n_79),
.B2(n_488),
.Y(n_487)
);

AOI22xp5_ASAP7_75t_L g514 ( 
.A1(n_55),
.A2(n_56),
.B1(n_152),
.B2(n_153),
.Y(n_514)
);

MAJx2_ASAP7_75t_L g517 ( 
.A(n_55),
.B(n_79),
.C(n_485),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_55),
.B(n_153),
.C(n_515),
.Y(n_536)
);

INVx4_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_57),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_58),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_64),
.B1(n_68),
.B2(n_69),
.Y(n_59)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_60),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g367 ( 
.A1(n_60),
.A2(n_68),
.B1(n_368),
.B2(n_369),
.Y(n_367)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_63),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_63),
.Y(n_324)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_64),
.Y(n_69)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_67),
.Y(n_222)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_67),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_68),
.B(n_410),
.C(n_411),
.Y(n_409)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

MAJx2_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_86),
.C(n_100),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_72),
.B(n_246),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_73),
.B(n_81),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

MAJx2_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_79),
.C(n_81),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_75),
.B(n_78),
.Y(n_74)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_77),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g208 ( 
.A(n_77),
.Y(n_208)
);

BUFx6f_ASAP7_75t_L g418 ( 
.A(n_77),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_78),
.B(n_266),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_79),
.B(n_402),
.Y(n_401)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_79),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_79),
.B(n_381),
.C(n_402),
.Y(n_491)
);

HB1xp67_ASAP7_75t_L g239 ( 
.A(n_80),
.Y(n_239)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_85),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_86),
.B(n_100),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_92),
.C(n_96),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_88),
.B(n_97),
.Y(n_285)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_92),
.B(n_285),
.Y(n_284)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

BUFx5_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx4_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_106),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_125),
.B2(n_130),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_107),
.B(n_126),
.C(n_129),
.Y(n_133)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_113),
.Y(n_108)
);

MAJx2_ASAP7_75t_L g160 ( 
.A(n_109),
.B(n_115),
.C(n_119),
.Y(n_160)
);

INVx5_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_112),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_119),
.B2(n_120),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_118),
.Y(n_274)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_121),
.B(n_123),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g486 ( 
.A(n_123),
.Y(n_486)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_125),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_158),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_132),
.B(n_159),
.C(n_174),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_134),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_133),
.B(n_135),
.C(n_147),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_147),
.Y(n_134)
);

XNOR2x2_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_146),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_137),
.B(n_142),
.Y(n_136)
);

NOR2xp67_ASAP7_75t_SL g186 ( 
.A(n_137),
.B(n_142),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_137),
.B(n_142),
.Y(n_187)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g185 ( 
.A1(n_146),
.A2(n_186),
.B(n_187),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g216 ( 
.A(n_148),
.B(n_152),
.C(n_154),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_148),
.A2(n_149),
.B1(n_415),
.B2(n_419),
.Y(n_414)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g490 ( 
.A(n_149),
.B(n_408),
.C(n_419),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_154),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g537 ( 
.A1(n_152),
.A2(n_153),
.B1(n_538),
.B2(n_539),
.Y(n_537)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_152),
.B(n_195),
.C(n_408),
.Y(n_551)
);

INVx2_ASAP7_75t_SL g152 ( 
.A(n_153),
.Y(n_152)
);

BUFx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_174),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_167),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_163),
.B(n_168),
.C(n_171),
.Y(n_198)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_171),
.B(n_235),
.Y(n_234)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

AOI21x1_ASAP7_75t_L g441 ( 
.A1(n_177),
.A2(n_442),
.B(n_443),
.Y(n_441)
);

AND2x2_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g443 ( 
.A(n_178),
.B(n_179),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_180),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_201),
.B2(n_202),
.Y(n_181)
);

HB1xp67_ASAP7_75t_L g436 ( 
.A(n_182),
.Y(n_436)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_200),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_188),
.Y(n_184)
);

HB1xp67_ASAP7_75t_L g429 ( 
.A(n_185),
.Y(n_429)
);

HB1xp67_ASAP7_75t_L g430 ( 
.A(n_188),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_198),
.B2(n_199),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_191),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g197 ( 
.A(n_191),
.Y(n_197)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_194),
.Y(n_193)
);

MAJx2_ASAP7_75t_L g351 ( 
.A(n_195),
.B(n_197),
.C(n_199),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g538 ( 
.A1(n_195),
.A2(n_196),
.B1(n_407),
.B2(n_408),
.Y(n_538)
);

OAI22xp5_ASAP7_75t_SL g553 ( 
.A1(n_195),
.A2(n_196),
.B1(n_379),
.B2(n_382),
.Y(n_553)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_198),
.Y(n_199)
);

INVxp33_ASAP7_75t_L g428 ( 
.A(n_200),
.Y(n_428)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

HB1xp67_ASAP7_75t_L g438 ( 
.A(n_202),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_203),
.B(n_215),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_204),
.B(n_348),
.C(n_349),
.Y(n_347)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_206),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_205),
.B(n_209),
.C(n_213),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_209),
.B1(n_213),
.B2(n_214),
.Y(n_206)
);

INVx1_ASAP7_75t_SL g213 ( 
.A(n_207),
.Y(n_213)
);

AOI22xp33_ASAP7_75t_L g463 ( 
.A1(n_207),
.A2(n_213),
.B1(n_464),
.B2(n_469),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g508 ( 
.A(n_207),
.B(n_469),
.C(n_509),
.Y(n_508)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_209),
.Y(n_214)
);

INVx4_ASAP7_75t_SL g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.Y(n_215)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_216),
.Y(n_349)
);

INVxp67_ASAP7_75t_SL g348 ( 
.A(n_217),
.Y(n_348)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_224),
.A2(n_250),
.B(n_342),
.Y(n_223)
);

NOR2xp67_ASAP7_75t_SL g224 ( 
.A(n_225),
.B(n_228),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_225),
.B(n_228),
.Y(n_342)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.Y(n_225)
);

A2O1A1Ixp33_ASAP7_75t_SL g228 ( 
.A1(n_229),
.A2(n_233),
.B(n_244),
.C(n_247),
.Y(n_228)
);

INVxp67_ASAP7_75t_SL g249 ( 
.A(n_229),
.Y(n_249)
);

HB1xp67_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_230),
.A2(n_233),
.B1(n_248),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_230),
.Y(n_340)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_231),
.Y(n_232)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_233),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.C(n_240),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_234),
.A2(n_237),
.B1(n_238),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_234),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_L g378 ( 
.A1(n_235),
.A2(n_379),
.B1(n_381),
.B2(n_382),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g381 ( 
.A(n_235),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_L g399 ( 
.A1(n_235),
.A2(n_381),
.B1(n_400),
.B2(n_401),
.Y(n_399)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_240),
.B(n_289),
.Y(n_288)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_241),
.Y(n_280)
);

INVx6_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_244),
.A2(n_245),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g250 ( 
.A1(n_251),
.A2(n_334),
.B(n_341),
.Y(n_250)
);

OAI21xp33_ASAP7_75t_L g251 ( 
.A1(n_252),
.A2(n_291),
.B(n_333),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_281),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_253),
.B(n_281),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_271),
.C(n_278),
.Y(n_253)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_254),
.A2(n_255),
.B1(n_303),
.B2(n_304),
.Y(n_302)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_265),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_261),
.B2(n_264),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_257),
.B(n_264),
.C(n_265),
.Y(n_283)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_261),
.Y(n_264)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx2_ASAP7_75t_SL g267 ( 
.A(n_268),
.Y(n_267)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_271),
.A2(n_278),
.B1(n_279),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_271),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_275),
.Y(n_294)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

BUFx4f_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_288),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_286),
.B2(n_287),
.Y(n_282)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_283),
.Y(n_286)
);

INVx1_ASAP7_75t_SL g287 ( 
.A(n_284),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_284),
.B(n_286),
.C(n_336),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_288),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_306),
.B(n_332),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_302),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_293),
.B(n_302),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.C(n_298),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_317),
.Y(n_316)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_295),
.A2(n_298),
.B1(n_299),
.B2(n_318),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_295),
.Y(n_318)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_307),
.A2(n_319),
.B(n_331),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_316),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_308),
.B(n_316),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_309),
.B(n_311),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_309),
.B(n_327),
.Y(n_326)
);

INVx3_ASAP7_75t_SL g312 ( 
.A(n_313),
.Y(n_312)
);

INVx8_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_315),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_326),
.B(n_330),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_325),
.Y(n_330)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

HB1xp67_ASAP7_75t_L g323 ( 
.A(n_324),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_337),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g341 ( 
.A(n_335),
.B(n_337),
.Y(n_341)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_431),
.Y(n_343)
);

NAND2xp33_ASAP7_75t_L g344 ( 
.A(n_345),
.B(n_420),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g445 ( 
.A1(n_345),
.A2(n_420),
.B1(n_432),
.B2(n_434),
.Y(n_445)
);

NOR2x1_ASAP7_75t_SL g446 ( 
.A(n_345),
.B(n_420),
.Y(n_446)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_364),
.Y(n_345)
);

INVxp33_ASAP7_75t_SL g454 ( 
.A(n_346),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_350),
.C(n_352),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_347),
.B(n_423),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_350),
.A2(n_351),
.B1(n_354),
.B2(n_355),
.Y(n_423)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_356),
.B(n_363),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_357),
.A2(n_358),
.B1(n_361),
.B2(n_362),
.Y(n_356)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_357),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_357),
.B(n_361),
.C(n_363),
.Y(n_385)
);

INVx2_ASAP7_75t_SL g361 ( 
.A(n_358),
.Y(n_361)
);

OAI22xp5_ASAP7_75t_SL g389 ( 
.A1(n_358),
.A2(n_361),
.B1(n_390),
.B2(n_391),
.Y(n_389)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_358),
.A2(n_361),
.B1(n_505),
.B2(n_506),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_358),
.B(n_505),
.C(n_510),
.Y(n_540)
);

BUFx6f_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx2_ASAP7_75t_L g468 ( 
.A(n_360),
.Y(n_468)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_361),
.B(n_388),
.C(n_476),
.Y(n_475)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_397),
.Y(n_364)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

XNOR2xp5_ASAP7_75t_L g365 ( 
.A(n_366),
.B(n_384),
.Y(n_365)
);

INVxp33_ASAP7_75t_SL g457 ( 
.A(n_366),
.Y(n_457)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_375),
.C(n_377),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_367),
.B(n_375),
.Y(n_425)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_374),
.Y(n_369)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_370),
.Y(n_411)
);

INVx4_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx2_ASAP7_75t_SL g372 ( 
.A(n_373),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_374),
.Y(n_410)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_377),
.B(n_425),
.Y(n_424)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_379),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g384 ( 
.A1(n_385),
.A2(n_386),
.B1(n_387),
.B2(n_396),
.Y(n_384)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_385),
.Y(n_396)
);

HB1xp67_ASAP7_75t_L g458 ( 
.A(n_386),
.Y(n_458)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

XOR2xp5_ASAP7_75t_L g387 ( 
.A(n_388),
.B(n_389),
.Y(n_387)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_391),
.Y(n_390)
);

BUFx2_ASAP7_75t_L g476 ( 
.A(n_391),
.Y(n_476)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_395),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_396),
.B(n_457),
.C(n_458),
.Y(n_456)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_397),
.Y(n_453)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_398),
.B(n_405),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

MAJx2_ASAP7_75t_L g479 ( 
.A(n_399),
.B(n_480),
.C(n_481),
.Y(n_479)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_401),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g403 ( 
.A(n_404),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_406),
.B(n_413),
.Y(n_405)
);

AOI22xp33_ASAP7_75t_L g406 ( 
.A1(n_407),
.A2(n_408),
.B1(n_409),
.B2(n_412),
.Y(n_406)
);

OAI22xp5_ASAP7_75t_L g480 ( 
.A1(n_407),
.A2(n_408),
.B1(n_413),
.B2(n_414),
.Y(n_480)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_408),
.Y(n_407)
);

INVxp67_ASAP7_75t_SL g412 ( 
.A(n_409),
.Y(n_412)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_409),
.Y(n_481)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_415),
.Y(n_419)
);

INVx2_ASAP7_75t_SL g416 ( 
.A(n_417),
.Y(n_416)
);

INVx3_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_424),
.C(n_426),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_422),
.B(n_424),
.Y(n_433)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_427),
.Y(n_426)
);

XNOR2xp5_ASAP7_75t_L g432 ( 
.A(n_427),
.B(n_433),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g427 ( 
.A(n_428),
.B(n_429),
.C(n_430),
.Y(n_427)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_434),
.Y(n_431)
);

NOR2xp67_ASAP7_75t_L g444 ( 
.A(n_432),
.B(n_434),
.Y(n_444)
);

MAJx2_ASAP7_75t_L g434 ( 
.A(n_435),
.B(n_437),
.C(n_439),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

O2A1O1Ixp33_ASAP7_75t_SL g440 ( 
.A1(n_441),
.A2(n_444),
.B(n_445),
.C(n_446),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_447),
.B(n_577),
.Y(n_576)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

OAI31xp33_ASAP7_75t_L g564 ( 
.A1(n_448),
.A2(n_546),
.A3(n_565),
.B(n_569),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_449),
.B(n_520),
.Y(n_448)
);

OA21x2_ASAP7_75t_SL g449 ( 
.A1(n_450),
.A2(n_492),
.B(n_518),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_451),
.B(n_455),
.Y(n_450)
);

OR2x2_ASAP7_75t_L g568 ( 
.A(n_451),
.B(n_455),
.Y(n_568)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_453),
.C(n_454),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_456),
.B(n_459),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_456),
.B(n_483),
.C(n_495),
.Y(n_494)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_482),
.Y(n_459)
);

INVxp67_ASAP7_75t_SL g495 ( 
.A(n_460),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_461),
.B(n_479),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_462),
.A2(n_475),
.B1(n_477),
.B2(n_478),
.Y(n_461)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_462),
.Y(n_477)
);

XOR2x2_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_470),
.Y(n_462)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_464),
.Y(n_469)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_466),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_468),
.Y(n_467)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_470),
.Y(n_509)
);

XOR2xp5_ASAP7_75t_L g552 ( 
.A(n_470),
.B(n_553),
.Y(n_552)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g472 ( 
.A(n_473),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

BUFx6f_ASAP7_75t_L g535 ( 
.A(n_474),
.Y(n_535)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_475),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_477),
.B(n_478),
.C(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_479),
.Y(n_498)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_489),
.Y(n_483)
);

MAJx2_ASAP7_75t_L g500 ( 
.A(n_484),
.B(n_490),
.C(n_491),
.Y(n_500)
);

XOR2x2_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_487),
.Y(n_484)
);

XNOR2xp5_ASAP7_75t_L g489 ( 
.A(n_490),
.B(n_491),
.Y(n_489)
);

INVxp67_ASAP7_75t_L g567 ( 
.A(n_492),
.Y(n_567)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_493),
.B(n_496),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_494),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_494),
.B(n_519),
.Y(n_518)
);

INVxp33_ASAP7_75t_SL g519 ( 
.A(n_496),
.Y(n_519)
);

XNOR2xp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_499),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_497),
.B(n_523),
.C(n_524),
.Y(n_522)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_500),
.B(n_501),
.Y(n_499)
);

INVxp33_ASAP7_75t_SL g523 ( 
.A(n_500),
.Y(n_523)
);

INVxp33_ASAP7_75t_SL g524 ( 
.A(n_501),
.Y(n_524)
);

XOR2x2_ASAP7_75t_L g501 ( 
.A(n_502),
.B(n_511),
.Y(n_501)
);

MAJx2_ASAP7_75t_L g543 ( 
.A(n_502),
.B(n_512),
.C(n_544),
.Y(n_543)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_503),
.A2(n_504),
.B1(n_508),
.B2(n_510),
.Y(n_502)
);

INVxp33_ASAP7_75t_SL g503 ( 
.A(n_504),
.Y(n_503)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_506),
.Y(n_505)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_508),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_L g511 ( 
.A(n_512),
.B(n_517),
.Y(n_511)
);

OAI22xp5_ASAP7_75t_L g512 ( 
.A1(n_513),
.A2(n_514),
.B1(n_515),
.B2(n_516),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_514),
.Y(n_513)
);

CKINVDCx16_ASAP7_75t_R g515 ( 
.A(n_516),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g544 ( 
.A(n_517),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g561 ( 
.A(n_520),
.B(n_562),
.Y(n_561)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_521),
.Y(n_520)
);

NOR2xp33_ASAP7_75t_L g521 ( 
.A(n_522),
.B(n_525),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g563 ( 
.A(n_522),
.B(n_525),
.Y(n_563)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_526),
.B(n_542),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_L g526 ( 
.A1(n_527),
.A2(n_528),
.B1(n_540),
.B2(n_541),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g555 ( 
.A(n_527),
.B(n_540),
.C(n_543),
.Y(n_555)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_528),
.Y(n_527)
);

XNOR2x1_ASAP7_75t_L g528 ( 
.A(n_529),
.B(n_537),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_530),
.B(n_536),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g554 ( 
.A(n_530),
.B(n_536),
.C(n_537),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_531),
.B(n_532),
.Y(n_530)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_533),
.Y(n_532)
);

INVx3_ASAP7_75t_L g533 ( 
.A(n_534),
.Y(n_533)
);

INVx6_ASAP7_75t_L g534 ( 
.A(n_535),
.Y(n_534)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_538),
.Y(n_539)
);

INVxp67_ASAP7_75t_SL g541 ( 
.A(n_540),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_543),
.Y(n_542)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_546),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g546 ( 
.A(n_547),
.B(n_557),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_547),
.B(n_558),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g547 ( 
.A(n_548),
.B(n_556),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_549),
.B(n_555),
.Y(n_548)
);

OR2x2_ASAP7_75t_L g556 ( 
.A(n_549),
.B(n_555),
.Y(n_556)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_550),
.B(n_554),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_551),
.B(n_552),
.Y(n_550)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_557),
.B(n_570),
.Y(n_569)
);

CKINVDCx20_ASAP7_75t_R g557 ( 
.A(n_558),
.Y(n_557)
);

NOR2xp33_ASAP7_75t_L g573 ( 
.A(n_560),
.B(n_574),
.Y(n_573)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_561),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g571 ( 
.A1(n_561),
.A2(n_572),
.B1(n_573),
.B2(n_576),
.Y(n_571)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_563),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_565),
.B(n_575),
.Y(n_574)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_566),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g566 ( 
.A(n_567),
.B(n_568),
.Y(n_566)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_575),
.Y(n_577)
);


endmodule