module fake_jpeg_6912_n_290 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_290);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_154;
wire n_127;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_155;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_7),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_11),
.Y(n_25)
);

CKINVDCx16_ASAP7_75t_R g26 ( 
.A(n_0),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_12),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_43),
.Y(n_65)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_20),
.B(n_0),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_34),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_39),
.Y(n_46)
);

INVx11_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_47)
);

OAI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_47),
.A2(n_64),
.B1(n_29),
.B2(n_45),
.Y(n_79)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_41),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_50),
.B(n_52),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_53),
.B(n_57),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_36),
.A2(n_19),
.B1(n_27),
.B2(n_25),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_54),
.A2(n_67),
.B1(n_26),
.B2(n_29),
.Y(n_78)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_34),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_35),
.Y(n_60)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_43),
.Y(n_62)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_40),
.A2(n_20),
.B1(n_32),
.B2(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_26),
.B1(n_32),
.B2(n_23),
.Y(n_67)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g83 ( 
.A(n_68),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_69),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_65),
.B(n_44),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_70),
.B(n_72),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_71),
.B(n_76),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_53),
.B(n_44),
.Y(n_72)
);

AND2x2_ASAP7_75t_SL g75 ( 
.A(n_48),
.B(n_44),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g92 ( 
.A(n_75),
.B(n_80),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_48),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_78),
.B(n_1),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g96 ( 
.A1(n_79),
.A2(n_66),
.B1(n_45),
.B2(n_49),
.Y(n_96)
);

NAND2x1_ASAP7_75t_SL g80 ( 
.A(n_55),
.B(n_44),
.Y(n_80)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_44),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_69),
.C(n_60),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_57),
.B(n_30),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_89),
.B(n_30),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_66),
.A2(n_30),
.B1(n_22),
.B2(n_21),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_94),
.Y(n_120)
);

BUFx24_ASAP7_75t_SL g94 ( 
.A(n_88),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_71),
.A2(n_49),
.B1(n_56),
.B2(n_50),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_100),
.B1(n_110),
.B2(n_112),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_96),
.A2(n_105),
.B1(n_81),
.B2(n_80),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_70),
.B(n_61),
.Y(n_97)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_55),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_99),
.B(n_102),
.C(n_113),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_79),
.A2(n_46),
.B1(n_51),
.B2(n_59),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_83),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_101),
.B(n_103),
.Y(n_137)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_75),
.Y(n_104)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_104),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_76),
.B(n_58),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_109),
.B(n_116),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_89),
.A2(n_51),
.B1(n_52),
.B2(n_33),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_74),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g128 ( 
.A(n_111),
.B(n_115),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_88),
.A2(n_33),
.B1(n_28),
.B2(n_24),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_75),
.B(n_38),
.C(n_30),
.Y(n_113)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_114),
.Y(n_134)
);

CKINVDCx14_ASAP7_75t_R g115 ( 
.A(n_83),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_88),
.B(n_22),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_119),
.A2(n_131),
.B1(n_140),
.B2(n_91),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g122 ( 
.A(n_97),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g150 ( 
.A(n_122),
.Y(n_150)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_124),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_95),
.Y(n_124)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_126),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_108),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g166 ( 
.A(n_130),
.B(n_86),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_92),
.A2(n_81),
.B1(n_75),
.B2(n_80),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_106),
.A2(n_81),
.B1(n_73),
.B2(n_91),
.Y(n_132)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_132),
.Y(n_143)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_92),
.A2(n_85),
.B(n_82),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g148 ( 
.A1(n_133),
.A2(n_136),
.B(n_138),
.Y(n_148)
);

MAJx2_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_106),
.C(n_116),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_135),
.B(n_102),
.C(n_112),
.Y(n_149)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_21),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_SL g138 ( 
.A1(n_92),
.A2(n_85),
.B(n_82),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_104),
.A2(n_73),
.B(n_87),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_139),
.A2(n_142),
.B(n_98),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_100),
.A2(n_91),
.B1(n_84),
.B2(n_87),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_109),
.B(n_113),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_141),
.B(n_28),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_98),
.A2(n_22),
.B(n_21),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_134),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_145),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_137),
.Y(n_145)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_147),
.B(n_152),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_149),
.B(n_151),
.C(n_162),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_129),
.B(n_110),
.C(n_111),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_132),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_123),
.B(n_103),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_153),
.B(n_154),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_127),
.B(n_101),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g188 ( 
.A1(n_155),
.A2(n_169),
.B(n_125),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_157),
.A2(n_122),
.B1(n_117),
.B2(n_136),
.Y(n_176)
);

NOR2x1_ASAP7_75t_L g158 ( 
.A(n_133),
.B(n_22),
.Y(n_158)
);

NOR2x1_ASAP7_75t_L g179 ( 
.A(n_158),
.B(n_136),
.Y(n_179)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_159),
.B(n_161),
.Y(n_174)
);

FAx1_ASAP7_75t_SL g160 ( 
.A(n_129),
.B(n_33),
.CI(n_28),
.CON(n_160),
.SN(n_160)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_160),
.B(n_167),
.Y(n_184)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_126),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_135),
.B(n_84),
.C(n_77),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g189 ( 
.A(n_163),
.B(n_168),
.C(n_1),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_139),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_164),
.Y(n_190)
);

BUFx24_ASAP7_75t_SL g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_165),
.Y(n_171)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_166),
.Y(n_181)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_131),
.B(n_86),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g169 ( 
.A1(n_138),
.A2(n_77),
.B(n_2),
.Y(n_169)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_180),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_176),
.A2(n_148),
.B1(n_155),
.B2(n_169),
.Y(n_196)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_146),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_177),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_179),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g180 ( 
.A(n_154),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_118),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_182),
.B(n_183),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_R g183 ( 
.A1(n_158),
.A2(n_121),
.B1(n_120),
.B2(n_118),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_162),
.B(n_121),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_185),
.B(n_189),
.C(n_151),
.Y(n_206)
);

AND2x2_ASAP7_75t_L g186 ( 
.A(n_149),
.B(n_142),
.Y(n_186)
);

AOI21xp5_ASAP7_75t_L g214 ( 
.A1(n_186),
.A2(n_191),
.B(n_9),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_188),
.A2(n_143),
.B(n_152),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_148),
.A2(n_2),
.B(n_3),
.Y(n_191)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_143),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_192),
.A2(n_159),
.B1(n_147),
.B2(n_167),
.Y(n_200)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_153),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_170),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_145),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_194),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_SL g217 ( 
.A(n_196),
.B(n_199),
.C(n_204),
.Y(n_217)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_200),
.Y(n_223)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_174),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_202),
.B(n_207),
.Y(n_226)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_203),
.Y(n_224)
);

MAJx2_ASAP7_75t_L g204 ( 
.A(n_182),
.B(n_163),
.C(n_160),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_185),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_178),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_190),
.A2(n_150),
.B1(n_160),
.B2(n_161),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g221 ( 
.A(n_208),
.B(n_214),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_146),
.B1(n_6),
.B2(n_7),
.Y(n_209)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_209),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_175),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_210),
.A2(n_211),
.B1(n_181),
.B2(n_173),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_180),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_170),
.B(n_8),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_213),
.Y(n_233)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_SL g219 ( 
.A(n_215),
.B(n_192),
.Y(n_219)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_179),
.B(n_9),
.Y(n_216)
);

AND2x2_ASAP7_75t_SL g220 ( 
.A(n_216),
.B(n_191),
.Y(n_220)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_219),
.Y(n_239)
);

BUFx12f_ASAP7_75t_SL g237 ( 
.A(n_220),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g222 ( 
.A(n_201),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_197),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_198),
.B(n_184),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_225),
.B(n_213),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_177),
.Y(n_227)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_227),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_228),
.B(n_230),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_195),
.B(n_172),
.Y(n_230)
);

INVxp67_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_205),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_195),
.B(n_172),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_206),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_204),
.B(n_189),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_234),
.B(n_188),
.C(n_208),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g236 ( 
.A(n_226),
.B(n_200),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_236),
.A2(n_244),
.B(n_246),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_238),
.B(n_234),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_240),
.Y(n_250)
);

AOI31xp67_ASAP7_75t_L g241 ( 
.A1(n_220),
.A2(n_199),
.A3(n_212),
.B(n_203),
.Y(n_241)
);

HAxp5_ASAP7_75t_SL g252 ( 
.A(n_241),
.B(n_224),
.CON(n_252),
.SN(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_242),
.B(n_243),
.C(n_230),
.Y(n_254)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_248),
.B(n_214),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_231),
.B(n_201),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_237),
.A2(n_223),
.B1(n_229),
.B2(n_220),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_238),
.B(n_232),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_251),
.B(n_242),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g266 ( 
.A(n_252),
.B(n_260),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_253),
.B(n_186),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_254),
.B(n_257),
.C(n_235),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_239),
.B(n_233),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_255),
.B(n_10),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_217),
.C(n_228),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_237),
.A2(n_217),
.B1(n_216),
.B2(n_186),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_258),
.A2(n_216),
.B1(n_245),
.B2(n_187),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g268 ( 
.A1(n_259),
.A2(n_211),
.B(n_210),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_241),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_261),
.B(n_268),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_250),
.B(n_256),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_269),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_266),
.B(n_260),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_272),
.B(n_273),
.C(n_276),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_253),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_262),
.B(n_257),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_275),
.B(n_266),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_249),
.Y(n_276)
);

NOR2xp67_ASAP7_75t_SL g277 ( 
.A(n_274),
.B(n_254),
.Y(n_277)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_277),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_278),
.A2(n_280),
.B(n_10),
.Y(n_283)
);

AO21x1_ASAP7_75t_SL g280 ( 
.A1(n_272),
.A2(n_252),
.B(n_270),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_171),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_281),
.B(n_16),
.C(n_13),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_283),
.B(n_284),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g286 ( 
.A(n_282),
.Y(n_286)
);

OAI321xp33_ASAP7_75t_L g287 ( 
.A1(n_286),
.A2(n_279),
.A3(n_14),
.B1(n_15),
.B2(n_16),
.C(n_12),
.Y(n_287)
);

OAI22xp33_ASAP7_75t_SL g288 ( 
.A1(n_287),
.A2(n_285),
.B1(n_14),
.B2(n_15),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_12),
.B1(n_15),
.B2(n_16),
.Y(n_289)
);

BUFx24_ASAP7_75t_SL g290 ( 
.A(n_289),
.Y(n_290)
);


endmodule