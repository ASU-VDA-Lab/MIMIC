module real_aes_9411_n_267 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_267);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_267;
wire n_476;
wire n_887;
wire n_599;
wire n_1279;
wire n_1314;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_503;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_571;
wire n_549;
wire n_1034;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_271;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1520;
wire n_1453;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_281;
wire n_962;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1224;
wire n_688;
wire n_1042;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_619;
wire n_1250;
wire n_1095;
wire n_1284;
wire n_360;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_488;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_1073;
wire n_404;
wire n_1301;
wire n_728;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1542;
wire n_1392;
wire n_665;
wire n_991;
wire n_667;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_278;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_277;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_676;
wire n_658;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_645;
wire n_1145;
wire n_1529;
wire n_557;
wire n_777;
wire n_985;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_720;
wire n_354;
wire n_1026;
wire n_492;
wire n_407;
wire n_1023;
wire n_419;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_268;
wire n_1194;
wire n_282;
wire n_389;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_679;
wire n_520;
wire n_926;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_1524;
wire n_762;
wire n_325;
wire n_1298;
wire n_442;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_1172;
wire n_459;
wire n_998;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_279;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_1185;
wire n_661;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_778;
wire n_1175;
wire n_1170;
wire n_522;
wire n_1475;
wire n_943;
wire n_977;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1113;
wire n_1268;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_274;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_273;
wire n_1482;
wire n_1038;
wire n_276;
wire n_1085;
wire n_295;
wire n_845;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1143;
wire n_929;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_650;
wire n_1211;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_1061;
wire n_849;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1381;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_280;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_372;
wire n_578;
wire n_938;
wire n_327;
wire n_774;
wire n_559;
wire n_1049;
wire n_466;
wire n_1277;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_1025;
wire n_532;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_879;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_269;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_275;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_272;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_270;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
INVxp33_ASAP7_75t_L g319 ( .A(n_0), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_0), .A2(n_40), .B1(n_420), .B2(n_425), .Y(n_419) );
INVx1_ASAP7_75t_L g1303 ( .A(n_1), .Y(n_1303) );
CKINVDCx5p33_ASAP7_75t_R g820 ( .A(n_2), .Y(n_820) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_3), .A2(n_242), .B1(n_426), .B2(n_539), .Y(n_1045) );
INVxp33_ASAP7_75t_L g1066 ( .A(n_3), .Y(n_1066) );
INVx1_ASAP7_75t_L g1089 ( .A(n_4), .Y(n_1089) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_5), .A2(n_191), .B1(n_894), .B2(n_1100), .Y(n_1160) );
AOI221xp5_ASAP7_75t_L g1186 ( .A1(n_5), .A2(n_141), .B1(n_321), .B2(n_356), .C(n_1187), .Y(n_1186) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_6), .Y(n_281) );
AND2x2_ASAP7_75t_L g306 ( .A(n_6), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_6), .B(n_216), .Y(n_335) );
INVx1_ASAP7_75t_L g387 ( .A(n_6), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_7), .Y(n_994) );
AOI22xp33_ASAP7_75t_L g1112 ( .A1(n_8), .A2(n_17), .B1(n_685), .B2(n_899), .Y(n_1112) );
INVx1_ASAP7_75t_L g1138 ( .A(n_8), .Y(n_1138) );
OA22x2_ASAP7_75t_L g1192 ( .A1(n_9), .A2(n_1193), .B1(n_1247), .B2(n_1248), .Y(n_1192) );
INVxp67_ASAP7_75t_SL g1248 ( .A(n_9), .Y(n_1248) );
INVxp67_ASAP7_75t_L g354 ( .A(n_10), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g451 ( .A1(n_10), .A2(n_91), .B1(n_425), .B2(n_452), .Y(n_451) );
OAI221xp5_ASAP7_75t_SL g791 ( .A1(n_11), .A2(n_66), .B1(n_792), .B2(n_794), .C(n_795), .Y(n_791) );
AOI221xp5_ASAP7_75t_L g823 ( .A1(n_11), .A2(n_111), .B1(n_416), .B2(n_824), .C(n_828), .Y(n_823) );
INVx1_ASAP7_75t_L g813 ( .A(n_12), .Y(n_813) );
INVx1_ASAP7_75t_L g1526 ( .A(n_13), .Y(n_1526) );
AOI22xp33_ASAP7_75t_L g1169 ( .A1(n_14), .A2(n_110), .B1(n_426), .B2(n_890), .Y(n_1169) );
INVx1_ASAP7_75t_L g1179 ( .A(n_14), .Y(n_1179) );
OAI332xp33_ASAP7_75t_L g1202 ( .A1(n_15), .A2(n_343), .A3(n_383), .B1(n_1203), .B2(n_1206), .B3(n_1210), .C1(n_1215), .C2(n_1218), .Y(n_1202) );
INVx1_ASAP7_75t_L g1243 ( .A(n_15), .Y(n_1243) );
INVx1_ASAP7_75t_L g854 ( .A(n_16), .Y(n_854) );
AOI221xp5_ASAP7_75t_L g1132 ( .A1(n_17), .A2(n_124), .B1(n_1133), .B2(n_1135), .C(n_1137), .Y(n_1132) );
INVx1_ASAP7_75t_L g1349 ( .A(n_18), .Y(n_1349) );
INVx1_ASAP7_75t_L g811 ( .A(n_19), .Y(n_811) );
INVx1_ASAP7_75t_L g626 ( .A(n_20), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_21), .A2(n_114), .B1(n_571), .B2(n_573), .Y(n_570) );
INVxp67_ASAP7_75t_SL g601 ( .A(n_21), .Y(n_601) );
INVxp33_ASAP7_75t_L g739 ( .A(n_22), .Y(n_739) );
AOI221xp5_ASAP7_75t_L g777 ( .A1(n_22), .A2(n_149), .B1(n_445), .B2(n_778), .C(n_779), .Y(n_777) );
INVx1_ASAP7_75t_L g577 ( .A(n_23), .Y(n_577) );
AOI22xp5_ASAP7_75t_L g900 ( .A1(n_24), .A2(n_238), .B1(n_901), .B2(n_902), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g960 ( .A1(n_24), .A2(n_238), .B1(n_961), .B2(n_963), .Y(n_960) );
AO221x2_ASAP7_75t_L g1293 ( .A1(n_25), .A2(n_70), .B1(n_1265), .B2(n_1273), .C(n_1294), .Y(n_1293) );
CKINVDCx5p33_ASAP7_75t_R g978 ( .A(n_26), .Y(n_978) );
INVx1_ASAP7_75t_L g1283 ( .A(n_27), .Y(n_1283) );
INVx2_ASAP7_75t_L g400 ( .A(n_28), .Y(n_400) );
OR2x2_ASAP7_75t_L g431 ( .A(n_28), .B(n_398), .Y(n_431) );
OAI22xp5_ASAP7_75t_L g619 ( .A1(n_29), .A2(n_115), .B1(n_564), .B2(n_620), .Y(n_619) );
OAI221xp5_ASAP7_75t_L g658 ( .A1(n_29), .A2(n_115), .B1(n_327), .B2(n_590), .C(n_659), .Y(n_658) );
INVx1_ASAP7_75t_L g784 ( .A(n_30), .Y(n_784) );
INVx1_ASAP7_75t_L g488 ( .A(n_31), .Y(n_488) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_32), .A2(n_54), .B1(n_684), .B2(n_685), .C(n_686), .Y(n_683) );
INVx1_ASAP7_75t_L g725 ( .A(n_32), .Y(n_725) );
OAI221xp5_ASAP7_75t_L g799 ( .A1(n_33), .A2(n_81), .B1(n_340), .B2(n_800), .C(n_801), .Y(n_799) );
OAI22xp5_ASAP7_75t_L g834 ( .A1(n_33), .A2(n_81), .B1(n_564), .B2(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g575 ( .A(n_34), .Y(n_575) );
AOI22xp33_ASAP7_75t_SL g560 ( .A1(n_35), .A2(n_146), .B1(n_425), .B2(n_561), .Y(n_560) );
INVxp33_ASAP7_75t_SL g588 ( .A(n_35), .Y(n_588) );
INVx1_ASAP7_75t_L g305 ( .A(n_36), .Y(n_305) );
OR2x2_ASAP7_75t_L g334 ( .A(n_36), .B(n_335), .Y(n_334) );
BUFx2_ASAP7_75t_L g346 ( .A(n_36), .Y(n_346) );
BUFx2_ASAP7_75t_L g394 ( .A(n_36), .Y(n_394) );
CKINVDCx5p33_ASAP7_75t_R g1002 ( .A(n_37), .Y(n_1002) );
CKINVDCx5p33_ASAP7_75t_R g1205 ( .A(n_38), .Y(n_1205) );
INVx1_ASAP7_75t_L g1347 ( .A(n_39), .Y(n_1347) );
INVxp33_ASAP7_75t_L g298 ( .A(n_40), .Y(n_298) );
INVx1_ASAP7_75t_L g643 ( .A(n_41), .Y(n_643) );
INVx1_ASAP7_75t_L g985 ( .A(n_42), .Y(n_985) );
AOI221xp5_ASAP7_75t_SL g1008 ( .A1(n_42), .A2(n_168), .B1(n_448), .B2(n_1009), .C(n_1011), .Y(n_1008) );
OAI22xp5_ASAP7_75t_L g1146 ( .A1(n_43), .A2(n_159), .B1(n_1023), .B2(n_1147), .Y(n_1146) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_43), .A2(n_148), .B1(n_500), .B2(n_723), .Y(n_1185) );
AOI221xp5_ASAP7_75t_L g1111 ( .A1(n_44), .A2(n_124), .B1(n_444), .B2(n_448), .C(n_635), .Y(n_1111) );
INVx1_ASAP7_75t_L g1139 ( .A(n_44), .Y(n_1139) );
INVx1_ASAP7_75t_L g979 ( .A(n_45), .Y(n_979) );
AOI221xp5_ASAP7_75t_L g1021 ( .A1(n_45), .A2(n_158), .B1(n_1022), .B2(n_1024), .C(n_1025), .Y(n_1021) );
INVxp67_ASAP7_75t_SL g804 ( .A(n_46), .Y(n_804) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_46), .A2(n_166), .B1(n_842), .B2(n_843), .Y(n_841) );
CKINVDCx16_ASAP7_75t_R g1094 ( .A(n_47), .Y(n_1094) );
INVx1_ASAP7_75t_L g1343 ( .A(n_48), .Y(n_1343) );
OAI221xp5_ASAP7_75t_SL g1042 ( .A1(n_49), .A2(n_235), .B1(n_519), .B2(n_564), .C(n_1043), .Y(n_1042) );
OAI221xp5_ASAP7_75t_L g1071 ( .A1(n_49), .A2(n_235), .B1(n_337), .B2(n_800), .C(n_1072), .Y(n_1071) );
INVx1_ASAP7_75t_L g757 ( .A(n_50), .Y(n_757) );
CKINVDCx5p33_ASAP7_75t_R g1038 ( .A(n_51), .Y(n_1038) );
OAI22xp33_ASAP7_75t_R g1528 ( .A1(n_52), .A2(n_251), .B1(n_564), .B2(n_1019), .Y(n_1528) );
OAI221xp5_ASAP7_75t_L g1545 ( .A1(n_52), .A2(n_251), .B1(n_340), .B2(n_800), .C(n_801), .Y(n_1545) );
AOI221xp5_ASAP7_75t_L g1049 ( .A1(n_53), .A2(n_153), .B1(n_1050), .B2(n_1052), .C(n_1055), .Y(n_1049) );
INVxp67_ASAP7_75t_SL g1080 ( .A(n_53), .Y(n_1080) );
INVx1_ASAP7_75t_L g728 ( .A(n_54), .Y(n_728) );
INVx1_ASAP7_75t_L g705 ( .A(n_55), .Y(n_705) );
CKINVDCx5p33_ASAP7_75t_R g976 ( .A(n_56), .Y(n_976) );
INVx1_ASAP7_75t_L g578 ( .A(n_57), .Y(n_578) );
INVx1_ASAP7_75t_L g989 ( .A(n_58), .Y(n_989) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_58), .A2(n_67), .B1(n_1014), .B2(n_1015), .Y(n_1013) );
INVx1_ASAP7_75t_L g1537 ( .A(n_59), .Y(n_1537) );
INVx1_ASAP7_75t_L g1517 ( .A(n_60), .Y(n_1517) );
AOI22xp33_ASAP7_75t_L g636 ( .A1(n_61), .A2(n_208), .B1(n_637), .B2(n_639), .Y(n_636) );
INVxp67_ASAP7_75t_SL g649 ( .A(n_61), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_62), .A2(n_105), .B1(n_499), .B2(n_502), .Y(n_498) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_62), .A2(n_201), .B1(n_425), .B2(n_541), .Y(n_540) );
AOI221xp5_ASAP7_75t_SL g1108 ( .A1(n_63), .A2(n_83), .B1(n_413), .B2(n_416), .C(n_535), .Y(n_1108) );
INVx1_ASAP7_75t_L g1123 ( .A(n_63), .Y(n_1123) );
INVx1_ASAP7_75t_L g1295 ( .A(n_64), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g888 ( .A1(n_65), .A2(n_85), .B1(n_889), .B2(n_891), .Y(n_888) );
INVxp67_ASAP7_75t_L g946 ( .A(n_65), .Y(n_946) );
AOI22xp33_ASAP7_75t_L g830 ( .A1(n_66), .A2(n_131), .B1(n_685), .B2(n_831), .Y(n_830) );
INVx1_ASAP7_75t_L g983 ( .A(n_67), .Y(n_983) );
INVx1_ASAP7_75t_L g633 ( .A(n_68), .Y(n_633) );
INVx1_ASAP7_75t_L g1105 ( .A(n_69), .Y(n_1105) );
INVx1_ASAP7_75t_L g1104 ( .A(n_71), .Y(n_1104) );
CKINVDCx5p33_ASAP7_75t_R g1214 ( .A(n_72), .Y(n_1214) );
INVx1_ASAP7_75t_L g1048 ( .A(n_73), .Y(n_1048) );
INVxp33_ASAP7_75t_SL g806 ( .A(n_74), .Y(n_806) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_74), .A2(n_227), .B1(n_838), .B2(n_839), .C(n_840), .Y(n_837) );
AOI221xp5_ASAP7_75t_L g1519 ( .A1(n_75), .A2(n_144), .B1(n_889), .B2(n_1520), .C(n_1522), .Y(n_1519) );
INVxp33_ASAP7_75t_L g1542 ( .A(n_75), .Y(n_1542) );
INVx1_ASAP7_75t_L g1358 ( .A(n_76), .Y(n_1358) );
AOI221xp5_ASAP7_75t_L g621 ( .A1(n_77), .A2(n_233), .B1(n_573), .B2(n_622), .C(n_624), .Y(n_621) );
INVxp33_ASAP7_75t_L g665 ( .A(n_77), .Y(n_665) );
CKINVDCx16_ASAP7_75t_R g1361 ( .A(n_78), .Y(n_1361) );
INVx1_ASAP7_75t_L g615 ( .A(n_79), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g1195 ( .A1(n_80), .A2(n_213), .B1(n_1196), .B2(n_1197), .Y(n_1195) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_80), .Y(n_1241) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_82), .Y(n_1151) );
INVx1_ASAP7_75t_L g1122 ( .A(n_83), .Y(n_1122) );
INVxp67_ASAP7_75t_L g348 ( .A(n_84), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g443 ( .A1(n_84), .A2(n_186), .B1(n_444), .B2(n_445), .C(n_448), .Y(n_443) );
INVxp67_ASAP7_75t_L g943 ( .A(n_85), .Y(n_943) );
XOR2x2_ASAP7_75t_L g1142 ( .A(n_86), .B(n_1143), .Y(n_1142) );
INVx1_ASAP7_75t_L g1304 ( .A(n_87), .Y(n_1304) );
AOI22xp33_ASAP7_75t_L g1534 ( .A1(n_88), .A2(n_244), .B1(n_828), .B2(n_1535), .Y(n_1534) );
INVxp67_ASAP7_75t_SL g1554 ( .A(n_88), .Y(n_1554) );
OAI221xp5_ASAP7_75t_L g1098 ( .A1(n_89), .A2(n_226), .B1(n_1027), .B2(n_1099), .C(n_1102), .Y(n_1098) );
INVx1_ASAP7_75t_L g1130 ( .A(n_89), .Y(n_1130) );
OAI22xp5_ASAP7_75t_L g1198 ( .A1(n_90), .A2(n_150), .B1(n_391), .B2(n_1199), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g1239 ( .A(n_90), .Y(n_1239) );
INVxp67_ASAP7_75t_L g360 ( .A(n_91), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g1363 ( .A(n_92), .Y(n_1363) );
OA22x2_ASAP7_75t_L g1509 ( .A1(n_92), .A2(n_1363), .B1(n_1510), .B2(n_1511), .Y(n_1509) );
AOI22xp33_ASAP7_75t_L g1562 ( .A1(n_92), .A2(n_1563), .B1(n_1567), .B2(n_1570), .Y(n_1562) );
INVx1_ASAP7_75t_L g1062 ( .A(n_93), .Y(n_1062) );
AOI22xp5_ASAP7_75t_L g1286 ( .A1(n_94), .A2(n_145), .B1(n_1287), .B2(n_1290), .Y(n_1286) );
INVx1_ASAP7_75t_L g398 ( .A(n_95), .Y(n_398) );
INVx1_ASAP7_75t_L g418 ( .A(n_95), .Y(n_418) );
INVx1_ASAP7_75t_L g609 ( .A(n_96), .Y(n_609) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_97), .Y(n_1514) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_98), .Y(n_998) );
INVx1_ASAP7_75t_L g874 ( .A(n_99), .Y(n_874) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_100), .A2(n_264), .B1(n_433), .B2(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g709 ( .A(n_100), .Y(n_709) );
OAI221xp5_ASAP7_75t_L g326 ( .A1(n_101), .A2(n_126), .B1(n_327), .B2(n_336), .C(n_340), .Y(n_326) );
OAI22xp5_ASAP7_75t_L g432 ( .A1(n_101), .A2(n_126), .B1(n_433), .B2(n_438), .Y(n_432) );
INVxp67_ASAP7_75t_SL g748 ( .A(n_102), .Y(n_748) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_102), .A2(n_218), .B1(n_448), .B2(n_635), .C(n_770), .Y(n_772) );
INVx1_ASAP7_75t_L g1103 ( .A(n_103), .Y(n_1103) );
AOI221xp5_ASAP7_75t_L g1125 ( .A1(n_103), .A2(n_226), .B1(n_1126), .B2(n_1128), .C(n_1129), .Y(n_1125) );
INVx1_ASAP7_75t_L g548 ( .A(n_104), .Y(n_548) );
AOI221xp5_ASAP7_75t_L g534 ( .A1(n_105), .A2(n_172), .B1(n_448), .B2(n_535), .C(n_537), .Y(n_534) );
INVxp33_ASAP7_75t_SL g736 ( .A(n_106), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g780 ( .A1(n_106), .A2(n_122), .B1(n_444), .B2(n_781), .Y(n_780) );
AOI22xp33_ASAP7_75t_L g509 ( .A1(n_107), .A2(n_248), .B1(n_502), .B2(n_510), .Y(n_509) );
INVxp67_ASAP7_75t_L g533 ( .A(n_107), .Y(n_533) );
INVxp33_ASAP7_75t_SL g490 ( .A(n_108), .Y(n_490) );
AOI21xp33_ASAP7_75t_L g527 ( .A1(n_108), .A2(n_528), .B(n_529), .Y(n_527) );
INVx1_ASAP7_75t_L g1280 ( .A(n_109), .Y(n_1280) );
OAI211xp5_ASAP7_75t_L g1171 ( .A1(n_110), .A2(n_1172), .B(n_1174), .C(n_1176), .Y(n_1171) );
INVxp33_ASAP7_75t_SL g797 ( .A(n_111), .Y(n_797) );
INVx1_ASAP7_75t_L g1115 ( .A(n_112), .Y(n_1115) );
AO221x2_ASAP7_75t_L g1300 ( .A1(n_113), .A2(n_195), .B1(n_1273), .B2(n_1301), .C(n_1302), .Y(n_1300) );
INVxp33_ASAP7_75t_L g593 ( .A(n_114), .Y(n_593) );
OAI221xp5_ASAP7_75t_L g980 ( .A1(n_116), .A2(n_143), .B1(n_327), .B2(n_590), .C(n_659), .Y(n_980) );
OAI22xp5_ASAP7_75t_L g1018 ( .A1(n_116), .A2(n_143), .B1(n_1019), .B2(n_1020), .Y(n_1018) );
INVx1_ASAP7_75t_L g562 ( .A(n_117), .Y(n_562) );
INVxp33_ASAP7_75t_SL g864 ( .A(n_118), .Y(n_864) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_118), .A2(n_157), .B1(n_510), .B2(n_722), .C(n_932), .Y(n_931) );
INVx1_ASAP7_75t_L g754 ( .A(n_119), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g773 ( .A1(n_119), .A2(n_179), .B1(n_425), .B2(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g1057 ( .A1(n_120), .A2(n_174), .B1(n_1058), .B2(n_1059), .Y(n_1057) );
INVx1_ASAP7_75t_L g1082 ( .A(n_120), .Y(n_1082) );
INVx1_ASAP7_75t_L g273 ( .A(n_121), .Y(n_273) );
INVxp33_ASAP7_75t_SL g740 ( .A(n_122), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g892 ( .A1(n_123), .A2(n_196), .B1(n_893), .B2(n_895), .Y(n_892) );
INVxp67_ASAP7_75t_SL g955 ( .A(n_123), .Y(n_955) );
XNOR2x1_ASAP7_75t_L g293 ( .A(n_125), .B(n_294), .Y(n_293) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_127), .Y(n_478) );
OAI221xp5_ASAP7_75t_L g518 ( .A1(n_127), .A2(n_206), .B1(n_438), .B2(n_519), .C(n_521), .Y(n_518) );
CKINVDCx5p33_ASAP7_75t_R g1166 ( .A(n_128), .Y(n_1166) );
INVx1_ASAP7_75t_L g369 ( .A(n_129), .Y(n_369) );
INVx1_ASAP7_75t_L g695 ( .A(n_130), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g719 ( .A1(n_130), .A2(n_169), .B1(n_720), .B2(n_722), .Y(n_719) );
INVxp33_ASAP7_75t_SL g796 ( .A(n_131), .Y(n_796) );
AOI22xp5_ASAP7_75t_L g1292 ( .A1(n_132), .A2(n_193), .B1(n_1265), .B2(n_1273), .Y(n_1292) );
AOI221xp5_ASAP7_75t_L g1531 ( .A1(n_133), .A2(n_220), .B1(n_1162), .B2(n_1532), .C(n_1533), .Y(n_1531) );
INVxp67_ASAP7_75t_SL g1549 ( .A(n_133), .Y(n_1549) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_134), .A2(n_224), .B1(n_504), .B2(n_507), .Y(n_506) );
INVxp33_ASAP7_75t_L g547 ( .A(n_134), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g701 ( .A1(n_135), .A2(n_249), .B1(n_637), .B2(n_639), .Y(n_701) );
AOI22xp33_ASAP7_75t_L g715 ( .A1(n_135), .A2(n_147), .B1(n_504), .B2(n_605), .Y(n_715) );
INVx1_ASAP7_75t_L g729 ( .A(n_136), .Y(n_729) );
OAI221xp5_ASAP7_75t_L g1201 ( .A1(n_137), .A2(n_231), .B1(n_590), .B2(n_659), .C(n_800), .Y(n_1201) );
OAI222xp33_ASAP7_75t_L g1225 ( .A1(n_137), .A2(n_150), .B1(n_231), .B2(n_1019), .C1(n_1020), .C2(n_1114), .Y(n_1225) );
XNOR2x1_ASAP7_75t_L g969 ( .A(n_138), .B(n_970), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g563 ( .A1(n_139), .A2(n_198), .B1(n_433), .B2(n_564), .Y(n_563) );
OAI221xp5_ASAP7_75t_L g589 ( .A1(n_139), .A2(n_198), .B1(n_327), .B2(n_336), .C(n_590), .Y(n_589) );
CKINVDCx5p33_ASAP7_75t_R g1005 ( .A(n_140), .Y(n_1005) );
AOI21xp33_ASAP7_75t_L g1161 ( .A1(n_141), .A2(n_1162), .B(n_1163), .Y(n_1161) );
INVx1_ASAP7_75t_L g1296 ( .A(n_142), .Y(n_1296) );
INVxp33_ASAP7_75t_L g1544 ( .A(n_144), .Y(n_1544) );
INVxp33_ASAP7_75t_L g583 ( .A(n_146), .Y(n_583) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_147), .A2(n_155), .B1(n_697), .B2(n_699), .C(n_700), .Y(n_696) );
OAI22xp33_ASAP7_75t_L g1148 ( .A1(n_148), .A2(n_161), .B1(n_640), .B2(n_1149), .Y(n_1148) );
INVxp33_ASAP7_75t_L g737 ( .A(n_149), .Y(n_737) );
INVx1_ASAP7_75t_L g380 ( .A(n_151), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_152), .Y(n_1000) );
INVx1_ASAP7_75t_L g1078 ( .A(n_153), .Y(n_1078) );
INVxp33_ASAP7_75t_SL g491 ( .A(n_154), .Y(n_491) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_154), .A2(n_217), .B1(n_426), .B2(n_526), .Y(n_525) );
AOI22xp33_ASAP7_75t_SL g711 ( .A1(n_155), .A2(n_249), .B1(n_500), .B2(n_712), .Y(n_711) );
INVx1_ASAP7_75t_L g704 ( .A(n_156), .Y(n_704) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_156), .A2(n_190), .B1(n_504), .B2(n_717), .Y(n_716) );
INVxp33_ASAP7_75t_SL g859 ( .A(n_157), .Y(n_859) );
INVx1_ASAP7_75t_L g974 ( .A(n_158), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g1183 ( .A1(n_159), .A2(n_161), .B1(n_300), .B2(n_1184), .Y(n_1183) );
AOI21xp5_ASAP7_75t_L g1170 ( .A1(n_160), .A2(n_778), .B(n_779), .Y(n_1170) );
INVx1_ASAP7_75t_L g1177 ( .A(n_160), .Y(n_1177) );
AOI22xp33_ASAP7_75t_SL g897 ( .A1(n_162), .A2(n_170), .B1(n_895), .B2(n_898), .Y(n_897) );
OAI211xp5_ASAP7_75t_SL g920 ( .A1(n_162), .A2(n_921), .B(n_926), .C(n_934), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_163), .A2(n_180), .B1(n_1287), .B2(n_1290), .Y(n_1309) );
INVx1_ASAP7_75t_L g579 ( .A(n_164), .Y(n_579) );
XNOR2xp5_ASAP7_75t_L g849 ( .A(n_165), .B(n_850), .Y(n_849) );
INVxp67_ASAP7_75t_SL g809 ( .A(n_166), .Y(n_809) );
OAI221xp5_ASAP7_75t_L g741 ( .A1(n_167), .A2(n_265), .B1(n_327), .B2(n_337), .C(n_340), .Y(n_741) );
OAI22xp33_ASAP7_75t_L g782 ( .A1(n_167), .A2(n_265), .B1(n_519), .B2(n_783), .Y(n_782) );
INVx1_ASAP7_75t_L g987 ( .A(n_168), .Y(n_987) );
INVx1_ASAP7_75t_L g703 ( .A(n_169), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g939 ( .A1(n_170), .A2(n_940), .B1(n_942), .B2(n_952), .C(n_958), .Y(n_939) );
INVx1_ASAP7_75t_L g1044 ( .A(n_171), .Y(n_1044) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_172), .A2(n_201), .B1(n_504), .B2(n_505), .Y(n_503) );
AOI221xp5_ASAP7_75t_L g634 ( .A1(n_173), .A2(n_255), .B1(n_444), .B2(n_448), .C(n_635), .Y(n_634) );
INVxp33_ASAP7_75t_SL g652 ( .A(n_173), .Y(n_652) );
INVx1_ASAP7_75t_L g1077 ( .A(n_174), .Y(n_1077) );
INVx1_ASAP7_75t_L g731 ( .A(n_175), .Y(n_731) );
INVx1_ASAP7_75t_L g618 ( .A(n_176), .Y(n_618) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_177), .Y(n_275) );
AND3x2_ASAP7_75t_L g1266 ( .A(n_177), .B(n_273), .C(n_1267), .Y(n_1266) );
NAND2xp5_ASAP7_75t_L g1277 ( .A(n_177), .B(n_273), .Y(n_1277) );
CKINVDCx5p33_ASAP7_75t_R g1158 ( .A(n_178), .Y(n_1158) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_179), .Y(n_747) );
AOI22xp5_ASAP7_75t_L g1310 ( .A1(n_181), .A2(n_221), .B1(n_1301), .B2(n_1311), .Y(n_1310) );
OAI221xp5_ASAP7_75t_L g1153 ( .A1(n_182), .A2(n_223), .B1(n_1149), .B2(n_1154), .C(n_1155), .Y(n_1153) );
INVx1_ASAP7_75t_L g1175 ( .A(n_182), .Y(n_1175) );
CKINVDCx5p33_ASAP7_75t_R g1211 ( .A(n_183), .Y(n_1211) );
INVx2_ASAP7_75t_L g286 ( .A(n_184), .Y(n_286) );
XOR2xp5_ASAP7_75t_L g612 ( .A(n_185), .B(n_613), .Y(n_612) );
INVxp33_ASAP7_75t_L g367 ( .A(n_186), .Y(n_367) );
INVx1_ASAP7_75t_L g629 ( .A(n_187), .Y(n_629) );
INVx1_ASAP7_75t_L g1106 ( .A(n_188), .Y(n_1106) );
INVx1_ASAP7_75t_L g815 ( .A(n_189), .Y(n_815) );
INVx1_ASAP7_75t_L g679 ( .A(n_190), .Y(n_679) );
INVx1_ASAP7_75t_L g1188 ( .A(n_191), .Y(n_1188) );
CKINVDCx5p33_ASAP7_75t_R g1216 ( .A(n_192), .Y(n_1216) );
AOI22xp5_ASAP7_75t_L g1328 ( .A1(n_194), .A2(n_203), .B1(n_1265), .B2(n_1273), .Y(n_1328) );
INVxp67_ASAP7_75t_SL g954 ( .A(n_196), .Y(n_954) );
INVx1_ASAP7_75t_L g788 ( .A(n_197), .Y(n_788) );
INVx1_ASAP7_75t_L g372 ( .A(n_199), .Y(n_372) );
INVx1_ASAP7_75t_L g1267 ( .A(n_200), .Y(n_1267) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_202), .A2(n_257), .B1(n_422), .B2(n_448), .C(n_568), .Y(n_567) );
INVxp67_ASAP7_75t_SL g599 ( .A(n_202), .Y(n_599) );
CKINVDCx16_ASAP7_75t_R g1271 ( .A(n_204), .Y(n_1271) );
XNOR2x1_ASAP7_75t_L g472 ( .A(n_205), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g1345 ( .A(n_205), .Y(n_1345) );
INVxp67_ASAP7_75t_SL g482 ( .A(n_206), .Y(n_482) );
INVx1_ASAP7_75t_L g1530 ( .A(n_207), .Y(n_1530) );
INVxp33_ASAP7_75t_L g651 ( .A(n_208), .Y(n_651) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_209), .Y(n_1204) );
INVx1_ASAP7_75t_L g644 ( .A(n_210), .Y(n_644) );
INVx1_ASAP7_75t_L g1524 ( .A(n_211), .Y(n_1524) );
INVx1_ASAP7_75t_L g760 ( .A(n_212), .Y(n_760) );
CKINVDCx5p33_ASAP7_75t_R g1237 ( .A(n_213), .Y(n_1237) );
CKINVDCx5p33_ASAP7_75t_R g1217 ( .A(n_214), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g1568 ( .A1(n_215), .A2(n_1510), .B1(n_1511), .B2(n_1569), .Y(n_1568) );
CKINVDCx5p33_ASAP7_75t_R g1569 ( .A(n_215), .Y(n_1569) );
INVx1_ASAP7_75t_L g288 ( .A(n_216), .Y(n_288) );
INVx2_ASAP7_75t_L g307 ( .A(n_216), .Y(n_307) );
INVxp33_ASAP7_75t_SL g486 ( .A(n_217), .Y(n_486) );
INVxp67_ASAP7_75t_SL g753 ( .A(n_218), .Y(n_753) );
AOI22xp5_ASAP7_75t_L g1327 ( .A1(n_219), .A2(n_243), .B1(n_1287), .B2(n_1290), .Y(n_1327) );
INVxp67_ASAP7_75t_SL g1553 ( .A(n_220), .Y(n_1553) );
INVxp33_ASAP7_75t_L g314 ( .A(n_222), .Y(n_314) );
AOI221xp5_ASAP7_75t_L g409 ( .A1(n_222), .A2(n_225), .B1(n_410), .B2(n_413), .C(n_416), .Y(n_409) );
INVx1_ASAP7_75t_L g1191 ( .A(n_223), .Y(n_1191) );
INVxp67_ASAP7_75t_L g517 ( .A(n_224), .Y(n_517) );
INVxp33_ASAP7_75t_L g308 ( .A(n_225), .Y(n_308) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_227), .Y(n_808) );
INVx1_ASAP7_75t_L g758 ( .A(n_228), .Y(n_758) );
INVx1_ASAP7_75t_L g816 ( .A(n_229), .Y(n_816) );
AOI22xp33_ASAP7_75t_L g1109 ( .A1(n_230), .A2(n_245), .B1(n_561), .B2(n_573), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1119 ( .A1(n_230), .A2(n_245), .B1(n_988), .B2(n_1120), .C(n_1121), .Y(n_1119) );
INVx1_ASAP7_75t_L g868 ( .A(n_232), .Y(n_868) );
INVxp33_ASAP7_75t_L g662 ( .A(n_233), .Y(n_662) );
CKINVDCx5p33_ASAP7_75t_R g1209 ( .A(n_234), .Y(n_1209) );
INVx1_ASAP7_75t_L g1359 ( .A(n_236), .Y(n_1359) );
INVx1_ASAP7_75t_L g376 ( .A(n_237), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g559 ( .A1(n_239), .A2(n_266), .B1(n_410), .B2(n_416), .C(n_452), .Y(n_559) );
INVxp33_ASAP7_75t_L g587 ( .A(n_239), .Y(n_587) );
INVx1_ASAP7_75t_L g1270 ( .A(n_240), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g1282 ( .A(n_240), .B(n_1279), .Y(n_1282) );
AOI21xp33_ASAP7_75t_L g1046 ( .A1(n_241), .A2(n_416), .B(n_691), .Y(n_1046) );
INVxp33_ASAP7_75t_L g1069 ( .A(n_241), .Y(n_1069) );
INVxp33_ASAP7_75t_L g1070 ( .A(n_242), .Y(n_1070) );
INVxp67_ASAP7_75t_SL g1548 ( .A(n_244), .Y(n_1548) );
INVx1_ASAP7_75t_L g880 ( .A(n_246), .Y(n_880) );
CKINVDCx5p33_ASAP7_75t_R g406 ( .A(n_247), .Y(n_406) );
INVxp33_ASAP7_75t_L g546 ( .A(n_248), .Y(n_546) );
INVx1_ASAP7_75t_L g1538 ( .A(n_250), .Y(n_1538) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_252), .A2(n_529), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g727 ( .A(n_252), .Y(n_727) );
INVx2_ASAP7_75t_L g285 ( .A(n_253), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g910 ( .A(n_254), .Y(n_910) );
INVxp67_ASAP7_75t_L g648 ( .A(n_255), .Y(n_648) );
INVx1_ASAP7_75t_L g1061 ( .A(n_256), .Y(n_1061) );
INVxp33_ASAP7_75t_SL g596 ( .A(n_257), .Y(n_596) );
INVx1_ASAP7_75t_L g762 ( .A(n_258), .Y(n_762) );
BUFx3_ASAP7_75t_L g403 ( .A(n_259), .Y(n_403) );
INVx1_ASAP7_75t_L g428 ( .A(n_259), .Y(n_428) );
BUFx3_ASAP7_75t_L g405 ( .A(n_260), .Y(n_405) );
INVx1_ASAP7_75t_L g424 ( .A(n_260), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g1207 ( .A(n_261), .Y(n_1207) );
CKINVDCx20_ASAP7_75t_R g1041 ( .A(n_262), .Y(n_1041) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_263), .Y(n_689) );
INVx1_ASAP7_75t_L g708 ( .A(n_264), .Y(n_708) );
INVxp33_ASAP7_75t_L g585 ( .A(n_266), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_268), .A2(n_289), .B(n_1256), .Y(n_267) );
HB1xp67_ASAP7_75t_L g268 ( .A(n_269), .Y(n_268) );
BUFx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
AND2x4_ASAP7_75t_L g270 ( .A(n_271), .B(n_276), .Y(n_270) );
AND2x4_ASAP7_75t_L g1561 ( .A(n_271), .B(n_277), .Y(n_1561) );
NOR2xp33_ASAP7_75t_SL g271 ( .A(n_272), .B(n_274), .Y(n_271) );
INVx1_ASAP7_75t_SL g1566 ( .A(n_272), .Y(n_1566) );
NAND2xp5_ASAP7_75t_L g1576 ( .A(n_272), .B(n_274), .Y(n_1576) );
HB1xp67_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x2_ASAP7_75t_L g1565 ( .A(n_274), .B(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
INVx1_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
NOR2xp33_ASAP7_75t_L g277 ( .A(n_278), .B(n_282), .Y(n_277) );
INVxp67_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
HB1xp67_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
AND2x2_ASAP7_75t_L g497 ( .A(n_280), .B(n_288), .Y(n_497) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g344 ( .A(n_281), .B(n_345), .Y(n_344) );
OR2x6_ASAP7_75t_L g282 ( .A(n_283), .B(n_287), .Y(n_282) );
INVx2_ASAP7_75t_SL g359 ( .A(n_283), .Y(n_359) );
INVx2_ASAP7_75t_SL g375 ( .A(n_283), .Y(n_375) );
OR2x2_ASAP7_75t_L g391 ( .A(n_283), .B(n_334), .Y(n_391) );
BUFx6f_ASAP7_75t_L g595 ( .A(n_283), .Y(n_595) );
INVx1_ASAP7_75t_L g1076 ( .A(n_283), .Y(n_1076) );
OAI22xp5_ASAP7_75t_L g1187 ( .A1(n_283), .A2(n_363), .B1(n_1158), .B2(n_1188), .Y(n_1187) );
BUFx6f_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AND2x4_ASAP7_75t_L g302 ( .A(n_285), .B(n_303), .Y(n_302) );
INVx1_ASAP7_75t_L g312 ( .A(n_285), .Y(n_312) );
AND2x2_ASAP7_75t_L g318 ( .A(n_285), .B(n_286), .Y(n_318) );
INVx2_ASAP7_75t_L g323 ( .A(n_285), .Y(n_323) );
INVx1_ASAP7_75t_L g366 ( .A(n_285), .Y(n_366) );
INVx2_ASAP7_75t_L g303 ( .A(n_286), .Y(n_303) );
INVx1_ASAP7_75t_L g325 ( .A(n_286), .Y(n_325) );
INVx1_ASAP7_75t_L g332 ( .A(n_286), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_286), .B(n_323), .Y(n_353) );
INVx1_ASAP7_75t_L g365 ( .A(n_286), .Y(n_365) );
INVx2_ASAP7_75t_SL g287 ( .A(n_288), .Y(n_287) );
XOR2xp5_ASAP7_75t_L g289 ( .A(n_290), .B(n_669), .Y(n_289) );
OAI22xp33_ASAP7_75t_L g290 ( .A1(n_291), .A2(n_551), .B1(n_552), .B2(n_668), .Y(n_290) );
INVxp67_ASAP7_75t_SL g668 ( .A(n_291), .Y(n_668) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_471), .B1(n_549), .B2(n_550), .Y(n_291) );
BUFx2_ASAP7_75t_SL g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g550 ( .A(n_293), .Y(n_550) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_388), .Y(n_294) );
NOR3xp33_ASAP7_75t_L g295 ( .A(n_296), .B(n_326), .C(n_342), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g296 ( .A(n_297), .B(n_313), .Y(n_296) );
AOI22xp33_ASAP7_75t_L g297 ( .A1(n_298), .A2(n_299), .B1(n_308), .B2(n_309), .Y(n_297) );
BUFx2_ASAP7_75t_L g487 ( .A(n_299), .Y(n_487) );
BUFx2_ASAP7_75t_L g584 ( .A(n_299), .Y(n_584) );
BUFx2_ASAP7_75t_L g663 ( .A(n_299), .Y(n_663) );
AOI22xp33_ASAP7_75t_L g795 ( .A1(n_299), .A2(n_796), .B1(n_797), .B2(n_798), .Y(n_795) );
BUFx2_ASAP7_75t_L g975 ( .A(n_299), .Y(n_975) );
BUFx2_ASAP7_75t_L g1067 ( .A(n_299), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1543 ( .A1(n_299), .A2(n_798), .B1(n_1524), .B2(n_1544), .Y(n_1543) );
AND2x4_ASAP7_75t_L g299 ( .A(n_300), .B(n_304), .Y(n_299) );
BUFx3_ASAP7_75t_L g605 ( .A(n_300), .Y(n_605) );
INVx1_ASAP7_75t_L g656 ( .A(n_300), .Y(n_656) );
INVx3_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx3_ASAP7_75t_L g371 ( .A(n_301), .Y(n_371) );
BUFx6f_ASAP7_75t_L g997 ( .A(n_301), .Y(n_997) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
BUFx6f_ASAP7_75t_L g356 ( .A(n_302), .Y(n_356) );
INVx1_ASAP7_75t_L g951 ( .A(n_302), .Y(n_951) );
AND2x4_ASAP7_75t_L g311 ( .A(n_303), .B(n_312), .Y(n_311) );
AND2x6_ASAP7_75t_L g309 ( .A(n_304), .B(n_310), .Y(n_309) );
AND2x4_ASAP7_75t_L g315 ( .A(n_304), .B(n_316), .Y(n_315) );
AND2x2_ASAP7_75t_L g320 ( .A(n_304), .B(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g492 ( .A(n_304), .B(n_321), .Y(n_492) );
AND2x2_ASAP7_75t_L g666 ( .A(n_304), .B(n_321), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g1118 ( .A1(n_304), .A2(n_512), .B1(n_1119), .B2(n_1125), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_304), .B(n_321), .Y(n_1173) );
AND2x2_ASAP7_75t_L g1178 ( .A(n_304), .B(n_918), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1180 ( .A(n_304), .B(n_371), .Y(n_1180) );
AND2x2_ASAP7_75t_L g1189 ( .A(n_304), .B(n_723), .Y(n_1189) );
AND2x4_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g384 ( .A(n_305), .Y(n_384) );
OR2x2_ASAP7_75t_L g858 ( .A(n_305), .B(n_431), .Y(n_858) );
INVx2_ASAP7_75t_L g924 ( .A(n_306), .Y(n_924) );
AND2x4_ASAP7_75t_L g941 ( .A(n_306), .B(n_501), .Y(n_941) );
AND2x2_ASAP7_75t_L g962 ( .A(n_306), .B(n_322), .Y(n_962) );
INVx1_ASAP7_75t_L g345 ( .A(n_307), .Y(n_345) );
INVx1_ASAP7_75t_L g386 ( .A(n_307), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g485 ( .A1(n_309), .A2(n_486), .B1(n_487), .B2(n_488), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_309), .A2(n_583), .B1(n_584), .B2(n_585), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_309), .A2(n_626), .B1(n_662), .B2(n_663), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g724 ( .A1(n_309), .A2(n_584), .B1(n_689), .B2(n_725), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g735 ( .A1(n_309), .A2(n_584), .B1(n_736), .B2(n_737), .Y(n_735) );
BUFx2_ASAP7_75t_L g798 ( .A(n_309), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g973 ( .A1(n_309), .A2(n_974), .B1(n_975), .B2(n_976), .Y(n_973) );
AOI22xp33_ASAP7_75t_L g1065 ( .A1(n_309), .A2(n_1044), .B1(n_1066), .B2(n_1067), .Y(n_1065) );
INVx1_ASAP7_75t_SL g1197 ( .A(n_309), .Y(n_1197) );
NAND2x1p5_ASAP7_75t_L g341 ( .A(n_310), .B(n_333), .Y(n_341) );
BUFx2_ASAP7_75t_L g502 ( .A(n_310), .Y(n_502) );
BUFx3_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
BUFx2_ASAP7_75t_L g484 ( .A(n_311), .Y(n_484) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_311), .Y(n_714) );
BUFx6f_ASAP7_75t_L g723 ( .A(n_311), .Y(n_723) );
BUFx3_ASAP7_75t_L g925 ( .A(n_311), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g313 ( .A1(n_314), .A2(n_315), .B1(n_319), .B2(n_320), .Y(n_313) );
AOI22xp33_ASAP7_75t_L g489 ( .A1(n_315), .A2(n_490), .B1(n_491), .B2(n_492), .Y(n_489) );
AOI22xp33_ASAP7_75t_L g586 ( .A1(n_315), .A2(n_492), .B1(n_587), .B2(n_588), .Y(n_586) );
AOI22xp33_ASAP7_75t_L g664 ( .A1(n_315), .A2(n_629), .B1(n_665), .B2(n_666), .Y(n_664) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_315), .A2(n_666), .B1(n_727), .B2(n_728), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_315), .A2(n_666), .B1(n_739), .B2(n_740), .Y(n_738) );
BUFx2_ASAP7_75t_L g793 ( .A(n_315), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g977 ( .A1(n_315), .A2(n_320), .B1(n_978), .B2(n_979), .Y(n_977) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_315), .A2(n_492), .B1(n_1069), .B2(n_1070), .Y(n_1068) );
INVx2_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g721 ( .A(n_317), .Y(n_721) );
INVx2_ASAP7_75t_SL g918 ( .A(n_317), .Y(n_918) );
INVx3_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx6f_ASAP7_75t_L g501 ( .A(n_318), .Y(n_501) );
INVx1_ASAP7_75t_L g794 ( .A(n_320), .Y(n_794) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_320), .A2(n_793), .B1(n_1526), .B2(n_1542), .Y(n_1541) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
BUFx2_ASAP7_75t_L g504 ( .A(n_322), .Y(n_504) );
INVx1_ASAP7_75t_L g1127 ( .A(n_322), .Y(n_1127) );
INVx1_ASAP7_75t_L g1134 ( .A(n_322), .Y(n_1134) );
BUFx6f_ASAP7_75t_L g1184 ( .A(n_322), .Y(n_1184) );
AND2x4_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx1_ASAP7_75t_L g339 ( .A(n_323), .Y(n_339) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx2_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx2_ASAP7_75t_L g800 ( .A(n_328), .Y(n_800) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
NAND2x1_ASAP7_75t_SL g329 ( .A(n_330), .B(n_333), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
HB1xp67_ASAP7_75t_L g477 ( .A(n_332), .Y(n_477) );
NAND2x1p5_ASAP7_75t_L g337 ( .A(n_333), .B(n_338), .Y(n_337) );
AND2x4_ASAP7_75t_L g476 ( .A(n_333), .B(n_477), .Y(n_476) );
AND2x4_ASAP7_75t_L g479 ( .A(n_333), .B(n_480), .Y(n_479) );
AND2x4_ASAP7_75t_L g483 ( .A(n_333), .B(n_484), .Y(n_483) );
INVx3_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g917 ( .A(n_335), .Y(n_917) );
BUFx4f_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
BUFx4f_ASAP7_75t_L g659 ( .A(n_337), .Y(n_659) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
OR2x6_ASAP7_75t_L g938 ( .A(n_339), .B(n_916), .Y(n_938) );
BUFx2_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
BUFx3_ASAP7_75t_L g590 ( .A(n_341), .Y(n_590) );
BUFx2_ASAP7_75t_L g1072 ( .A(n_341), .Y(n_1072) );
OAI33xp33_ASAP7_75t_L g342 ( .A1(n_343), .A2(n_347), .A3(n_357), .B1(n_368), .B2(n_373), .B3(n_381), .Y(n_342) );
OAI33xp33_ASAP7_75t_L g591 ( .A1(n_343), .A2(n_381), .A3(n_592), .B1(n_598), .B2(n_603), .B3(n_606), .Y(n_591) );
OAI33xp33_ASAP7_75t_L g646 ( .A1(n_343), .A2(n_381), .A3(n_647), .B1(n_650), .B2(n_655), .B3(n_657), .Y(n_646) );
HB1xp67_ASAP7_75t_L g743 ( .A(n_343), .Y(n_743) );
OAI33xp33_ASAP7_75t_L g802 ( .A1(n_343), .A2(n_803), .A3(n_807), .B1(n_810), .B2(n_814), .B3(n_817), .Y(n_802) );
OAI33xp33_ASAP7_75t_L g981 ( .A1(n_343), .A2(n_381), .A3(n_982), .B1(n_986), .B2(n_991), .B3(n_999), .Y(n_981) );
OAI33xp33_ASAP7_75t_L g1073 ( .A1(n_343), .A2(n_381), .A3(n_1074), .B1(n_1079), .B2(n_1083), .B3(n_1086), .Y(n_1073) );
OAI33xp33_ASAP7_75t_L g1546 ( .A1(n_343), .A2(n_1547), .A3(n_1550), .B1(n_1555), .B2(n_1556), .B3(n_1557), .Y(n_1546) );
OR2x6_ASAP7_75t_L g343 ( .A(n_344), .B(n_346), .Y(n_343) );
BUFx2_ASAP7_75t_L g470 ( .A(n_346), .Y(n_470) );
INVx2_ASAP7_75t_L g496 ( .A(n_346), .Y(n_496) );
OAI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_349), .B1(n_354), .B2(n_355), .Y(n_347) );
OAI22xp5_ASAP7_75t_L g368 ( .A1(n_349), .A2(n_369), .B1(n_370), .B2(n_372), .Y(n_368) );
OAI22xp5_ASAP7_75t_L g647 ( .A1(n_349), .A2(n_604), .B1(n_648), .B2(n_649), .Y(n_647) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx2_ASAP7_75t_L g600 ( .A(n_350), .Y(n_600) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g756 ( .A(n_351), .Y(n_756) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
BUFx3_ASAP7_75t_L g930 ( .A(n_352), .Y(n_930) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g752 ( .A(n_353), .Y(n_752) );
BUFx2_ASAP7_75t_L g993 ( .A(n_353), .Y(n_993) );
OAI22xp5_ASAP7_75t_L g749 ( .A1(n_355), .A2(n_750), .B1(n_753), .B2(n_754), .Y(n_749) );
OAI22xp5_ASAP7_75t_L g755 ( .A1(n_355), .A2(n_756), .B1(n_757), .B2(n_758), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g1203 ( .A1(n_355), .A2(n_929), .B1(n_1204), .B2(n_1205), .Y(n_1203) );
INVx4_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
BUFx3_ASAP7_75t_L g505 ( .A(n_356), .Y(n_505) );
INVx2_ASAP7_75t_SL g602 ( .A(n_356), .Y(n_602) );
INVx2_ASAP7_75t_SL g1120 ( .A(n_356), .Y(n_1120) );
INVx2_ASAP7_75t_SL g1136 ( .A(n_356), .Y(n_1136) );
OAI22xp33_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_360), .B1(n_361), .B2(n_367), .Y(n_357) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_358), .A2(n_953), .B1(n_954), .B2(n_955), .C(n_956), .Y(n_952) );
BUFx2_ASAP7_75t_L g984 ( .A(n_358), .Y(n_984) );
OAI22xp33_ASAP7_75t_L g1547 ( .A1(n_358), .A2(n_761), .B1(n_1548), .B2(n_1549), .Y(n_1547) );
OAI22xp33_ASAP7_75t_L g1555 ( .A1(n_358), .A2(n_944), .B1(n_1517), .B2(n_1537), .Y(n_1555) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g761 ( .A(n_362), .Y(n_761) );
INVx2_ASAP7_75t_L g1001 ( .A(n_362), .Y(n_1001) );
INVx2_ASAP7_75t_L g362 ( .A(n_363), .Y(n_362) );
BUFx3_ASAP7_75t_L g805 ( .A(n_363), .Y(n_805) );
BUFx6f_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g379 ( .A(n_365), .B(n_366), .Y(n_379) );
INVx1_ASAP7_75t_L g481 ( .A(n_366), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g408 ( .A1(n_369), .A2(n_409), .B1(n_419), .B2(n_429), .C(n_432), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_370), .A2(n_1211), .B1(n_1212), .B2(n_1214), .Y(n_1210) );
INVx2_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g508 ( .A(n_371), .Y(n_508) );
INVx2_ASAP7_75t_L g718 ( .A(n_371), .Y(n_718) );
INVx2_ASAP7_75t_L g1085 ( .A(n_371), .Y(n_1085) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_372), .A2(n_376), .B1(n_460), .B2(n_465), .Y(n_459) );
OAI22xp33_ASAP7_75t_L g373 ( .A1(n_374), .A2(n_376), .B1(n_377), .B2(n_380), .Y(n_373) );
OAI22xp33_ASAP7_75t_L g657 ( .A1(n_374), .A2(n_377), .B1(n_633), .B2(n_643), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g803 ( .A1(n_374), .A2(n_804), .B1(n_805), .B2(n_806), .Y(n_803) );
OAI22xp33_ASAP7_75t_L g814 ( .A1(n_374), .A2(n_805), .B1(n_815), .B2(n_816), .Y(n_814) );
INVx3_ASAP7_75t_L g374 ( .A(n_375), .Y(n_374) );
OAI22xp33_ASAP7_75t_L g744 ( .A1(n_377), .A2(n_745), .B1(n_747), .B2(n_748), .Y(n_744) );
OAI22xp33_ASAP7_75t_L g1086 ( .A1(n_377), .A2(n_1048), .B1(n_1061), .B2(n_1087), .Y(n_1086) );
BUFx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g654 ( .A(n_378), .Y(n_654) );
OAI22xp33_ASAP7_75t_L g1129 ( .A1(n_378), .A2(n_595), .B1(n_1104), .B2(n_1130), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1137 ( .A1(n_378), .A2(n_595), .B1(n_1138), .B2(n_1139), .Y(n_1137) );
INVx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx2_ASAP7_75t_L g597 ( .A(n_379), .Y(n_597) );
BUFx2_ASAP7_75t_L g608 ( .A(n_379), .Y(n_608) );
INVx2_ASAP7_75t_L g959 ( .A(n_379), .Y(n_959) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_380), .A2(n_443), .B1(n_451), .B2(n_454), .C(n_456), .Y(n_442) );
OAI33xp33_ASAP7_75t_L g742 ( .A1(n_381), .A2(n_743), .A3(n_744), .B1(n_749), .B2(n_755), .B3(n_759), .Y(n_742) );
INVx1_ASAP7_75t_L g818 ( .A(n_381), .Y(n_818) );
CKINVDCx8_ASAP7_75t_R g381 ( .A(n_382), .Y(n_381) );
INVx5_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx6_ASAP7_75t_L g512 ( .A(n_383), .Y(n_512) );
OR2x6_ASAP7_75t_L g383 ( .A(n_384), .B(n_385), .Y(n_383) );
NAND2x1p5_ASAP7_75t_L g879 ( .A(n_384), .B(n_396), .Y(n_879) );
INVx2_ASAP7_75t_L g933 ( .A(n_385), .Y(n_933) );
NAND2x1p5_ASAP7_75t_L g385 ( .A(n_386), .B(n_387), .Y(n_385) );
AOI21xp33_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_406), .B(n_407), .Y(n_388) );
AOI22xp5_ASAP7_75t_L g513 ( .A1(n_389), .A2(n_514), .B1(n_515), .B2(n_548), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_389), .A2(n_514), .B1(n_557), .B2(n_579), .Y(n_556) );
AOI21xp33_ASAP7_75t_L g614 ( .A1(n_389), .A2(n_615), .B(n_616), .Y(n_614) );
AOI22xp5_ASAP7_75t_L g675 ( .A1(n_389), .A2(n_676), .B1(n_677), .B2(n_705), .Y(n_675) );
AOI21xp33_ASAP7_75t_SL g1037 ( .A1(n_389), .A2(n_1038), .B(n_1039), .Y(n_1037) );
INVx5_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g785 ( .A(n_390), .Y(n_785) );
INVx1_ASAP7_75t_L g1004 ( .A(n_390), .Y(n_1004) );
INVx2_ASAP7_75t_L g1513 ( .A(n_390), .Y(n_1513) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx2_ASAP7_75t_L g1140 ( .A(n_391), .Y(n_1140) );
INVx2_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
OR2x6_ASAP7_75t_L g911 ( .A(n_393), .B(n_912), .Y(n_911) );
AND2x4_ASAP7_75t_L g393 ( .A(n_394), .B(n_395), .Y(n_393) );
AND2x4_ASAP7_75t_L g904 ( .A(n_394), .B(n_417), .Y(n_904) );
INVx2_ASAP7_75t_L g1114 ( .A(n_395), .Y(n_1114) );
AND2x2_ASAP7_75t_L g395 ( .A(n_396), .B(n_401), .Y(n_395) );
AND2x4_ASAP7_75t_L g434 ( .A(n_396), .B(n_435), .Y(n_434) );
AND2x4_ASAP7_75t_L g439 ( .A(n_396), .B(n_440), .Y(n_439) );
INVx1_ASAP7_75t_L g458 ( .A(n_396), .Y(n_458) );
AND2x4_ASAP7_75t_L g520 ( .A(n_396), .B(n_435), .Y(n_520) );
BUFx2_ASAP7_75t_L g544 ( .A(n_396), .Y(n_544) );
AND2x2_ASAP7_75t_L g565 ( .A(n_396), .B(n_440), .Y(n_565) );
AND2x2_ASAP7_75t_L g682 ( .A(n_396), .B(n_440), .Y(n_682) );
AND2x4_ASAP7_75t_L g396 ( .A(n_397), .B(n_399), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g417 ( .A(n_399), .B(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
AND2x2_ASAP7_75t_L g450 ( .A(n_400), .B(n_418), .Y(n_450) );
INVx6_ASAP7_75t_L g415 ( .A(n_401), .Y(n_415) );
INVx2_ASAP7_75t_L g572 ( .A(n_401), .Y(n_572) );
BUFx2_ASAP7_75t_L g778 ( .A(n_401), .Y(n_778) );
AND2x4_ASAP7_75t_L g401 ( .A(n_402), .B(n_404), .Y(n_401) );
INVx1_ASAP7_75t_L g441 ( .A(n_402), .Y(n_441) );
INVx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g412 ( .A(n_403), .B(n_405), .Y(n_412) );
AND2x4_ASAP7_75t_L g423 ( .A(n_403), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g437 ( .A(n_404), .Y(n_437) );
INVx2_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
AND2x4_ASAP7_75t_L g427 ( .A(n_405), .B(n_428), .Y(n_427) );
AOI31xp33_ASAP7_75t_L g407 ( .A1(n_408), .A2(n_442), .A3(n_459), .B(n_468), .Y(n_407) );
BUFx2_ASAP7_75t_L g1532 ( .A(n_410), .Y(n_1532) );
BUFx4f_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
AND2x4_ASAP7_75t_L g455 ( .A(n_411), .B(n_430), .Y(n_455) );
INVx2_ASAP7_75t_SL g536 ( .A(n_411), .Y(n_536) );
AND2x4_ASAP7_75t_L g543 ( .A(n_411), .B(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g635 ( .A(n_411), .Y(n_635) );
BUFx6f_ASAP7_75t_L g896 ( .A(n_411), .Y(n_896) );
BUFx6f_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_412), .Y(n_447) );
HB1xp67_ASAP7_75t_L g842 ( .A(n_413), .Y(n_842) );
BUFx6f_ASAP7_75t_L g413 ( .A(n_414), .Y(n_413) );
INVx1_ASAP7_75t_L g638 ( .A(n_414), .Y(n_638) );
INVx2_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_415), .Y(n_453) );
INVx2_ASAP7_75t_SL g528 ( .A(n_415), .Y(n_528) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_415), .Y(n_542) );
INVx2_ASAP7_75t_L g691 ( .A(n_415), .Y(n_691) );
INVx1_ASAP7_75t_L g894 ( .A(n_415), .Y(n_894) );
INVx1_ASAP7_75t_L g899 ( .A(n_415), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g529 ( .A(n_417), .Y(n_529) );
INVx2_ASAP7_75t_SL g631 ( .A(n_417), .Y(n_631) );
INVx1_ASAP7_75t_L g779 ( .A(n_417), .Y(n_779) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g901 ( .A(n_421), .Y(n_901) );
INVx2_ASAP7_75t_SL g421 ( .A(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g429 ( .A(n_422), .B(n_430), .Y(n_429) );
BUFx3_ASAP7_75t_L g561 ( .A(n_422), .Y(n_561) );
BUFx6f_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
BUFx2_ASAP7_75t_L g444 ( .A(n_423), .Y(n_444) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_423), .Y(n_526) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_423), .Y(n_539) );
BUFx6f_ASAP7_75t_L g770 ( .A(n_423), .Y(n_770) );
BUFx2_ASAP7_75t_L g838 ( .A(n_423), .Y(n_838) );
INVx2_ASAP7_75t_SL g871 ( .A(n_423), .Y(n_871) );
BUFx3_ASAP7_75t_L g890 ( .A(n_423), .Y(n_890) );
INVx1_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
INVx1_ASAP7_75t_L g1230 ( .A(n_425), .Y(n_1230) );
BUFx6f_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
BUFx3_ASAP7_75t_L g902 ( .A(n_426), .Y(n_902) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx2_ASAP7_75t_L g467 ( .A(n_427), .Y(n_467) );
INVx1_ASAP7_75t_L g574 ( .A(n_427), .Y(n_574) );
BUFx6f_ASAP7_75t_L g641 ( .A(n_427), .Y(n_641) );
INVx1_ASAP7_75t_L g857 ( .A(n_427), .Y(n_857) );
INVx1_ASAP7_75t_L g463 ( .A(n_428), .Y(n_463) );
AOI21xp33_ASAP7_75t_L g516 ( .A1(n_429), .A2(n_517), .B(n_518), .Y(n_516) );
AOI221xp5_ASAP7_75t_L g558 ( .A1(n_429), .A2(n_559), .B1(n_560), .B2(n_562), .C(n_563), .Y(n_558) );
AOI211xp5_ASAP7_75t_L g617 ( .A1(n_429), .A2(n_618), .B(n_619), .C(n_621), .Y(n_617) );
AOI22xp33_ASAP7_75t_L g702 ( .A1(n_429), .A2(n_460), .B1(n_703), .B2(n_704), .Y(n_702) );
INVx1_ASAP7_75t_L g833 ( .A(n_429), .Y(n_833) );
AOI211xp5_ASAP7_75t_L g1017 ( .A1(n_429), .A2(n_994), .B(n_1018), .C(n_1021), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1040 ( .A1(n_429), .A2(n_1041), .B(n_1042), .Y(n_1040) );
HB1xp67_ASAP7_75t_L g1518 ( .A(n_429), .Y(n_1518) );
AND2x2_ASAP7_75t_L g769 ( .A(n_430), .B(n_770), .Y(n_769) );
AOI222xp33_ASAP7_75t_L g1097 ( .A1(n_430), .A2(n_434), .B1(n_565), .B2(n_1098), .C1(n_1105), .C2(n_1106), .Y(n_1097) );
OAI21xp5_ASAP7_75t_L g1145 ( .A1(n_430), .A2(n_1146), .B(n_1148), .Y(n_1145) );
INVx2_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g461 ( .A(n_431), .B(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g466 ( .A(n_431), .B(n_467), .Y(n_466) );
A2O1A1Ixp33_ASAP7_75t_SL g1220 ( .A1(n_431), .A2(n_1221), .B(n_1222), .C(n_1224), .Y(n_1220) );
INVx2_ASAP7_75t_SL g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g620 ( .A(n_434), .Y(n_620) );
INVx1_ASAP7_75t_L g835 ( .A(n_434), .Y(n_835) );
INVx2_ASAP7_75t_SL g1019 ( .A(n_434), .Y(n_1019) );
INVxp67_ASAP7_75t_L g1154 ( .A(n_435), .Y(n_1154) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g877 ( .A(n_436), .Y(n_877) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx2_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g783 ( .A(n_439), .Y(n_783) );
INVx2_ASAP7_75t_L g883 ( .A(n_440), .Y(n_883) );
INVx1_ASAP7_75t_L g1155 ( .A(n_440), .Y(n_1155) );
BUFx3_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_445), .Y(n_839) );
BUFx6f_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AND2x4_ASAP7_75t_L g456 ( .A(n_446), .B(n_457), .Y(n_456) );
INVx1_ASAP7_75t_L g569 ( .A(n_446), .Y(n_569) );
INVx1_ASAP7_75t_L g1010 ( .A(n_446), .Y(n_1010) );
AOI22xp5_ASAP7_75t_L g1102 ( .A1(n_446), .A2(n_770), .B1(n_1103), .B2(n_1104), .Y(n_1102) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g827 ( .A(n_447), .Y(n_827) );
INVx1_ASAP7_75t_L g1054 ( .A(n_447), .Y(n_1054) );
INVx3_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g840 ( .A(n_449), .Y(n_840) );
OAI221xp5_ASAP7_75t_L g1231 ( .A1(n_449), .A2(n_1204), .B1(n_1209), .B2(n_1232), .C(n_1234), .Y(n_1231) );
BUFx3_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
INVx2_ASAP7_75t_SL g700 ( .A(n_450), .Y(n_700) );
INVx2_ASAP7_75t_L g887 ( .A(n_450), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g1221 ( .A1(n_452), .A2(n_1024), .B1(n_1214), .B2(n_1216), .Y(n_1221) );
INVx4_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g829 ( .A(n_453), .Y(n_829) );
INVx1_ASAP7_75t_L g1152 ( .A(n_453), .Y(n_1152) );
AOI221xp5_ASAP7_75t_L g1007 ( .A1(n_454), .A2(n_456), .B1(n_1002), .B2(n_1008), .C(n_1013), .Y(n_1007) );
AOI221xp5_ASAP7_75t_L g1047 ( .A1(n_454), .A2(n_456), .B1(n_1048), .B2(n_1049), .C(n_1057), .Y(n_1047) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g532 ( .A(n_455), .Y(n_532) );
AOI221xp5_ASAP7_75t_L g566 ( .A1(n_455), .A2(n_456), .B1(n_567), .B2(n_570), .C(n_575), .Y(n_566) );
INVx2_ASAP7_75t_SL g694 ( .A(n_455), .Y(n_694) );
INVx1_ASAP7_75t_L g845 ( .A(n_455), .Y(n_845) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_456), .A2(n_531), .B1(n_633), .B2(n_634), .C(n_636), .Y(n_632) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_456), .A2(n_693), .B1(n_695), .B2(n_696), .C(n_701), .Y(n_692) );
AOI221xp5_ASAP7_75t_L g771 ( .A1(n_456), .A2(n_693), .B1(n_762), .B2(n_772), .C(n_773), .Y(n_771) );
HB1xp67_ASAP7_75t_L g846 ( .A(n_456), .Y(n_846) );
AOI21xp33_ASAP7_75t_L g1107 ( .A1(n_456), .A2(n_1108), .B(n_1109), .Y(n_1107) );
INVx1_ASAP7_75t_L g1224 ( .A(n_456), .Y(n_1224) );
AOI221xp5_ASAP7_75t_L g1529 ( .A1(n_456), .A2(n_531), .B1(n_1530), .B2(n_1531), .C(n_1534), .Y(n_1529) );
INVx1_ASAP7_75t_SL g457 ( .A(n_458), .Y(n_457) );
OR2x2_ASAP7_75t_L g1020 ( .A(n_458), .B(n_883), .Y(n_1020) );
AOI22xp33_ASAP7_75t_L g545 ( .A1(n_460), .A2(n_465), .B1(n_546), .B2(n_547), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_460), .A2(n_465), .B1(n_577), .B2(n_578), .Y(n_576) );
AOI22xp33_ASAP7_75t_SL g642 ( .A1(n_460), .A2(n_465), .B1(n_643), .B2(n_644), .Y(n_642) );
AOI22xp5_ASAP7_75t_L g766 ( .A1(n_460), .A2(n_757), .B1(n_760), .B2(n_767), .Y(n_766) );
AOI22xp33_ASAP7_75t_L g847 ( .A1(n_460), .A2(n_465), .B1(n_813), .B2(n_815), .Y(n_847) );
AOI22xp33_ASAP7_75t_SL g1030 ( .A1(n_460), .A2(n_465), .B1(n_998), .B2(n_1000), .Y(n_1030) );
AOI22xp33_ASAP7_75t_L g1060 ( .A1(n_460), .A2(n_465), .B1(n_1061), .B2(n_1062), .Y(n_1060) );
AOI22xp33_ASAP7_75t_L g1536 ( .A1(n_460), .A2(n_465), .B1(n_1537), .B2(n_1538), .Y(n_1536) );
INVx6_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g628 ( .A(n_462), .Y(n_628) );
INVx2_ASAP7_75t_L g1028 ( .A(n_462), .Y(n_1028) );
BUFx2_ASAP7_75t_L g1525 ( .A(n_462), .Y(n_1525) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AND2x2_ASAP7_75t_L g524 ( .A(n_463), .B(n_464), .Y(n_524) );
AOI211xp5_ASAP7_75t_L g678 ( .A1(n_465), .A2(n_679), .B(n_680), .C(n_683), .Y(n_678) );
AOI221xp5_ASAP7_75t_L g776 ( .A1(n_465), .A2(n_758), .B1(n_777), .B2(n_780), .C(n_782), .Y(n_776) );
INVx4_ASAP7_75t_L g465 ( .A(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g781 ( .A(n_467), .Y(n_781) );
INVx2_ASAP7_75t_L g1101 ( .A(n_467), .Y(n_1101) );
AOI31xp33_ASAP7_75t_L g616 ( .A1(n_468), .A2(n_617), .A3(n_632), .B(n_642), .Y(n_616) );
INVx5_ASAP7_75t_L g764 ( .A(n_468), .Y(n_764) );
BUFx8_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
INVx2_ASAP7_75t_L g514 ( .A(n_469), .Y(n_514) );
OAI31xp33_ASAP7_75t_L g919 ( .A1(n_469), .A2(n_920), .A3(n_939), .B(n_960), .Y(n_919) );
AOI31xp33_ASAP7_75t_L g1515 ( .A1(n_469), .A2(n_1516), .A3(n_1529), .B(n_1536), .Y(n_1515) );
INVx2_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
BUFx2_ASAP7_75t_L g676 ( .A(n_470), .Y(n_676) );
INVx1_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
HB1xp67_ASAP7_75t_L g549 ( .A(n_472), .Y(n_549) );
AND2x2_ASAP7_75t_L g473 ( .A(n_474), .B(n_513), .Y(n_473) );
AND4x1_ASAP7_75t_L g474 ( .A(n_475), .B(n_485), .C(n_489), .D(n_493), .Y(n_474) );
AOI221xp5_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_478), .B1(n_479), .B2(n_482), .C(n_483), .Y(n_475) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_476), .A2(n_479), .B1(n_483), .B2(n_708), .C(n_709), .Y(n_707) );
AOI221xp5_ASAP7_75t_L g1141 ( .A1(n_476), .A2(n_479), .B1(n_483), .B2(n_1105), .C(n_1106), .Y(n_1141) );
AOI21xp5_ASAP7_75t_L g1190 ( .A1(n_476), .A2(n_483), .B(n_1191), .Y(n_1190) );
AND2x2_ASAP7_75t_L g936 ( .A(n_477), .B(n_915), .Y(n_936) );
AOI22xp33_ASAP7_75t_L g1174 ( .A1(n_479), .A2(n_1140), .B1(n_1151), .B2(n_1175), .Y(n_1174) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
OAI211xp5_ASAP7_75t_L g521 ( .A1(n_488), .A2(n_522), .B(n_525), .C(n_527), .Y(n_521) );
AOI33xp33_ASAP7_75t_L g493 ( .A1(n_494), .A2(n_498), .A3(n_503), .B1(n_506), .B2(n_509), .B3(n_512), .Y(n_493) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
AOI33xp33_ASAP7_75t_L g710 ( .A1(n_495), .A2(n_512), .A3(n_711), .B1(n_715), .B2(n_716), .B3(n_719), .Y(n_710) );
AOI22xp5_ASAP7_75t_L g1131 ( .A1(n_495), .A2(n_1115), .B1(n_1132), .B2(n_1140), .Y(n_1131) );
AOI322xp5_ASAP7_75t_L g1182 ( .A1(n_495), .A2(n_512), .A3(n_1166), .B1(n_1183), .B2(n_1185), .C1(n_1186), .C2(n_1189), .Y(n_1182) );
AND2x4_ASAP7_75t_L g495 ( .A(n_496), .B(n_497), .Y(n_495) );
OR2x6_ASAP7_75t_L g886 ( .A(n_496), .B(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g913 ( .A(n_496), .Y(n_913) );
BUFx2_ASAP7_75t_L g1246 ( .A(n_496), .Y(n_1246) );
INVx1_ASAP7_75t_L g957 ( .A(n_497), .Y(n_957) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g511 ( .A(n_500), .Y(n_511) );
AOI22xp5_ASAP7_75t_L g1121 ( .A1(n_500), .A2(n_1122), .B1(n_1123), .B2(n_1124), .Y(n_1121) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx1_ASAP7_75t_L g812 ( .A(n_505), .Y(n_812) );
INVx1_ASAP7_75t_L g1081 ( .A(n_505), .Y(n_1081) );
INVx2_ASAP7_75t_SL g990 ( .A(n_507), .Y(n_990) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
INVx1_ASAP7_75t_L g1128 ( .A(n_508), .Y(n_1128) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx1_ASAP7_75t_L g1557 ( .A(n_512), .Y(n_1557) );
NAND3xp33_ASAP7_75t_L g515 ( .A(n_516), .B(n_530), .C(n_545), .Y(n_515) );
INVx2_ASAP7_75t_L g519 ( .A(n_520), .Y(n_519) );
OAI211xp5_ASAP7_75t_L g1043 ( .A1(n_522), .A2(n_1044), .B(n_1045), .C(n_1046), .Y(n_1043) );
INVx2_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_SL g1149 ( .A(n_523), .Y(n_1149) );
INVx1_ASAP7_75t_L g1523 ( .A(n_523), .Y(n_1523) );
BUFx4f_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g625 ( .A(n_524), .Y(n_625) );
BUFx2_ASAP7_75t_L g688 ( .A(n_524), .Y(n_688) );
INVx2_ASAP7_75t_L g862 ( .A(n_524), .Y(n_862) );
INVx1_ASAP7_75t_L g1233 ( .A(n_524), .Y(n_1233) );
INVx2_ASAP7_75t_L g623 ( .A(n_526), .Y(n_623) );
INVx2_ASAP7_75t_SL g698 ( .A(n_526), .Y(n_698) );
BUFx3_ASAP7_75t_L g1235 ( .A(n_526), .Y(n_1235) );
INVx1_ASAP7_75t_L g775 ( .A(n_528), .Y(n_775) );
INVx1_ASAP7_75t_L g1527 ( .A(n_529), .Y(n_1527) );
AOI221xp5_ASAP7_75t_L g530 ( .A1(n_531), .A2(n_533), .B1(n_534), .B2(n_540), .C(n_543), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx2_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
INVx1_ASAP7_75t_L g684 ( .A(n_538), .Y(n_684) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
BUFx3_ASAP7_75t_L g1156 ( .A(n_544), .Y(n_1156) );
INVx1_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AO22x1_ASAP7_75t_L g552 ( .A1(n_553), .A2(n_610), .B1(n_611), .B2(n_667), .Y(n_552) );
BUFx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g667 ( .A(n_554), .Y(n_667) );
XOR2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_609), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_580), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_558), .B(n_566), .C(n_576), .Y(n_557) );
INVxp67_ASAP7_75t_L g1238 ( .A(n_561), .Y(n_1238) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_562), .A2(n_578), .B1(n_600), .B2(n_604), .Y(n_603) );
INVx3_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
INVx1_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g699 ( .A(n_569), .Y(n_699) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx2_ASAP7_75t_SL g866 ( .A(n_572), .Y(n_866) );
INVx1_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g685 ( .A(n_574), .Y(n_685) );
INVx1_ASAP7_75t_L g1535 ( .A(n_574), .Y(n_1535) );
OAI22xp33_ASAP7_75t_L g606 ( .A1(n_575), .A2(n_577), .B1(n_594), .B2(n_607), .Y(n_606) );
NOR3xp33_ASAP7_75t_L g580 ( .A(n_581), .B(n_589), .C(n_591), .Y(n_580) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_582), .B(n_586), .Y(n_581) );
OAI22xp33_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B1(n_596), .B2(n_597), .Y(n_592) );
OAI22xp33_ASAP7_75t_L g650 ( .A1(n_594), .A2(n_651), .B1(n_652), .B2(n_653), .Y(n_650) );
BUFx2_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx1_ASAP7_75t_L g746 ( .A(n_595), .Y(n_746) );
INVx1_ASAP7_75t_L g1088 ( .A(n_595), .Y(n_1088) );
OAI22xp5_ASAP7_75t_SL g1215 ( .A1(n_595), .A2(n_761), .B1(n_1216), .B2(n_1217), .Y(n_1215) );
OAI22xp5_ASAP7_75t_SL g598 ( .A1(n_599), .A2(n_600), .B1(n_601), .B2(n_602), .Y(n_598) );
OAI22xp5_ASAP7_75t_L g655 ( .A1(n_600), .A2(n_618), .B1(n_644), .B2(n_656), .Y(n_655) );
OAI221xp5_ASAP7_75t_L g926 ( .A1(n_602), .A2(n_854), .B1(n_868), .B2(n_927), .C(n_931), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g1550 ( .A1(n_602), .A2(n_1551), .B1(n_1553), .B2(n_1554), .Y(n_1550) );
OAI22xp33_ASAP7_75t_L g1556 ( .A1(n_602), .A2(n_761), .B1(n_1530), .B2(n_1538), .Y(n_1556) );
OAI22xp5_ASAP7_75t_L g807 ( .A1(n_604), .A2(n_756), .B1(n_808), .B2(n_809), .Y(n_807) );
CKINVDCx5p33_ASAP7_75t_R g604 ( .A(n_605), .Y(n_604) );
OAI22xp33_ASAP7_75t_L g1074 ( .A1(n_607), .A2(n_1075), .B1(n_1077), .B2(n_1078), .Y(n_1074) );
INVx2_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_614), .B(n_645), .Y(n_613) );
INVx2_ASAP7_75t_SL g622 ( .A(n_623), .Y(n_622) );
OAI221xp5_ASAP7_75t_L g624 ( .A1(n_625), .A2(n_626), .B1(n_627), .B2(n_629), .C(n_630), .Y(n_624) );
INVx2_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g1029 ( .A(n_631), .Y(n_1029) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
INVx1_ASAP7_75t_L g843 ( .A(n_640), .Y(n_843) );
OAI22xp5_ASAP7_75t_L g1236 ( .A1(n_640), .A2(n_1237), .B1(n_1238), .B2(n_1239), .Y(n_1236) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
BUFx6f_ASAP7_75t_L g1016 ( .A(n_641), .Y(n_1016) );
BUFx6f_ASAP7_75t_L g1059 ( .A(n_641), .Y(n_1059) );
NOR3xp33_ASAP7_75t_L g645 ( .A(n_646), .B(n_658), .C(n_660), .Y(n_645) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
HB1xp67_ASAP7_75t_L g801 ( .A(n_659), .Y(n_801) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_664), .Y(n_660) );
BUFx3_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
OAI22xp5_ASAP7_75t_L g670 ( .A1(n_671), .A2(n_967), .B1(n_1253), .B2(n_1254), .Y(n_670) );
INVx1_ASAP7_75t_L g1253 ( .A(n_671), .Y(n_1253) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_786), .B1(n_965), .B2(n_966), .Y(n_671) );
INVx1_ASAP7_75t_L g965 ( .A(n_672), .Y(n_965) );
XOR2x2_ASAP7_75t_L g672 ( .A(n_673), .B(n_730), .Y(n_672) );
XNOR2xp5_ASAP7_75t_L g673 ( .A(n_674), .B(n_729), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_675), .B(n_706), .Y(n_674) );
INVx2_ASAP7_75t_L g1031 ( .A(n_676), .Y(n_1031) );
NAND3xp33_ASAP7_75t_SL g677 ( .A(n_678), .B(n_692), .C(n_702), .Y(n_677) );
INVx2_ASAP7_75t_SL g681 ( .A(n_682), .Y(n_681) );
OAI21xp5_ASAP7_75t_SL g686 ( .A1(n_687), .A2(n_689), .B(n_690), .Y(n_686) );
INVx2_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g1026 ( .A(n_688), .Y(n_1026) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_691), .Y(n_1014) );
BUFx3_ASAP7_75t_L g1058 ( .A(n_691), .Y(n_1058) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g1056 ( .A(n_700), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1533 ( .A(n_700), .Y(n_1533) );
AND4x1_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .C(n_724), .D(n_726), .Y(n_706) );
INVx2_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
INVx2_ASAP7_75t_L g1124 ( .A(n_713), .Y(n_1124) );
INVx2_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
INVx2_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
BUFx3_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_723), .Y(n_722) );
XNOR2x1_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
AND2x2_ASAP7_75t_L g732 ( .A(n_733), .B(n_763), .Y(n_732) );
NOR3xp33_ASAP7_75t_L g733 ( .A(n_734), .B(n_741), .C(n_742), .Y(n_733) );
NAND2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_738), .Y(n_734) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_745), .A2(n_760), .B1(n_761), .B2(n_762), .Y(n_759) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
BUFx2_ASAP7_75t_L g750 ( .A(n_751), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g1079 ( .A1(n_751), .A2(n_1080), .B1(n_1081), .B2(n_1082), .Y(n_1079) );
INVx2_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
HB1xp67_ASAP7_75t_L g1552 ( .A(n_752), .Y(n_1552) );
OAI22xp5_ASAP7_75t_L g810 ( .A1(n_756), .A2(n_811), .B1(n_812), .B2(n_813), .Y(n_810) );
AOI22xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B1(n_784), .B2(n_785), .Y(n_763) );
INVx1_ASAP7_75t_SL g848 ( .A(n_764), .Y(n_848) );
NAND3xp33_ASAP7_75t_L g765 ( .A(n_766), .B(n_771), .C(n_776), .Y(n_765) );
INVx1_ASAP7_75t_L g767 ( .A(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g768 ( .A(n_769), .Y(n_768) );
BUFx2_ASAP7_75t_L g831 ( .A(n_770), .Y(n_831) );
INVx1_ASAP7_75t_L g1023 ( .A(n_770), .Y(n_1023) );
INVx1_ASAP7_75t_L g1051 ( .A(n_770), .Y(n_1051) );
INVx2_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_L g1244 ( .A(n_779), .Y(n_1244) );
AOI21xp5_ASAP7_75t_L g819 ( .A1(n_785), .A2(n_820), .B(n_821), .Y(n_819) );
INVx1_ASAP7_75t_L g966 ( .A(n_786), .Y(n_966) );
XOR2xp5_ASAP7_75t_L g786 ( .A(n_787), .B(n_849), .Y(n_786) );
XNOR2xp5_ASAP7_75t_L g787 ( .A(n_788), .B(n_789), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_819), .Y(n_789) );
NOR3xp33_ASAP7_75t_SL g790 ( .A(n_791), .B(n_799), .C(n_802), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
BUFx3_ASAP7_75t_L g953 ( .A(n_805), .Y(n_953) );
OAI22xp5_ASAP7_75t_L g1206 ( .A1(n_805), .A2(n_1207), .B1(n_1208), .B2(n_1209), .Y(n_1206) );
AOI221xp5_ASAP7_75t_SL g822 ( .A1(n_811), .A2(n_823), .B1(n_830), .B2(n_832), .C(n_834), .Y(n_822) );
AOI221xp5_ASAP7_75t_L g836 ( .A1(n_816), .A2(n_837), .B1(n_841), .B2(n_844), .C(n_846), .Y(n_836) );
INVx1_ASAP7_75t_L g817 ( .A(n_818), .Y(n_817) );
AOI31xp33_ASAP7_75t_L g821 ( .A1(n_822), .A2(n_836), .A3(n_847), .B(n_848), .Y(n_821) );
INVx1_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
INVx3_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
HB1xp67_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
CKINVDCx5p33_ASAP7_75t_R g844 ( .A(n_845), .Y(n_844) );
AND3x1_ASAP7_75t_L g850 ( .A(n_851), .B(n_909), .C(n_919), .Y(n_850) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_872), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_853), .B(n_863), .Y(n_852) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_854), .A2(n_855), .B1(n_859), .B2(n_860), .Y(n_853) );
CKINVDCx6p67_ASAP7_75t_R g855 ( .A(n_856), .Y(n_855) );
OR2x6_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
INVx2_ASAP7_75t_L g891 ( .A(n_857), .Y(n_891) );
OR2x6_ASAP7_75t_L g861 ( .A(n_858), .B(n_862), .Y(n_861) );
INVx1_ASAP7_75t_L g867 ( .A(n_858), .Y(n_867) );
CKINVDCx6p67_ASAP7_75t_R g860 ( .A(n_861), .Y(n_860) );
BUFx3_ASAP7_75t_L g1159 ( .A(n_862), .Y(n_1159) );
INVx1_ASAP7_75t_L g1168 ( .A(n_862), .Y(n_1168) );
AOI22xp33_ASAP7_75t_L g863 ( .A1(n_864), .A2(n_865), .B1(n_868), .B2(n_869), .Y(n_863) );
AND2x2_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .Y(n_865) );
AND2x2_ASAP7_75t_L g869 ( .A(n_867), .B(n_870), .Y(n_869) );
INVx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx2_ASAP7_75t_SL g1162 ( .A(n_871), .Y(n_1162) );
NAND3xp33_ASAP7_75t_SL g872 ( .A(n_873), .B(n_884), .C(n_905), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g873 ( .A1(n_874), .A2(n_875), .B1(n_880), .B2(n_881), .Y(n_873) );
AOI22xp33_ASAP7_75t_L g934 ( .A1(n_874), .A2(n_880), .B1(n_935), .B2(n_937), .Y(n_934) );
INVx2_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
NAND2x1p5_ASAP7_75t_L g876 ( .A(n_877), .B(n_878), .Y(n_876) );
INVx2_ASAP7_75t_SL g878 ( .A(n_879), .Y(n_878) );
OR2x6_ASAP7_75t_L g882 ( .A(n_879), .B(n_883), .Y(n_882) );
INVx1_ASAP7_75t_L g908 ( .A(n_879), .Y(n_908) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
AOI33xp33_ASAP7_75t_L g884 ( .A1(n_885), .A2(n_888), .A3(n_892), .B1(n_897), .B2(n_900), .B3(n_903), .Y(n_884) );
CKINVDCx5p33_ASAP7_75t_R g885 ( .A(n_886), .Y(n_885) );
INVx1_ASAP7_75t_L g1164 ( .A(n_887), .Y(n_1164) );
BUFx3_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
INVx2_ASAP7_75t_SL g1012 ( .A(n_890), .Y(n_1012) );
BUFx2_ASAP7_75t_L g1024 ( .A(n_891), .Y(n_1024) );
HB1xp67_ASAP7_75t_L g893 ( .A(n_894), .Y(n_893) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g907 ( .A(n_896), .B(n_908), .Y(n_907) );
BUFx2_ASAP7_75t_SL g1223 ( .A(n_896), .Y(n_1223) );
BUFx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
BUFx4f_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g905 ( .A(n_906), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_910), .B(n_911), .Y(n_909) );
NOR2xp67_ASAP7_75t_L g912 ( .A(n_913), .B(n_914), .Y(n_912) );
INVx2_ASAP7_75t_L g1116 ( .A(n_913), .Y(n_1116) );
AOI211xp5_ASAP7_75t_L g1143 ( .A1(n_913), .A2(n_1144), .B(n_1171), .C(n_1181), .Y(n_1143) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_918), .Y(n_914) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
OR2x2_ASAP7_75t_L g958 ( .A(n_916), .B(n_959), .Y(n_958) );
INVx2_ASAP7_75t_L g916 ( .A(n_917), .Y(n_916) );
INVx8_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
AND2x4_ASAP7_75t_L g922 ( .A(n_923), .B(n_925), .Y(n_922) );
AND2x4_ASAP7_75t_L g964 ( .A(n_923), .B(n_950), .Y(n_964) );
INVx1_ASAP7_75t_L g923 ( .A(n_924), .Y(n_923) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx2_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
OAI22xp5_ASAP7_75t_L g1083 ( .A1(n_929), .A2(n_1041), .B1(n_1062), .B2(n_1084), .Y(n_1083) );
INVx2_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_SL g945 ( .A(n_930), .Y(n_945) );
INVx2_ASAP7_75t_L g988 ( .A(n_930), .Y(n_988) );
INVx2_ASAP7_75t_SL g932 ( .A(n_933), .Y(n_932) );
HB1xp67_ASAP7_75t_L g935 ( .A(n_936), .Y(n_935) );
CKINVDCx11_ASAP7_75t_R g937 ( .A(n_938), .Y(n_937) );
CKINVDCx6p67_ASAP7_75t_R g940 ( .A(n_941), .Y(n_940) );
OAI22xp5_ASAP7_75t_SL g942 ( .A1(n_943), .A2(n_944), .B1(n_946), .B2(n_947), .Y(n_942) );
BUFx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_949), .Y(n_948) );
INVx1_ASAP7_75t_L g949 ( .A(n_950), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
OAI22xp33_ASAP7_75t_L g982 ( .A1(n_953), .A2(n_983), .B1(n_984), .B2(n_985), .Y(n_982) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
INVx3_ASAP7_75t_L g961 ( .A(n_962), .Y(n_961) );
INVx3_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
AOI22xp33_ASAP7_75t_L g967 ( .A1(n_968), .A2(n_1032), .B1(n_1250), .B2(n_1252), .Y(n_967) );
INVx2_ASAP7_75t_L g968 ( .A(n_969), .Y(n_968) );
HB1xp67_ASAP7_75t_L g1252 ( .A(n_969), .Y(n_1252) );
AOI22xp33_ASAP7_75t_L g1254 ( .A1(n_969), .A2(n_1032), .B1(n_1033), .B2(n_1255), .Y(n_1254) );
AND2x2_ASAP7_75t_L g970 ( .A(n_971), .B(n_1003), .Y(n_970) );
NOR3xp33_ASAP7_75t_SL g971 ( .A(n_972), .B(n_980), .C(n_981), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g972 ( .A(n_973), .B(n_977), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g1025 ( .A1(n_976), .A2(n_978), .B1(n_1026), .B2(n_1027), .C(n_1029), .Y(n_1025) );
OAI22xp33_ASAP7_75t_L g999 ( .A1(n_984), .A2(n_1000), .B1(n_1001), .B2(n_1002), .Y(n_999) );
OAI22xp5_ASAP7_75t_L g986 ( .A1(n_987), .A2(n_988), .B1(n_989), .B2(n_990), .Y(n_986) );
OAI22xp5_ASAP7_75t_L g991 ( .A1(n_992), .A2(n_994), .B1(n_995), .B2(n_998), .Y(n_991) );
BUFx2_ASAP7_75t_L g992 ( .A(n_993), .Y(n_992) );
INVx2_ASAP7_75t_L g1213 ( .A(n_993), .Y(n_1213) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVx2_ASAP7_75t_L g996 ( .A(n_997), .Y(n_996) );
AOI21xp5_ASAP7_75t_L g1003 ( .A1(n_1004), .A2(n_1005), .B(n_1006), .Y(n_1003) );
AOI31xp33_ASAP7_75t_L g1006 ( .A1(n_1007), .A2(n_1017), .A3(n_1030), .B(n_1031), .Y(n_1006) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1010), .Y(n_1009) );
AOI22xp33_ASAP7_75t_L g1222 ( .A1(n_1011), .A2(n_1211), .B1(n_1217), .B2(n_1223), .Y(n_1222) );
INVx1_ASAP7_75t_L g1011 ( .A(n_1012), .Y(n_1011) );
HB1xp67_ASAP7_75t_L g1015 ( .A(n_1016), .Y(n_1015) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx2_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx2_ASAP7_75t_L g1147 ( .A(n_1028), .Y(n_1147) );
HB1xp67_ASAP7_75t_L g1229 ( .A(n_1028), .Y(n_1229) );
INVx2_ASAP7_75t_L g1242 ( .A(n_1028), .Y(n_1242) );
AOI31xp33_ASAP7_75t_L g1039 ( .A1(n_1031), .A2(n_1040), .A3(n_1047), .B(n_1060), .Y(n_1039) );
INVx2_ASAP7_75t_L g1032 ( .A(n_1033), .Y(n_1032) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1033), .Y(n_1251) );
XNOR2x1_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1090), .Y(n_1033) );
INVx1_ASAP7_75t_L g1034 ( .A(n_1035), .Y(n_1034) );
XNOR2x1_ASAP7_75t_L g1035 ( .A(n_1036), .B(n_1089), .Y(n_1035) );
AND2x2_ASAP7_75t_L g1036 ( .A(n_1037), .B(n_1063), .Y(n_1036) );
INVx1_ASAP7_75t_L g1050 ( .A(n_1051), .Y(n_1050) );
HB1xp67_ASAP7_75t_L g1052 ( .A(n_1053), .Y(n_1052) );
INVx1_ASAP7_75t_L g1053 ( .A(n_1054), .Y(n_1053) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NOR3xp33_ASAP7_75t_SL g1063 ( .A(n_1064), .B(n_1071), .C(n_1073), .Y(n_1063) );
NAND2xp5_ASAP7_75t_L g1064 ( .A(n_1065), .B(n_1068), .Y(n_1064) );
INVx1_ASAP7_75t_L g1075 ( .A(n_1076), .Y(n_1075) );
INVx2_ASAP7_75t_L g1208 ( .A(n_1076), .Y(n_1208) );
HB1xp67_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
INVx1_ASAP7_75t_L g1087 ( .A(n_1088), .Y(n_1087) );
OAI22x1_ASAP7_75t_L g1090 ( .A1(n_1091), .A2(n_1092), .B1(n_1192), .B2(n_1249), .Y(n_1090) );
INVx1_ASAP7_75t_L g1091 ( .A(n_1092), .Y(n_1091) );
XNOR2x1_ASAP7_75t_L g1092 ( .A(n_1093), .B(n_1142), .Y(n_1092) );
XNOR2x1_ASAP7_75t_L g1093 ( .A(n_1094), .B(n_1095), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1263 ( .A1(n_1094), .A2(n_1264), .B1(n_1271), .B2(n_1272), .Y(n_1263) );
OR2x2_ASAP7_75t_L g1095 ( .A(n_1096), .B(n_1117), .Y(n_1095) );
AOI31xp33_ASAP7_75t_SL g1096 ( .A1(n_1097), .A2(n_1107), .A3(n_1110), .B(n_1116), .Y(n_1096) );
INVx1_ASAP7_75t_L g1099 ( .A(n_1100), .Y(n_1099) );
BUFx2_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
INVx2_ASAP7_75t_L g1521 ( .A(n_1101), .Y(n_1521) );
AOI22xp5_ASAP7_75t_L g1110 ( .A1(n_1111), .A2(n_1112), .B1(n_1113), .B2(n_1115), .Y(n_1110) );
INVx2_ASAP7_75t_L g1113 ( .A(n_1114), .Y(n_1113) );
NAND3xp33_ASAP7_75t_L g1117 ( .A(n_1118), .B(n_1131), .C(n_1141), .Y(n_1117) );
INVx2_ASAP7_75t_L g1126 ( .A(n_1127), .Y(n_1126) );
INVx1_ASAP7_75t_L g1133 ( .A(n_1134), .Y(n_1133) );
INVxp67_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
NAND4xp25_ASAP7_75t_L g1144 ( .A(n_1145), .B(n_1150), .C(n_1157), .D(n_1165), .Y(n_1144) );
A2O1A1Ixp33_ASAP7_75t_L g1150 ( .A1(n_1151), .A2(n_1152), .B(n_1153), .C(n_1156), .Y(n_1150) );
OAI211xp5_ASAP7_75t_L g1157 ( .A1(n_1158), .A2(n_1159), .B(n_1160), .C(n_1161), .Y(n_1157) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
OAI211xp5_ASAP7_75t_L g1165 ( .A1(n_1166), .A2(n_1167), .B(n_1169), .C(n_1170), .Y(n_1165) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1168), .Y(n_1167) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1196 ( .A(n_1173), .Y(n_1196) );
AOI22xp5_ASAP7_75t_L g1176 ( .A1(n_1177), .A2(n_1178), .B1(n_1179), .B2(n_1180), .Y(n_1176) );
INVx1_ASAP7_75t_L g1218 ( .A(n_1178), .Y(n_1218) );
INVx2_ASAP7_75t_L g1199 ( .A(n_1180), .Y(n_1199) );
NAND2xp5_ASAP7_75t_L g1181 ( .A(n_1182), .B(n_1190), .Y(n_1181) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1192), .Y(n_1249) );
INVx1_ASAP7_75t_L g1247 ( .A(n_1193), .Y(n_1247) );
NAND3xp33_ASAP7_75t_L g1193 ( .A(n_1194), .B(n_1200), .C(n_1219), .Y(n_1193) );
NOR2xp33_ASAP7_75t_L g1194 ( .A(n_1195), .B(n_1198), .Y(n_1194) );
NOR2xp33_ASAP7_75t_L g1200 ( .A(n_1201), .B(n_1202), .Y(n_1200) );
OAI22xp5_ASAP7_75t_L g1227 ( .A1(n_1205), .A2(n_1207), .B1(n_1228), .B2(n_1230), .Y(n_1227) );
INVx2_ASAP7_75t_L g1212 ( .A(n_1213), .Y(n_1212) );
OAI31xp33_ASAP7_75t_L g1219 ( .A1(n_1220), .A2(n_1225), .A3(n_1226), .B(n_1245), .Y(n_1219) );
OAI22xp5_ASAP7_75t_L g1226 ( .A1(n_1227), .A2(n_1231), .B1(n_1236), .B2(n_1240), .Y(n_1226) );
INVx1_ASAP7_75t_L g1228 ( .A(n_1229), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1240 ( .A1(n_1232), .A2(n_1241), .B1(n_1242), .B2(n_1243), .C(n_1244), .Y(n_1240) );
BUFx2_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
CKINVDCx8_ASAP7_75t_R g1245 ( .A(n_1246), .Y(n_1245) );
INVx1_ASAP7_75t_L g1250 ( .A(n_1251), .Y(n_1250) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1252), .Y(n_1255) );
OAI221xp5_ASAP7_75t_L g1256 ( .A1(n_1257), .A2(n_1506), .B1(n_1508), .B2(n_1558), .C(n_1562), .Y(n_1256) );
NOR2x1_ASAP7_75t_L g1257 ( .A(n_1258), .B(n_1443), .Y(n_1257) );
NAND3xp33_ASAP7_75t_L g1258 ( .A(n_1259), .B(n_1364), .C(n_1403), .Y(n_1258) );
OAI21xp5_ASAP7_75t_L g1259 ( .A1(n_1260), .A2(n_1320), .B(n_1338), .Y(n_1259) );
AOI22xp5_ASAP7_75t_L g1260 ( .A1(n_1261), .A2(n_1297), .B1(n_1314), .B2(n_1316), .Y(n_1260) );
NOR2xp33_ASAP7_75t_L g1429 ( .A(n_1261), .B(n_1324), .Y(n_1429) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1262), .B(n_1284), .Y(n_1261) );
CKINVDCx6p67_ASAP7_75t_R g1313 ( .A(n_1262), .Y(n_1313) );
OAI222xp33_ASAP7_75t_L g1320 ( .A1(n_1262), .A2(n_1321), .B1(n_1324), .B2(n_1329), .C1(n_1333), .C2(n_1337), .Y(n_1320) );
AND2x2_ASAP7_75t_L g1323 ( .A(n_1262), .B(n_1285), .Y(n_1323) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1262), .B(n_1336), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1395 ( .A(n_1262), .B(n_1318), .Y(n_1395) );
AND2x2_ASAP7_75t_L g1402 ( .A(n_1262), .B(n_1335), .Y(n_1402) );
AND2x2_ASAP7_75t_L g1407 ( .A(n_1262), .B(n_1383), .Y(n_1407) );
OR2x2_ASAP7_75t_L g1427 ( .A(n_1262), .B(n_1336), .Y(n_1427) );
AND2x2_ASAP7_75t_L g1437 ( .A(n_1262), .B(n_1306), .Y(n_1437) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1262), .B(n_1442), .Y(n_1441) );
AND2x2_ASAP7_75t_L g1449 ( .A(n_1262), .B(n_1410), .Y(n_1449) );
OR2x6_ASAP7_75t_SL g1262 ( .A(n_1263), .B(n_1274), .Y(n_1262) );
INVx1_ASAP7_75t_L g1264 ( .A(n_1265), .Y(n_1264) );
AND2x2_ASAP7_75t_L g1265 ( .A(n_1266), .B(n_1268), .Y(n_1265) );
AND2x4_ASAP7_75t_L g1273 ( .A(n_1266), .B(n_1269), .Y(n_1273) );
AND2x4_ASAP7_75t_L g1301 ( .A(n_1266), .B(n_1268), .Y(n_1301) );
INVx1_ASAP7_75t_L g1279 ( .A(n_1267), .Y(n_1279) );
HB1xp67_ASAP7_75t_L g1573 ( .A(n_1268), .Y(n_1573) );
INVx1_ASAP7_75t_L g1268 ( .A(n_1269), .Y(n_1268) );
INVx1_ASAP7_75t_L g1269 ( .A(n_1270), .Y(n_1269) );
NAND2xp5_ASAP7_75t_L g1278 ( .A(n_1270), .B(n_1279), .Y(n_1278) );
OAI22xp5_ASAP7_75t_L g1360 ( .A1(n_1272), .A2(n_1361), .B1(n_1362), .B2(n_1363), .Y(n_1360) );
INVx1_ASAP7_75t_SL g1272 ( .A(n_1273), .Y(n_1272) );
INVx2_ASAP7_75t_L g1312 ( .A(n_1273), .Y(n_1312) );
OAI22xp5_ASAP7_75t_L g1274 ( .A1(n_1275), .A2(n_1280), .B1(n_1281), .B2(n_1283), .Y(n_1274) );
OAI22xp33_ASAP7_75t_L g1302 ( .A1(n_1275), .A2(n_1281), .B1(n_1303), .B2(n_1304), .Y(n_1302) );
BUFx3_ASAP7_75t_L g1348 ( .A(n_1275), .Y(n_1348) );
OAI22xp33_ASAP7_75t_L g1357 ( .A1(n_1275), .A2(n_1351), .B1(n_1358), .B2(n_1359), .Y(n_1357) );
BUFx6f_ASAP7_75t_L g1275 ( .A(n_1276), .Y(n_1275) );
OAI22xp5_ASAP7_75t_L g1294 ( .A1(n_1276), .A2(n_1281), .B1(n_1295), .B2(n_1296), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1276 ( .A(n_1277), .B(n_1278), .Y(n_1276) );
OR2x2_ASAP7_75t_L g1281 ( .A(n_1277), .B(n_1282), .Y(n_1281) );
INVx1_ASAP7_75t_L g1289 ( .A(n_1277), .Y(n_1289) );
INVx1_ASAP7_75t_L g1288 ( .A(n_1278), .Y(n_1288) );
HB1xp67_ASAP7_75t_L g1575 ( .A(n_1279), .Y(n_1575) );
INVx1_ASAP7_75t_L g1352 ( .A(n_1281), .Y(n_1352) );
INVx1_ASAP7_75t_L g1291 ( .A(n_1282), .Y(n_1291) );
INVx1_ASAP7_75t_L g1383 ( .A(n_1284), .Y(n_1383) );
OAI221xp5_ASAP7_75t_L g1404 ( .A1(n_1284), .A2(n_1405), .B1(n_1411), .B2(n_1414), .C(n_1416), .Y(n_1404) );
NOR2xp33_ASAP7_75t_L g1442 ( .A(n_1284), .B(n_1319), .Y(n_1442) );
OR2x2_ASAP7_75t_L g1284 ( .A(n_1285), .B(n_1293), .Y(n_1284) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1285), .B(n_1293), .Y(n_1306) );
INVx1_ASAP7_75t_L g1336 ( .A(n_1285), .Y(n_1336) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1285), .B(n_1367), .Y(n_1410) );
NOR2xp33_ASAP7_75t_SL g1481 ( .A(n_1285), .B(n_1482), .Y(n_1481) );
AND2x2_ASAP7_75t_L g1285 ( .A(n_1286), .B(n_1292), .Y(n_1285) );
AND2x4_ASAP7_75t_L g1287 ( .A(n_1288), .B(n_1289), .Y(n_1287) );
AND2x4_ASAP7_75t_L g1290 ( .A(n_1289), .B(n_1291), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1293), .B(n_1336), .Y(n_1335) );
INVx1_ASAP7_75t_L g1367 ( .A(n_1293), .Y(n_1367) );
AND2x2_ASAP7_75t_L g1461 ( .A(n_1293), .B(n_1313), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1305), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1492 ( .A(n_1298), .B(n_1447), .Y(n_1492) );
NAND2xp5_ASAP7_75t_L g1498 ( .A(n_1298), .B(n_1499), .Y(n_1498) );
INVx1_ASAP7_75t_L g1298 ( .A(n_1299), .Y(n_1298) );
INVx1_ASAP7_75t_L g1315 ( .A(n_1299), .Y(n_1315) );
INVx1_ASAP7_75t_L g1380 ( .A(n_1299), .Y(n_1380) );
NAND2xp5_ASAP7_75t_L g1420 ( .A(n_1299), .B(n_1421), .Y(n_1420) );
NAND2xp5_ASAP7_75t_L g1457 ( .A(n_1299), .B(n_1407), .Y(n_1457) );
HB1xp67_ASAP7_75t_L g1299 ( .A(n_1300), .Y(n_1299) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1300), .B(n_1326), .Y(n_1325) );
INVx2_ASAP7_75t_SL g1332 ( .A(n_1300), .Y(n_1332) );
OR2x2_ASAP7_75t_L g1387 ( .A(n_1300), .B(n_1326), .Y(n_1387) );
INVx1_ASAP7_75t_L g1344 ( .A(n_1301), .Y(n_1344) );
INVx1_ASAP7_75t_L g1362 ( .A(n_1301), .Y(n_1362) );
NAND2xp5_ASAP7_75t_L g1305 ( .A(n_1306), .B(n_1307), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1318 ( .A(n_1306), .B(n_1319), .Y(n_1318) );
AOI322xp5_ASAP7_75t_L g1493 ( .A1(n_1306), .A2(n_1354), .A3(n_1367), .B1(n_1393), .B2(n_1470), .C1(n_1494), .C2(n_1495), .Y(n_1493) );
NAND2xp5_ASAP7_75t_L g1375 ( .A(n_1307), .B(n_1335), .Y(n_1375) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1307), .B(n_1383), .Y(n_1500) );
AND2x2_ASAP7_75t_L g1307 ( .A(n_1308), .B(n_1313), .Y(n_1307) );
INVx4_ASAP7_75t_L g1319 ( .A(n_1308), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1308), .B(n_1331), .Y(n_1330) );
NOR2xp33_ASAP7_75t_L g1384 ( .A(n_1308), .B(n_1313), .Y(n_1384) );
INVx2_ASAP7_75t_L g1400 ( .A(n_1308), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1428 ( .A(n_1308), .B(n_1332), .Y(n_1428) );
NAND2xp5_ASAP7_75t_L g1451 ( .A(n_1308), .B(n_1449), .Y(n_1451) );
AND2x2_ASAP7_75t_L g1470 ( .A(n_1308), .B(n_1356), .Y(n_1470) );
A2O1A1Ixp33_ASAP7_75t_SL g1477 ( .A1(n_1308), .A2(n_1478), .B(n_1479), .C(n_1486), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1308), .B(n_1393), .Y(n_1482) );
OR2x2_ASAP7_75t_L g1485 ( .A(n_1308), .B(n_1401), .Y(n_1485) );
AND2x6_ASAP7_75t_L g1308 ( .A(n_1309), .B(n_1310), .Y(n_1308) );
INVx2_ASAP7_75t_L g1311 ( .A(n_1312), .Y(n_1311) );
OAI22xp5_ASAP7_75t_L g1342 ( .A1(n_1312), .A2(n_1343), .B1(n_1344), .B2(n_1345), .Y(n_1342) );
INVx1_ASAP7_75t_L g1507 ( .A(n_1312), .Y(n_1507) );
AND2x2_ASAP7_75t_L g1317 ( .A(n_1313), .B(n_1318), .Y(n_1317) );
AND2x2_ASAP7_75t_L g1334 ( .A(n_1313), .B(n_1335), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1313), .B(n_1410), .Y(n_1409) );
AND2x2_ASAP7_75t_L g1421 ( .A(n_1313), .B(n_1367), .Y(n_1421) );
NOR3xp33_ASAP7_75t_SL g1462 ( .A(n_1313), .B(n_1319), .C(n_1463), .Y(n_1462) );
OR2x2_ASAP7_75t_L g1474 ( .A(n_1313), .B(n_1367), .Y(n_1474) );
AND2x2_ASAP7_75t_L g1491 ( .A(n_1313), .B(n_1336), .Y(n_1491) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1315), .Y(n_1314) );
INVx1_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1322 ( .A(n_1319), .Y(n_1322) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1319), .B(n_1331), .Y(n_1369) );
AND2x2_ASAP7_75t_L g1370 ( .A(n_1319), .B(n_1371), .Y(n_1370) );
NAND2xp5_ASAP7_75t_L g1436 ( .A(n_1319), .B(n_1334), .Y(n_1436) );
AND2x2_ASAP7_75t_L g1447 ( .A(n_1319), .B(n_1409), .Y(n_1447) );
AND2x2_ASAP7_75t_L g1475 ( .A(n_1319), .B(n_1476), .Y(n_1475) );
NAND2xp5_ASAP7_75t_L g1321 ( .A(n_1322), .B(n_1323), .Y(n_1321) );
OAI211xp5_ASAP7_75t_L g1430 ( .A1(n_1324), .A2(n_1431), .B(n_1434), .C(n_1438), .Y(n_1430) );
INVx1_ASAP7_75t_L g1324 ( .A(n_1325), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1331 ( .A(n_1326), .B(n_1332), .Y(n_1331) );
OR2x2_ASAP7_75t_L g1337 ( .A(n_1326), .B(n_1332), .Y(n_1337) );
AOI22xp5_ASAP7_75t_L g1366 ( .A1(n_1326), .A2(n_1367), .B1(n_1368), .B2(n_1370), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1326), .B(n_1356), .Y(n_1378) );
OR2x2_ASAP7_75t_L g1389 ( .A(n_1326), .B(n_1355), .Y(n_1389) );
INVx2_ASAP7_75t_L g1413 ( .A(n_1326), .Y(n_1413) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1326), .B(n_1426), .Y(n_1425) );
OAI21xp5_ASAP7_75t_L g1445 ( .A1(n_1326), .A2(n_1446), .B(n_1448), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1456 ( .A(n_1326), .B(n_1355), .Y(n_1456) );
O2A1O1Ixp33_ASAP7_75t_L g1496 ( .A1(n_1326), .A2(n_1440), .B(n_1497), .C(n_1498), .Y(n_1496) );
AND2x4_ASAP7_75t_L g1326 ( .A(n_1327), .B(n_1328), .Y(n_1326) );
INVx1_ASAP7_75t_L g1329 ( .A(n_1330), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1373 ( .A(n_1331), .B(n_1374), .Y(n_1373) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1331), .B(n_1449), .Y(n_1448) );
INVx2_ASAP7_75t_SL g1393 ( .A(n_1332), .Y(n_1393) );
AND2x2_ASAP7_75t_L g1502 ( .A(n_1332), .B(n_1355), .Y(n_1502) );
INVx1_ASAP7_75t_L g1333 ( .A(n_1334), .Y(n_1333) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_1334), .B(n_1392), .Y(n_1418) );
INVx1_ASAP7_75t_L g1467 ( .A(n_1335), .Y(n_1467) );
INVx2_ASAP7_75t_L g1415 ( .A(n_1337), .Y(n_1415) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1353), .Y(n_1339) );
OAI21xp5_ASAP7_75t_L g1403 ( .A1(n_1340), .A2(n_1404), .B(n_1430), .Y(n_1403) );
NAND2xp5_ASAP7_75t_L g1453 ( .A(n_1340), .B(n_1413), .Y(n_1453) );
CKINVDCx5p33_ASAP7_75t_R g1340 ( .A(n_1341), .Y(n_1340) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1341), .B(n_1354), .Y(n_1376) );
AOI221xp5_ASAP7_75t_L g1444 ( .A1(n_1341), .A2(n_1445), .B1(n_1450), .B2(n_1452), .C(n_1454), .Y(n_1444) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1341), .Y(n_1487) );
OR2x6_ASAP7_75t_SL g1341 ( .A(n_1342), .B(n_1346), .Y(n_1341) );
OAI22xp5_ASAP7_75t_L g1346 ( .A1(n_1347), .A2(n_1348), .B1(n_1349), .B2(n_1350), .Y(n_1346) );
HB1xp67_ASAP7_75t_L g1350 ( .A(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1352), .Y(n_1351) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1353), .B(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_SL g1353 ( .A(n_1354), .Y(n_1353) );
NOR3xp33_ASAP7_75t_L g1484 ( .A(n_1354), .B(n_1432), .C(n_1485), .Y(n_1484) );
INVx3_ASAP7_75t_L g1354 ( .A(n_1355), .Y(n_1354) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1355), .Y(n_1394) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1355), .B(n_1413), .Y(n_1464) );
INVx3_ASAP7_75t_L g1355 ( .A(n_1356), .Y(n_1355) );
OR2x2_ASAP7_75t_L g1386 ( .A(n_1356), .B(n_1387), .Y(n_1386) );
OR2x2_ASAP7_75t_L g1356 ( .A(n_1357), .B(n_1360), .Y(n_1356) );
NOR2xp33_ASAP7_75t_L g1364 ( .A(n_1365), .B(n_1388), .Y(n_1364) );
A2O1A1Ixp33_ASAP7_75t_L g1365 ( .A1(n_1366), .A2(n_1372), .B(n_1376), .C(n_1377), .Y(n_1365) );
INVx1_ASAP7_75t_L g1368 ( .A(n_1369), .Y(n_1368) );
AOI22xp5_ASAP7_75t_L g1377 ( .A1(n_1370), .A2(n_1378), .B1(n_1379), .B2(n_1385), .Y(n_1377) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1371), .B(n_1423), .Y(n_1422) );
INVxp67_ASAP7_75t_L g1372 ( .A(n_1373), .Y(n_1372) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
INVx1_ASAP7_75t_L g1424 ( .A(n_1378), .Y(n_1424) );
AND2x2_ASAP7_75t_L g1459 ( .A(n_1378), .B(n_1393), .Y(n_1459) );
AND2x2_ASAP7_75t_L g1379 ( .A(n_1380), .B(n_1381), .Y(n_1379) );
INVx1_ASAP7_75t_L g1503 ( .A(n_1381), .Y(n_1503) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1382), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1383), .B(n_1384), .Y(n_1382) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1384), .Y(n_1433) );
INVx1_ASAP7_75t_L g1385 ( .A(n_1386), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1478 ( .A(n_1386), .B(n_1467), .Y(n_1478) );
INVx1_ASAP7_75t_L g1476 ( .A(n_1387), .Y(n_1476) );
A2O1A1Ixp33_ASAP7_75t_L g1388 ( .A1(n_1389), .A2(n_1390), .B(n_1395), .C(n_1396), .Y(n_1388) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1389), .Y(n_1417) );
INVxp67_ASAP7_75t_SL g1390 ( .A(n_1391), .Y(n_1390) );
OAI21xp5_ASAP7_75t_L g1434 ( .A1(n_1391), .A2(n_1435), .B(n_1437), .Y(n_1434) );
AND2x2_ASAP7_75t_L g1391 ( .A(n_1392), .B(n_1394), .Y(n_1391) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1393), .Y(n_1401) );
INVx1_ASAP7_75t_L g1440 ( .A(n_1393), .Y(n_1440) );
NAND2xp5_ASAP7_75t_L g1414 ( .A(n_1394), .B(n_1415), .Y(n_1414) );
AND2x2_ASAP7_75t_L g1495 ( .A(n_1394), .B(n_1476), .Y(n_1495) );
OAI22xp5_ASAP7_75t_L g1501 ( .A1(n_1395), .A2(n_1502), .B1(n_1503), .B2(n_1504), .Y(n_1501) );
AND2x2_ASAP7_75t_L g1397 ( .A(n_1398), .B(n_1402), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1399), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1494 ( .A(n_1399), .B(n_1432), .Y(n_1494) );
NAND2xp5_ASAP7_75t_L g1399 ( .A(n_1400), .B(n_1401), .Y(n_1399) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_1400), .B(n_1413), .Y(n_1412) );
INVx2_ASAP7_75t_L g1423 ( .A(n_1400), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1460 ( .A(n_1400), .B(n_1461), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1406), .B(n_1408), .Y(n_1405) );
INVx1_ASAP7_75t_L g1406 ( .A(n_1407), .Y(n_1406) );
OAI221xp5_ASAP7_75t_L g1479 ( .A1(n_1408), .A2(n_1455), .B1(n_1463), .B2(n_1480), .C(n_1483), .Y(n_1479) );
INVx1_ASAP7_75t_L g1408 ( .A(n_1409), .Y(n_1408) );
OAI21xp5_ASAP7_75t_SL g1472 ( .A1(n_1409), .A2(n_1473), .B(n_1475), .Y(n_1472) );
INVx1_ASAP7_75t_L g1432 ( .A(n_1410), .Y(n_1432) );
INVxp67_ASAP7_75t_SL g1411 ( .A(n_1412), .Y(n_1411) );
INVx1_ASAP7_75t_L g1505 ( .A(n_1413), .Y(n_1505) );
OAI211xp5_ASAP7_75t_L g1489 ( .A1(n_1414), .A2(n_1490), .B(n_1492), .C(n_1493), .Y(n_1489) );
NAND3xp33_ASAP7_75t_L g1469 ( .A(n_1415), .B(n_1470), .C(n_1471), .Y(n_1469) );
AOI211xp5_ASAP7_75t_L g1416 ( .A1(n_1417), .A2(n_1418), .B(n_1419), .C(n_1429), .Y(n_1416) );
A2O1A1Ixp33_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1422), .B(n_1424), .C(n_1425), .Y(n_1419) );
NOR2xp33_ASAP7_75t_L g1426 ( .A(n_1427), .B(n_1428), .Y(n_1426) );
INVx1_ASAP7_75t_L g1471 ( .A(n_1427), .Y(n_1471) );
OR2x2_ASAP7_75t_L g1431 ( .A(n_1432), .B(n_1433), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1466 ( .A(n_1432), .B(n_1467), .Y(n_1466) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1497 ( .A(n_1437), .Y(n_1497) );
INVx1_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
NOR2xp33_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
NAND3xp33_ASAP7_75t_L g1443 ( .A(n_1444), .B(n_1477), .C(n_1488), .Y(n_1443) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1447), .Y(n_1446) );
INVx1_ASAP7_75t_L g1450 ( .A(n_1451), .Y(n_1450) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OAI211xp5_ASAP7_75t_L g1454 ( .A1(n_1455), .A2(n_1457), .B(n_1458), .C(n_1472), .Y(n_1454) );
INVx1_ASAP7_75t_L g1455 ( .A(n_1456), .Y(n_1455) );
AOI221xp5_ASAP7_75t_L g1458 ( .A1(n_1459), .A2(n_1460), .B1(n_1462), .B2(n_1465), .C(n_1468), .Y(n_1458) );
INVx1_ASAP7_75t_L g1463 ( .A(n_1464), .Y(n_1463) );
INVx1_ASAP7_75t_L g1465 ( .A(n_1466), .Y(n_1465) );
INVx1_ASAP7_75t_SL g1468 ( .A(n_1469), .Y(n_1468) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1474), .Y(n_1473) );
INVxp67_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
OAI31xp33_ASAP7_75t_SL g1488 ( .A1(n_1486), .A2(n_1489), .A3(n_1496), .B(n_1501), .Y(n_1488) );
CKINVDCx14_ASAP7_75t_R g1486 ( .A(n_1487), .Y(n_1486) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1499 ( .A(n_1500), .Y(n_1499) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
HB1xp67_ASAP7_75t_L g1508 ( .A(n_1509), .Y(n_1508) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1511), .Y(n_1510) );
AND2x2_ASAP7_75t_L g1511 ( .A(n_1512), .B(n_1539), .Y(n_1511) );
AOI21xp5_ASAP7_75t_L g1512 ( .A1(n_1513), .A2(n_1514), .B(n_1515), .Y(n_1512) );
AOI211xp5_ASAP7_75t_L g1516 ( .A1(n_1517), .A2(n_1518), .B(n_1519), .C(n_1528), .Y(n_1516) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
OAI221xp5_ASAP7_75t_L g1522 ( .A1(n_1523), .A2(n_1524), .B1(n_1525), .B2(n_1526), .C(n_1527), .Y(n_1522) );
NOR3xp33_ASAP7_75t_L g1539 ( .A(n_1540), .B(n_1545), .C(n_1546), .Y(n_1539) );
NAND2xp5_ASAP7_75t_L g1540 ( .A(n_1541), .B(n_1543), .Y(n_1540) );
INVx1_ASAP7_75t_L g1551 ( .A(n_1552), .Y(n_1551) );
INVx4_ASAP7_75t_SL g1558 ( .A(n_1559), .Y(n_1558) );
BUFx3_ASAP7_75t_L g1559 ( .A(n_1560), .Y(n_1559) );
BUFx2_ASAP7_75t_L g1560 ( .A(n_1561), .Y(n_1560) );
INVx2_ASAP7_75t_L g1563 ( .A(n_1564), .Y(n_1563) );
CKINVDCx5p33_ASAP7_75t_R g1564 ( .A(n_1565), .Y(n_1564) );
A2O1A1Ixp33_ASAP7_75t_L g1571 ( .A1(n_1566), .A2(n_1572), .B(n_1574), .C(n_1576), .Y(n_1571) );
INVxp33_ASAP7_75t_SL g1567 ( .A(n_1568), .Y(n_1567) );
HB1xp67_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1573), .Y(n_1572) );
INVx1_ASAP7_75t_L g1574 ( .A(n_1575), .Y(n_1574) );
endmodule