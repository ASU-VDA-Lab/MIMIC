module fake_jpeg_6055_n_105 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_105);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_105;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_33),
.Y(n_44)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_8),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_14),
.Y(n_48)
);

BUFx4f_ASAP7_75t_L g49 ( 
.A(n_7),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_3),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_12),
.Y(n_51)
);

INVx13_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_39),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_19),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_25),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_40),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_22),
.Y(n_60)
);

BUFx12f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

CKINVDCx14_ASAP7_75t_R g62 ( 
.A(n_23),
.Y(n_62)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

INVx5_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_64),
.B(n_65),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_48),
.Y(n_65)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_52),
.Y(n_66)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_66),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_53),
.A2(n_21),
.B(n_42),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_67),
.Y(n_71)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_68),
.Y(n_74)
);

OAI22xp33_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_49),
.B1(n_51),
.B2(n_57),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_50),
.B1(n_55),
.B2(n_62),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_66),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_75),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_69),
.A2(n_45),
.B1(n_46),
.B2(n_59),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_76),
.A2(n_60),
.B1(n_58),
.B2(n_43),
.Y(n_88)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_78),
.B(n_79),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_70),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_80),
.A2(n_56),
.B1(n_70),
.B2(n_74),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_83),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_88),
.B1(n_61),
.B2(n_0),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_77),
.A2(n_74),
.B1(n_47),
.B2(n_54),
.Y(n_83)
);

A2O1A1Ixp33_ASAP7_75t_L g85 ( 
.A1(n_77),
.A2(n_71),
.B(n_1),
.C(n_2),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_86),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_80),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_87),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_61),
.C(n_24),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_92),
.B(n_93),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_91),
.A2(n_84),
.B(n_75),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_94),
.A2(n_89),
.B1(n_90),
.B2(n_0),
.Y(n_96)
);

A2O1A1O1Ixp25_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_95),
.B(n_1),
.C(n_5),
.D(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_98),
.B(n_4),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_99),
.A2(n_9),
.B(n_13),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_15),
.C(n_16),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_17),
.Y(n_102)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_102),
.A2(n_18),
.A3(n_20),
.B1(n_26),
.B2(n_27),
.C1(n_28),
.C2(n_29),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_103),
.A2(n_30),
.B1(n_31),
.B2(n_35),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_104),
.B(n_37),
.Y(n_105)
);


endmodule