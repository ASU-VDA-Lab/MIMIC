module real_jpeg_30035_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_271;
wire n_131;
wire n_281;
wire n_276;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_160;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_262;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_195;
wire n_61;
wire n_110;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_277;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_191;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_279;
wire n_59;
wire n_169;
wire n_216;
wire n_128;
wire n_167;
wire n_179;
wire n_202;
wire n_213;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;

OAI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_0),
.A2(n_27),
.B1(n_29),
.B2(n_42),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_0),
.Y(n_42)
);

AOI22xp33_ASAP7_75t_L g87 ( 
.A1(n_0),
.A2(n_42),
.B1(n_80),
.B2(n_81),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g94 ( 
.A1(n_0),
.A2(n_32),
.B1(n_35),
.B2(n_42),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_L g101 ( 
.A1(n_0),
.A2(n_42),
.B1(n_48),
.B2(n_49),
.Y(n_101)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_1),
.Y(n_65)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_1),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g123 ( 
.A(n_1),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_2),
.A2(n_48),
.B1(n_49),
.B2(n_55),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_2),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_2),
.A2(n_27),
.B1(n_29),
.B2(n_55),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_2),
.A2(n_32),
.B1(n_35),
.B2(n_55),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_3),
.A2(n_80),
.B1(n_81),
.B2(n_133),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_3),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_3),
.A2(n_48),
.B1(n_49),
.B2(n_133),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_3),
.A2(n_27),
.B1(n_29),
.B2(n_133),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_3),
.A2(n_32),
.B1(n_35),
.B2(n_133),
.Y(n_231)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_4),
.A2(n_48),
.B1(n_49),
.B2(n_57),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_4),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_4),
.A2(n_27),
.B1(n_29),
.B2(n_57),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_4),
.A2(n_32),
.B1(n_35),
.B2(n_57),
.Y(n_119)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_6),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_6),
.B(n_83),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_6),
.B(n_48),
.Y(n_191)
);

AOI21xp33_ASAP7_75t_L g195 ( 
.A1(n_6),
.A2(n_48),
.B(n_191),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g215 ( 
.A1(n_6),
.A2(n_27),
.B1(n_29),
.B2(n_151),
.Y(n_215)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_6),
.A2(n_32),
.B(n_36),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_6),
.B(n_99),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_6),
.A2(n_62),
.B1(n_65),
.B2(n_239),
.Y(n_241)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_8),
.A2(n_80),
.B1(n_81),
.B2(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_8),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_8),
.A2(n_48),
.B1(n_49),
.B2(n_106),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_8),
.A2(n_27),
.B1(n_29),
.B2(n_106),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_8),
.A2(n_32),
.B1(n_35),
.B2(n_106),
.Y(n_226)
);

INVx13_ASAP7_75t_L g81 ( 
.A(n_9),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_10),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_10),
.A2(n_28),
.B1(n_32),
.B2(n_35),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_10),
.A2(n_28),
.B1(n_80),
.B2(n_81),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_10),
.A2(n_28),
.B1(n_48),
.B2(n_49),
.Y(n_128)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_11),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_12),
.A2(n_80),
.B1(n_81),
.B2(n_153),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_12),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_12),
.A2(n_48),
.B1(n_49),
.B2(n_153),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_12),
.A2(n_27),
.B1(n_29),
.B2(n_153),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_12),
.A2(n_32),
.B1(n_35),
.B2(n_153),
.Y(n_239)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_13),
.Y(n_50)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_14),
.Y(n_47)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_15),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_135),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_134),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_19),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_20),
.B(n_109),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_20),
.B(n_109),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_89),
.B2(n_108),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_59),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_43),
.B(n_58),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_24),
.B(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_37),
.Y(n_24)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_25),
.A2(n_39),
.B(n_199),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_30),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_26),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_27),
.Y(n_29)
);

OAI22xp33_ASAP7_75t_L g40 ( 
.A1(n_27),
.A2(n_29),
.B1(n_34),
.B2(n_36),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_27),
.A2(n_29),
.B1(n_46),
.B2(n_51),
.Y(n_52)
);

NAND2xp33_ASAP7_75t_SL g192 ( 
.A(n_27),
.B(n_46),
.Y(n_192)
);

A2O1A1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_27),
.A2(n_34),
.B(n_151),
.C(n_218),
.Y(n_217)
);

AOI32xp33_ASAP7_75t_L g189 ( 
.A1(n_29),
.A2(n_49),
.A3(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g73 ( 
.A(n_30),
.B(n_41),
.Y(n_73)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_31),
.A2(n_39),
.B1(n_72),
.B2(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_31),
.A2(n_37),
.B(n_97),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_31),
.A2(n_39),
.B1(n_198),
.B2(n_199),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_31),
.A2(n_39),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_31),
.A2(n_39),
.B1(n_198),
.B2(n_216),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_31),
.B(n_151),
.Y(n_237)
);

OA22x2_ASAP7_75t_L g31 ( 
.A1(n_32),
.A2(n_34),
.B1(n_35),
.B2(n_36),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_32),
.Y(n_35)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_35),
.B(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_SL g37 ( 
.A(n_38),
.B(n_41),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_72),
.B(n_73),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_SL g143 ( 
.A1(n_39),
.A2(n_73),
.B(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_44),
.A2(n_52),
.B1(n_53),
.B2(n_56),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_44),
.B(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_44),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_44),
.A2(n_52),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_44),
.A2(n_52),
.B1(n_147),
.B2(n_177),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_44),
.A2(n_52),
.B1(n_177),
.B2(n_195),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_45),
.B(n_52),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B1(n_49),
.B2(n_51),
.Y(n_45)
);

INVx6_ASAP7_75t_L g190 ( 
.A(n_46),
.Y(n_190)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_48),
.A2(n_49),
.B1(n_78),
.B2(n_79),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_48),
.B(n_78),
.Y(n_165)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_49),
.A2(n_82),
.B1(n_150),
.B2(n_165),
.Y(n_164)
);

INVx11_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_52),
.B(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_52),
.B(n_128),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g53 ( 
.A(n_54),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_54),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_74),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_71),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_61),
.A2(n_75),
.B1(n_76),
.B2(n_88),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_61),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_61),
.A2(n_71),
.B1(n_88),
.B2(n_115),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_66),
.B(n_69),
.Y(n_61)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_62),
.A2(n_119),
.B(n_120),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_62),
.A2(n_119),
.B1(n_167),
.B2(n_168),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_62),
.A2(n_95),
.B(n_226),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_62),
.A2(n_65),
.B1(n_231),
.B2(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_63),
.B(n_93),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_63),
.A2(n_70),
.B(n_121),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_63),
.A2(n_67),
.B1(n_230),
.B2(n_232),
.Y(n_229)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_65),
.B(n_151),
.Y(n_243)
);

INVx5_ASAP7_75t_SL g66 ( 
.A(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_67),
.B(n_70),
.Y(n_95)
);

INVx11_ASAP7_75t_L g168 ( 
.A(n_67),
.Y(n_168)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_71),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_L g76 ( 
.A1(n_77),
.A2(n_84),
.B(n_85),
.Y(n_76)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_77),
.A2(n_83),
.B1(n_150),
.B2(n_152),
.Y(n_149)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_78),
.A2(n_80),
.B(n_82),
.C(n_83),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_78),
.B(n_80),
.Y(n_82)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

HAxp5_ASAP7_75t_SL g150 ( 
.A(n_80),
.B(n_151),
.CON(n_150),
.SN(n_150)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_83),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_83),
.B(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_86),
.B(n_87),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_86),
.A2(n_104),
.B1(n_105),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_86),
.A2(n_104),
.B1(n_132),
.B2(n_158),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_89),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_98),
.C(n_102),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_90),
.B(n_112),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_96),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_91),
.B(n_96),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_95),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_92),
.A2(n_167),
.B(n_168),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_122),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_98),
.A2(n_102),
.B1(n_103),
.B2(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_98),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_104),
.A2(n_105),
.B(n_107),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_114),
.C(n_116),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_110),
.A2(n_111),
.B1(n_114),
.B2(n_280),
.Y(n_279)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_114),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_116),
.B(n_279),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_125),
.C(n_130),
.Y(n_116)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_117),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_124),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_124),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_121),
.Y(n_120)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g271 ( 
.A1(n_125),
.A2(n_130),
.B1(n_131),
.B2(n_272),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_125),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B(n_129),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_126),
.A2(n_161),
.B(n_162),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_276),
.B(n_281),
.Y(n_135)
);

O2A1O1Ixp33_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_181),
.B(n_262),
.C(n_275),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_169),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_138),
.B(n_169),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_154),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_140),
.B(n_141),
.C(n_154),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_145),
.C(n_149),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_142),
.A2(n_143),
.B1(n_145),
.B2(n_146),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_146),
.Y(n_145)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_148),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_SL g171 ( 
.A(n_149),
.B(n_172),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_152),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g154 ( 
.A(n_155),
.B(n_163),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_156),
.A2(n_157),
.B1(n_159),
.B2(n_160),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_156),
.B(n_160),
.C(n_163),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_164),
.B(n_166),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_173),
.C(n_175),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_170),
.A2(n_171),
.B1(n_257),
.B2(n_259),
.Y(n_256)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g257 ( 
.A1(n_173),
.A2(n_174),
.B1(n_175),
.B2(n_258),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_174),
.Y(n_173)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_175),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_178),
.C(n_180),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_176),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_204),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_180),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_182),
.B(n_261),
.Y(n_181)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_183),
.A2(n_254),
.B(n_260),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_209),
.B(n_253),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_200),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_185),
.B(n_200),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_193),
.C(n_196),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_186),
.A2(n_187),
.B1(n_250),
.B2(n_251),
.Y(n_249)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_189),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_193),
.A2(n_194),
.B1(n_196),
.B2(n_197),
.Y(n_251)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_194),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_255)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_210),
.A2(n_247),
.B(n_252),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_227),
.B(n_246),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_219),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_212),
.B(n_219),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_213),
.A2(n_214),
.B1(n_217),
.B2(n_234),
.Y(n_233)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_217),
.Y(n_234)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_221),
.A2(n_222),
.B1(n_223),
.B2(n_224),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_221),
.B(n_224),
.C(n_225),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g223 ( 
.A(n_224),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_226),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_235),
.B(n_245),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_233),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_229),
.B(n_233),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_240),
.B(n_244),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_238),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_237),
.B(n_238),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_248),
.B(n_249),
.Y(n_252)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_SL g260 ( 
.A(n_255),
.B(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_257),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_263),
.B(n_264),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_265),
.A2(n_266),
.B1(n_273),
.B2(n_274),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_269),
.B2(n_270),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_270),
.C(n_274),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_277),
.B(n_278),
.Y(n_281)
);


endmodule