module fake_jpeg_15546_n_22 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_22);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_22;

wire n_13;
wire n_21;
wire n_10;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_16;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

AOI22xp33_ASAP7_75t_L g10 ( 
.A1(n_5),
.A2(n_8),
.B1(n_2),
.B2(n_0),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_6),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_1),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_16),
.C(n_12),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g15 ( 
.A1(n_10),
.A2(n_0),
.B(n_1),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_15),
.A2(n_13),
.B1(n_11),
.B2(n_10),
.Y(n_17)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_12),
.B(n_2),
.C(n_3),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_17),
.A2(n_11),
.B1(n_4),
.B2(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g19 ( 
.A(n_18),
.B(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_20),
.Y(n_21)
);

MAJx2_ASAP7_75t_L g22 ( 
.A(n_21),
.B(n_20),
.C(n_9),
.Y(n_22)
);


endmodule