module fake_jpeg_20386_n_100 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_91;
wire n_54;
wire n_93;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_28),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_30),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_2),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_25),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_24),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_34),
.Y(n_41)
);

INVx8_ASAP7_75t_SL g42 ( 
.A(n_20),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_27),
.Y(n_43)
);

AOI21xp33_ASAP7_75t_L g44 ( 
.A1(n_13),
.A2(n_3),
.B(n_6),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_47),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_39),
.B1(n_44),
.B2(n_6),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_41),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_49),
.B(n_50),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g50 ( 
.A(n_36),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_0),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_51),
.B(n_52),
.Y(n_56)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_3),
.Y(n_53)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_53),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_4),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_54),
.Y(n_63)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_57),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_41),
.B1(n_39),
.B2(n_38),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_58),
.B(n_62),
.Y(n_74)
);

BUFx24_ASAP7_75t_L g60 ( 
.A(n_50),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g77 ( 
.A(n_60),
.Y(n_77)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_64),
.B(n_37),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_65),
.Y(n_69)
);

NOR2x1_ASAP7_75t_SL g79 ( 
.A(n_66),
.B(n_5),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_55),
.B(n_63),
.C(n_60),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_72),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_56),
.Y(n_70)
);

NAND3xp33_ASAP7_75t_L g81 ( 
.A(n_70),
.B(n_71),
.C(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_64),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_73),
.B(n_76),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_4),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_63),
.B(n_43),
.Y(n_76)
);

OAI22xp33_ASAP7_75t_SL g78 ( 
.A1(n_69),
.A2(n_40),
.B1(n_35),
.B2(n_5),
.Y(n_78)
);

INVxp67_ASAP7_75t_L g88 ( 
.A(n_78),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_79),
.B(n_83),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g80 ( 
.A(n_74),
.Y(n_80)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g83 ( 
.A1(n_74),
.A2(n_17),
.B1(n_8),
.B2(n_10),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_76),
.A2(n_19),
.B1(n_11),
.B2(n_12),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_66),
.C(n_67),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_84),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_87),
.A2(n_90),
.B1(n_77),
.B2(n_85),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_89),
.A2(n_80),
.B1(n_82),
.B2(n_81),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_91),
.B(n_92),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_91),
.C(n_86),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_88),
.B(n_14),
.Y(n_96)
);

AOI322xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_88),
.A3(n_15),
.B1(n_16),
.B2(n_18),
.C1(n_21),
.C2(n_23),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_26),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_29),
.B(n_31),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_33),
.C(n_7),
.Y(n_100)
);


endmodule