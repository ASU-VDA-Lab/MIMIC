module real_jpeg_26106_n_11 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_10, n_9, n_11);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_11;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_78;
wire n_83;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_208;
wire n_62;
wire n_239;
wire n_162;
wire n_245;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_203;
wire n_198;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_12;
wire n_124;
wire n_24;
wire n_92;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_169;
wire n_88;
wire n_59;
wire n_128;
wire n_244;
wire n_202;
wire n_179;
wire n_167;
wire n_213;
wire n_133;
wire n_216;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_1),
.A2(n_20),
.B1(n_24),
.B2(n_46),
.Y(n_45)
);

CKINVDCx16_ASAP7_75t_R g46 ( 
.A(n_1),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_1),
.A2(n_37),
.B1(n_38),
.B2(n_46),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_1),
.A2(n_46),
.B1(n_54),
.B2(n_55),
.Y(n_117)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_2),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_60),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_5),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_5),
.A2(n_54),
.B1(n_55),
.B2(n_60),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_5),
.A2(n_20),
.B1(n_24),
.B2(n_60),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_6),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_6),
.A2(n_20),
.B1(n_24),
.B2(n_30),
.Y(n_43)
);

OAI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_6),
.A2(n_30),
.B1(n_37),
.B2(n_38),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_6),
.A2(n_30),
.B1(n_54),
.B2(n_55),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_6),
.B(n_20),
.C(n_23),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_6),
.B(n_171),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_6),
.B(n_36),
.C(n_38),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_6),
.B(n_52),
.C(n_55),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_6),
.B(n_95),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_6),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_6),
.B(n_71),
.Y(n_206)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_10),
.Y(n_82)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_10),
.Y(n_83)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_10),
.Y(n_118)
);

XOR2xp5_ASAP7_75t_L g11 ( 
.A(n_12),
.B(n_101),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_99),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_87),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_14),
.B(n_87),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_62),
.C(n_73),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_15),
.A2(n_62),
.B1(n_63),
.B2(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_15),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_17),
.B1(n_31),
.B2(n_32),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_16),
.B(n_33),
.C(n_48),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_16),
.A2(n_17),
.B1(n_90),
.B2(n_98),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_16),
.A2(n_17),
.B1(n_91),
.B2(n_97),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_16),
.A2(n_17),
.B1(n_76),
.B2(n_77),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_16),
.B(n_64),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_16),
.A2(n_17),
.B1(n_64),
.B2(n_65),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_16),
.A2(n_17),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI21xp5_ASAP7_75t_L g73 ( 
.A1(n_17),
.A2(n_74),
.B(n_77),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_17),
.B(n_65),
.Y(n_120)
);

AOI211xp5_ASAP7_75t_L g150 ( 
.A1(n_17),
.A2(n_119),
.B(n_122),
.C(n_151),
.Y(n_150)
);

AND2x2_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_29),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_25),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_SL g25 ( 
.A(n_19),
.B(n_26),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_19),
.Y(n_171)
);

OA22x2_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_20),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_20),
.A2(n_24),
.B1(n_36),
.B2(n_40),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_20),
.B(n_182),
.Y(n_181)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_22),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_26)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_27),
.Y(n_28)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_27),
.Y(n_158)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_47),
.B1(n_48),
.B2(n_61),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_34),
.A2(n_35),
.B1(n_42),
.B2(n_44),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_34),
.B(n_35),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_34),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_41),
.Y(n_34)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_35),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_35)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_L g58 ( 
.A1(n_37),
.A2(n_38),
.B1(n_52),
.B2(n_53),
.Y(n_58)
);

INVx5_ASAP7_75t_SL g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_38),
.B(n_193),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVxp67_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_43),
.B(n_66),
.Y(n_65)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g93 ( 
.A1(n_45),
.A2(n_94),
.B1(n_95),
.B2(n_96),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_47),
.A2(n_48),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_59),
.Y(n_48)
);

INVxp33_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g119 ( 
.A(n_50),
.B(n_86),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_51),
.B(n_58),
.Y(n_57)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_51),
.A2(n_57),
.B1(n_69),
.B2(n_85),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_53),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_55),
.B(n_203),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_64),
.B(n_67),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_64),
.B(n_149),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_64),
.A2(n_65),
.B1(n_119),
.B2(n_149),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_64),
.A2(n_65),
.B1(n_177),
.B2(n_178),
.Y(n_176)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_65),
.B(n_154),
.C(n_169),
.Y(n_168)
);

O2A1O1Ixp33_ASAP7_75t_L g217 ( 
.A1(n_65),
.A2(n_119),
.B(n_151),
.C(n_214),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_73),
.B(n_243),
.Y(n_242)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_74),
.A2(n_75),
.B1(n_109),
.B2(n_110),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_76),
.B(n_84),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_76),
.A2(n_77),
.B1(n_84),
.B2(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_79),
.A2(n_81),
.B1(n_117),
.B2(n_118),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_137),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_81),
.B(n_83),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_81),
.A2(n_117),
.B1(n_136),
.B2(n_138),
.Y(n_135)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_83),
.Y(n_204)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_84),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

XNOR2xp5_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_89),
.Y(n_87)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_93),
.Y(n_92)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_240),
.B(n_246),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_141),
.B(n_239),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_105),
.B(n_124),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_105),
.B(n_124),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_106),
.A2(n_113),
.B1(n_114),
.B2(n_123),
.Y(n_105)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_106),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_108),
.B1(n_111),
.B2(n_112),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_108),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_108),
.B(n_111),
.C(n_113),
.Y(n_245)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_112),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_115),
.A2(n_120),
.B(n_121),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_115),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_115),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_116),
.B(n_119),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_116),
.A2(n_119),
.B1(n_149),
.B2(n_230),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_116),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_119),
.B(n_135),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_119),
.A2(n_135),
.B1(n_148),
.B2(n_149),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_119),
.B(n_191),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_119),
.A2(n_149),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_119),
.A2(n_149),
.B1(n_191),
.B2(n_192),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_119),
.A2(n_149),
.B1(n_179),
.B2(n_220),
.Y(n_219)
);

CKINVDCx14_ASAP7_75t_R g140 ( 
.A(n_120),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_120),
.A2(n_121),
.B(n_153),
.Y(n_231)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g132 ( 
.A1(n_122),
.A2(n_133),
.B(n_140),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_130),
.C(n_132),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_125),
.A2(n_126),
.B1(n_130),
.B2(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_127),
.A2(n_128),
.B1(n_153),
.B2(n_160),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_127),
.A2(n_128),
.B1(n_133),
.B2(n_134),
.Y(n_228)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_130),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_132),
.B(n_235),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_135),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_233),
.B(n_238),
.Y(n_141)
);

A2O1A1Ixp33_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_172),
.B(n_224),
.C(n_232),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_162),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_144),
.B(n_162),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_145),
.A2(n_146),
.B1(n_152),
.B2(n_161),
.Y(n_144)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_150),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_147),
.B(n_150),
.C(n_161),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_149),
.B(n_176),
.C(n_179),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_149),
.B(n_155),
.C(n_198),
.Y(n_211)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_152),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_156),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_154),
.A2(n_155),
.B1(n_156),
.B2(n_157),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_154),
.A2(n_155),
.B1(n_169),
.B2(n_170),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_154),
.B(n_180),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_154),
.A2(n_155),
.B1(n_195),
.B2(n_196),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_154),
.B(n_208),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_154),
.A2(n_155),
.B1(n_180),
.B2(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_155),
.B(n_202),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_155),
.B(n_206),
.Y(n_205)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_159),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.C(n_167),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_184),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_164),
.A2(n_165),
.B1(n_213),
.B2(n_214),
.Y(n_212)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_185),
.Y(n_184)
);

CKINVDCx14_ASAP7_75t_R g185 ( 
.A(n_166),
.Y(n_185)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_173),
.B(n_223),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_186),
.B(n_222),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_183),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g222 ( 
.A(n_175),
.B(n_183),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g218 ( 
.A(n_176),
.B(n_219),
.Y(n_218)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_179),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_181),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_216),
.B(n_221),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_188),
.A2(n_210),
.B(n_215),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_199),
.B(n_209),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_194),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_190),
.B(n_194),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_207),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_212),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_211),
.B(n_212),
.Y(n_215)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_217),
.B(n_218),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_217),
.B(n_218),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_226),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_231),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_228),
.B(n_229),
.C(n_231),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_237),
.Y(n_238)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_241),
.Y(n_240)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_242),
.B(n_245),
.Y(n_246)
);


endmodule