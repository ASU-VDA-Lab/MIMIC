module fake_jpeg_7887_n_279 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_279);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_279;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_57;
wire n_21;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_122;
wire n_75;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

INVx1_ASAP7_75t_L g17 ( 
.A(n_16),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_2),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

INVx11_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx10_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

INVx3_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_7),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_7),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_31),
.B(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_35),
.B(n_41),
.Y(n_51)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_36),
.Y(n_69)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_19),
.Y(n_37)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_24),
.B(n_0),
.C(n_1),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_38),
.B(n_17),
.C(n_28),
.Y(n_70)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_39),
.B(n_23),
.Y(n_63)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_19),
.Y(n_40)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_31),
.B(n_16),
.Y(n_41)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g53 ( 
.A(n_43),
.Y(n_53)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_44),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_23),
.B(n_16),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_45),
.B(n_17),
.Y(n_64)
);

BUFx4f_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_49),
.Y(n_74)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_50),
.B(n_52),
.Y(n_86)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_54),
.A2(n_68),
.B1(n_42),
.B2(n_20),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g72 ( 
.A(n_55),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_35),
.B(n_18),
.Y(n_56)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_56),
.Y(n_91)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_33),
.B1(n_23),
.B2(n_25),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_58),
.A2(n_20),
.B1(n_28),
.B2(n_34),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_41),
.B(n_18),
.Y(n_59)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_60),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_45),
.B(n_32),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_61),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

BUFx2_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_63),
.A2(n_66),
.B(n_24),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_64),
.B(n_65),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_30),
.Y(n_65)
);

OR2x4_ASAP7_75t_L g66 ( 
.A(n_38),
.B(n_24),
.Y(n_66)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_44),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_67),
.B(n_49),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_44),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_70),
.B(n_17),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_63),
.B(n_70),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_71),
.A2(n_73),
.B(n_80),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_48),
.A2(n_42),
.B1(n_33),
.B2(n_22),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_79),
.A2(n_81),
.B1(n_82),
.B2(n_90),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_48),
.A2(n_33),
.B1(n_25),
.B2(n_22),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_54),
.A2(n_22),
.B1(n_25),
.B2(n_20),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_83),
.A2(n_84),
.B1(n_57),
.B2(n_52),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_47),
.A2(n_28),
.B1(n_34),
.B2(n_32),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_64),
.B(n_29),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_85),
.B(n_87),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_51),
.B(n_29),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_47),
.A2(n_43),
.B1(n_36),
.B2(n_39),
.Y(n_90)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_86),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g140 ( 
.A(n_94),
.B(n_96),
.Y(n_140)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_86),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_85),
.B(n_51),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_97),
.B(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_34),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_76),
.B(n_30),
.Y(n_100)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_100),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_0),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_101),
.B(n_102),
.Y(n_130)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_90),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_80),
.B(n_49),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_112),
.Y(n_123)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_105),
.B(n_106),
.Y(n_131)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_78),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_107),
.B(n_110),
.Y(n_134)
);

AOI32xp33_ASAP7_75t_L g108 ( 
.A1(n_71),
.A2(n_53),
.A3(n_67),
.B1(n_43),
.B2(n_36),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g133 ( 
.A1(n_108),
.A2(n_118),
.B(n_74),
.C(n_88),
.Y(n_133)
);

AOI21xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_73),
.B(n_93),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g143 ( 
.A1(n_109),
.A2(n_117),
.B(n_88),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_89),
.B(n_2),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_81),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_111),
.B(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_73),
.B(n_50),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_78),
.A2(n_69),
.B1(n_53),
.B2(n_39),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_78),
.B1(n_69),
.B2(n_74),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_89),
.B(n_3),
.Y(n_116)
);

AOI32xp33_ASAP7_75t_L g118 ( 
.A1(n_73),
.A2(n_67),
.A3(n_60),
.B1(n_62),
.B2(n_29),
.Y(n_118)
);

OAI21xp33_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_92),
.B(n_91),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_SL g149 ( 
.A(n_119),
.B(n_125),
.C(n_133),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_120),
.A2(n_137),
.B1(n_141),
.B2(n_143),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_106),
.A2(n_46),
.B1(n_74),
.B2(n_91),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_121),
.A2(n_128),
.B1(n_98),
.B2(n_104),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_114),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_122),
.B(n_136),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_113),
.B(n_67),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_112),
.Y(n_146)
);

NOR2x1_ASAP7_75t_R g125 ( 
.A(n_108),
.B(n_29),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_95),
.B(n_99),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_127),
.B(n_132),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_105),
.A2(n_102),
.B1(n_111),
.B2(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_92),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g135 ( 
.A(n_118),
.B(n_4),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_135),
.A2(n_139),
.B(n_116),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_97),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_96),
.B(n_4),
.Y(n_139)
);

INVx4_ASAP7_75t_SL g141 ( 
.A(n_107),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_142),
.B(n_46),
.Y(n_168)
);

INVx13_ASAP7_75t_L g144 ( 
.A(n_115),
.Y(n_144)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_144),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_146),
.B(n_21),
.C(n_27),
.Y(n_195)
);

AOI21xp5_ASAP7_75t_SL g147 ( 
.A1(n_143),
.A2(n_113),
.B(n_109),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_SL g194 ( 
.A(n_147),
.B(n_155),
.Y(n_194)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_148),
.B(n_150),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_140),
.Y(n_150)
);

AOI21xp33_ASAP7_75t_L g152 ( 
.A1(n_135),
.A2(n_100),
.B(n_101),
.Y(n_152)
);

NAND3xp33_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_139),
.C(n_126),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_154),
.A2(n_161),
.B1(n_168),
.B2(n_26),
.Y(n_188)
);

A2O1A1Ixp33_ASAP7_75t_L g156 ( 
.A1(n_123),
.A2(n_109),
.B(n_94),
.C(n_115),
.Y(n_156)
);

AOI21xp5_ASAP7_75t_L g183 ( 
.A1(n_156),
.A2(n_123),
.B(n_129),
.Y(n_183)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_131),
.Y(n_157)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

INVx13_ASAP7_75t_L g158 ( 
.A(n_141),
.Y(n_158)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_158),
.Y(n_174)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_126),
.B(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_160),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_142),
.A2(n_98),
.B1(n_104),
.B2(n_88),
.Y(n_161)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_163),
.Y(n_181)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_132),
.Y(n_164)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_164),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_129),
.B(n_4),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g187 ( 
.A(n_165),
.B(n_170),
.Y(n_187)
);

XOR2x1_ASAP7_75t_L g166 ( 
.A(n_125),
.B(n_21),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_166),
.A2(n_136),
.B1(n_137),
.B2(n_144),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_138),
.Y(n_167)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_167),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_127),
.B(n_27),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_124),
.Y(n_177)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_134),
.Y(n_170)
);

A2O1A1Ixp33_ASAP7_75t_SL g171 ( 
.A1(n_122),
.A2(n_62),
.B(n_60),
.C(n_68),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_171),
.A2(n_75),
.B(n_27),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_172),
.B(n_154),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g175 ( 
.A(n_163),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_175),
.Y(n_209)
);

NAND3xp33_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_149),
.C(n_155),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_177),
.B(n_185),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_153),
.A2(n_128),
.B1(n_133),
.B2(n_135),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g211 ( 
.A1(n_178),
.A2(n_186),
.B1(n_170),
.B2(n_171),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g200 ( 
.A1(n_183),
.A2(n_188),
.B(n_190),
.Y(n_200)
);

AO22x1_ASAP7_75t_SL g184 ( 
.A1(n_166),
.A2(n_130),
.B1(n_139),
.B2(n_26),
.Y(n_184)
);

AO21x1_ASAP7_75t_L g202 ( 
.A1(n_184),
.A2(n_169),
.B(n_171),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g185 ( 
.A(n_168),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_148),
.A2(n_26),
.B1(n_19),
.B2(n_21),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_147),
.B(n_75),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_192),
.B(n_195),
.C(n_146),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_158),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_193),
.B(n_167),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_174),
.B(n_145),
.Y(n_196)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_196),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_189),
.B(n_162),
.Y(n_197)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_197),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_184),
.A2(n_149),
.B1(n_159),
.B2(n_151),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_198),
.A2(n_190),
.B(n_172),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_202),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_201),
.B(n_195),
.C(n_192),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_145),
.Y(n_203)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

OAI21xp5_ASAP7_75t_SL g232 ( 
.A1(n_204),
.A2(n_206),
.B(n_214),
.Y(n_232)
);

OA21x2_ASAP7_75t_SL g206 ( 
.A1(n_184),
.A2(n_156),
.B(n_162),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_207),
.B(n_208),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_194),
.B(n_161),
.Y(n_210)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_210),
.B(n_213),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_211),
.A2(n_215),
.B1(n_180),
.B2(n_191),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_179),
.A2(n_171),
.B1(n_165),
.B2(n_26),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_212),
.A2(n_187),
.B1(n_21),
.B2(n_8),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g213 ( 
.A(n_194),
.B(n_171),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_175),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_178),
.A2(n_75),
.B1(n_21),
.B2(n_7),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_182),
.B(n_5),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_216),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_224),
.C(n_225),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_221),
.A2(n_222),
.B1(n_202),
.B2(n_200),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_177),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_201),
.B(n_173),
.C(n_186),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_226),
.Y(n_236)
);

BUFx24_ASAP7_75t_SL g227 ( 
.A(n_205),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_225),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_199),
.B(n_187),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_200),
.C(n_213),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_211),
.A2(n_215),
.B(n_197),
.Y(n_233)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_233),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_229),
.B(n_198),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_239),
.C(n_240),
.Y(n_248)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_235),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_209),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_216),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_241),
.B(n_242),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_218),
.A2(n_209),
.B1(n_214),
.B2(n_21),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_218),
.B(n_5),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_244),
.B(n_221),
.C(n_222),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_217),
.B(n_5),
.C(n_6),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_245),
.B(n_230),
.C(n_232),
.Y(n_246)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_249),
.B(n_250),
.C(n_251),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_238),
.B(n_219),
.C(n_224),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_237),
.A2(n_228),
.B(n_220),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_238),
.B(n_220),
.C(n_8),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_252),
.B(n_253),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_236),
.A2(n_6),
.B(n_9),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_255),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g257 ( 
.A(n_247),
.B(n_240),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_257),
.B(n_262),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_248),
.B(n_234),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_259),
.B(n_6),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_244),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_261),
.B(n_246),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g263 ( 
.A(n_254),
.B(n_245),
.Y(n_263)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_263),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_264),
.B(n_267),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_257),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_265),
.B(n_268),
.Y(n_271)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_260),
.Y(n_268)
);

OR2x2_ASAP7_75t_L g272 ( 
.A(n_269),
.B(n_11),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_266),
.A2(n_256),
.B1(n_13),
.B2(n_14),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g275 ( 
.A(n_270),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_272),
.A2(n_256),
.B(n_267),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_273),
.B(n_271),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_275),
.B(n_14),
.Y(n_277)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_277),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_13),
.Y(n_279)
);


endmodule