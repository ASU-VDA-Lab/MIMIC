module fake_netlist_1_7405_n_1468 (n_117, n_44, n_185, n_22, n_57, n_26, n_284, n_278, n_60, n_114, n_41, n_94, n_125, n_9, n_161, n_177, n_130, n_189, n_311, n_19, n_292, n_309, n_160, n_154, n_7, n_29, n_328, n_229, n_252, n_152, n_113, n_206, n_17, n_288, n_6, n_296, n_157, n_79, n_202, n_38, n_142, n_232, n_316, n_31, n_211, n_275, n_0, n_131, n_112, n_205, n_162, n_163, n_105, n_227, n_231, n_298, n_144, n_27, n_53, n_183, n_199, n_83, n_28, n_48, n_100, n_305, n_228, n_236, n_150, n_3, n_18, n_301, n_66, n_222, n_234, n_286, n_15, n_190, n_246, n_321, n_324, n_39, n_279, n_303, n_326, n_289, n_249, n_244, n_50, n_73, n_49, n_119, n_141, n_97, n_167, n_171, n_65, n_196, n_192, n_312, n_137, n_277, n_45, n_85, n_250, n_314, n_237, n_181, n_101, n_62, n_255, n_36, n_37, n_91, n_108, n_116, n_230, n_209, n_274, n_16, n_282, n_319, n_241, n_95, n_238, n_318, n_293, n_135, n_42, n_24, n_247, n_304, n_294, n_313, n_210, n_184, n_322, n_310, n_191, n_307, n_46, n_32, n_235, n_243, n_268, n_174, n_248, n_72, n_299, n_43, n_89, n_256, n_67, n_77, n_20, n_54, n_172, n_329, n_251, n_59, n_218, n_1, n_271, n_302, n_270, n_153, n_61, n_259, n_308, n_93, n_140, n_207, n_224, n_96, n_219, n_133, n_149, n_81, n_69, n_214, n_204, n_88, n_33, n_107, n_254, n_262, n_10, n_239, n_87, n_98, n_276, n_320, n_285, n_195, n_165, n_34, n_5, n_23, n_8, n_217, n_139, n_193, n_273, n_120, n_70, n_245, n_90, n_260, n_78, n_197, n_201, n_317, n_4, n_40, n_111, n_64, n_265, n_264, n_200, n_208, n_126, n_178, n_118, n_179, n_315, n_86, n_143, n_295, n_263, n_166, n_186, n_75, n_136, n_283, n_76, n_216, n_147, n_148, n_212, n_92, n_11, n_168, n_134, n_233, n_82, n_106, n_173, n_327, n_325, n_51, n_225, n_220, n_267, n_221, n_203, n_52, n_102, n_115, n_80, n_300, n_158, n_121, n_35, n_240, n_103, n_180, n_104, n_74, n_272, n_146, n_306, n_47, n_215, n_242, n_155, n_13, n_198, n_169, n_156, n_124, n_297, n_128, n_129, n_63, n_14, n_71, n_56, n_188, n_127, n_291, n_170, n_281, n_58, n_122, n_187, n_138, n_323, n_258, n_253, n_84, n_266, n_55, n_12, n_213, n_182, n_226, n_159, n_176, n_68, n_2, n_123, n_223, n_25, n_30, n_194, n_287, n_110, n_261, n_164, n_175, n_145, n_290, n_280, n_21, n_99, n_109, n_132, n_151, n_257, n_269, n_1468);
input n_117;
input n_44;
input n_185;
input n_22;
input n_57;
input n_26;
input n_284;
input n_278;
input n_60;
input n_114;
input n_41;
input n_94;
input n_125;
input n_9;
input n_161;
input n_177;
input n_130;
input n_189;
input n_311;
input n_19;
input n_292;
input n_309;
input n_160;
input n_154;
input n_7;
input n_29;
input n_328;
input n_229;
input n_252;
input n_152;
input n_113;
input n_206;
input n_17;
input n_288;
input n_6;
input n_296;
input n_157;
input n_79;
input n_202;
input n_38;
input n_142;
input n_232;
input n_316;
input n_31;
input n_211;
input n_275;
input n_0;
input n_131;
input n_112;
input n_205;
input n_162;
input n_163;
input n_105;
input n_227;
input n_231;
input n_298;
input n_144;
input n_27;
input n_53;
input n_183;
input n_199;
input n_83;
input n_28;
input n_48;
input n_100;
input n_305;
input n_228;
input n_236;
input n_150;
input n_3;
input n_18;
input n_301;
input n_66;
input n_222;
input n_234;
input n_286;
input n_15;
input n_190;
input n_246;
input n_321;
input n_324;
input n_39;
input n_279;
input n_303;
input n_326;
input n_289;
input n_249;
input n_244;
input n_50;
input n_73;
input n_49;
input n_119;
input n_141;
input n_97;
input n_167;
input n_171;
input n_65;
input n_196;
input n_192;
input n_312;
input n_137;
input n_277;
input n_45;
input n_85;
input n_250;
input n_314;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_37;
input n_91;
input n_108;
input n_116;
input n_230;
input n_209;
input n_274;
input n_16;
input n_282;
input n_319;
input n_241;
input n_95;
input n_238;
input n_318;
input n_293;
input n_135;
input n_42;
input n_24;
input n_247;
input n_304;
input n_294;
input n_313;
input n_210;
input n_184;
input n_322;
input n_310;
input n_191;
input n_307;
input n_46;
input n_32;
input n_235;
input n_243;
input n_268;
input n_174;
input n_248;
input n_72;
input n_299;
input n_43;
input n_89;
input n_256;
input n_67;
input n_77;
input n_20;
input n_54;
input n_172;
input n_329;
input n_251;
input n_59;
input n_218;
input n_1;
input n_271;
input n_302;
input n_270;
input n_153;
input n_61;
input n_259;
input n_308;
input n_93;
input n_140;
input n_207;
input n_224;
input n_96;
input n_219;
input n_133;
input n_149;
input n_81;
input n_69;
input n_214;
input n_204;
input n_88;
input n_33;
input n_107;
input n_254;
input n_262;
input n_10;
input n_239;
input n_87;
input n_98;
input n_276;
input n_320;
input n_285;
input n_195;
input n_165;
input n_34;
input n_5;
input n_23;
input n_8;
input n_217;
input n_139;
input n_193;
input n_273;
input n_120;
input n_70;
input n_245;
input n_90;
input n_260;
input n_78;
input n_197;
input n_201;
input n_317;
input n_4;
input n_40;
input n_111;
input n_64;
input n_265;
input n_264;
input n_200;
input n_208;
input n_126;
input n_178;
input n_118;
input n_179;
input n_315;
input n_86;
input n_143;
input n_295;
input n_263;
input n_166;
input n_186;
input n_75;
input n_136;
input n_283;
input n_76;
input n_216;
input n_147;
input n_148;
input n_212;
input n_92;
input n_11;
input n_168;
input n_134;
input n_233;
input n_82;
input n_106;
input n_173;
input n_327;
input n_325;
input n_51;
input n_225;
input n_220;
input n_267;
input n_221;
input n_203;
input n_52;
input n_102;
input n_115;
input n_80;
input n_300;
input n_158;
input n_121;
input n_35;
input n_240;
input n_103;
input n_180;
input n_104;
input n_74;
input n_272;
input n_146;
input n_306;
input n_47;
input n_215;
input n_242;
input n_155;
input n_13;
input n_198;
input n_169;
input n_156;
input n_124;
input n_297;
input n_128;
input n_129;
input n_63;
input n_14;
input n_71;
input n_56;
input n_188;
input n_127;
input n_291;
input n_170;
input n_281;
input n_58;
input n_122;
input n_187;
input n_138;
input n_323;
input n_258;
input n_253;
input n_84;
input n_266;
input n_55;
input n_12;
input n_213;
input n_182;
input n_226;
input n_159;
input n_176;
input n_68;
input n_2;
input n_123;
input n_223;
input n_25;
input n_30;
input n_194;
input n_287;
input n_110;
input n_261;
input n_164;
input n_175;
input n_145;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_132;
input n_151;
input n_257;
input n_269;
output n_1468;
wire n_1309;
wire n_963;
wire n_1034;
wire n_949;
wire n_1277;
wire n_1312;
wire n_858;
wire n_646;
wire n_1334;
wire n_829;
wire n_1198;
wire n_1382;
wire n_667;
wire n_988;
wire n_1363;
wire n_655;
wire n_1298;
wire n_1391;
wire n_903;
wire n_965;
wire n_918;
wire n_770;
wire n_1211;
wire n_878;
wire n_637;
wire n_564;
wire n_779;
wire n_528;
wire n_1128;
wire n_850;
wire n_672;
wire n_627;
wire n_1118;
wire n_1161;
wire n_1030;
wire n_807;
wire n_877;
wire n_1445;
wire n_545;
wire n_896;
wire n_334;
wire n_588;
wire n_1019;
wire n_940;
wire n_789;
wire n_1197;
wire n_1163;
wire n_1404;
wire n_387;
wire n_452;
wire n_518;
wire n_1336;
wire n_411;
wire n_1341;
wire n_1381;
wire n_860;
wire n_1208;
wire n_1201;
wire n_1342;
wire n_340;
wire n_373;
wire n_1194;
wire n_922;
wire n_465;
wire n_636;
wire n_914;
wire n_1352;
wire n_1005;
wire n_1097;
wire n_1125;
wire n_1017;
wire n_773;
wire n_847;
wire n_668;
wire n_437;
wire n_680;
wire n_642;
wire n_1267;
wire n_830;
wire n_1112;
wire n_517;
wire n_1295;
wire n_1297;
wire n_502;
wire n_543;
wire n_1159;
wire n_1250;
wire n_1002;
wire n_1355;
wire n_915;
wire n_367;
wire n_999;
wire n_769;
wire n_624;
wire n_725;
wire n_1407;
wire n_1018;
wire n_979;
wire n_499;
wire n_1349;
wire n_1033;
wire n_1063;
wire n_1010;
wire n_533;
wire n_490;
wire n_648;
wire n_613;
wire n_892;
wire n_571;
wire n_610;
wire n_771;
wire n_1337;
wire n_474;
wire n_402;
wire n_413;
wire n_676;
wire n_950;
wire n_995;
wire n_938;
wire n_331;
wire n_746;
wire n_1307;
wire n_619;
wire n_501;
wire n_699;
wire n_338;
wire n_551;
wire n_404;
wire n_1061;
wire n_509;
wire n_849;
wire n_864;
wire n_961;
wire n_1448;
wire n_1140;
wire n_611;
wire n_990;
wire n_800;
wire n_626;
wire n_1414;
wire n_1209;
wire n_1399;
wire n_1441;
wire n_926;
wire n_1274;
wire n_537;
wire n_660;
wire n_839;
wire n_1210;
wire n_1001;
wire n_1129;
wire n_450;
wire n_1406;
wire n_1099;
wire n_1328;
wire n_1369;
wire n_556;
wire n_1214;
wire n_379;
wire n_641;
wire n_966;
wire n_527;
wire n_797;
wire n_666;
wire n_1443;
wire n_1313;
wire n_954;
wire n_574;
wire n_823;
wire n_706;
wire n_822;
wire n_1181;
wire n_1438;
wire n_390;
wire n_514;
wire n_486;
wire n_568;
wire n_716;
wire n_899;
wire n_1066;
wire n_1251;
wire n_1199;
wire n_883;
wire n_573;
wire n_1308;
wire n_673;
wire n_1071;
wire n_1323;
wire n_1377;
wire n_1079;
wire n_409;
wire n_1321;
wire n_677;
wire n_1354;
wire n_1242;
wire n_756;
wire n_1385;
wire n_1240;
wire n_1139;
wire n_577;
wire n_1394;
wire n_870;
wire n_1324;
wire n_790;
wire n_761;
wire n_1287;
wire n_472;
wire n_1100;
wire n_419;
wire n_1193;
wire n_1119;
wire n_825;
wire n_477;
wire n_815;
wire n_908;
wire n_429;
wire n_488;
wire n_821;
wire n_745;
wire n_684;
wire n_1281;
wire n_1388;
wire n_1102;
wire n_723;
wire n_972;
wire n_1437;
wire n_997;
wire n_1387;
wire n_1244;
wire n_1464;
wire n_1184;
wire n_947;
wire n_620;
wire n_1141;
wire n_1213;
wire n_1452;
wire n_359;
wire n_1402;
wire n_1189;
wire n_1316;
wire n_923;
wire n_1205;
wire n_1172;
wire n_741;
wire n_1142;
wire n_1447;
wire n_1228;
wire n_831;
wire n_859;
wire n_1165;
wire n_1300;
wire n_1467;
wire n_930;
wire n_994;
wire n_1413;
wire n_410;
wire n_774;
wire n_1207;
wire n_1463;
wire n_377;
wire n_510;
wire n_1075;
wire n_1282;
wire n_493;
wire n_855;
wire n_722;
wire n_1083;
wire n_690;
wire n_1365;
wire n_1164;
wire n_451;
wire n_487;
wire n_748;
wire n_1373;
wire n_824;
wire n_793;
wire n_753;
wire n_355;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_1461;
wire n_1226;
wire n_1233;
wire n_1067;
wire n_866;
wire n_1108;
wire n_350;
wire n_433;
wire n_1311;
wire n_483;
wire n_395;
wire n_992;
wire n_361;
wire n_1077;
wire n_838;
wire n_705;
wire n_964;
wire n_590;
wire n_407;
wire n_1229;
wire n_792;
wire n_1412;
wire n_925;
wire n_1289;
wire n_957;
wire n_808;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_1306;
wire n_958;
wire n_468;
wire n_1453;
wire n_917;
wire n_523;
wire n_920;
wire n_1202;
wire n_1333;
wire n_1361;
wire n_911;
wire n_980;
wire n_817;
wire n_1056;
wire n_856;
wire n_1345;
wire n_661;
wire n_890;
wire n_787;
wire n_1015;
wire n_548;
wire n_1048;
wire n_973;
wire n_587;
wire n_476;
wire n_434;
wire n_489;
wire n_752;
wire n_1098;
wire n_1012;
wire n_461;
wire n_857;
wire n_1090;
wire n_786;
wire n_1121;
wire n_576;
wire n_1179;
wire n_1435;
wire n_796;
wire n_1216;
wire n_927;
wire n_1405;
wire n_1433;
wire n_840;
wire n_846;
wire n_968;
wire n_512;
wire n_1330;
wire n_586;
wire n_1246;
wire n_1276;
wire n_560;
wire n_697;
wire n_780;
wire n_447;
wire n_897;
wire n_1188;
wire n_580;
wire n_1009;
wire n_921;
wire n_854;
wire n_1011;
wire n_1155;
wire n_511;
wire n_467;
wire n_692;
wire n_1415;
wire n_644;
wire n_1116;
wire n_818;
wire n_738;
wire n_1225;
wire n_575;
wire n_711;
wire n_977;
wire n_884;
wire n_767;
wire n_393;
wire n_550;
wire n_826;
wire n_399;
wire n_1235;
wire n_1171;
wire n_459;
wire n_907;
wire n_1062;
wire n_708;
wire n_1271;
wire n_634;
wire n_696;
wire n_1203;
wire n_1013;
wire n_1000;
wire n_1370;
wire n_939;
wire n_953;
wire n_391;
wire n_478;
wire n_482;
wire n_394;
wire n_442;
wire n_485;
wire n_1248;
wire n_519;
wire n_1465;
wire n_1020;
wire n_1106;
wire n_635;
wire n_731;
wire n_986;
wire n_507;
wire n_605;
wire n_704;
wire n_633;
wire n_873;
wire n_1322;
wire n_751;
wire n_1147;
wire n_466;
wire n_900;
wire n_952;
wire n_685;
wire n_565;
wire n_1035;
wire n_475;
wire n_578;
wire n_542;
wire n_430;
wire n_943;
wire n_1326;
wire n_557;
wire n_842;
wire n_1269;
wire n_439;
wire n_614;
wire n_1346;
wire n_1107;
wire n_446;
wire n_423;
wire n_342;
wire n_799;
wire n_1427;
wire n_1050;
wire n_643;
wire n_874;
wire n_1049;
wire n_454;
wire n_687;
wire n_970;
wire n_984;
wire n_720;
wire n_806;
wire n_1157;
wire n_539;
wire n_1153;
wire n_816;
wire n_522;
wire n_898;
wire n_1135;
wire n_669;
wire n_541;
wire n_363;
wire n_733;
wire n_894;
wire n_376;
wire n_744;
wire n_520;
wire n_681;
wire n_942;
wire n_1029;
wire n_508;
wire n_721;
wire n_1060;
wire n_438;
wire n_640;
wire n_1037;
wire n_686;
wire n_944;
wire n_1110;
wire n_498;
wire n_1069;
wire n_1123;
wire n_811;
wire n_530;
wire n_737;
wire n_1266;
wire n_795;
wire n_1232;
wire n_449;
wire n_734;
wire n_919;
wire n_763;
wire n_1174;
wire n_657;
wire n_583;
wire n_841;
wire n_582;
wire n_1440;
wire n_1397;
wire n_1356;
wire n_836;
wire n_561;
wire n_1096;
wire n_594;
wire n_531;
wire n_1136;
wire n_1007;
wire n_1117;
wire n_1408;
wire n_424;
wire n_714;
wire n_932;
wire n_837;
wire n_1339;
wire n_1315;
wire n_1432;
wire n_867;
wire n_1070;
wire n_1270;
wire n_675;
wire n_504;
wire n_581;
wire n_698;
wire n_555;
wire n_901;
wire n_834;
wire n_727;
wire n_1038;
wire n_1162;
wire n_1103;
wire n_785;
wire n_375;
wire n_688;
wire n_347;
wire n_515;
wire n_1290;
wire n_1234;
wire n_592;
wire n_1045;
wire n_1449;
wire n_1115;
wire n_521;
wire n_625;
wire n_585;
wire n_1190;
wire n_1237;
wire n_713;
wire n_457;
wire n_736;
wire n_606;
wire n_332;
wire n_1292;
wire n_1425;
wire n_421;
wire n_1148;
wire n_739;
wire n_1166;
wire n_987;
wire n_1086;
wire n_406;
wire n_1416;
wire n_1236;
wire n_791;
wire n_707;
wire n_603;
wire n_1261;
wire n_885;
wire n_500;
wire n_607;
wire n_496;
wire n_1362;
wire n_801;
wire n_1059;
wire n_701;
wire n_612;
wire n_1418;
wire n_1032;
wire n_1284;
wire n_1358;
wire n_336;
wire n_464;
wire n_1243;
wire n_1196;
wire n_1338;
wire n_814;
wire n_985;
wire n_1191;
wire n_971;
wire n_904;
wire n_1301;
wire n_532;
wire n_400;
wire n_1455;
wire n_386;
wire n_432;
wire n_659;
wire n_1329;
wire n_1185;
wire n_389;
wire n_436;
wire n_1217;
wire n_715;
wire n_330;
wire n_1087;
wire n_662;
wire n_1372;
wire n_1460;
wire n_1451;
wire n_617;
wire n_598;
wire n_732;
wire n_724;
wire n_599;
wire n_1459;
wire n_609;
wire n_909;
wire n_1273;
wire n_366;
wire n_1319;
wire n_596;
wire n_1215;
wire n_951;
wire n_1024;
wire n_1016;
wire n_652;
wire n_333;
wire n_1417;
wire n_1357;
wire n_638;
wire n_563;
wire n_479;
wire n_623;
wire n_1222;
wire n_593;
wire n_872;
wire n_809;
wire n_1101;
wire n_1072;
wire n_865;
wire n_1064;
wire n_1380;
wire n_1254;
wire n_764;
wire n_426;
wire n_1375;
wire n_969;
wire n_417;
wire n_1253;
wire n_632;
wire n_1182;
wire n_828;
wire n_1138;
wire n_506;
wire n_1458;
wire n_381;
wire n_1255;
wire n_1299;
wire n_1450;
wire n_1332;
wire n_427;
wire n_703;
wire n_415;
wire n_1272;
wire n_928;
wire n_352;
wire n_882;
wire n_871;
wire n_803;
wire n_1429;
wire n_729;
wire n_805;
wire n_693;
wire n_1036;
wire n_1145;
wire n_651;
wire n_1303;
wire n_1320;
wire n_747;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_959;
wire n_719;
wire n_1206;
wire n_1257;
wire n_710;
wire n_1178;
wire n_546;
wire n_412;
wire n_664;
wire n_1249;
wire n_788;
wire n_1454;
wire n_1383;
wire n_403;
wire n_516;
wire n_549;
wire n_832;
wire n_996;
wire n_420;
wire n_1089;
wire n_1434;
wire n_1058;
wire n_388;
wire n_1396;
wire n_1400;
wire n_1082;
wire n_1052;
wire n_1055;
wire n_974;
wire n_591;
wire n_933;
wire n_1252;
wire n_416;
wire n_536;
wire n_1256;
wire n_1259;
wire n_1351;
wire n_1318;
wire n_956;
wire n_989;
wire n_754;
wire n_775;
wire n_616;
wire n_1227;
wire n_365;
wire n_495;
wire n_364;
wire n_566;
wire n_1144;
wire n_344;
wire n_503;
wire n_1279;
wire n_1152;
wire n_1068;
wire n_1149;
wire n_1430;
wire n_615;
wire n_1386;
wire n_1170;
wire n_804;
wire n_570;
wire n_1133;
wire n_1317;
wire n_440;
wire n_422;
wire n_679;
wire n_1131;
wire n_597;
wire n_1039;
wire n_1395;
wire n_835;
wire n_778;
wire n_1156;
wire n_1288;
wire n_1340;
wire n_1042;
wire n_1130;
wire n_584;
wire n_912;
wire n_1325;
wire n_1043;
wire n_1283;
wire n_346;
wire n_397;
wire n_1008;
wire n_1109;
wire n_1026;
wire n_1027;
wire n_1040;
wire n_1367;
wire n_569;
wire n_946;
wire n_960;
wire n_1168;
wire n_343;
wire n_458;
wire n_1084;
wire n_618;
wire n_341;
wire n_470;
wire n_1085;
wire n_1073;
wire n_868;
wire n_1466;
wire n_473;
wire n_991;
wire n_843;
wire n_1263;
wire n_1393;
wire n_538;
wire n_492;
wire n_1426;
wire n_1150;
wire n_1462;
wire n_1327;
wire n_368;
wire n_1444;
wire n_650;
wire n_469;
wire n_1187;
wire n_742;
wire n_913;
wire n_845;
wire n_891;
wire n_1134;
wire n_494;
wire n_372;
wire n_631;
wire n_934;
wire n_425;
wire n_562;
wire n_1436;
wire n_1192;
wire n_983;
wire n_781;
wire n_709;
wire n_1105;
wire n_408;
wire n_1378;
wire n_385;
wire n_1127;
wire n_1348;
wire n_1173;
wire n_663;
wire n_513;
wire n_1092;
wire n_1124;
wire n_1278;
wire n_998;
wire n_604;
wire n_1260;
wire n_755;
wire n_1409;
wire n_848;
wire n_1031;
wire n_1293;
wire n_1280;
wire n_1158;
wire n_743;
wire n_757;
wire n_750;
wire n_448;
wire n_645;
wire n_348;
wire n_1022;
wire n_802;
wire n_353;
wire n_993;
wire n_1122;
wire n_1224;
wire n_383;
wire n_762;
wire n_1422;
wire n_981;
wire n_1095;
wire n_758;
wire n_544;
wire n_1175;
wire n_853;
wire n_1376;
wire n_765;
wire n_1177;
wire n_1310;
wire n_462;
wire n_1347;
wire n_1384;
wire n_783;
wire n_1074;
wire n_1374;
wire n_463;
wire n_1379;
wire n_1003;
wire n_678;
wire n_1200;
wire n_384;
wire n_978;
wire n_547;
wire n_1247;
wire n_628;
wire n_812;
wire n_777;
wire n_351;
wire n_401;
wire n_345;
wire n_360;
wire n_481;
wire n_443;
wire n_694;
wire n_1262;
wire n_1360;
wire n_1078;
wire n_702;
wire n_572;
wire n_1094;
wire n_1204;
wire n_392;
wire n_1169;
wire n_975;
wire n_1081;
wire n_1457;
wire n_671;
wire n_540;
wire n_937;
wire n_1093;
wire n_1275;
wire n_955;
wire n_945;
wire n_554;
wire n_726;
wire n_712;
wire n_608;
wire n_567;
wire n_888;
wire n_529;
wire n_455;
wire n_1025;
wire n_1389;
wire n_1132;
wire n_630;
wire n_1180;
wire n_647;
wire n_1364;
wire n_1350;
wire n_844;
wire n_1403;
wire n_1160;
wire n_1420;
wire n_1245;
wire n_1195;
wire n_1241;
wire n_1302;
wire n_895;
wire n_798;
wire n_887;
wire n_471;
wire n_1014;
wire n_1410;
wire n_1442;
wire n_665;
wire n_1154;
wire n_863;
wire n_1265;
wire n_730;
wire n_1212;
wire n_735;
wire n_1091;
wire n_784;
wire n_354;
wire n_1220;
wire n_893;
wire n_1028;
wire n_910;
wire n_935;
wire n_1046;
wire n_1183;
wire n_460;
wire n_813;
wire n_1076;
wire n_369;
wire n_1186;
wire n_1167;
wire n_674;
wire n_810;
wire n_982;
wire n_889;
wire n_689;
wire n_902;
wire n_1423;
wire n_1113;
wire n_1264;
wire n_760;
wire n_941;
wire n_1368;
wire n_362;
wire n_931;
wire n_827;
wire n_1218;
wire n_1343;
wire n_1041;
wire n_1080;
wire n_1126;
wire n_1151;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_1065;
wire n_622;
wire n_601;
wire n_1331;
wire n_1176;
wire n_649;
wire n_526;
wire n_1047;
wire n_768;
wire n_869;
wire n_880;
wire n_621;
wire n_370;
wire n_589;
wire n_505;
wire n_682;
wire n_906;
wire n_357;
wire n_653;
wire n_881;
wire n_1439;
wire n_374;
wire n_718;
wire n_1411;
wire n_1238;
wire n_1114;
wire n_1286;
wire n_948;
wire n_1304;
wire n_1314;
wire n_717;
wire n_861;
wire n_654;
wire n_1221;
wire n_428;
wire n_794;
wire n_1268;
wire n_639;
wire n_1305;
wire n_552;
wire n_1023;
wire n_1057;
wire n_435;
wire n_1359;
wire n_1294;
wire n_1051;
wire n_1088;
wire n_851;
wire n_396;
wire n_398;
wire n_445;
wire n_656;
wire n_1230;
wire n_553;
wire n_1431;
wire n_349;
wire n_1021;
wire n_1456;
wire n_749;
wire n_535;
wire n_1006;
wire n_1054;
wire n_1353;
wire n_1231;
wire n_358;
wire n_456;
wire n_962;
wire n_1424;
wire n_782;
wire n_524;
wire n_1044;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_1239;
wire n_1335;
wire n_924;
wire n_378;
wire n_441;
wire n_1285;
wire n_1344;
wire n_335;
wire n_700;
wire n_534;
wire n_1401;
wire n_1296;
wire n_1428;
wire n_766;
wire n_602;
wire n_1143;
wire n_629;
wire n_1053;
wire n_1223;
wire n_1421;
wire n_1390;
wire n_967;
wire n_1419;
wire n_1258;
wire n_418;
wire n_380;
wire n_356;
wire n_600;
wire n_371;
wire n_820;
wire n_558;
wire n_670;
wire n_1004;
wire n_683;
wire n_1371;
wire n_929;
wire n_1111;
wire n_976;
wire n_1446;
wire n_695;
wire n_1104;
wire n_1392;
wire n_1120;
wire n_1219;
wire n_595;
wire n_759;
wire n_559;
wire n_1366;
wire n_480;
wire n_453;
wire n_833;
wire n_1146;
wire n_414;
wire n_1137;
wire n_916;
wire n_740;
wire n_772;
wire n_819;
wire n_405;
wire n_1398;
wire n_491;
wire n_1291;
INVx1_ASAP7_75t_L g330 ( .A(n_293), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_38), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_327), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_201), .Y(n_333) );
CKINVDCx16_ASAP7_75t_R g334 ( .A(n_241), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_99), .Y(n_335) );
CKINVDCx5p33_ASAP7_75t_R g336 ( .A(n_314), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_295), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_73), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_3), .Y(n_339) );
CKINVDCx5p33_ASAP7_75t_R g340 ( .A(n_126), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_196), .Y(n_341) );
HB1xp67_ASAP7_75t_L g342 ( .A(n_197), .Y(n_342) );
CKINVDCx20_ASAP7_75t_R g343 ( .A(n_16), .Y(n_343) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_238), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_51), .Y(n_345) );
CKINVDCx5p33_ASAP7_75t_R g346 ( .A(n_145), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_300), .Y(n_347) );
CKINVDCx16_ASAP7_75t_R g348 ( .A(n_164), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_140), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_229), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_184), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_142), .Y(n_352) );
CKINVDCx5p33_ASAP7_75t_R g353 ( .A(n_174), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_209), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_104), .Y(n_355) );
CKINVDCx20_ASAP7_75t_R g356 ( .A(n_325), .Y(n_356) );
BUFx5_ASAP7_75t_L g357 ( .A(n_110), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_218), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_257), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_132), .Y(n_360) );
CKINVDCx5p33_ASAP7_75t_R g361 ( .A(n_262), .Y(n_361) );
NOR2xp67_ASAP7_75t_L g362 ( .A(n_141), .B(n_60), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_170), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g364 ( .A(n_298), .Y(n_364) );
CKINVDCx5p33_ASAP7_75t_R g365 ( .A(n_19), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_322), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_161), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_276), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_59), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_263), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_269), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_165), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_166), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_90), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_131), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_70), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_74), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_284), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_37), .Y(n_379) );
INVx2_ASAP7_75t_SL g380 ( .A(n_90), .Y(n_380) );
CKINVDCx5p33_ASAP7_75t_R g381 ( .A(n_5), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_162), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_281), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_212), .Y(n_384) );
CKINVDCx20_ASAP7_75t_R g385 ( .A(n_272), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_242), .Y(n_386) );
CKINVDCx5p33_ASAP7_75t_R g387 ( .A(n_228), .Y(n_387) );
CKINVDCx5p33_ASAP7_75t_R g388 ( .A(n_63), .Y(n_388) );
INVx1_ASAP7_75t_L g389 ( .A(n_243), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_302), .Y(n_390) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_156), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_294), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_329), .Y(n_393) );
HB1xp67_ASAP7_75t_L g394 ( .A(n_136), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_61), .Y(n_395) );
BUFx3_ASAP7_75t_L g396 ( .A(n_188), .Y(n_396) );
AND2x4_ASAP7_75t_L g397 ( .A(n_65), .B(n_4), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_220), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_40), .Y(n_399) );
CKINVDCx20_ASAP7_75t_R g400 ( .A(n_5), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_155), .Y(n_401) );
BUFx2_ASAP7_75t_L g402 ( .A(n_168), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_303), .Y(n_403) );
BUFx3_ASAP7_75t_L g404 ( .A(n_66), .Y(n_404) );
CKINVDCx5p33_ASAP7_75t_R g405 ( .A(n_259), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_58), .Y(n_406) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_12), .Y(n_407) );
OR2x2_ASAP7_75t_L g408 ( .A(n_282), .B(n_318), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_251), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_46), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_316), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_204), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_185), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_19), .Y(n_414) );
BUFx3_ASAP7_75t_L g415 ( .A(n_198), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_163), .Y(n_416) );
CKINVDCx16_ASAP7_75t_R g417 ( .A(n_157), .Y(n_417) );
BUFx6f_ASAP7_75t_L g418 ( .A(n_248), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_290), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_11), .Y(n_420) );
CKINVDCx5p33_ASAP7_75t_R g421 ( .A(n_171), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_178), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_27), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_91), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_191), .Y(n_425) );
CKINVDCx5p33_ASAP7_75t_R g426 ( .A(n_58), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_187), .Y(n_427) );
BUFx10_ASAP7_75t_L g428 ( .A(n_138), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_177), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_192), .Y(n_430) );
INVxp67_ASAP7_75t_SL g431 ( .A(n_47), .Y(n_431) );
BUFx6f_ASAP7_75t_L g432 ( .A(n_53), .Y(n_432) );
BUFx6f_ASAP7_75t_L g433 ( .A(n_216), .Y(n_433) );
CKINVDCx5p33_ASAP7_75t_R g434 ( .A(n_96), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_214), .Y(n_435) );
CKINVDCx5p33_ASAP7_75t_R g436 ( .A(n_182), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_217), .Y(n_437) );
BUFx5_ASAP7_75t_L g438 ( .A(n_292), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_249), .Y(n_439) );
INVxp67_ASAP7_75t_SL g440 ( .A(n_63), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_321), .Y(n_441) );
CKINVDCx5p33_ASAP7_75t_R g442 ( .A(n_167), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_219), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g444 ( .A(n_260), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_289), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_224), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_175), .Y(n_447) );
CKINVDCx5p33_ASAP7_75t_R g448 ( .A(n_245), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_144), .Y(n_449) );
INVx1_ASAP7_75t_L g450 ( .A(n_274), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_73), .Y(n_451) );
INVx2_ASAP7_75t_L g452 ( .A(n_70), .Y(n_452) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_176), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_147), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_34), .Y(n_455) );
BUFx2_ASAP7_75t_L g456 ( .A(n_137), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_98), .Y(n_457) );
INVx1_ASAP7_75t_SL g458 ( .A(n_288), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_160), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_306), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_151), .Y(n_461) );
INVx2_ASAP7_75t_SL g462 ( .A(n_85), .Y(n_462) );
HB1xp67_ASAP7_75t_L g463 ( .A(n_119), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_102), .Y(n_464) );
HB1xp67_ASAP7_75t_L g465 ( .A(n_181), .Y(n_465) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_320), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_10), .Y(n_467) );
NOR2xp67_ASAP7_75t_L g468 ( .A(n_301), .B(n_80), .Y(n_468) );
CKINVDCx16_ASAP7_75t_R g469 ( .A(n_116), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_221), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_315), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_252), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_41), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_172), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_89), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_273), .Y(n_476) );
CKINVDCx5p33_ASAP7_75t_R g477 ( .A(n_107), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_169), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_50), .B(n_77), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_77), .Y(n_480) );
BUFx2_ASAP7_75t_L g481 ( .A(n_126), .Y(n_481) );
CKINVDCx5p33_ASAP7_75t_R g482 ( .A(n_234), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_239), .Y(n_483) );
CKINVDCx5p33_ASAP7_75t_R g484 ( .A(n_213), .Y(n_484) );
BUFx2_ASAP7_75t_L g485 ( .A(n_124), .Y(n_485) );
CKINVDCx20_ASAP7_75t_R g486 ( .A(n_230), .Y(n_486) );
INVx1_ASAP7_75t_L g487 ( .A(n_231), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_296), .Y(n_488) );
HB1xp67_ASAP7_75t_L g489 ( .A(n_258), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_62), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_299), .Y(n_491) );
INVx2_ASAP7_75t_L g492 ( .A(n_183), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_215), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_49), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_235), .Y(n_495) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_55), .B(n_134), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_247), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_190), .Y(n_498) );
CKINVDCx5p33_ASAP7_75t_R g499 ( .A(n_246), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_44), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_123), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_202), .Y(n_502) );
CKINVDCx5p33_ASAP7_75t_R g503 ( .A(n_154), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_180), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_115), .B(n_34), .Y(n_505) );
BUFx2_ASAP7_75t_L g506 ( .A(n_150), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g507 ( .A(n_93), .Y(n_507) );
CKINVDCx5p33_ASAP7_75t_R g508 ( .A(n_107), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_275), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_146), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_10), .Y(n_511) );
CKINVDCx5p33_ASAP7_75t_R g512 ( .A(n_67), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_250), .Y(n_513) );
BUFx6f_ASAP7_75t_L g514 ( .A(n_418), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_438), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_357), .Y(n_516) );
INVx3_ASAP7_75t_L g517 ( .A(n_357), .Y(n_517) );
AND2x2_ASAP7_75t_SL g518 ( .A(n_342), .B(n_129), .Y(n_518) );
AND2x6_ASAP7_75t_L g519 ( .A(n_396), .B(n_130), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_438), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_342), .B(n_0), .Y(n_521) );
AND2x6_ASAP7_75t_L g522 ( .A(n_396), .B(n_133), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_463), .B(n_0), .Y(n_523) );
INVx1_ASAP7_75t_L g524 ( .A(n_357), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_391), .B(n_1), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_438), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_438), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_463), .B(n_1), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_357), .Y(n_529) );
INVx2_ASAP7_75t_L g530 ( .A(n_438), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_391), .B(n_2), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_357), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_357), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g534 ( .A1(n_400), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_534) );
AND2x2_ASAP7_75t_SL g535 ( .A(n_394), .B(n_135), .Y(n_535) );
OA21x2_ASAP7_75t_L g536 ( .A1(n_352), .A2(n_143), .B(n_139), .Y(n_536) );
INVx3_ASAP7_75t_L g537 ( .A(n_404), .Y(n_537) );
INVx5_ASAP7_75t_L g538 ( .A(n_418), .Y(n_538) );
INVx2_ASAP7_75t_L g539 ( .A(n_438), .Y(n_539) );
CKINVDCx20_ASAP7_75t_R g540 ( .A(n_374), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_394), .Y(n_541) );
NOR2xp33_ASAP7_75t_SL g542 ( .A(n_334), .B(n_328), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_338), .B(n_6), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_418), .Y(n_544) );
AND2x4_ASAP7_75t_L g545 ( .A(n_465), .B(n_6), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_481), .B(n_7), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_418), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_433), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_433), .Y(n_549) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_447), .B(n_7), .Y(n_550) );
INVx5_ASAP7_75t_L g551 ( .A(n_433), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_433), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_465), .Y(n_553) );
HB1xp67_ASAP7_75t_L g554 ( .A(n_485), .Y(n_554) );
INVxp67_ASAP7_75t_L g555 ( .A(n_380), .Y(n_555) );
BUFx6f_ASAP7_75t_L g556 ( .A(n_453), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_453), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_489), .Y(n_558) );
NOR2x1p5_ASAP7_75t_L g559 ( .A(n_541), .B(n_431), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_540), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_517), .Y(n_561) );
NOR2x1p5_ASAP7_75t_L g562 ( .A(n_541), .B(n_431), .Y(n_562) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_555), .B(n_402), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_517), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_517), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_517), .Y(n_566) );
INVx2_ASAP7_75t_L g567 ( .A(n_515), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_553), .B(n_456), .Y(n_568) );
NAND3xp33_ASAP7_75t_L g569 ( .A(n_516), .B(n_489), .C(n_333), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_515), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_553), .B(n_506), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_520), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_520), .Y(n_573) );
AOI22xp5_ASAP7_75t_L g574 ( .A1(n_518), .A2(n_535), .B1(n_523), .B2(n_528), .Y(n_574) );
INVx1_ASAP7_75t_SL g575 ( .A(n_554), .Y(n_575) );
AND2x4_ASAP7_75t_L g576 ( .A(n_521), .B(n_397), .Y(n_576) );
NAND2xp5_ASAP7_75t_SL g577 ( .A(n_558), .B(n_348), .Y(n_577) );
OR2x2_ASAP7_75t_L g578 ( .A(n_558), .B(n_469), .Y(n_578) );
INVx6_ASAP7_75t_L g579 ( .A(n_538), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_520), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_526), .Y(n_581) );
CKINVDCx6p67_ASAP7_75t_R g582 ( .A(n_518), .Y(n_582) );
AND2x6_ASAP7_75t_L g583 ( .A(n_521), .B(n_415), .Y(n_583) );
INVx4_ASAP7_75t_L g584 ( .A(n_519), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_537), .B(n_417), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_526), .Y(n_586) );
INVx3_ASAP7_75t_L g587 ( .A(n_527), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_527), .Y(n_588) );
INVx5_ASAP7_75t_L g589 ( .A(n_519), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_527), .Y(n_590) );
INVxp67_ASAP7_75t_SL g591 ( .A(n_525), .Y(n_591) );
INVx1_ASAP7_75t_L g592 ( .A(n_530), .Y(n_592) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_514), .Y(n_593) );
AND3x1_ASAP7_75t_L g594 ( .A(n_523), .B(n_462), .C(n_335), .Y(n_594) );
INVx2_ASAP7_75t_SL g595 ( .A(n_521), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_537), .B(n_466), .Y(n_596) );
NOR2xp33_ASAP7_75t_L g597 ( .A(n_537), .B(n_368), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_530), .Y(n_598) );
INVx3_ASAP7_75t_L g599 ( .A(n_539), .Y(n_599) );
NAND2xp5_ASAP7_75t_SL g600 ( .A(n_584), .B(n_518), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_591), .Y(n_601) );
OAI21xp33_ASAP7_75t_L g602 ( .A1(n_574), .A2(n_545), .B(n_521), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_575), .B(n_546), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_576), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_582), .A2(n_535), .B1(n_545), .B2(n_529), .Y(n_605) );
INVx4_ASAP7_75t_L g606 ( .A(n_583), .Y(n_606) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_582), .A2(n_535), .B1(n_545), .B2(n_529), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_581), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g609 ( .A(n_585), .B(n_545), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_596), .B(n_528), .Y(n_610) );
INVx2_ASAP7_75t_SL g611 ( .A(n_559), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_574), .A2(n_546), .B1(n_542), .B2(n_543), .Y(n_612) );
NOR2xp33_ASAP7_75t_L g613 ( .A(n_568), .B(n_525), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g614 ( .A(n_571), .B(n_531), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_581), .Y(n_615) );
BUFx3_ASAP7_75t_L g616 ( .A(n_583), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_576), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_576), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g619 ( .A1(n_595), .A2(n_532), .B(n_524), .Y(n_619) );
OAI22xp5_ASAP7_75t_SL g620 ( .A1(n_560), .A2(n_534), .B1(n_400), .B2(n_343), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_571), .B(n_531), .Y(n_621) );
NOR2xp33_ASAP7_75t_SL g622 ( .A(n_584), .B(n_356), .Y(n_622) );
INVx2_ASAP7_75t_L g623 ( .A(n_581), .Y(n_623) );
NOR2xp33_ASAP7_75t_L g624 ( .A(n_577), .B(n_550), .Y(n_624) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_578), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g626 ( .A(n_578), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_562), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_583), .B(n_542), .Y(n_628) );
INVx2_ASAP7_75t_SL g629 ( .A(n_583), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_594), .Y(n_630) );
AND2x6_ASAP7_75t_SL g631 ( .A(n_563), .B(n_331), .Y(n_631) );
INVx2_ASAP7_75t_L g632 ( .A(n_587), .Y(n_632) );
NAND2xp5_ASAP7_75t_SL g633 ( .A(n_584), .B(n_539), .Y(n_633) );
OR2x6_ASAP7_75t_L g634 ( .A(n_584), .B(n_479), .Y(n_634) );
AND2x2_ASAP7_75t_L g635 ( .A(n_569), .B(n_440), .Y(n_635) );
OAI22xp5_ASAP7_75t_L g636 ( .A1(n_569), .A2(n_358), .B1(n_370), .B2(n_356), .Y(n_636) );
AOI21xp5_ASAP7_75t_L g637 ( .A1(n_566), .A2(n_532), .B(n_524), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_597), .B(n_533), .Y(n_638) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_566), .B(n_533), .Y(n_639) );
AOI22xp5_ASAP7_75t_L g640 ( .A1(n_570), .A2(n_370), .B1(n_385), .B2(n_358), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_561), .B(n_332), .Y(n_641) );
OR2x6_ASAP7_75t_L g642 ( .A(n_561), .B(n_505), .Y(n_642) );
OR2x2_ASAP7_75t_L g643 ( .A(n_570), .B(n_339), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_561), .B(n_336), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_564), .B(n_344), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g646 ( .A(n_564), .B(n_428), .Y(n_646) );
NAND2xp5_ASAP7_75t_L g647 ( .A(n_564), .B(n_346), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_580), .A2(n_385), .B1(n_486), .B2(n_444), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_565), .B(n_353), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_587), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_589), .B(n_330), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_580), .A2(n_444), .B1(n_495), .B2(n_486), .Y(n_652) );
AOI22xp5_ASAP7_75t_L g653 ( .A1(n_586), .A2(n_495), .B1(n_509), .B2(n_364), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_565), .B(n_361), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_565), .B(n_363), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_586), .A2(n_522), .B1(n_519), .B2(n_376), .Y(n_656) );
NAND2xp5_ASAP7_75t_SL g657 ( .A(n_589), .B(n_337), .Y(n_657) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_590), .B(n_371), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_587), .Y(n_659) );
AND2x2_ASAP7_75t_L g660 ( .A(n_590), .B(n_340), .Y(n_660) );
NOR3xp33_ASAP7_75t_L g661 ( .A(n_587), .B(n_365), .C(n_345), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_599), .Y(n_662) );
OAI22xp5_ASAP7_75t_SL g663 ( .A1(n_592), .A2(n_509), .B1(n_388), .B2(n_407), .Y(n_663) );
AOI22xp5_ASAP7_75t_L g664 ( .A1(n_592), .A2(n_426), .B1(n_434), .B2(n_381), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_598), .B(n_387), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_599), .Y(n_666) );
HB1xp67_ASAP7_75t_L g667 ( .A(n_599), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_567), .B(n_405), .Y(n_668) );
INVx2_ASAP7_75t_L g669 ( .A(n_567), .Y(n_669) );
A2O1A1Ixp33_ASAP7_75t_L g670 ( .A1(n_572), .A2(n_378), .B(n_379), .C(n_355), .Y(n_670) );
INVx1_ASAP7_75t_L g671 ( .A(n_572), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_573), .A2(n_378), .B(n_410), .C(n_395), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_573), .B(n_421), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_588), .B(n_436), .Y(n_674) );
INVx4_ASAP7_75t_L g675 ( .A(n_589), .Y(n_675) );
NAND2xp5_ASAP7_75t_SL g676 ( .A(n_589), .B(n_341), .Y(n_676) );
NAND2xp33_ASAP7_75t_L g677 ( .A(n_589), .B(n_519), .Y(n_677) );
INVx2_ASAP7_75t_L g678 ( .A(n_588), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_614), .B(n_475), .Y(n_679) );
AND2x2_ASAP7_75t_L g680 ( .A(n_603), .B(n_477), .Y(n_680) );
OR2x2_ASAP7_75t_L g681 ( .A(n_626), .B(n_507), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g682 ( .A(n_621), .B(n_508), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_613), .B(n_512), .Y(n_683) );
INVx2_ASAP7_75t_L g684 ( .A(n_604), .Y(n_684) );
BUFx6f_ASAP7_75t_L g685 ( .A(n_606), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g686 ( .A1(n_605), .A2(n_420), .B1(n_423), .B2(n_414), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_601), .B(n_424), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g688 ( .A1(n_633), .A2(n_536), .B(n_349), .Y(n_688) );
AOI21xp5_ASAP7_75t_L g689 ( .A1(n_619), .A2(n_536), .B(n_350), .Y(n_689) );
AOI21xp5_ASAP7_75t_L g690 ( .A1(n_638), .A2(n_536), .B(n_351), .Y(n_690) );
AOI21xp5_ASAP7_75t_L g691 ( .A1(n_609), .A2(n_354), .B(n_347), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_617), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_605), .A2(n_455), .B1(n_464), .B2(n_451), .Y(n_693) );
OAI22xp5_ASAP7_75t_L g694 ( .A1(n_607), .A2(n_473), .B1(n_480), .B2(n_467), .Y(n_694) );
AOI22xp5_ASAP7_75t_L g695 ( .A1(n_607), .A2(n_500), .B1(n_501), .B2(n_490), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_618), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_669), .Y(n_697) );
NAND2xp5_ASAP7_75t_SL g698 ( .A(n_606), .B(n_442), .Y(n_698) );
OAI22xp5_ASAP7_75t_L g699 ( .A1(n_612), .A2(n_511), .B1(n_377), .B2(n_406), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_610), .A2(n_360), .B(n_359), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_660), .B(n_369), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_643), .B(n_377), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_627), .B(n_406), .Y(n_703) );
BUFx8_ASAP7_75t_SL g704 ( .A(n_634), .Y(n_704) );
CKINVDCx5p33_ASAP7_75t_R g705 ( .A(n_663), .Y(n_705) );
AND2x4_ASAP7_75t_L g706 ( .A(n_661), .B(n_611), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_667), .Y(n_707) );
O2A1O1Ixp5_ASAP7_75t_L g708 ( .A1(n_600), .A2(n_496), .B(n_393), .C(n_401), .Y(n_708) );
OAI22xp5_ASAP7_75t_L g709 ( .A1(n_600), .A2(n_457), .B1(n_494), .B2(n_452), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_630), .A2(n_452), .B1(n_494), .B2(n_457), .C(n_496), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_616), .B(n_362), .Y(n_711) );
AOI21xp5_ASAP7_75t_L g712 ( .A1(n_677), .A2(n_367), .B(n_366), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_640), .B(n_428), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_624), .B(n_458), .Y(n_714) );
INVx1_ASAP7_75t_L g715 ( .A(n_667), .Y(n_715) );
AOI21xp5_ASAP7_75t_L g716 ( .A1(n_639), .A2(n_373), .B(n_372), .Y(n_716) );
AOI21xp5_ASAP7_75t_L g717 ( .A1(n_637), .A2(n_382), .B(n_375), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_635), .B(n_448), .Y(n_718) );
O2A1O1Ixp5_ASAP7_75t_L g719 ( .A1(n_628), .A2(n_393), .B(n_401), .C(n_352), .Y(n_719) );
AND2x4_ASAP7_75t_SL g720 ( .A(n_648), .B(n_399), .Y(n_720) );
INVx2_ASAP7_75t_L g721 ( .A(n_669), .Y(n_721) );
A2O1A1Ixp33_ASAP7_75t_L g722 ( .A1(n_624), .A2(n_468), .B(n_384), .C(n_386), .Y(n_722) );
INVx1_ASAP7_75t_L g723 ( .A(n_642), .Y(n_723) );
OR2x2_ASAP7_75t_L g724 ( .A(n_652), .B(n_8), .Y(n_724) );
AND2x2_ASAP7_75t_L g725 ( .A(n_653), .B(n_399), .Y(n_725) );
AND2x2_ASAP7_75t_L g726 ( .A(n_636), .B(n_399), .Y(n_726) );
AND2x4_ASAP7_75t_L g727 ( .A(n_634), .B(n_383), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_642), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g729 ( .A1(n_641), .A2(n_390), .B(n_389), .Y(n_729) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_642), .B(n_471), .Y(n_730) );
INVx2_ASAP7_75t_L g731 ( .A(n_678), .Y(n_731) );
OAI22xp33_ASAP7_75t_L g732 ( .A1(n_622), .A2(n_432), .B1(n_399), .B2(n_482), .Y(n_732) );
NAND2xp5_ASAP7_75t_SL g733 ( .A(n_629), .B(n_484), .Y(n_733) );
OAI21xp33_ASAP7_75t_L g734 ( .A1(n_664), .A2(n_503), .B(n_499), .Y(n_734) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_634), .Y(n_735) );
AOI21xp5_ASAP7_75t_L g736 ( .A1(n_644), .A2(n_398), .B(n_392), .Y(n_736) );
OAI22xp5_ASAP7_75t_L g737 ( .A1(n_670), .A2(n_408), .B1(n_409), .B2(n_403), .Y(n_737) );
AOI21xp5_ASAP7_75t_L g738 ( .A1(n_645), .A2(n_412), .B(n_411), .Y(n_738) );
INVx1_ASAP7_75t_L g739 ( .A(n_650), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_678), .Y(n_740) );
BUFx8_ASAP7_75t_L g741 ( .A(n_620), .Y(n_741) );
NAND3xp33_ASAP7_75t_L g742 ( .A(n_670), .B(n_432), .C(n_416), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_659), .Y(n_743) );
NOR2x1_ASAP7_75t_L g744 ( .A(n_672), .B(n_413), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g745 ( .A1(n_647), .A2(n_422), .B(n_419), .Y(n_745) );
OAI21xp5_ASAP7_75t_L g746 ( .A1(n_672), .A2(n_522), .B(n_519), .Y(n_746) );
AOI21xp5_ASAP7_75t_L g747 ( .A1(n_649), .A2(n_427), .B(n_425), .Y(n_747) );
AOI21xp5_ASAP7_75t_L g748 ( .A1(n_654), .A2(n_435), .B(n_430), .Y(n_748) );
AOI21xp5_ASAP7_75t_L g749 ( .A1(n_655), .A2(n_439), .B(n_437), .Y(n_749) );
O2A1O1Ixp33_ASAP7_75t_SL g750 ( .A1(n_651), .A2(n_441), .B(n_445), .C(n_443), .Y(n_750) );
OAI22xp5_ASAP7_75t_L g751 ( .A1(n_671), .A2(n_432), .B1(n_449), .B2(n_446), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_646), .B(n_519), .Y(n_752) );
O2A1O1Ixp33_ASAP7_75t_L g753 ( .A1(n_658), .A2(n_454), .B(n_459), .C(n_450), .Y(n_753) );
AOI21xp5_ASAP7_75t_L g754 ( .A1(n_665), .A2(n_461), .B(n_460), .Y(n_754) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_668), .A2(n_472), .B(n_474), .C(n_470), .Y(n_755) );
INVx2_ASAP7_75t_SL g756 ( .A(n_623), .Y(n_756) );
AOI21xp5_ASAP7_75t_L g757 ( .A1(n_673), .A2(n_478), .B(n_476), .Y(n_757) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_674), .B(n_487), .C(n_483), .Y(n_758) );
BUFx2_ASAP7_75t_L g759 ( .A(n_631), .Y(n_759) );
INVx2_ASAP7_75t_L g760 ( .A(n_623), .Y(n_760) );
BUFx3_ASAP7_75t_L g761 ( .A(n_632), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_632), .B(n_522), .Y(n_762) );
OAI22xp5_ASAP7_75t_L g763 ( .A1(n_656), .A2(n_491), .B1(n_493), .B2(n_488), .Y(n_763) );
OR2x6_ASAP7_75t_SL g764 ( .A(n_608), .B(n_497), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_615), .B(n_522), .Y(n_765) );
AND2x4_ASAP7_75t_L g766 ( .A(n_662), .B(n_498), .Y(n_766) );
AOI21xp5_ASAP7_75t_L g767 ( .A1(n_656), .A2(n_504), .B(n_502), .Y(n_767) );
AOI21xp5_ASAP7_75t_L g768 ( .A1(n_666), .A2(n_513), .B(n_510), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g769 ( .A1(n_651), .A2(n_522), .B1(n_429), .B2(n_492), .Y(n_769) );
NOR2xp33_ASAP7_75t_R g770 ( .A(n_675), .B(n_8), .Y(n_770) );
INVx1_ASAP7_75t_SL g771 ( .A(n_657), .Y(n_771) );
NOR2xp33_ASAP7_75t_L g772 ( .A(n_676), .B(n_9), .Y(n_772) );
AOI221xp5_ASAP7_75t_SL g773 ( .A1(n_602), .A2(n_544), .B1(n_549), .B2(n_548), .C(n_547), .Y(n_773) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_603), .Y(n_774) );
OAI22xp5_ASAP7_75t_L g775 ( .A1(n_605), .A2(n_544), .B1(n_548), .B2(n_547), .Y(n_775) );
NAND2xp5_ASAP7_75t_L g776 ( .A(n_614), .B(n_11), .Y(n_776) );
O2A1O1Ixp33_ASAP7_75t_L g777 ( .A1(n_625), .A2(n_552), .B(n_549), .C(n_14), .Y(n_777) );
INVx1_ASAP7_75t_L g778 ( .A(n_601), .Y(n_778) );
INVx2_ASAP7_75t_L g779 ( .A(n_604), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_614), .B(n_13), .Y(n_780) );
AND2x2_ASAP7_75t_L g781 ( .A(n_603), .B(n_13), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_614), .B(n_14), .Y(n_782) );
BUFx4f_ASAP7_75t_L g783 ( .A(n_634), .Y(n_783) );
OAI22xp5_ASAP7_75t_SL g784 ( .A1(n_620), .A2(n_453), .B1(n_17), .B2(n_15), .Y(n_784) );
NAND2xp33_ASAP7_75t_SL g785 ( .A(n_606), .B(n_514), .Y(n_785) );
INVx1_ASAP7_75t_L g786 ( .A(n_601), .Y(n_786) );
NOR2x1_ASAP7_75t_L g787 ( .A(n_614), .B(n_514), .Y(n_787) );
BUFx6f_ASAP7_75t_L g788 ( .A(n_606), .Y(n_788) );
BUFx6f_ASAP7_75t_L g789 ( .A(n_606), .Y(n_789) );
NAND2xp33_ASAP7_75t_L g790 ( .A(n_602), .B(n_514), .Y(n_790) );
INVx4_ASAP7_75t_L g791 ( .A(n_606), .Y(n_791) );
INVx1_ASAP7_75t_SL g792 ( .A(n_603), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_604), .Y(n_793) );
OAI22xp5_ASAP7_75t_L g794 ( .A1(n_605), .A2(n_579), .B1(n_551), .B2(n_556), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g795 ( .A(n_614), .B(n_18), .Y(n_795) );
O2A1O1Ixp33_ASAP7_75t_L g796 ( .A1(n_625), .A2(n_22), .B(n_20), .C(n_21), .Y(n_796) );
AND2x4_ASAP7_75t_L g797 ( .A(n_735), .B(n_21), .Y(n_797) );
INVx5_ASAP7_75t_L g798 ( .A(n_704), .Y(n_798) );
OAI22x1_ASAP7_75t_L g799 ( .A1(n_705), .A2(n_24), .B1(n_22), .B2(n_23), .Y(n_799) );
AOI21xp5_ASAP7_75t_L g800 ( .A1(n_690), .A2(n_752), .B(n_762), .Y(n_800) );
BUFx12f_ASAP7_75t_L g801 ( .A(n_741), .Y(n_801) );
AOI21xp5_ASAP7_75t_L g802 ( .A1(n_689), .A2(n_593), .B(n_557), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_792), .B(n_24), .Y(n_803) );
OAI21xp5_ASAP7_75t_L g804 ( .A1(n_719), .A2(n_579), .B(n_557), .Y(n_804) );
AOI21xp5_ASAP7_75t_L g805 ( .A1(n_765), .A2(n_593), .B(n_557), .Y(n_805) );
INVx2_ASAP7_75t_L g806 ( .A(n_778), .Y(n_806) );
INVx3_ASAP7_75t_SL g807 ( .A(n_735), .Y(n_807) );
NAND3xp33_ASAP7_75t_L g808 ( .A(n_722), .B(n_557), .C(n_556), .Y(n_808) );
INVx3_ASAP7_75t_SL g809 ( .A(n_735), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_792), .B(n_25), .Y(n_810) );
AO21x1_ASAP7_75t_L g811 ( .A1(n_790), .A2(n_557), .B(n_556), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g812 ( .A1(n_783), .A2(n_556), .B1(n_579), .B2(n_27), .Y(n_812) );
BUFx6f_ASAP7_75t_L g813 ( .A(n_783), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_786), .Y(n_814) );
A2O1A1Ixp33_ASAP7_75t_L g815 ( .A1(n_777), .A2(n_593), .B(n_28), .C(n_25), .Y(n_815) );
BUFx6f_ASAP7_75t_L g816 ( .A(n_685), .Y(n_816) );
AO32x2_ASAP7_75t_L g817 ( .A1(n_709), .A2(n_26), .A3(n_28), .B1(n_29), .B2(n_30), .Y(n_817) );
AOI21xp5_ASAP7_75t_L g818 ( .A1(n_688), .A2(n_149), .B(n_148), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_774), .B(n_31), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_741), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g821 ( .A(n_686), .B(n_31), .Y(n_821) );
INVx2_ASAP7_75t_L g822 ( .A(n_697), .Y(n_822) );
AO31x2_ASAP7_75t_L g823 ( .A1(n_709), .A2(n_35), .A3(n_32), .B(n_33), .Y(n_823) );
OAI21xp5_ASAP7_75t_L g824 ( .A1(n_708), .A2(n_153), .B(n_152), .Y(n_824) );
INVx1_ASAP7_75t_L g825 ( .A(n_776), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g826 ( .A(n_681), .B(n_713), .Y(n_826) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_695), .B(n_32), .Y(n_827) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_706), .B(n_33), .Y(n_828) );
AOI21xp5_ASAP7_75t_L g829 ( .A1(n_721), .A2(n_740), .B(n_731), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_680), .B(n_35), .Y(n_830) );
OAI21x1_ASAP7_75t_L g831 ( .A1(n_787), .A2(n_159), .B(n_158), .Y(n_831) );
INVx2_ASAP7_75t_SL g832 ( .A(n_727), .Y(n_832) );
BUFx12f_ASAP7_75t_L g833 ( .A(n_759), .Y(n_833) );
AO32x2_ASAP7_75t_L g834 ( .A1(n_699), .A2(n_36), .A3(n_37), .B1(n_38), .B2(n_39), .Y(n_834) );
AND2x4_ASAP7_75t_L g835 ( .A(n_706), .B(n_36), .Y(n_835) );
CKINVDCx20_ASAP7_75t_R g836 ( .A(n_770), .Y(n_836) );
OAI21xp33_ASAP7_75t_L g837 ( .A1(n_683), .A2(n_40), .B(n_41), .Y(n_837) );
A2O1A1Ixp33_ASAP7_75t_L g838 ( .A1(n_753), .A2(n_45), .B(n_42), .C(n_43), .Y(n_838) );
A2O1A1Ixp33_ASAP7_75t_L g839 ( .A1(n_755), .A2(n_50), .B(n_48), .C(n_49), .Y(n_839) );
AO21x1_ASAP7_75t_L g840 ( .A1(n_746), .A2(n_179), .B(n_173), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g841 ( .A1(n_724), .A2(n_53), .B1(n_51), .B2(n_52), .Y(n_841) );
INVx2_ASAP7_75t_SL g842 ( .A(n_781), .Y(n_842) );
INVx2_ASAP7_75t_L g843 ( .A(n_684), .Y(n_843) );
AO31x2_ASAP7_75t_L g844 ( .A1(n_763), .A2(n_54), .A3(n_56), .B(n_57), .Y(n_844) );
AO32x2_ASAP7_75t_L g845 ( .A1(n_737), .A2(n_56), .A3(n_57), .B1(n_59), .B2(n_60), .Y(n_845) );
INVx3_ASAP7_75t_L g846 ( .A(n_720), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g847 ( .A1(n_691), .A2(n_189), .B(n_186), .Y(n_847) );
INVx2_ASAP7_75t_SL g848 ( .A(n_725), .Y(n_848) );
AND2x4_ASAP7_75t_L g849 ( .A(n_707), .B(n_61), .Y(n_849) );
AOI21xp33_ASAP7_75t_L g850 ( .A1(n_730), .A2(n_62), .B(n_64), .Y(n_850) );
OAI21x1_ASAP7_75t_L g851 ( .A1(n_712), .A2(n_194), .B(n_193), .Y(n_851) );
INVx2_ASAP7_75t_L g852 ( .A(n_779), .Y(n_852) );
NOR2xp33_ASAP7_75t_L g853 ( .A(n_679), .B(n_64), .Y(n_853) );
O2A1O1Ixp33_ASAP7_75t_L g854 ( .A1(n_693), .A2(n_65), .B(n_66), .C(n_67), .Y(n_854) );
CKINVDCx16_ASAP7_75t_R g855 ( .A(n_764), .Y(n_855) );
BUFx6f_ASAP7_75t_L g856 ( .A(n_685), .Y(n_856) );
OAI22xp5_ASAP7_75t_SL g857 ( .A1(n_784), .A2(n_68), .B1(n_69), .B2(n_71), .Y(n_857) );
AOI21xp5_ASAP7_75t_L g858 ( .A1(n_754), .A2(n_199), .B(n_195), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g859 ( .A1(n_746), .A2(n_203), .B(n_200), .Y(n_859) );
AOI21xp5_ASAP7_75t_L g860 ( .A1(n_729), .A2(n_206), .B(n_205), .Y(n_860) );
AO31x2_ASAP7_75t_L g861 ( .A1(n_763), .A2(n_68), .A3(n_69), .B(n_71), .Y(n_861) );
INVx1_ASAP7_75t_L g862 ( .A(n_780), .Y(n_862) );
AOI21xp5_ASAP7_75t_L g863 ( .A1(n_736), .A2(n_208), .B(n_207), .Y(n_863) );
AO32x2_ASAP7_75t_L g864 ( .A1(n_694), .A2(n_72), .A3(n_74), .B1(n_75), .B2(n_76), .Y(n_864) );
O2A1O1Ixp33_ASAP7_75t_L g865 ( .A1(n_796), .A2(n_72), .B(n_75), .C(n_76), .Y(n_865) );
A2O1A1Ixp33_ASAP7_75t_L g866 ( .A1(n_700), .A2(n_78), .B(n_79), .C(n_81), .Y(n_866) );
INVx1_ASAP7_75t_SL g867 ( .A(n_766), .Y(n_867) );
O2A1O1Ixp33_ASAP7_75t_L g868 ( .A1(n_737), .A2(n_78), .B(n_81), .C(n_82), .Y(n_868) );
AOI21xp5_ASAP7_75t_L g869 ( .A1(n_738), .A2(n_211), .B(n_210), .Y(n_869) );
AND2x4_ASAP7_75t_L g870 ( .A(n_715), .B(n_82), .Y(n_870) );
AOI21xp33_ASAP7_75t_L g871 ( .A1(n_723), .A2(n_83), .B(n_84), .Y(n_871) );
CKINVDCx8_ASAP7_75t_R g872 ( .A(n_711), .Y(n_872) );
A2O1A1Ixp33_ASAP7_75t_L g873 ( .A1(n_745), .A2(n_83), .B(n_84), .C(n_86), .Y(n_873) );
AND2x2_ASAP7_75t_L g874 ( .A(n_682), .B(n_86), .Y(n_874) );
AND2x2_ASAP7_75t_SL g875 ( .A(n_791), .B(n_87), .Y(n_875) );
HB1xp67_ASAP7_75t_L g876 ( .A(n_728), .Y(n_876) );
AO31x2_ASAP7_75t_L g877 ( .A1(n_775), .A2(n_88), .A3(n_89), .B(n_91), .Y(n_877) );
AND2x6_ASAP7_75t_L g878 ( .A(n_788), .B(n_92), .Y(n_878) );
INVx4_ASAP7_75t_L g879 ( .A(n_788), .Y(n_879) );
AO32x2_ASAP7_75t_L g880 ( .A1(n_751), .A2(n_92), .A3(n_93), .B1(n_94), .B2(n_95), .Y(n_880) );
NOR2xp33_ASAP7_75t_L g881 ( .A(n_714), .B(n_94), .Y(n_881) );
INVxp67_ASAP7_75t_L g882 ( .A(n_782), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_702), .B(n_95), .Y(n_883) );
NAND2x1p5_ASAP7_75t_L g884 ( .A(n_791), .B(n_96), .Y(n_884) );
AOI21xp5_ASAP7_75t_L g885 ( .A1(n_747), .A2(n_261), .B(n_326), .Y(n_885) );
INVx3_ASAP7_75t_L g886 ( .A(n_793), .Y(n_886) );
AND2x2_ASAP7_75t_L g887 ( .A(n_701), .B(n_97), .Y(n_887) );
AO31x2_ASAP7_75t_L g888 ( .A1(n_794), .A2(n_97), .A3(n_98), .B(n_99), .Y(n_888) );
NAND2xp33_ASAP7_75t_SL g889 ( .A(n_788), .B(n_100), .Y(n_889) );
NAND2xp5_ASAP7_75t_L g890 ( .A(n_692), .B(n_101), .Y(n_890) );
BUFx8_ASAP7_75t_SL g891 ( .A(n_726), .Y(n_891) );
AO31x2_ASAP7_75t_L g892 ( .A1(n_767), .A2(n_103), .A3(n_105), .B(n_106), .Y(n_892) );
INVx3_ASAP7_75t_L g893 ( .A(n_766), .Y(n_893) );
AOI21xp5_ASAP7_75t_L g894 ( .A1(n_748), .A2(n_266), .B(n_324), .Y(n_894) );
AO32x2_ASAP7_75t_L g895 ( .A1(n_756), .A2(n_108), .A3(n_109), .B1(n_110), .B2(n_111), .Y(n_895) );
AO21x1_ASAP7_75t_L g896 ( .A1(n_732), .A2(n_267), .B(n_323), .Y(n_896) );
INVx3_ASAP7_75t_L g897 ( .A(n_761), .Y(n_897) );
A2O1A1Ixp33_ASAP7_75t_L g898 ( .A1(n_749), .A2(n_111), .B(n_112), .C(n_113), .Y(n_898) );
OAI22xp33_ASAP7_75t_SL g899 ( .A1(n_795), .A2(n_112), .B1(n_113), .B2(n_114), .Y(n_899) );
AND2x4_ASAP7_75t_L g900 ( .A(n_696), .B(n_114), .Y(n_900) );
AND2x2_ASAP7_75t_L g901 ( .A(n_758), .B(n_117), .Y(n_901) );
INVx5_ASAP7_75t_L g902 ( .A(n_789), .Y(n_902) );
AO31x2_ASAP7_75t_L g903 ( .A1(n_717), .A2(n_118), .A3(n_119), .B(n_120), .Y(n_903) );
AOI22xp5_ASAP7_75t_L g904 ( .A1(n_744), .A2(n_118), .B1(n_120), .B2(n_121), .Y(n_904) );
BUFx3_ASAP7_75t_L g905 ( .A(n_743), .Y(n_905) );
BUFx2_ASAP7_75t_L g906 ( .A(n_789), .Y(n_906) );
NAND3xp33_ASAP7_75t_L g907 ( .A(n_710), .B(n_121), .C(n_122), .Y(n_907) );
AO21x1_ASAP7_75t_L g908 ( .A1(n_772), .A2(n_271), .B(n_319), .Y(n_908) );
INVx1_ASAP7_75t_L g909 ( .A(n_687), .Y(n_909) );
BUFx3_ASAP7_75t_L g910 ( .A(n_739), .Y(n_910) );
BUFx2_ASAP7_75t_L g911 ( .A(n_760), .Y(n_911) );
AOI21xp5_ASAP7_75t_L g912 ( .A1(n_757), .A2(n_270), .B(n_317), .Y(n_912) );
INVx1_ASAP7_75t_L g913 ( .A(n_703), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_718), .B(n_125), .Y(n_914) );
AND2x2_ASAP7_75t_L g915 ( .A(n_734), .B(n_127), .Y(n_915) );
O2A1O1Ixp33_ASAP7_75t_SL g916 ( .A1(n_771), .A2(n_698), .B(n_733), .C(n_742), .Y(n_916) );
AO31x2_ASAP7_75t_L g917 ( .A1(n_716), .A2(n_127), .A3(n_128), .B(n_222), .Y(n_917) );
INVx5_ASAP7_75t_L g918 ( .A(n_785), .Y(n_918) );
AO31x2_ASAP7_75t_L g919 ( .A1(n_768), .A2(n_128), .A3(n_223), .B(n_225), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_742), .B(n_226), .Y(n_920) );
BUFx2_ASAP7_75t_L g921 ( .A(n_771), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_750), .B(n_227), .Y(n_922) );
BUFx2_ASAP7_75t_L g923 ( .A(n_769), .Y(n_923) );
INVx6_ASAP7_75t_SL g924 ( .A(n_727), .Y(n_924) );
AO21x2_ASAP7_75t_L g925 ( .A1(n_690), .A2(n_232), .B(n_233), .Y(n_925) );
AOI221xp5_ASAP7_75t_SL g926 ( .A1(n_699), .A2(n_236), .B1(n_237), .B2(n_240), .C(n_244), .Y(n_926) );
A2O1A1Ixp33_ASAP7_75t_L g927 ( .A1(n_777), .A2(n_253), .B(n_254), .C(n_255), .Y(n_927) );
NAND2xp5_ASAP7_75t_L g928 ( .A(n_792), .B(n_256), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_778), .Y(n_929) );
AOI22xp33_ASAP7_75t_L g930 ( .A1(n_783), .A2(n_264), .B1(n_265), .B2(n_268), .Y(n_930) );
INVx4_ASAP7_75t_L g931 ( .A(n_704), .Y(n_931) );
INVx1_ASAP7_75t_L g932 ( .A(n_778), .Y(n_932) );
BUFx6f_ASAP7_75t_L g933 ( .A(n_735), .Y(n_933) );
AOI221xp5_ASAP7_75t_L g934 ( .A1(n_792), .A2(n_277), .B1(n_278), .B2(n_279), .C(n_280), .Y(n_934) );
AND2x2_ASAP7_75t_L g935 ( .A(n_792), .B(n_283), .Y(n_935) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_792), .A2(n_285), .B1(n_286), .B2(n_287), .C(n_291), .Y(n_936) );
INVx2_ASAP7_75t_SL g937 ( .A(n_783), .Y(n_937) );
BUFx12f_ASAP7_75t_L g938 ( .A(n_798), .Y(n_938) );
AND2x2_ASAP7_75t_L g939 ( .A(n_855), .B(n_297), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_814), .Y(n_940) );
BUFx12f_ASAP7_75t_L g941 ( .A(n_798), .Y(n_941) );
BUFx6f_ASAP7_75t_L g942 ( .A(n_902), .Y(n_942) );
INVx2_ASAP7_75t_L g943 ( .A(n_806), .Y(n_943) );
INVx2_ASAP7_75t_L g944 ( .A(n_929), .Y(n_944) );
NAND2xp5_ASAP7_75t_L g945 ( .A(n_909), .B(n_932), .Y(n_945) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_911), .Y(n_946) );
INVx2_ASAP7_75t_L g947 ( .A(n_843), .Y(n_947) );
OAI22x1_ASAP7_75t_L g948 ( .A1(n_835), .A2(n_304), .B1(n_305), .B2(n_307), .Y(n_948) );
OA21x2_ASAP7_75t_L g949 ( .A1(n_926), .A2(n_308), .B(n_309), .Y(n_949) );
INVx1_ASAP7_75t_L g950 ( .A(n_900), .Y(n_950) );
INVx1_ASAP7_75t_L g951 ( .A(n_900), .Y(n_951) );
OAI221xp5_ASAP7_75t_L g952 ( .A1(n_826), .A2(n_310), .B1(n_311), .B2(n_312), .C(n_313), .Y(n_952) );
BUFx8_ASAP7_75t_L g953 ( .A(n_801), .Y(n_953) );
INVx2_ASAP7_75t_SL g954 ( .A(n_798), .Y(n_954) );
INVxp33_ASAP7_75t_L g955 ( .A(n_813), .Y(n_955) );
INVx1_ASAP7_75t_L g956 ( .A(n_849), .Y(n_956) );
AND2x4_ASAP7_75t_L g957 ( .A(n_937), .B(n_813), .Y(n_957) );
HB1xp67_ASAP7_75t_L g958 ( .A(n_911), .Y(n_958) );
NOR2xp33_ASAP7_75t_L g959 ( .A(n_832), .B(n_882), .Y(n_959) );
INVx2_ASAP7_75t_L g960 ( .A(n_852), .Y(n_960) );
AOI21xp5_ASAP7_75t_L g961 ( .A1(n_805), .A2(n_804), .B(n_824), .Y(n_961) );
AND2x4_ASAP7_75t_L g962 ( .A(n_910), .B(n_902), .Y(n_962) );
AND2x2_ASAP7_75t_L g963 ( .A(n_875), .B(n_835), .Y(n_963) );
AND2x4_ASAP7_75t_L g964 ( .A(n_902), .B(n_913), .Y(n_964) );
NAND2xp5_ASAP7_75t_L g965 ( .A(n_825), .B(n_862), .Y(n_965) );
BUFx2_ASAP7_75t_L g966 ( .A(n_924), .Y(n_966) );
BUFx3_ASAP7_75t_L g967 ( .A(n_807), .Y(n_967) );
AOI21xp5_ASAP7_75t_L g968 ( .A1(n_829), .A2(n_818), .B(n_916), .Y(n_968) );
INVx1_ASAP7_75t_SL g969 ( .A(n_867), .Y(n_969) );
AND2x2_ASAP7_75t_L g970 ( .A(n_901), .B(n_870), .Y(n_970) );
BUFx3_ASAP7_75t_L g971 ( .A(n_809), .Y(n_971) );
NOR2xp33_ASAP7_75t_L g972 ( .A(n_842), .B(n_872), .Y(n_972) );
OA21x2_ASAP7_75t_L g973 ( .A1(n_840), .A2(n_831), .B(n_859), .Y(n_973) );
OR2x6_ASAP7_75t_L g974 ( .A(n_931), .B(n_884), .Y(n_974) );
INVx1_ASAP7_75t_L g975 ( .A(n_803), .Y(n_975) );
INVx1_ASAP7_75t_L g976 ( .A(n_810), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_876), .Y(n_977) );
INVx1_ASAP7_75t_L g978 ( .A(n_819), .Y(n_978) );
INVx1_ASAP7_75t_SL g979 ( .A(n_921), .Y(n_979) );
OA21x2_ASAP7_75t_L g980 ( .A1(n_920), .A2(n_908), .B(n_851), .Y(n_980) );
BUFx3_ASAP7_75t_L g981 ( .A(n_933), .Y(n_981) );
BUFx3_ASAP7_75t_L g982 ( .A(n_833), .Y(n_982) );
AND2x4_ASAP7_75t_L g983 ( .A(n_905), .B(n_886), .Y(n_983) );
OAI21xp5_ASAP7_75t_L g984 ( .A1(n_815), .A2(n_927), .B(n_890), .Y(n_984) );
INVx1_ASAP7_75t_L g985 ( .A(n_883), .Y(n_985) );
NAND2xp5_ASAP7_75t_L g986 ( .A(n_874), .B(n_887), .Y(n_986) );
BUFx3_ASAP7_75t_L g987 ( .A(n_836), .Y(n_987) );
INVx3_ASAP7_75t_L g988 ( .A(n_879), .Y(n_988) );
AO31x2_ASAP7_75t_L g989 ( .A1(n_923), .A2(n_839), .A3(n_838), .B(n_921), .Y(n_989) );
INVx1_ASAP7_75t_L g990 ( .A(n_797), .Y(n_990) );
INVx3_ASAP7_75t_L g991 ( .A(n_816), .Y(n_991) );
AND2x4_ASAP7_75t_L g992 ( .A(n_846), .B(n_897), .Y(n_992) );
INVx1_ASAP7_75t_L g993 ( .A(n_823), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_823), .Y(n_994) );
NAND2xp5_ASAP7_75t_L g995 ( .A(n_853), .B(n_822), .Y(n_995) );
AND2x2_ASAP7_75t_L g996 ( .A(n_828), .B(n_893), .Y(n_996) );
HB1xp67_ASAP7_75t_L g997 ( .A(n_906), .Y(n_997) );
AO31x2_ASAP7_75t_L g998 ( .A1(n_923), .A2(n_866), .A3(n_922), .B(n_873), .Y(n_998) );
INVx1_ASAP7_75t_L g999 ( .A(n_830), .Y(n_999) );
AOI21xp5_ASAP7_75t_L g1000 ( .A1(n_925), .A2(n_928), .B(n_808), .Y(n_1000) );
OAI21x1_ASAP7_75t_L g1001 ( .A1(n_860), .A2(n_894), .B(n_885), .Y(n_1001) );
CKINVDCx6p67_ASAP7_75t_R g1002 ( .A(n_820), .Y(n_1002) );
INVx3_ASAP7_75t_L g1003 ( .A(n_816), .Y(n_1003) );
AO31x2_ASAP7_75t_L g1004 ( .A1(n_898), .A2(n_881), .A3(n_847), .B(n_863), .Y(n_1004) );
NOR2xp33_ASAP7_75t_L g1005 ( .A(n_891), .B(n_924), .Y(n_1005) );
AND2x4_ASAP7_75t_L g1006 ( .A(n_935), .B(n_856), .Y(n_1006) );
NAND2xp5_ASAP7_75t_L g1007 ( .A(n_848), .B(n_914), .Y(n_1007) );
CKINVDCx12_ASAP7_75t_R g1008 ( .A(n_857), .Y(n_1008) );
AOI21xp5_ASAP7_75t_L g1009 ( .A1(n_858), .A2(n_869), .B(n_912), .Y(n_1009) );
NAND2x1p5_ASAP7_75t_L g1010 ( .A(n_856), .B(n_918), .Y(n_1010) );
INVx1_ASAP7_75t_L g1011 ( .A(n_844), .Y(n_1011) );
BUFx2_ASAP7_75t_L g1012 ( .A(n_878), .Y(n_1012) );
INVx1_ASAP7_75t_L g1013 ( .A(n_861), .Y(n_1013) );
AOI22xp33_ASAP7_75t_L g1014 ( .A1(n_841), .A2(n_907), .B1(n_827), .B2(n_821), .Y(n_1014) );
CKINVDCx5p33_ASAP7_75t_R g1015 ( .A(n_799), .Y(n_1015) );
NOR2xp33_ASAP7_75t_L g1016 ( .A(n_865), .B(n_850), .Y(n_1016) );
NOR2xp33_ASAP7_75t_L g1017 ( .A(n_899), .B(n_868), .Y(n_1017) );
AOI21xp5_ASAP7_75t_L g1018 ( .A1(n_837), .A2(n_854), .B(n_889), .Y(n_1018) );
A2O1A1Ixp33_ASAP7_75t_L g1019 ( .A1(n_904), .A2(n_915), .B(n_871), .C(n_812), .Y(n_1019) );
OAI21x1_ASAP7_75t_L g1020 ( .A1(n_930), .A2(n_936), .B(n_934), .Y(n_1020) );
INVxp67_ASAP7_75t_SL g1021 ( .A(n_878), .Y(n_1021) );
BUFx8_ASAP7_75t_L g1022 ( .A(n_878), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_892), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_892), .Y(n_1024) );
OR2x2_ASAP7_75t_L g1025 ( .A(n_877), .B(n_903), .Y(n_1025) );
AND2x2_ASAP7_75t_L g1026 ( .A(n_845), .B(n_834), .Y(n_1026) );
CKINVDCx20_ASAP7_75t_R g1027 ( .A(n_895), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_895), .Y(n_1028) );
CKINVDCx20_ASAP7_75t_R g1029 ( .A(n_845), .Y(n_1029) );
INVx1_ASAP7_75t_L g1030 ( .A(n_834), .Y(n_1030) );
AND2x2_ASAP7_75t_L g1031 ( .A(n_834), .B(n_864), .Y(n_1031) );
AO21x2_ASAP7_75t_L g1032 ( .A1(n_919), .A2(n_917), .B(n_888), .Y(n_1032) );
INVx1_ASAP7_75t_L g1033 ( .A(n_817), .Y(n_1033) );
OA21x2_ASAP7_75t_L g1034 ( .A1(n_817), .A2(n_864), .B(n_880), .Y(n_1034) );
OAI21x1_ASAP7_75t_SL g1035 ( .A1(n_817), .A2(n_864), .B(n_880), .Y(n_1035) );
AOI21xp5_ASAP7_75t_L g1036 ( .A1(n_802), .A2(n_800), .B(n_790), .Y(n_1036) );
A2O1A1Ixp33_ASAP7_75t_L g1037 ( .A1(n_881), .A2(n_602), .B(n_853), .C(n_574), .Y(n_1037) );
INVx2_ASAP7_75t_L g1038 ( .A(n_806), .Y(n_1038) );
AO31x2_ASAP7_75t_L g1039 ( .A1(n_840), .A2(n_811), .A3(n_908), .B(n_896), .Y(n_1039) );
NAND2xp5_ASAP7_75t_L g1040 ( .A(n_909), .B(n_574), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1041 ( .A(n_798), .Y(n_1041) );
INVx1_ASAP7_75t_L g1042 ( .A(n_814), .Y(n_1042) );
AND2x2_ASAP7_75t_L g1043 ( .A(n_855), .B(n_792), .Y(n_1043) );
OA21x2_ASAP7_75t_L g1044 ( .A1(n_802), .A2(n_926), .B(n_773), .Y(n_1044) );
AOI21xp5_ASAP7_75t_L g1045 ( .A1(n_802), .A2(n_800), .B(n_790), .Y(n_1045) );
INVx2_ASAP7_75t_L g1046 ( .A(n_806), .Y(n_1046) );
INVx2_ASAP7_75t_L g1047 ( .A(n_806), .Y(n_1047) );
INVx2_ASAP7_75t_L g1048 ( .A(n_806), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1049 ( .A(n_855), .B(n_792), .Y(n_1049) );
OR2x2_ASAP7_75t_L g1050 ( .A(n_855), .B(n_792), .Y(n_1050) );
AO31x2_ASAP7_75t_L g1051 ( .A1(n_840), .A2(n_811), .A3(n_908), .B(n_896), .Y(n_1051) );
AND2x4_ASAP7_75t_L g1052 ( .A(n_937), .B(n_813), .Y(n_1052) );
A2O1A1Ixp33_ASAP7_75t_L g1053 ( .A1(n_881), .A2(n_602), .B(n_853), .C(n_574), .Y(n_1053) );
INVx4_ASAP7_75t_L g1054 ( .A(n_798), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_911), .Y(n_1055) );
NAND2x1p5_ASAP7_75t_L g1056 ( .A(n_902), .B(n_783), .Y(n_1056) );
OAI22xp5_ASAP7_75t_L g1057 ( .A1(n_875), .A2(n_574), .B1(n_582), .B2(n_605), .Y(n_1057) );
A2O1A1Ixp33_ASAP7_75t_L g1058 ( .A1(n_881), .A2(n_602), .B(n_853), .C(n_574), .Y(n_1058) );
INVx2_ASAP7_75t_SL g1059 ( .A(n_798), .Y(n_1059) );
NAND2xp5_ASAP7_75t_L g1060 ( .A(n_909), .B(n_574), .Y(n_1060) );
AND2x2_ASAP7_75t_L g1061 ( .A(n_855), .B(n_792), .Y(n_1061) );
NAND2xp5_ASAP7_75t_L g1062 ( .A(n_909), .B(n_574), .Y(n_1062) );
INVx2_ASAP7_75t_L g1063 ( .A(n_806), .Y(n_1063) );
INVx2_ASAP7_75t_L g1064 ( .A(n_806), .Y(n_1064) );
INVx3_ASAP7_75t_L g1065 ( .A(n_902), .Y(n_1065) );
AOI21xp33_ASAP7_75t_L g1066 ( .A1(n_865), .A2(n_881), .B(n_808), .Y(n_1066) );
INVx1_ASAP7_75t_L g1067 ( .A(n_814), .Y(n_1067) );
AOI22xp33_ASAP7_75t_L g1068 ( .A1(n_875), .A2(n_582), .B1(n_574), .B2(n_826), .Y(n_1068) );
INVx3_ASAP7_75t_L g1069 ( .A(n_902), .Y(n_1069) );
INVx1_ASAP7_75t_L g1070 ( .A(n_814), .Y(n_1070) );
INVx2_ASAP7_75t_L g1071 ( .A(n_806), .Y(n_1071) );
OR2x2_ASAP7_75t_L g1072 ( .A(n_855), .B(n_792), .Y(n_1072) );
AOI21xp5_ASAP7_75t_L g1073 ( .A1(n_802), .A2(n_800), .B(n_790), .Y(n_1073) );
INVx1_ASAP7_75t_L g1074 ( .A(n_814), .Y(n_1074) );
NAND2xp5_ASAP7_75t_L g1075 ( .A(n_909), .B(n_574), .Y(n_1075) );
NAND2xp5_ASAP7_75t_L g1076 ( .A(n_909), .B(n_574), .Y(n_1076) );
INVx1_ASAP7_75t_L g1077 ( .A(n_993), .Y(n_1077) );
HB1xp67_ASAP7_75t_L g1078 ( .A(n_946), .Y(n_1078) );
AO21x2_ASAP7_75t_L g1079 ( .A1(n_1036), .A2(n_1073), .B(n_1045), .Y(n_1079) );
INVx1_ASAP7_75t_L g1080 ( .A(n_940), .Y(n_1080) );
INVx1_ASAP7_75t_L g1081 ( .A(n_1042), .Y(n_1081) );
INVx3_ASAP7_75t_L g1082 ( .A(n_942), .Y(n_1082) );
OR2x2_ASAP7_75t_L g1083 ( .A(n_958), .B(n_1055), .Y(n_1083) );
OAI21xp5_ASAP7_75t_L g1084 ( .A1(n_1037), .A2(n_1058), .B(n_1053), .Y(n_1084) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_1056), .Y(n_1085) );
AND2x2_ASAP7_75t_L g1086 ( .A(n_943), .B(n_1038), .Y(n_1086) );
INVx1_ASAP7_75t_SL g1087 ( .A(n_967), .Y(n_1087) );
INVx2_ASAP7_75t_L g1088 ( .A(n_944), .Y(n_1088) );
INVx3_ASAP7_75t_L g1089 ( .A(n_942), .Y(n_1089) );
AND2x4_ASAP7_75t_L g1090 ( .A(n_1021), .B(n_1012), .Y(n_1090) );
AND2x2_ASAP7_75t_L g1091 ( .A(n_1046), .B(n_1047), .Y(n_1091) );
BUFx2_ASAP7_75t_L g1092 ( .A(n_997), .Y(n_1092) );
CKINVDCx20_ASAP7_75t_R g1093 ( .A(n_953), .Y(n_1093) );
OR2x2_ASAP7_75t_L g1094 ( .A(n_958), .B(n_1055), .Y(n_1094) );
INVx1_ASAP7_75t_L g1095 ( .A(n_1067), .Y(n_1095) );
AND2x2_ASAP7_75t_L g1096 ( .A(n_1048), .B(n_1063), .Y(n_1096) );
INVx1_ASAP7_75t_L g1097 ( .A(n_994), .Y(n_1097) );
NAND2x1p5_ASAP7_75t_L g1098 ( .A(n_942), .B(n_1065), .Y(n_1098) );
OAI21xp5_ASAP7_75t_L g1099 ( .A1(n_1016), .A2(n_1019), .B(n_1018), .Y(n_1099) );
AND2x2_ASAP7_75t_L g1100 ( .A(n_1064), .B(n_1071), .Y(n_1100) );
INVxp67_ASAP7_75t_L g1101 ( .A(n_1043), .Y(n_1101) );
NAND3xp33_ASAP7_75t_SL g1102 ( .A(n_1015), .B(n_1068), .C(n_963), .Y(n_1102) );
INVx3_ASAP7_75t_L g1103 ( .A(n_1056), .Y(n_1103) );
NAND2xp5_ASAP7_75t_L g1104 ( .A(n_1040), .B(n_1060), .Y(n_1104) );
AO21x2_ASAP7_75t_L g1105 ( .A1(n_961), .A2(n_1035), .B(n_1000), .Y(n_1105) );
NAND2xp5_ASAP7_75t_L g1106 ( .A(n_1040), .B(n_1060), .Y(n_1106) );
INVx1_ASAP7_75t_L g1107 ( .A(n_1011), .Y(n_1107) );
INVx1_ASAP7_75t_L g1108 ( .A(n_1013), .Y(n_1108) );
AND2x2_ASAP7_75t_L g1109 ( .A(n_947), .B(n_960), .Y(n_1109) );
BUFx2_ASAP7_75t_L g1110 ( .A(n_979), .Y(n_1110) );
INVx1_ASAP7_75t_L g1111 ( .A(n_1028), .Y(n_1111) );
CKINVDCx20_ASAP7_75t_R g1112 ( .A(n_953), .Y(n_1112) );
AO21x2_ASAP7_75t_L g1113 ( .A1(n_1023), .A2(n_1024), .B(n_968), .Y(n_1113) );
INVx2_ASAP7_75t_L g1114 ( .A(n_1044), .Y(n_1114) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_962), .Y(n_1115) );
INVx1_ASAP7_75t_L g1116 ( .A(n_1070), .Y(n_1116) );
HB1xp67_ASAP7_75t_L g1117 ( .A(n_962), .Y(n_1117) );
OR2x2_ASAP7_75t_L g1118 ( .A(n_945), .B(n_965), .Y(n_1118) );
AND2x2_ASAP7_75t_L g1119 ( .A(n_1074), .B(n_945), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_977), .Y(n_1120) );
AND2x4_ASAP7_75t_L g1121 ( .A(n_1006), .B(n_990), .Y(n_1121) );
INVx1_ASAP7_75t_L g1122 ( .A(n_956), .Y(n_1122) );
HB1xp67_ASAP7_75t_L g1123 ( .A(n_964), .Y(n_1123) );
BUFx3_ASAP7_75t_L g1124 ( .A(n_971), .Y(n_1124) );
CKINVDCx20_ASAP7_75t_R g1125 ( .A(n_1002), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g1126 ( .A1(n_1068), .A2(n_1057), .B1(n_1027), .B2(n_1029), .Y(n_1126) );
OR2x2_ASAP7_75t_L g1127 ( .A(n_1050), .B(n_1072), .Y(n_1127) );
AND2x4_ASAP7_75t_L g1128 ( .A(n_964), .B(n_1065), .Y(n_1128) );
INVx1_ASAP7_75t_L g1129 ( .A(n_1033), .Y(n_1129) );
OR2x2_ASAP7_75t_L g1130 ( .A(n_969), .B(n_1025), .Y(n_1130) );
INVxp67_ASAP7_75t_L g1131 ( .A(n_1049), .Y(n_1131) );
AOI21xp5_ASAP7_75t_SL g1132 ( .A1(n_948), .A2(n_952), .B(n_949), .Y(n_1132) );
AND2x2_ASAP7_75t_L g1133 ( .A(n_970), .B(n_1017), .Y(n_1133) );
INVxp67_ASAP7_75t_L g1134 ( .A(n_1061), .Y(n_1134) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1030), .Y(n_1135) );
AND2x2_ASAP7_75t_L g1136 ( .A(n_1017), .B(n_999), .Y(n_1136) );
AO21x2_ASAP7_75t_L g1137 ( .A1(n_1032), .A2(n_1018), .B(n_984), .Y(n_1137) );
AND2x2_ASAP7_75t_L g1138 ( .A(n_1031), .B(n_1026), .Y(n_1138) );
OA21x2_ASAP7_75t_L g1139 ( .A1(n_984), .A2(n_1009), .B(n_1001), .Y(n_1139) );
INVx1_ASAP7_75t_L g1140 ( .A(n_1034), .Y(n_1140) );
AND2x2_ASAP7_75t_L g1141 ( .A(n_975), .B(n_976), .Y(n_1141) );
AND2x4_ASAP7_75t_L g1142 ( .A(n_1069), .B(n_950), .Y(n_1142) );
INVx3_ASAP7_75t_L g1143 ( .A(n_1069), .Y(n_1143) );
INVx1_ASAP7_75t_L g1144 ( .A(n_959), .Y(n_1144) );
INVx1_ASAP7_75t_L g1145 ( .A(n_959), .Y(n_1145) );
INVx1_ASAP7_75t_L g1146 ( .A(n_985), .Y(n_1146) );
HB1xp67_ASAP7_75t_L g1147 ( .A(n_969), .Y(n_1147) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1034), .Y(n_1148) );
BUFx2_ASAP7_75t_L g1149 ( .A(n_1022), .Y(n_1149) );
INVx1_ASAP7_75t_L g1150 ( .A(n_951), .Y(n_1150) );
CKINVDCx5p33_ASAP7_75t_R g1151 ( .A(n_1022), .Y(n_1151) );
OAI21xp5_ASAP7_75t_L g1152 ( .A1(n_1016), .A2(n_1014), .B(n_1066), .Y(n_1152) );
INVx2_ASAP7_75t_L g1153 ( .A(n_1039), .Y(n_1153) );
AND2x2_ASAP7_75t_L g1154 ( .A(n_978), .B(n_1076), .Y(n_1154) );
BUFx2_ASAP7_75t_L g1155 ( .A(n_1010), .Y(n_1155) );
INVx3_ASAP7_75t_L g1156 ( .A(n_1010), .Y(n_1156) );
NAND2xp5_ASAP7_75t_L g1157 ( .A(n_1062), .B(n_1076), .Y(n_1157) );
INVx2_ASAP7_75t_L g1158 ( .A(n_1039), .Y(n_1158) );
INVx2_ASAP7_75t_L g1159 ( .A(n_1051), .Y(n_1159) );
NAND2xp5_ASAP7_75t_L g1160 ( .A(n_1062), .B(n_1075), .Y(n_1160) );
BUFx4f_ASAP7_75t_L g1161 ( .A(n_974), .Y(n_1161) );
INVx1_ASAP7_75t_L g1162 ( .A(n_998), .Y(n_1162) );
HB1xp67_ASAP7_75t_L g1163 ( .A(n_983), .Y(n_1163) );
INVx1_ASAP7_75t_L g1164 ( .A(n_998), .Y(n_1164) );
OAI21xp5_ASAP7_75t_L g1165 ( .A1(n_1014), .A2(n_995), .B(n_986), .Y(n_1165) );
INVx1_ASAP7_75t_L g1166 ( .A(n_998), .Y(n_1166) );
INVx2_ASAP7_75t_L g1167 ( .A(n_1051), .Y(n_1167) );
AO21x2_ASAP7_75t_L g1168 ( .A1(n_1020), .A2(n_995), .B(n_986), .Y(n_1168) );
INVx1_ASAP7_75t_L g1169 ( .A(n_989), .Y(n_1169) );
INVx2_ASAP7_75t_L g1170 ( .A(n_1051), .Y(n_1170) );
HB1xp67_ASAP7_75t_L g1171 ( .A(n_988), .Y(n_1171) );
AOI21x1_ASAP7_75t_L g1172 ( .A1(n_980), .A2(n_973), .B(n_1007), .Y(n_1172) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_1138), .B(n_989), .Y(n_1173) );
BUFx3_ASAP7_75t_L g1174 ( .A(n_1124), .Y(n_1174) );
OR2x2_ASAP7_75t_L g1175 ( .A(n_1130), .B(n_989), .Y(n_1175) );
AND2x2_ASAP7_75t_L g1176 ( .A(n_1138), .B(n_1003), .Y(n_1176) );
INVx1_ASAP7_75t_L g1177 ( .A(n_1120), .Y(n_1177) );
INVx4_ASAP7_75t_L g1178 ( .A(n_1161), .Y(n_1178) );
AND2x2_ASAP7_75t_L g1179 ( .A(n_1136), .B(n_991), .Y(n_1179) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1146), .Y(n_1180) );
OR2x2_ASAP7_75t_L g1181 ( .A(n_1130), .B(n_996), .Y(n_1181) );
AND2x2_ASAP7_75t_L g1182 ( .A(n_1099), .B(n_1004), .Y(n_1182) );
AND2x4_ASAP7_75t_SL g1183 ( .A(n_1103), .B(n_1054), .Y(n_1183) );
AND2x2_ASAP7_75t_L g1184 ( .A(n_1119), .B(n_1004), .Y(n_1184) );
AND2x2_ASAP7_75t_L g1185 ( .A(n_1119), .B(n_1004), .Y(n_1185) );
INVx1_ASAP7_75t_L g1186 ( .A(n_1080), .Y(n_1186) );
BUFx4f_ASAP7_75t_L g1187 ( .A(n_1103), .Y(n_1187) );
AND2x2_ASAP7_75t_L g1188 ( .A(n_1133), .B(n_939), .Y(n_1188) );
AND2x4_ASAP7_75t_L g1189 ( .A(n_1077), .B(n_1097), .Y(n_1189) );
AND2x2_ASAP7_75t_L g1190 ( .A(n_1133), .B(n_981), .Y(n_1190) );
INVx1_ASAP7_75t_L g1191 ( .A(n_1081), .Y(n_1191) );
AND2x2_ASAP7_75t_L g1192 ( .A(n_1088), .B(n_973), .Y(n_1192) );
NAND2xp5_ASAP7_75t_L g1193 ( .A(n_1154), .B(n_972), .Y(n_1193) );
AND2x4_ASAP7_75t_L g1194 ( .A(n_1077), .B(n_1054), .Y(n_1194) );
INVx1_ASAP7_75t_L g1195 ( .A(n_1095), .Y(n_1195) );
INVx3_ASAP7_75t_L g1196 ( .A(n_1090), .Y(n_1196) );
HB1xp67_ASAP7_75t_L g1197 ( .A(n_1110), .Y(n_1197) );
AND2x2_ASAP7_75t_SL g1198 ( .A(n_1161), .B(n_1005), .Y(n_1198) );
NAND2xp5_ASAP7_75t_L g1199 ( .A(n_1154), .B(n_972), .Y(n_1199) );
OR2x2_ASAP7_75t_L g1200 ( .A(n_1083), .B(n_1059), .Y(n_1200) );
BUFx2_ASAP7_75t_L g1201 ( .A(n_1161), .Y(n_1201) );
INVx1_ASAP7_75t_L g1202 ( .A(n_1116), .Y(n_1202) );
OAI33xp33_ASAP7_75t_L g1203 ( .A1(n_1126), .A2(n_1008), .A3(n_938), .B1(n_941), .B2(n_1041), .B3(n_954), .Y(n_1203) );
INVx1_ASAP7_75t_L g1204 ( .A(n_1141), .Y(n_1204) );
AND2x4_ASAP7_75t_L g1205 ( .A(n_1097), .B(n_992), .Y(n_1205) );
AND2x2_ASAP7_75t_L g1206 ( .A(n_1135), .B(n_1052), .Y(n_1206) );
NAND3xp33_ASAP7_75t_SL g1207 ( .A(n_1093), .B(n_1005), .C(n_966), .Y(n_1207) );
AND2x2_ASAP7_75t_L g1208 ( .A(n_1135), .B(n_957), .Y(n_1208) );
INVxp67_ASAP7_75t_L g1209 ( .A(n_1124), .Y(n_1209) );
AND2x2_ASAP7_75t_L g1210 ( .A(n_1140), .B(n_957), .Y(n_1210) );
AND2x2_ASAP7_75t_L g1211 ( .A(n_1140), .B(n_992), .Y(n_1211) );
INVx2_ASAP7_75t_SL g1212 ( .A(n_1128), .Y(n_1212) );
INVx1_ASAP7_75t_L g1213 ( .A(n_1141), .Y(n_1213) );
NAND2xp5_ASAP7_75t_SL g1214 ( .A(n_1152), .B(n_982), .Y(n_1214) );
AND2x2_ASAP7_75t_L g1215 ( .A(n_1148), .B(n_955), .Y(n_1215) );
AND2x2_ASAP7_75t_L g1216 ( .A(n_1148), .B(n_987), .Y(n_1216) );
AND2x2_ASAP7_75t_L g1217 ( .A(n_1129), .B(n_1086), .Y(n_1217) );
BUFx4f_ASAP7_75t_L g1218 ( .A(n_1149), .Y(n_1218) );
AND2x2_ASAP7_75t_L g1219 ( .A(n_1129), .B(n_1086), .Y(n_1219) );
AND2x4_ASAP7_75t_L g1220 ( .A(n_1107), .B(n_1108), .Y(n_1220) );
HB1xp67_ASAP7_75t_L g1221 ( .A(n_1110), .Y(n_1221) );
AND2x2_ASAP7_75t_L g1222 ( .A(n_1091), .B(n_1096), .Y(n_1222) );
INVx2_ASAP7_75t_SL g1223 ( .A(n_1128), .Y(n_1223) );
INVx2_ASAP7_75t_L g1224 ( .A(n_1114), .Y(n_1224) );
AND2x2_ASAP7_75t_L g1225 ( .A(n_1100), .B(n_1109), .Y(n_1225) );
AND2x2_ASAP7_75t_L g1226 ( .A(n_1109), .B(n_1111), .Y(n_1226) );
AND2x2_ASAP7_75t_L g1227 ( .A(n_1111), .B(n_1168), .Y(n_1227) );
AND2x2_ASAP7_75t_L g1228 ( .A(n_1168), .B(n_1169), .Y(n_1228) );
AND2x2_ASAP7_75t_L g1229 ( .A(n_1168), .B(n_1169), .Y(n_1229) );
INVx1_ASAP7_75t_L g1230 ( .A(n_1118), .Y(n_1230) );
AND2x2_ASAP7_75t_L g1231 ( .A(n_1162), .B(n_1164), .Y(n_1231) );
CKINVDCx8_ASAP7_75t_R g1232 ( .A(n_1149), .Y(n_1232) );
NAND2xp5_ASAP7_75t_L g1233 ( .A(n_1118), .B(n_1165), .Y(n_1233) );
NAND2xp5_ASAP7_75t_L g1234 ( .A(n_1144), .B(n_1145), .Y(n_1234) );
AOI22xp33_ASAP7_75t_L g1235 ( .A1(n_1102), .A2(n_1084), .B1(n_1101), .B2(n_1134), .Y(n_1235) );
AND2x2_ASAP7_75t_L g1236 ( .A(n_1162), .B(n_1164), .Y(n_1236) );
NAND2xp5_ASAP7_75t_L g1237 ( .A(n_1104), .B(n_1106), .Y(n_1237) );
INVx1_ASAP7_75t_L g1238 ( .A(n_1122), .Y(n_1238) );
AND2x2_ASAP7_75t_L g1239 ( .A(n_1166), .B(n_1137), .Y(n_1239) );
OR2x2_ASAP7_75t_L g1240 ( .A(n_1083), .B(n_1094), .Y(n_1240) );
OR2x2_ASAP7_75t_L g1241 ( .A(n_1094), .B(n_1092), .Y(n_1241) );
AND2x2_ASAP7_75t_L g1242 ( .A(n_1166), .B(n_1137), .Y(n_1242) );
AND2x2_ASAP7_75t_L g1243 ( .A(n_1137), .B(n_1092), .Y(n_1243) );
OR2x2_ASAP7_75t_L g1244 ( .A(n_1127), .B(n_1078), .Y(n_1244) );
AND2x2_ASAP7_75t_L g1245 ( .A(n_1172), .B(n_1150), .Y(n_1245) );
NAND2xp5_ASAP7_75t_L g1246 ( .A(n_1157), .B(n_1160), .Y(n_1246) );
OR2x2_ASAP7_75t_L g1247 ( .A(n_1127), .B(n_1147), .Y(n_1247) );
INVxp67_ASAP7_75t_SL g1248 ( .A(n_1171), .Y(n_1248) );
OR2x2_ASAP7_75t_L g1249 ( .A(n_1131), .B(n_1123), .Y(n_1249) );
OR2x2_ASAP7_75t_L g1250 ( .A(n_1240), .B(n_1105), .Y(n_1250) );
INVx2_ASAP7_75t_L g1251 ( .A(n_1224), .Y(n_1251) );
AND2x2_ASAP7_75t_L g1252 ( .A(n_1184), .B(n_1105), .Y(n_1252) );
NAND2xp5_ASAP7_75t_L g1253 ( .A(n_1204), .B(n_1115), .Y(n_1253) );
OR2x2_ASAP7_75t_L g1254 ( .A(n_1240), .B(n_1105), .Y(n_1254) );
AND2x2_ASAP7_75t_L g1255 ( .A(n_1184), .B(n_1153), .Y(n_1255) );
NAND2xp5_ASAP7_75t_L g1256 ( .A(n_1213), .B(n_1117), .Y(n_1256) );
HB1xp67_ASAP7_75t_L g1257 ( .A(n_1197), .Y(n_1257) );
AND2x2_ASAP7_75t_L g1258 ( .A(n_1185), .B(n_1153), .Y(n_1258) );
AND2x2_ASAP7_75t_L g1259 ( .A(n_1173), .B(n_1158), .Y(n_1259) );
INVx3_ASAP7_75t_L g1260 ( .A(n_1189), .Y(n_1260) );
OR2x2_ASAP7_75t_L g1261 ( .A(n_1241), .B(n_1159), .Y(n_1261) );
AND2x2_ASAP7_75t_L g1262 ( .A(n_1173), .B(n_1159), .Y(n_1262) );
INVx1_ASAP7_75t_L g1263 ( .A(n_1189), .Y(n_1263) );
INVxp67_ASAP7_75t_SL g1264 ( .A(n_1248), .Y(n_1264) );
INVx1_ASAP7_75t_L g1265 ( .A(n_1189), .Y(n_1265) );
AND2x2_ASAP7_75t_L g1266 ( .A(n_1182), .B(n_1167), .Y(n_1266) );
INVx1_ASAP7_75t_L g1267 ( .A(n_1220), .Y(n_1267) );
INVxp67_ASAP7_75t_SL g1268 ( .A(n_1221), .Y(n_1268) );
HB1xp67_ASAP7_75t_L g1269 ( .A(n_1176), .Y(n_1269) );
NOR2xp33_ASAP7_75t_L g1270 ( .A(n_1203), .B(n_1087), .Y(n_1270) );
INVx1_ASAP7_75t_L g1271 ( .A(n_1220), .Y(n_1271) );
HB1xp67_ASAP7_75t_L g1272 ( .A(n_1176), .Y(n_1272) );
INVx2_ASAP7_75t_SL g1273 ( .A(n_1194), .Y(n_1273) );
BUFx3_ASAP7_75t_L g1274 ( .A(n_1174), .Y(n_1274) );
AND2x4_ASAP7_75t_L g1275 ( .A(n_1239), .B(n_1242), .Y(n_1275) );
AND2x2_ASAP7_75t_L g1276 ( .A(n_1182), .B(n_1167), .Y(n_1276) );
INVx1_ASAP7_75t_L g1277 ( .A(n_1220), .Y(n_1277) );
INVx1_ASAP7_75t_L g1278 ( .A(n_1245), .Y(n_1278) );
AND2x2_ASAP7_75t_L g1279 ( .A(n_1245), .B(n_1170), .Y(n_1279) );
INVx3_ASAP7_75t_L g1280 ( .A(n_1194), .Y(n_1280) );
NAND2xp5_ASAP7_75t_L g1281 ( .A(n_1222), .B(n_1163), .Y(n_1281) );
INVx1_ASAP7_75t_L g1282 ( .A(n_1231), .Y(n_1282) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1231), .Y(n_1283) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_1225), .Y(n_1284) );
INVx1_ASAP7_75t_L g1285 ( .A(n_1236), .Y(n_1285) );
NAND2xp5_ASAP7_75t_L g1286 ( .A(n_1225), .B(n_1230), .Y(n_1286) );
AND2x2_ASAP7_75t_L g1287 ( .A(n_1217), .B(n_1170), .Y(n_1287) );
OAI22xp5_ASAP7_75t_SL g1288 ( .A1(n_1232), .A2(n_1093), .B1(n_1112), .B2(n_1125), .Y(n_1288) );
NAND2x1p5_ASAP7_75t_L g1289 ( .A(n_1178), .B(n_1090), .Y(n_1289) );
AND2x2_ASAP7_75t_L g1290 ( .A(n_1217), .B(n_1172), .Y(n_1290) );
AND2x2_ASAP7_75t_L g1291 ( .A(n_1219), .B(n_1113), .Y(n_1291) );
AND2x2_ASAP7_75t_L g1292 ( .A(n_1219), .B(n_1113), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1293 ( .A(n_1200), .Y(n_1293) );
AND2x2_ASAP7_75t_L g1294 ( .A(n_1242), .B(n_1113), .Y(n_1294) );
OR2x2_ASAP7_75t_L g1295 ( .A(n_1241), .B(n_1079), .Y(n_1295) );
AND2x2_ASAP7_75t_L g1296 ( .A(n_1226), .B(n_1139), .Y(n_1296) );
INVx1_ASAP7_75t_L g1297 ( .A(n_1236), .Y(n_1297) );
INVx3_ASAP7_75t_L g1298 ( .A(n_1194), .Y(n_1298) );
NAND3xp33_ASAP7_75t_L g1299 ( .A(n_1214), .B(n_1235), .C(n_1232), .Y(n_1299) );
NAND2xp5_ASAP7_75t_L g1300 ( .A(n_1226), .B(n_1121), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1301 ( .A(n_1227), .B(n_1139), .Y(n_1301) );
AND2x2_ASAP7_75t_L g1302 ( .A(n_1275), .B(n_1243), .Y(n_1302) );
AND2x2_ASAP7_75t_L g1303 ( .A(n_1275), .B(n_1243), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1304 ( .A(n_1284), .B(n_1216), .Y(n_1304) );
AND2x2_ASAP7_75t_L g1305 ( .A(n_1275), .B(n_1227), .Y(n_1305) );
AND2x2_ASAP7_75t_L g1306 ( .A(n_1275), .B(n_1228), .Y(n_1306) );
INVx1_ASAP7_75t_L g1307 ( .A(n_1257), .Y(n_1307) );
NOR2xp33_ASAP7_75t_L g1308 ( .A(n_1288), .B(n_1207), .Y(n_1308) );
INVx1_ASAP7_75t_L g1309 ( .A(n_1293), .Y(n_1309) );
INVx1_ASAP7_75t_L g1310 ( .A(n_1264), .Y(n_1310) );
INVx1_ASAP7_75t_L g1311 ( .A(n_1282), .Y(n_1311) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1252), .B(n_1228), .Y(n_1312) );
INVx1_ASAP7_75t_L g1313 ( .A(n_1282), .Y(n_1313) );
AND2x2_ASAP7_75t_L g1314 ( .A(n_1252), .B(n_1229), .Y(n_1314) );
NAND2xp5_ASAP7_75t_L g1315 ( .A(n_1283), .B(n_1216), .Y(n_1315) );
INVx3_ASAP7_75t_L g1316 ( .A(n_1280), .Y(n_1316) );
INVx1_ASAP7_75t_L g1317 ( .A(n_1283), .Y(n_1317) );
INVx1_ASAP7_75t_L g1318 ( .A(n_1285), .Y(n_1318) );
NAND2xp5_ASAP7_75t_L g1319 ( .A(n_1285), .B(n_1247), .Y(n_1319) );
INVx1_ASAP7_75t_L g1320 ( .A(n_1297), .Y(n_1320) );
INVx1_ASAP7_75t_L g1321 ( .A(n_1278), .Y(n_1321) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1296), .B(n_1229), .Y(n_1322) );
AND2x4_ASAP7_75t_SL g1323 ( .A(n_1280), .B(n_1178), .Y(n_1323) );
NOR2xp33_ASAP7_75t_L g1324 ( .A(n_1288), .B(n_1209), .Y(n_1324) );
AND2x2_ASAP7_75t_L g1325 ( .A(n_1296), .B(n_1192), .Y(n_1325) );
INVxp33_ASAP7_75t_SL g1326 ( .A(n_1269), .Y(n_1326) );
INVx1_ASAP7_75t_L g1327 ( .A(n_1297), .Y(n_1327) );
INVx2_ASAP7_75t_L g1328 ( .A(n_1278), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1329 ( .A(n_1291), .B(n_1192), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1291), .B(n_1211), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1331 ( .A(n_1286), .B(n_1247), .Y(n_1331) );
INVx1_ASAP7_75t_L g1332 ( .A(n_1268), .Y(n_1332) );
INVx2_ASAP7_75t_L g1333 ( .A(n_1251), .Y(n_1333) );
INVx1_ASAP7_75t_L g1334 ( .A(n_1272), .Y(n_1334) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1292), .B(n_1211), .Y(n_1335) );
OAI221xp5_ASAP7_75t_L g1336 ( .A1(n_1299), .A2(n_1218), .B1(n_1199), .B2(n_1193), .C(n_1246), .Y(n_1336) );
OR2x2_ASAP7_75t_L g1337 ( .A(n_1250), .B(n_1175), .Y(n_1337) );
HB1xp67_ASAP7_75t_L g1338 ( .A(n_1274), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1339 ( .A(n_1292), .B(n_1233), .Y(n_1339) );
NAND2xp5_ASAP7_75t_L g1340 ( .A(n_1290), .B(n_1244), .Y(n_1340) );
OR2x2_ASAP7_75t_L g1341 ( .A(n_1250), .B(n_1175), .Y(n_1341) );
OR2x2_ASAP7_75t_L g1342 ( .A(n_1254), .B(n_1181), .Y(n_1342) );
OR2x2_ASAP7_75t_L g1343 ( .A(n_1254), .B(n_1181), .Y(n_1343) );
OR2x2_ASAP7_75t_L g1344 ( .A(n_1295), .B(n_1215), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1290), .B(n_1215), .Y(n_1345) );
NAND2xp5_ASAP7_75t_L g1346 ( .A(n_1287), .B(n_1186), .Y(n_1346) );
NAND2xp5_ASAP7_75t_L g1347 ( .A(n_1287), .B(n_1191), .Y(n_1347) );
OR2x2_ASAP7_75t_L g1348 ( .A(n_1295), .B(n_1210), .Y(n_1348) );
AND2x4_ASAP7_75t_L g1349 ( .A(n_1260), .B(n_1196), .Y(n_1349) );
INVx1_ASAP7_75t_L g1350 ( .A(n_1310), .Y(n_1350) );
AND2x2_ASAP7_75t_L g1351 ( .A(n_1322), .B(n_1294), .Y(n_1351) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1322), .B(n_1294), .Y(n_1352) );
INVx1_ASAP7_75t_L g1353 ( .A(n_1321), .Y(n_1353) );
INVx1_ASAP7_75t_L g1354 ( .A(n_1342), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1355 ( .A(n_1339), .B(n_1301), .Y(n_1355) );
INVxp67_ASAP7_75t_L g1356 ( .A(n_1338), .Y(n_1356) );
HB1xp67_ASAP7_75t_L g1357 ( .A(n_1326), .Y(n_1357) );
INVx1_ASAP7_75t_L g1358 ( .A(n_1342), .Y(n_1358) );
HB1xp67_ASAP7_75t_L g1359 ( .A(n_1326), .Y(n_1359) );
NOR2x1_ASAP7_75t_L g1360 ( .A(n_1308), .B(n_1274), .Y(n_1360) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1312), .B(n_1259), .Y(n_1361) );
INVx2_ASAP7_75t_SL g1362 ( .A(n_1323), .Y(n_1362) );
OR2x2_ASAP7_75t_L g1363 ( .A(n_1340), .B(n_1261), .Y(n_1363) );
AND2x2_ASAP7_75t_L g1364 ( .A(n_1314), .B(n_1259), .Y(n_1364) );
OR2x2_ASAP7_75t_L g1365 ( .A(n_1344), .B(n_1261), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1366 ( .A(n_1314), .B(n_1262), .Y(n_1366) );
INVxp67_ASAP7_75t_L g1367 ( .A(n_1324), .Y(n_1367) );
NOR2xp33_ASAP7_75t_L g1368 ( .A(n_1336), .B(n_1270), .Y(n_1368) );
OR2x2_ASAP7_75t_L g1369 ( .A(n_1343), .B(n_1344), .Y(n_1369) );
INVx2_ASAP7_75t_L g1370 ( .A(n_1333), .Y(n_1370) );
AND2x2_ASAP7_75t_L g1371 ( .A(n_1305), .B(n_1262), .Y(n_1371) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1343), .Y(n_1372) );
NOR2x1_ASAP7_75t_L g1373 ( .A(n_1332), .B(n_1112), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1311), .Y(n_1374) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1305), .B(n_1255), .Y(n_1375) );
OR2x2_ASAP7_75t_L g1376 ( .A(n_1345), .B(n_1279), .Y(n_1376) );
OR2x2_ASAP7_75t_L g1377 ( .A(n_1337), .B(n_1255), .Y(n_1377) );
AND2x2_ASAP7_75t_L g1378 ( .A(n_1306), .B(n_1258), .Y(n_1378) );
NAND2xp5_ASAP7_75t_L g1379 ( .A(n_1309), .B(n_1266), .Y(n_1379) );
NAND4xp25_ASAP7_75t_L g1380 ( .A(n_1307), .B(n_1188), .C(n_1256), .D(n_1253), .Y(n_1380) );
INVx1_ASAP7_75t_L g1381 ( .A(n_1313), .Y(n_1381) );
NAND2xp5_ASAP7_75t_L g1382 ( .A(n_1334), .B(n_1266), .Y(n_1382) );
NAND2xp5_ASAP7_75t_L g1383 ( .A(n_1330), .B(n_1276), .Y(n_1383) );
INVx1_ASAP7_75t_L g1384 ( .A(n_1317), .Y(n_1384) );
NAND2x1_ASAP7_75t_L g1385 ( .A(n_1362), .B(n_1316), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1386 ( .A(n_1351), .B(n_1306), .Y(n_1386) );
INVx1_ASAP7_75t_L g1387 ( .A(n_1369), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1388 ( .A(n_1367), .B(n_1331), .Y(n_1388) );
NOR2xp67_ASAP7_75t_SL g1389 ( .A(n_1362), .B(n_1151), .Y(n_1389) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1353), .Y(n_1390) );
INVx2_ASAP7_75t_L g1391 ( .A(n_1370), .Y(n_1391) );
OAI21xp33_ASAP7_75t_L g1392 ( .A1(n_1368), .A2(n_1303), .B(n_1302), .Y(n_1392) );
AOI21xp5_ASAP7_75t_L g1393 ( .A1(n_1360), .A2(n_1273), .B(n_1198), .Y(n_1393) );
NAND2xp5_ASAP7_75t_L g1394 ( .A(n_1354), .B(n_1330), .Y(n_1394) );
AOI21xp33_ASAP7_75t_L g1395 ( .A1(n_1368), .A2(n_1234), .B(n_1200), .Y(n_1395) );
NAND2xp5_ASAP7_75t_L g1396 ( .A(n_1358), .B(n_1335), .Y(n_1396) );
AOI21xp5_ASAP7_75t_L g1397 ( .A1(n_1380), .A2(n_1198), .B(n_1280), .Y(n_1397) );
INVx1_ASAP7_75t_L g1398 ( .A(n_1372), .Y(n_1398) );
NAND2xp5_ASAP7_75t_SL g1399 ( .A(n_1357), .B(n_1316), .Y(n_1399) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1351), .B(n_1302), .Y(n_1400) );
INVx1_ASAP7_75t_L g1401 ( .A(n_1365), .Y(n_1401) );
INVx1_ASAP7_75t_L g1402 ( .A(n_1365), .Y(n_1402) );
INVx2_ASAP7_75t_L g1403 ( .A(n_1370), .Y(n_1403) );
INVx2_ASAP7_75t_L g1404 ( .A(n_1350), .Y(n_1404) );
OR2x2_ASAP7_75t_L g1405 ( .A(n_1377), .B(n_1337), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1406 ( .A(n_1352), .B(n_1335), .Y(n_1406) );
A2O1A1Ixp33_ASAP7_75t_L g1407 ( .A1(n_1373), .A2(n_1201), .B(n_1298), .C(n_1187), .Y(n_1407) );
INVxp67_ASAP7_75t_L g1408 ( .A(n_1359), .Y(n_1408) );
OAI321xp33_ASAP7_75t_L g1409 ( .A1(n_1356), .A2(n_1341), .A3(n_1289), .B1(n_1277), .B2(n_1263), .C(n_1267), .Y(n_1409) );
OAI21xp5_ASAP7_75t_SL g1410 ( .A1(n_1393), .A2(n_1183), .B(n_1289), .Y(n_1410) );
NAND2xp5_ASAP7_75t_L g1411 ( .A(n_1401), .B(n_1352), .Y(n_1411) );
OAI22xp33_ASAP7_75t_L g1412 ( .A1(n_1385), .A2(n_1298), .B1(n_1376), .B2(n_1383), .Y(n_1412) );
INVx1_ASAP7_75t_L g1413 ( .A(n_1404), .Y(n_1413) );
INVx1_ASAP7_75t_L g1414 ( .A(n_1404), .Y(n_1414) );
OAI221xp5_ASAP7_75t_SL g1415 ( .A1(n_1392), .A2(n_1363), .B1(n_1348), .B2(n_1341), .C(n_1304), .Y(n_1415) );
INVx1_ASAP7_75t_L g1416 ( .A(n_1405), .Y(n_1416) );
A2O1A1Ixp33_ASAP7_75t_L g1417 ( .A1(n_1389), .A2(n_1183), .B(n_1366), .C(n_1364), .Y(n_1417) );
AOI221xp5_ASAP7_75t_L g1418 ( .A1(n_1395), .A2(n_1379), .B1(n_1382), .B2(n_1381), .C(n_1384), .Y(n_1418) );
INVxp67_ASAP7_75t_L g1419 ( .A(n_1408), .Y(n_1419) );
AOI222xp33_ASAP7_75t_L g1420 ( .A1(n_1388), .A2(n_1188), .B1(n_1319), .B2(n_1347), .C1(n_1346), .C2(n_1320), .Y(n_1420) );
AOI21xp5_ASAP7_75t_L g1421 ( .A1(n_1399), .A2(n_1355), .B(n_1363), .Y(n_1421) );
AOI322xp5_ASAP7_75t_L g1422 ( .A1(n_1387), .A2(n_1361), .A3(n_1371), .B1(n_1375), .B2(n_1378), .C1(n_1303), .C2(n_1325), .Y(n_1422) );
OAI22xp33_ASAP7_75t_L g1423 ( .A1(n_1409), .A2(n_1376), .B1(n_1289), .B2(n_1260), .Y(n_1423) );
NOR2xp33_ASAP7_75t_L g1424 ( .A(n_1402), .B(n_1125), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1398), .B(n_1318), .Y(n_1425) );
INVxp67_ASAP7_75t_L g1426 ( .A(n_1399), .Y(n_1426) );
NAND2xp5_ASAP7_75t_L g1427 ( .A(n_1386), .B(n_1406), .Y(n_1427) );
OAI22xp5_ASAP7_75t_L g1428 ( .A1(n_1407), .A2(n_1348), .B1(n_1315), .B2(n_1281), .Y(n_1428) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1390), .Y(n_1429) );
OAI211xp5_ASAP7_75t_SL g1430 ( .A1(n_1397), .A2(n_1249), .B(n_1237), .C(n_1374), .Y(n_1430) );
AOI22xp5_ASAP7_75t_L g1431 ( .A1(n_1386), .A2(n_1327), .B1(n_1349), .B2(n_1329), .Y(n_1431) );
O2A1O1Ixp33_ASAP7_75t_SL g1432 ( .A1(n_1394), .A2(n_1223), .B(n_1212), .C(n_1300), .Y(n_1432) );
NAND2xp5_ASAP7_75t_L g1433 ( .A(n_1396), .B(n_1328), .Y(n_1433) );
NAND2xp5_ASAP7_75t_L g1434 ( .A(n_1400), .B(n_1328), .Y(n_1434) );
NAND4xp25_ASAP7_75t_L g1435 ( .A(n_1391), .B(n_1190), .C(n_1249), .D(n_1179), .Y(n_1435) );
AOI221xp5_ASAP7_75t_L g1436 ( .A1(n_1403), .A2(n_1271), .B1(n_1267), .B2(n_1265), .C(n_1277), .Y(n_1436) );
XOR2x2_ASAP7_75t_L g1437 ( .A(n_1403), .B(n_1190), .Y(n_1437) );
A2O1A1Ixp33_ASAP7_75t_L g1438 ( .A1(n_1389), .A2(n_1187), .B(n_1349), .C(n_1329), .Y(n_1438) );
NAND2xp33_ASAP7_75t_SL g1439 ( .A(n_1428), .B(n_1410), .Y(n_1439) );
OAI221xp5_ASAP7_75t_L g1440 ( .A1(n_1426), .A2(n_1417), .B1(n_1419), .B2(n_1430), .C(n_1415), .Y(n_1440) );
AND2x2_ASAP7_75t_L g1441 ( .A(n_1419), .B(n_1422), .Y(n_1441) );
NAND4xp25_ASAP7_75t_L g1442 ( .A(n_1438), .B(n_1424), .C(n_1420), .D(n_1418), .Y(n_1442) );
NAND2xp5_ASAP7_75t_L g1443 ( .A(n_1416), .B(n_1421), .Y(n_1443) );
NAND2xp5_ASAP7_75t_SL g1444 ( .A(n_1423), .B(n_1412), .Y(n_1444) );
NAND2xp5_ASAP7_75t_L g1445 ( .A(n_1427), .B(n_1436), .Y(n_1445) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1429), .Y(n_1446) );
INVx1_ASAP7_75t_L g1447 ( .A(n_1425), .Y(n_1447) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1443), .Y(n_1448) );
AND3x2_ASAP7_75t_L g1449 ( .A(n_1441), .B(n_1155), .C(n_1413), .Y(n_1449) );
NAND4xp25_ASAP7_75t_L g1450 ( .A(n_1439), .B(n_1435), .C(n_1432), .D(n_1431), .Y(n_1450) );
NAND3xp33_ASAP7_75t_SL g1451 ( .A(n_1444), .B(n_1411), .C(n_1098), .Y(n_1451) );
NAND4xp25_ASAP7_75t_SL g1452 ( .A(n_1440), .B(n_1434), .C(n_1433), .D(n_1414), .Y(n_1452) );
NAND4xp25_ASAP7_75t_L g1453 ( .A(n_1442), .B(n_1205), .C(n_1132), .D(n_1179), .Y(n_1453) );
AND2x2_ASAP7_75t_L g1454 ( .A(n_1448), .B(n_1447), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1455 ( .A(n_1453), .B(n_1445), .Y(n_1455) );
OR4x2_ASAP7_75t_L g1456 ( .A(n_1451), .B(n_1437), .C(n_1446), .D(n_1187), .Y(n_1456) );
AOI21xp5_ASAP7_75t_L g1457 ( .A1(n_1452), .A2(n_1132), .B(n_1177), .Y(n_1457) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1454), .Y(n_1458) );
XNOR2xp5_ASAP7_75t_L g1459 ( .A(n_1455), .B(n_1450), .Y(n_1459) );
INVx4_ASAP7_75t_L g1460 ( .A(n_1456), .Y(n_1460) );
INVx1_ASAP7_75t_L g1461 ( .A(n_1458), .Y(n_1461) );
OAI22x1_ASAP7_75t_L g1462 ( .A1(n_1459), .A2(n_1449), .B1(n_1457), .B2(n_1085), .Y(n_1462) );
AO221x2_ASAP7_75t_L g1463 ( .A1(n_1461), .A2(n_1460), .B1(n_1180), .B2(n_1202), .C(n_1195), .Y(n_1463) );
AO221x1_ASAP7_75t_L g1464 ( .A1(n_1462), .A2(n_1143), .B1(n_1156), .B2(n_1082), .C(n_1089), .Y(n_1464) );
OAI21xp5_ASAP7_75t_L g1465 ( .A1(n_1464), .A2(n_1463), .B(n_1098), .Y(n_1465) );
AOI21xp5_ASAP7_75t_L g1466 ( .A1(n_1465), .A2(n_1142), .B(n_1238), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1466), .B(n_1142), .Y(n_1467) );
AOI22xp33_ASAP7_75t_SL g1468 ( .A1(n_1467), .A2(n_1121), .B1(n_1206), .B2(n_1208), .Y(n_1468) );
endmodule