module fake_jpeg_2299_n_100 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_100);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_100;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

INVxp67_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx6_ASAP7_75t_L g28 ( 
.A(n_17),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx2_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx24_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx10_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_28),
.B(n_26),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_40),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_27),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_42),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_42),
.A2(n_27),
.B1(n_33),
.B2(n_31),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_44),
.A2(n_50),
.B1(n_32),
.B2(n_30),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g45 ( 
.A1(n_39),
.A2(n_33),
.B1(n_34),
.B2(n_36),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_38),
.B1(n_41),
.B2(n_37),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_38),
.A2(n_36),
.B1(n_29),
.B2(n_30),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g60 ( 
.A(n_52),
.B(n_58),
.Y(n_60)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_43),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_0),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_55),
.B(n_2),
.Y(n_69)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_57),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g57 ( 
.A(n_49),
.B(n_32),
.Y(n_57)
);

AO22x2_ASAP7_75t_L g59 ( 
.A1(n_47),
.A2(n_19),
.B1(n_23),
.B2(n_22),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g61 ( 
.A(n_59),
.B(n_1),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_3),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_54),
.Y(n_62)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_59),
.B(n_1),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_64),
.B(n_59),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_58),
.A2(n_49),
.B1(n_47),
.B2(n_4),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_66),
.B(n_49),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_69),
.B(n_25),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_47),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_72),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_73),
.A2(n_74),
.B1(n_78),
.B2(n_79),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_47),
.B1(n_3),
.B2(n_4),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_63),
.B(n_2),
.Y(n_75)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g81 ( 
.A1(n_76),
.A2(n_61),
.B(n_68),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_65),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_77),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_67),
.B(n_12),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g88 ( 
.A1(n_81),
.A2(n_6),
.B(n_7),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_78),
.B(n_66),
.C(n_62),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_83),
.B(n_86),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_73),
.A2(n_71),
.B1(n_70),
.B2(n_8),
.Y(n_85)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_85),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_20),
.C(n_16),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_89),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_82),
.A2(n_6),
.B(n_7),
.Y(n_89)
);

OAI322xp33_ASAP7_75t_L g93 ( 
.A1(n_91),
.A2(n_87),
.A3(n_84),
.B1(n_83),
.B2(n_80),
.C1(n_86),
.C2(n_15),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_93),
.B(n_90),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_94),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_92),
.B1(n_9),
.B2(n_10),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_96),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g98 ( 
.A(n_97),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_8),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g100 ( 
.A(n_99),
.B(n_9),
.Y(n_100)
);


endmodule