module real_aes_8128_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_178;
wire n_409;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_725;
wire n_504;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_502;
wire n_434;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_713;
wire n_598;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_721;
wire n_446;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_719;
wire n_473;
wire n_465;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
A2O1A1Ixp33_ASAP7_75t_SL g174 ( .A1(n_0), .A2(n_175), .B(n_176), .C(n_180), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_1), .B(n_169), .Y(n_182) );
INVx1_ASAP7_75t_L g113 ( .A(n_2), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g153 ( .A(n_3), .B(n_154), .Y(n_153) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_4), .A2(n_163), .B(n_475), .Y(n_474) );
A2O1A1Ixp33_ASAP7_75t_L g518 ( .A1(n_5), .A2(n_143), .B(n_160), .C(n_519), .Y(n_518) );
AOI21xp5_ASAP7_75t_L g248 ( .A1(n_6), .A2(n_163), .B(n_249), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_7), .B(n_169), .Y(n_481) );
AO21x2_ASAP7_75t_L g256 ( .A1(n_8), .A2(n_135), .B(n_257), .Y(n_256) );
AND2x6_ASAP7_75t_L g160 ( .A(n_9), .B(n_161), .Y(n_160) );
A2O1A1Ixp33_ASAP7_75t_L g226 ( .A1(n_10), .A2(n_143), .B(n_160), .C(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g572 ( .A(n_11), .Y(n_572) );
NOR2xp33_ASAP7_75t_L g114 ( .A(n_12), .B(n_40), .Y(n_114) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_13), .B(n_179), .Y(n_521) );
INVx1_ASAP7_75t_L g140 ( .A(n_14), .Y(n_140) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_15), .B(n_154), .Y(n_263) );
A2O1A1Ixp33_ASAP7_75t_L g529 ( .A1(n_16), .A2(n_155), .B(n_530), .C(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_17), .B(n_169), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_18), .B(n_197), .Y(n_495) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_19), .A2(n_143), .B(n_189), .C(n_196), .Y(n_188) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_20), .A2(n_178), .B(n_231), .C(n_539), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_21), .B(n_441), .Y(n_440) );
NAND2xp5_ASAP7_75t_SL g503 ( .A(n_22), .B(n_179), .Y(n_503) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_23), .B(n_179), .Y(n_470) );
CKINVDCx16_ASAP7_75t_R g499 ( .A(n_24), .Y(n_499) );
INVx1_ASAP7_75t_L g469 ( .A(n_25), .Y(n_469) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_26), .A2(n_143), .B(n_196), .C(n_260), .Y(n_259) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_27), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g517 ( .A(n_28), .Y(n_517) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_29), .A2(n_104), .B1(n_115), .B2(n_727), .Y(n_103) );
INVx1_ASAP7_75t_L g493 ( .A(n_30), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g170 ( .A1(n_31), .A2(n_163), .B(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g145 ( .A(n_32), .Y(n_145) );
A2O1A1Ixp33_ASAP7_75t_L g211 ( .A1(n_33), .A2(n_158), .B(n_212), .C(n_213), .Y(n_211) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_34), .Y(n_523) );
A2O1A1Ixp33_ASAP7_75t_L g477 ( .A1(n_35), .A2(n_178), .B(n_478), .C(n_480), .Y(n_477) );
INVxp67_ASAP7_75t_L g494 ( .A(n_36), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_37), .B(n_262), .Y(n_261) );
CKINVDCx14_ASAP7_75t_R g476 ( .A(n_38), .Y(n_476) );
A2O1A1Ixp33_ASAP7_75t_L g467 ( .A1(n_39), .A2(n_143), .B(n_196), .C(n_468), .Y(n_467) );
A2O1A1Ixp33_ASAP7_75t_L g569 ( .A1(n_41), .A2(n_180), .B(n_570), .C(n_571), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g186 ( .A(n_42), .B(n_187), .Y(n_186) );
CKINVDCx20_ASAP7_75t_R g234 ( .A(n_43), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_44), .B(n_154), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_45), .B(n_163), .Y(n_258) );
CKINVDCx20_ASAP7_75t_R g472 ( .A(n_46), .Y(n_472) );
CKINVDCx20_ASAP7_75t_R g490 ( .A(n_47), .Y(n_490) );
A2O1A1Ixp33_ASAP7_75t_L g239 ( .A1(n_48), .A2(n_158), .B(n_212), .C(n_240), .Y(n_239) );
INVx1_ASAP7_75t_L g177 ( .A(n_49), .Y(n_177) );
AOI22xp33_ASAP7_75t_L g123 ( .A1(n_50), .A2(n_124), .B1(n_438), .B2(n_439), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_50), .Y(n_438) );
INVx1_ASAP7_75t_L g241 ( .A(n_51), .Y(n_241) );
INVx1_ASAP7_75t_L g537 ( .A(n_52), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_53), .B(n_163), .Y(n_238) );
OAI22xp5_ASAP7_75t_SL g125 ( .A1(n_54), .A2(n_72), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_54), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g201 ( .A(n_55), .Y(n_201) );
AOI222xp33_ASAP7_75t_SL g444 ( .A1(n_56), .A2(n_445), .B1(n_451), .B2(n_721), .C1(n_722), .C2(n_723), .Y(n_444) );
CKINVDCx14_ASAP7_75t_R g568 ( .A(n_57), .Y(n_568) );
INVx1_ASAP7_75t_L g161 ( .A(n_58), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_59), .B(n_163), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_60), .B(n_169), .Y(n_254) );
A2O1A1Ixp33_ASAP7_75t_L g251 ( .A1(n_61), .A2(n_150), .B(n_195), .C(n_252), .Y(n_251) );
OAI22xp5_ASAP7_75t_L g448 ( .A1(n_62), .A2(n_71), .B1(n_449), .B2(n_450), .Y(n_448) );
CKINVDCx20_ASAP7_75t_R g449 ( .A(n_62), .Y(n_449) );
INVx1_ASAP7_75t_L g139 ( .A(n_63), .Y(n_139) );
INVx1_ASAP7_75t_SL g479 ( .A(n_64), .Y(n_479) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_65), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_66), .B(n_154), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g541 ( .A(n_67), .B(n_169), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g228 ( .A(n_68), .B(n_155), .Y(n_228) );
INVx1_ASAP7_75t_L g502 ( .A(n_69), .Y(n_502) );
CKINVDCx16_ASAP7_75t_R g172 ( .A(n_70), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g450 ( .A(n_71), .Y(n_450) );
INVx1_ASAP7_75t_L g127 ( .A(n_72), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_73), .B(n_191), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g142 ( .A1(n_74), .A2(n_143), .B(n_148), .C(n_158), .Y(n_142) );
CKINVDCx16_ASAP7_75t_R g250 ( .A(n_75), .Y(n_250) );
INVx1_ASAP7_75t_L g108 ( .A(n_76), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g566 ( .A1(n_77), .A2(n_163), .B(n_567), .Y(n_566) );
CKINVDCx20_ASAP7_75t_R g506 ( .A(n_78), .Y(n_506) );
AOI21xp5_ASAP7_75t_L g526 ( .A1(n_79), .A2(n_163), .B(n_527), .Y(n_526) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_80), .A2(n_187), .B(n_489), .Y(n_488) );
CKINVDCx16_ASAP7_75t_R g466 ( .A(n_81), .Y(n_466) );
AOI22xp5_ASAP7_75t_L g445 ( .A1(n_82), .A2(n_446), .B1(n_447), .B2(n_448), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g446 ( .A(n_82), .Y(n_446) );
INVx1_ASAP7_75t_L g528 ( .A(n_83), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g192 ( .A(n_84), .B(n_193), .Y(n_192) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_85), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g535 ( .A1(n_86), .A2(n_163), .B(n_536), .Y(n_535) );
INVx1_ASAP7_75t_L g531 ( .A(n_87), .Y(n_531) );
INVx2_ASAP7_75t_L g137 ( .A(n_88), .Y(n_137) );
INVx1_ASAP7_75t_L g520 ( .A(n_89), .Y(n_520) );
CKINVDCx20_ASAP7_75t_R g167 ( .A(n_90), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g229 ( .A(n_91), .B(n_179), .Y(n_229) );
OR2x2_ASAP7_75t_L g110 ( .A(n_92), .B(n_111), .Y(n_110) );
OR2x2_ASAP7_75t_L g455 ( .A(n_92), .B(n_112), .Y(n_455) );
INVx2_ASAP7_75t_L g720 ( .A(n_92), .Y(n_720) );
A2O1A1Ixp33_ASAP7_75t_L g500 ( .A1(n_93), .A2(n_143), .B(n_158), .C(n_501), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_94), .B(n_163), .Y(n_210) );
INVx1_ASAP7_75t_L g214 ( .A(n_95), .Y(n_214) );
INVxp67_ASAP7_75t_L g253 ( .A(n_96), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_97), .B(n_135), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g107 ( .A(n_98), .B(n_108), .Y(n_107) );
INVx1_ASAP7_75t_L g149 ( .A(n_99), .Y(n_149) );
INVx1_ASAP7_75t_L g224 ( .A(n_100), .Y(n_224) );
INVx2_ASAP7_75t_L g540 ( .A(n_101), .Y(n_540) );
AND2x2_ASAP7_75t_L g243 ( .A(n_102), .B(n_199), .Y(n_243) );
CKINVDCx6p67_ASAP7_75t_R g104 ( .A(n_105), .Y(n_104) );
INVx1_ASAP7_75t_L g728 ( .A(n_105), .Y(n_728) );
NAND2xp5_ASAP7_75t_L g105 ( .A(n_106), .B(n_109), .Y(n_105) );
INVx1_ASAP7_75t_SL g106 ( .A(n_107), .Y(n_106) );
INVx1_ASAP7_75t_SL g109 ( .A(n_110), .Y(n_109) );
INVx2_ASAP7_75t_L g122 ( .A(n_110), .Y(n_122) );
HB1xp67_ASAP7_75t_L g442 ( .A(n_110), .Y(n_442) );
NOR2x2_ASAP7_75t_L g721 ( .A(n_111), .B(n_720), .Y(n_721) );
INVx2_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
OR2x2_ASAP7_75t_L g719 ( .A(n_112), .B(n_720), .Y(n_719) );
AND2x2_ASAP7_75t_L g112 ( .A(n_113), .B(n_114), .Y(n_112) );
OA21x2_ASAP7_75t_L g115 ( .A1(n_116), .A2(n_121), .B(n_443), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_117), .Y(n_116) );
NAND3xp33_ASAP7_75t_L g443 ( .A(n_117), .B(n_440), .C(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_118), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OAI21xp5_ASAP7_75t_L g121 ( .A1(n_122), .A2(n_123), .B(n_440), .Y(n_121) );
INVx1_ASAP7_75t_L g439 ( .A(n_124), .Y(n_439) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_125), .B(n_128), .Y(n_124) );
INVx1_ASAP7_75t_L g452 ( .A(n_128), .Y(n_452) );
OAI22xp5_ASAP7_75t_L g723 ( .A1(n_128), .A2(n_457), .B1(n_724), .B2(n_725), .Y(n_723) );
OR3x1_ASAP7_75t_L g128 ( .A(n_129), .B(n_346), .C(n_395), .Y(n_128) );
NAND5xp2_ASAP7_75t_L g129 ( .A(n_130), .B(n_280), .C(n_309), .D(n_317), .E(n_332), .Y(n_129) );
O2A1O1Ixp33_ASAP7_75t_L g130 ( .A1(n_131), .A2(n_203), .B(n_219), .C(n_264), .Y(n_130) );
NOR2xp33_ASAP7_75t_L g131 ( .A(n_132), .B(n_183), .Y(n_131) );
AND2x2_ASAP7_75t_L g275 ( .A(n_132), .B(n_272), .Y(n_275) );
AND2x2_ASAP7_75t_L g308 ( .A(n_132), .B(n_184), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_132), .B(n_207), .Y(n_401) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_168), .Y(n_132) );
INVx2_ASAP7_75t_L g206 ( .A(n_133), .Y(n_206) );
BUFx2_ASAP7_75t_L g375 ( .A(n_133), .Y(n_375) );
AO21x2_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_141), .B(n_166), .Y(n_133) );
NOR2xp33_ASAP7_75t_L g166 ( .A(n_134), .B(n_167), .Y(n_166) );
INVx3_ASAP7_75t_L g169 ( .A(n_134), .Y(n_169) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_134), .B(n_218), .Y(n_217) );
AO21x2_ASAP7_75t_L g222 ( .A1(n_134), .A2(n_223), .B(n_233), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g471 ( .A(n_134), .B(n_472), .Y(n_471) );
AO21x2_ASAP7_75t_L g497 ( .A1(n_134), .A2(n_498), .B(n_505), .Y(n_497) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_134), .B(n_523), .Y(n_522) );
INVx4_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
HB1xp67_ASAP7_75t_L g247 ( .A(n_135), .Y(n_247) );
AOI21xp5_ASAP7_75t_L g257 ( .A1(n_135), .A2(n_258), .B(n_259), .Y(n_257) );
BUFx6f_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g235 ( .A(n_136), .Y(n_235) );
AND2x2_ASAP7_75t_L g136 ( .A(n_137), .B(n_138), .Y(n_136) );
AND2x2_ASAP7_75t_SL g199 ( .A(n_137), .B(n_138), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_139), .B(n_140), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_142), .B(n_162), .Y(n_141) );
INVx5_ASAP7_75t_L g173 ( .A(n_143), .Y(n_173) );
AND2x6_ASAP7_75t_L g143 ( .A(n_144), .B(n_146), .Y(n_143) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_144), .Y(n_157) );
BUFx3_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
INVx2_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
INVx1_ASAP7_75t_L g165 ( .A(n_145), .Y(n_165) );
INVx1_ASAP7_75t_L g232 ( .A(n_145), .Y(n_232) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_147), .Y(n_152) );
INVx3_ASAP7_75t_L g155 ( .A(n_147), .Y(n_155) );
AND2x2_ASAP7_75t_L g164 ( .A(n_147), .B(n_165), .Y(n_164) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_147), .Y(n_179) );
INVx1_ASAP7_75t_L g262 ( .A(n_147), .Y(n_262) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_153), .C(n_156), .Y(n_148) );
INVx1_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
OAI22xp33_ASAP7_75t_L g492 ( .A1(n_151), .A2(n_154), .B1(n_493), .B2(n_494), .Y(n_492) );
NOR2xp33_ASAP7_75t_L g530 ( .A(n_151), .B(n_531), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g539 ( .A(n_151), .B(n_540), .Y(n_539) );
INVx4_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g191 ( .A(n_152), .Y(n_191) );
INVx2_ASAP7_75t_L g175 ( .A(n_154), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g252 ( .A(n_154), .B(n_253), .Y(n_252) );
O2A1O1Ixp33_ASAP7_75t_L g468 ( .A1(n_154), .A2(n_194), .B(n_469), .C(n_470), .Y(n_468) );
INVx5_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_155), .B(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx3_ASAP7_75t_L g480 ( .A(n_157), .Y(n_480) );
INVx1_ASAP7_75t_L g158 ( .A(n_159), .Y(n_158) );
O2A1O1Ixp33_ASAP7_75t_SL g171 ( .A1(n_159), .A2(n_172), .B(n_173), .C(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_L g249 ( .A1(n_159), .A2(n_173), .B(n_250), .C(n_251), .Y(n_249) );
O2A1O1Ixp33_ASAP7_75t_L g475 ( .A1(n_159), .A2(n_173), .B(n_476), .C(n_477), .Y(n_475) );
O2A1O1Ixp33_ASAP7_75t_SL g489 ( .A1(n_159), .A2(n_173), .B(n_490), .C(n_491), .Y(n_489) );
O2A1O1Ixp33_ASAP7_75t_SL g527 ( .A1(n_159), .A2(n_173), .B(n_528), .C(n_529), .Y(n_527) );
O2A1O1Ixp33_ASAP7_75t_SL g536 ( .A1(n_159), .A2(n_173), .B(n_537), .C(n_538), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g567 ( .A1(n_159), .A2(n_173), .B(n_568), .C(n_569), .Y(n_567) );
INVx4_ASAP7_75t_SL g159 ( .A(n_160), .Y(n_159) );
AND2x4_ASAP7_75t_L g163 ( .A(n_160), .B(n_164), .Y(n_163) );
BUFx3_ASAP7_75t_L g196 ( .A(n_160), .Y(n_196) );
NAND2x1p5_ASAP7_75t_L g225 ( .A(n_160), .B(n_164), .Y(n_225) );
BUFx2_ASAP7_75t_L g187 ( .A(n_163), .Y(n_187) );
INVx1_ASAP7_75t_L g195 ( .A(n_165), .Y(n_195) );
AND2x2_ASAP7_75t_L g183 ( .A(n_168), .B(n_184), .Y(n_183) );
INVx2_ASAP7_75t_L g273 ( .A(n_168), .Y(n_273) );
AND2x2_ASAP7_75t_L g359 ( .A(n_168), .B(n_272), .Y(n_359) );
AND2x2_ASAP7_75t_L g414 ( .A(n_168), .B(n_206), .Y(n_414) );
OA21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_170), .B(n_182), .Y(n_168) );
INVx2_ASAP7_75t_L g212 ( .A(n_173), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_177), .B(n_178), .Y(n_176) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_178), .B(n_479), .Y(n_478) );
INVx4_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx2_ASAP7_75t_L g570 ( .A(n_179), .Y(n_570) );
INVx2_ASAP7_75t_L g504 ( .A(n_180), .Y(n_504) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
HB1xp67_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
INVx1_ASAP7_75t_L g532 ( .A(n_181), .Y(n_532) );
INVx1_ASAP7_75t_L g331 ( .A(n_183), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_183), .B(n_207), .Y(n_378) );
INVx5_ASAP7_75t_L g272 ( .A(n_184), .Y(n_272) );
AND2x4_ASAP7_75t_L g293 ( .A(n_184), .B(n_273), .Y(n_293) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_184), .Y(n_315) );
AND2x2_ASAP7_75t_L g390 ( .A(n_184), .B(n_375), .Y(n_390) );
AND2x2_ASAP7_75t_L g393 ( .A(n_184), .B(n_208), .Y(n_393) );
OR2x6_ASAP7_75t_L g184 ( .A(n_185), .B(n_200), .Y(n_184) );
AOI21xp5_ASAP7_75t_SL g185 ( .A1(n_186), .A2(n_188), .B(n_197), .Y(n_185) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_190), .A2(n_192), .B(n_194), .Y(n_189) );
INVx2_ASAP7_75t_L g193 ( .A(n_191), .Y(n_193) );
O2A1O1Ixp33_ASAP7_75t_L g213 ( .A1(n_193), .A2(n_214), .B(n_215), .C(n_216), .Y(n_213) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_193), .A2(n_216), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_193), .A2(n_502), .B(n_503), .C(n_504), .Y(n_501) );
O2A1O1Ixp5_ASAP7_75t_L g519 ( .A1(n_193), .A2(n_504), .B(n_520), .C(n_521), .Y(n_519) );
INVx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g491 ( .A(n_195), .B(n_492), .Y(n_491) );
INVx1_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
NOR2xp33_ASAP7_75t_L g505 ( .A(n_198), .B(n_506), .Y(n_505) );
INVx2_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
INVx1_ASAP7_75t_L g202 ( .A(n_199), .Y(n_202) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_199), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g237 ( .A1(n_199), .A2(n_238), .B(n_239), .Y(n_237) );
O2A1O1Ixp33_ASAP7_75t_L g465 ( .A1(n_199), .A2(n_225), .B(n_466), .C(n_467), .Y(n_465) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_199), .A2(n_566), .B(n_573), .Y(n_565) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_201), .B(n_202), .Y(n_200) );
AO21x2_ASAP7_75t_L g515 ( .A1(n_202), .A2(n_516), .B(n_522), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_203), .B(n_273), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_203), .B(n_404), .Y(n_403) );
INVx2_ASAP7_75t_SL g203 ( .A(n_204), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_205), .B(n_207), .Y(n_204) );
AND2x2_ASAP7_75t_L g298 ( .A(n_205), .B(n_273), .Y(n_298) );
AND2x2_ASAP7_75t_L g316 ( .A(n_205), .B(n_208), .Y(n_316) );
INVx1_ASAP7_75t_L g336 ( .A(n_205), .Y(n_336) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_205), .B(n_272), .Y(n_381) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_205), .Y(n_423) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g292 ( .A(n_206), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_207), .B(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g325 ( .A(n_207), .Y(n_325) );
O2A1O1Ixp33_ASAP7_75t_L g328 ( .A1(n_207), .A2(n_268), .B(n_329), .C(n_331), .Y(n_328) );
AND2x2_ASAP7_75t_L g335 ( .A(n_207), .B(n_336), .Y(n_335) );
OR2x2_ASAP7_75t_L g344 ( .A(n_207), .B(n_345), .Y(n_344) );
AND2x2_ASAP7_75t_L g348 ( .A(n_207), .B(n_272), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_207), .B(n_359), .Y(n_358) );
AND2x2_ASAP7_75t_L g363 ( .A(n_207), .B(n_273), .Y(n_363) );
AND2x2_ASAP7_75t_L g413 ( .A(n_207), .B(n_414), .Y(n_413) );
INVx5_ASAP7_75t_L g207 ( .A(n_208), .Y(n_207) );
BUFx2_ASAP7_75t_L g277 ( .A(n_208), .Y(n_277) );
AND2x2_ASAP7_75t_L g318 ( .A(n_208), .B(n_271), .Y(n_318) );
AND2x2_ASAP7_75t_L g330 ( .A(n_208), .B(n_305), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_208), .B(n_359), .Y(n_377) );
OR2x6_ASAP7_75t_L g208 ( .A(n_209), .B(n_217), .Y(n_208) );
AND2x2_ASAP7_75t_L g219 ( .A(n_220), .B(n_244), .Y(n_219) );
INVx1_ASAP7_75t_L g266 ( .A(n_220), .Y(n_266) );
AND2x2_ASAP7_75t_L g220 ( .A(n_221), .B(n_236), .Y(n_220) );
OR2x2_ASAP7_75t_L g268 ( .A(n_221), .B(n_236), .Y(n_268) );
NAND3xp33_ASAP7_75t_L g274 ( .A(n_221), .B(n_275), .C(n_276), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_221), .B(n_246), .Y(n_285) );
OR2x2_ASAP7_75t_L g300 ( .A(n_221), .B(n_288), .Y(n_300) );
AND2x2_ASAP7_75t_L g306 ( .A(n_221), .B(n_255), .Y(n_306) );
NOR2xp33_ASAP7_75t_L g436 ( .A(n_221), .B(n_437), .Y(n_436) );
INVx5_ASAP7_75t_SL g221 ( .A(n_222), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_222), .B(n_246), .Y(n_303) );
AND2x2_ASAP7_75t_L g342 ( .A(n_222), .B(n_256), .Y(n_342) );
NAND2xp5_ASAP7_75t_SL g370 ( .A(n_222), .B(n_255), .Y(n_370) );
OR2x2_ASAP7_75t_L g373 ( .A(n_222), .B(n_255), .Y(n_373) );
OAI21xp5_ASAP7_75t_L g223 ( .A1(n_224), .A2(n_225), .B(n_226), .Y(n_223) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_225), .A2(n_499), .B(n_500), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g516 ( .A1(n_225), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g227 ( .A1(n_228), .A2(n_229), .B(n_230), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g260 ( .A1(n_230), .A2(n_261), .B(n_263), .Y(n_260) );
INVx2_ASAP7_75t_L g230 ( .A(n_231), .Y(n_230) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g233 ( .A(n_234), .B(n_235), .Y(n_233) );
INVx2_ASAP7_75t_L g487 ( .A(n_235), .Y(n_487) );
INVx5_ASAP7_75t_SL g288 ( .A(n_236), .Y(n_288) );
OR2x2_ASAP7_75t_L g294 ( .A(n_236), .B(n_245), .Y(n_294) );
AND2x2_ASAP7_75t_L g310 ( .A(n_236), .B(n_311), .Y(n_310) );
AOI321xp33_ASAP7_75t_L g317 ( .A1(n_236), .A2(n_318), .A3(n_319), .B1(n_320), .B2(n_326), .C(n_328), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_236), .B(n_244), .Y(n_327) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_236), .Y(n_340) );
OR2x2_ASAP7_75t_L g387 ( .A(n_236), .B(n_285), .Y(n_387) );
AND2x2_ASAP7_75t_L g409 ( .A(n_236), .B(n_306), .Y(n_409) );
AND2x2_ASAP7_75t_L g428 ( .A(n_236), .B(n_246), .Y(n_428) );
OR2x6_ASAP7_75t_L g236 ( .A(n_237), .B(n_243), .Y(n_236) );
INVx1_ASAP7_75t_SL g244 ( .A(n_245), .Y(n_244) );
OR2x2_ASAP7_75t_L g245 ( .A(n_246), .B(n_255), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_246), .B(n_255), .Y(n_269) );
AND2x2_ASAP7_75t_L g278 ( .A(n_246), .B(n_279), .Y(n_278) );
INVx3_ASAP7_75t_L g305 ( .A(n_246), .Y(n_305) );
AND2x2_ASAP7_75t_L g311 ( .A(n_246), .B(n_306), .Y(n_311) );
INVxp67_ASAP7_75t_L g341 ( .A(n_246), .Y(n_341) );
OR2x2_ASAP7_75t_L g383 ( .A(n_246), .B(n_288), .Y(n_383) );
OA21x2_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_248), .B(n_254), .Y(n_246) );
OA21x2_ASAP7_75t_L g473 ( .A1(n_247), .A2(n_474), .B(n_481), .Y(n_473) );
OA21x2_ASAP7_75t_L g525 ( .A1(n_247), .A2(n_526), .B(n_533), .Y(n_525) );
OA21x2_ASAP7_75t_L g534 ( .A1(n_247), .A2(n_535), .B(n_541), .Y(n_534) );
OR2x2_ASAP7_75t_L g265 ( .A(n_255), .B(n_266), .Y(n_265) );
INVx1_ASAP7_75t_SL g279 ( .A(n_255), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_255), .B(n_268), .Y(n_312) );
AND2x2_ASAP7_75t_L g361 ( .A(n_255), .B(n_305), .Y(n_361) );
AND2x2_ASAP7_75t_L g399 ( .A(n_255), .B(n_288), .Y(n_399) );
INVx2_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_256), .B(n_288), .Y(n_287) );
A2O1A1Ixp33_ASAP7_75t_L g264 ( .A1(n_265), .A2(n_267), .B(n_270), .C(n_274), .Y(n_264) );
OAI22xp5_ASAP7_75t_L g391 ( .A1(n_265), .A2(n_267), .B1(n_392), .B2(n_394), .Y(n_391) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_267), .A2(n_290), .B1(n_345), .B2(n_431), .Y(n_430) );
OR2x2_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
INVx1_ASAP7_75t_SL g419 ( .A(n_268), .Y(n_419) );
INVx1_ASAP7_75t_SL g319 ( .A(n_269), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_271), .B(n_291), .Y(n_321) );
AOI222xp33_ASAP7_75t_L g332 ( .A1(n_271), .A2(n_312), .B1(n_319), .B2(n_333), .C1(n_337), .C2(n_343), .Y(n_332) );
AND2x2_ASAP7_75t_L g422 ( .A(n_271), .B(n_423), .Y(n_422) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_273), .Y(n_271) );
INVx2_ASAP7_75t_L g297 ( .A(n_272), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g367 ( .A(n_272), .B(n_292), .Y(n_367) );
HB1xp67_ASAP7_75t_L g404 ( .A(n_272), .Y(n_404) );
AND2x2_ASAP7_75t_L g407 ( .A(n_272), .B(n_316), .Y(n_407) );
NOR2xp33_ASAP7_75t_L g433 ( .A(n_272), .B(n_423), .Y(n_433) );
INVx1_ASAP7_75t_L g324 ( .A(n_273), .Y(n_324) );
HB1xp67_ASAP7_75t_L g352 ( .A(n_273), .Y(n_352) );
O2A1O1Ixp33_ASAP7_75t_L g415 ( .A1(n_275), .A2(n_416), .B(n_417), .C(n_420), .Y(n_415) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_278), .Y(n_276) );
NAND3xp33_ASAP7_75t_L g338 ( .A(n_277), .B(n_339), .C(n_342), .Y(n_338) );
OR2x2_ASAP7_75t_L g366 ( .A(n_277), .B(n_367), .Y(n_366) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_277), .B(n_293), .Y(n_394) );
OR2x2_ASAP7_75t_L g299 ( .A(n_279), .B(n_300), .Y(n_299) );
AOI211xp5_ASAP7_75t_L g280 ( .A1(n_281), .A2(n_283), .B(n_289), .C(n_301), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g410 ( .A(n_282), .B(n_411), .Y(n_410) );
AND2x2_ASAP7_75t_L g388 ( .A(n_283), .B(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_286), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g398 ( .A(n_284), .B(n_399), .Y(n_398) );
INVx1_ASAP7_75t_SL g284 ( .A(n_285), .Y(n_284) );
INVx1_ASAP7_75t_SL g286 ( .A(n_287), .Y(n_286) );
OR2x2_ASAP7_75t_L g302 ( .A(n_287), .B(n_303), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_288), .B(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g356 ( .A(n_288), .B(n_306), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_288), .B(n_361), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_288), .B(n_305), .Y(n_371) );
OAI22xp5_ASAP7_75t_L g289 ( .A1(n_290), .A2(n_294), .B1(n_295), .B2(n_299), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_293), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_291), .B(n_363), .Y(n_362) );
BUFx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_293), .B(n_335), .Y(n_334) );
OAI221xp5_ASAP7_75t_SL g357 ( .A1(n_294), .A2(n_358), .B1(n_360), .B2(n_362), .C(n_364), .Y(n_357) );
INVx1_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_297), .B(n_298), .Y(n_296) );
AND2x2_ASAP7_75t_L g412 ( .A(n_297), .B(n_413), .Y(n_412) );
AND2x2_ASAP7_75t_L g425 ( .A(n_297), .B(n_414), .Y(n_425) );
INVx1_ASAP7_75t_L g345 ( .A(n_298), .Y(n_345) );
INVx1_ASAP7_75t_L g416 ( .A(n_299), .Y(n_416) );
AOI21xp5_ASAP7_75t_L g405 ( .A1(n_300), .A2(n_383), .B(n_406), .Y(n_405) );
AOI21xp33_ASAP7_75t_L g301 ( .A1(n_302), .A2(n_304), .B(n_307), .Y(n_301) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
OAI21xp5_ASAP7_75t_SL g309 ( .A1(n_310), .A2(n_312), .B(n_313), .Y(n_309) );
INVx1_ASAP7_75t_L g349 ( .A(n_310), .Y(n_349) );
AOI221xp5_ASAP7_75t_L g396 ( .A1(n_311), .A2(n_397), .B1(n_400), .B2(n_402), .C(n_405), .Y(n_396) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_315), .B(n_316), .Y(n_314) );
AOI22xp5_ASAP7_75t_L g408 ( .A1(n_319), .A2(n_409), .B1(n_410), .B2(n_412), .Y(n_408) );
NAND2xp5_ASAP7_75t_SL g320 ( .A(n_321), .B(n_322), .Y(n_320) );
INVx1_ASAP7_75t_L g385 ( .A(n_321), .Y(n_385) );
INVx1_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2xp67_ASAP7_75t_SL g323 ( .A(n_324), .B(n_325), .Y(n_323) );
AND2x2_ASAP7_75t_L g389 ( .A(n_325), .B(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g354 ( .A(n_330), .Y(n_354) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_335), .B(n_359), .Y(n_411) );
INVxp67_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g339 ( .A(n_340), .B(n_341), .Y(n_339) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_341), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g427 ( .A(n_342), .B(n_428), .Y(n_427) );
AND2x4_ASAP7_75t_L g434 ( .A(n_342), .B(n_435), .Y(n_434) );
INVx1_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
OAI211xp5_ASAP7_75t_SL g346 ( .A1(n_347), .A2(n_349), .B(n_350), .C(n_384), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
AOI211xp5_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_353), .B(n_357), .C(n_376), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx1_ASAP7_75t_SL g437 ( .A(n_361), .Y(n_437) );
AND2x2_ASAP7_75t_L g374 ( .A(n_363), .B(n_375), .Y(n_374) );
AOI22xp5_ASAP7_75t_L g364 ( .A1(n_365), .A2(n_368), .B1(n_372), .B2(n_374), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
OR2x2_ASAP7_75t_L g369 ( .A(n_370), .B(n_371), .Y(n_369) );
OR2x2_ASAP7_75t_L g382 ( .A(n_370), .B(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g435 ( .A(n_371), .Y(n_435) );
INVxp67_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
AOI31xp33_ASAP7_75t_L g376 ( .A1(n_377), .A2(n_378), .A3(n_379), .B(n_382), .Y(n_376) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
AOI211xp5_ASAP7_75t_L g384 ( .A1(n_385), .A2(n_386), .B(n_388), .C(n_391), .Y(n_384) );
INVx1_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
CKINVDCx16_ASAP7_75t_R g392 ( .A(n_393), .Y(n_392) );
NAND5xp2_ASAP7_75t_L g395 ( .A(n_396), .B(n_408), .C(n_415), .D(n_429), .E(n_432), .Y(n_395) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_407), .A2(n_433), .B1(n_434), .B2(n_436), .Y(n_432) );
INVx1_ASAP7_75t_SL g431 ( .A(n_409), .Y(n_431) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AOI21xp33_ASAP7_75t_L g420 ( .A1(n_421), .A2(n_424), .B(n_426), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVxp67_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx1_ASAP7_75t_SL g441 ( .A(n_442), .Y(n_441) );
CKINVDCx16_ASAP7_75t_R g722 ( .A(n_445), .Y(n_722) );
INVx1_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
OAI22xp5_ASAP7_75t_SL g451 ( .A1(n_452), .A2(n_453), .B1(n_456), .B2(n_719), .Y(n_451) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g724 ( .A(n_454), .Y(n_724) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR3x1_ASAP7_75t_L g457 ( .A(n_458), .B(n_630), .C(n_677), .Y(n_457) );
NAND3xp33_ASAP7_75t_SL g458 ( .A(n_459), .B(n_576), .C(n_601), .Y(n_458) );
AOI221xp5_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_514), .B1(n_542), .B2(n_545), .C(n_553), .Y(n_459) );
OAI21xp5_ASAP7_75t_L g460 ( .A1(n_461), .A2(n_482), .B(n_507), .Y(n_460) );
INVx1_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_462), .B(n_555), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_462), .B(n_558), .Y(n_674) );
AND2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_473), .Y(n_462) );
AND2x2_ASAP7_75t_L g544 ( .A(n_463), .B(n_513), .Y(n_544) );
AND2x2_ASAP7_75t_L g594 ( .A(n_463), .B(n_512), .Y(n_594) );
AND2x2_ASAP7_75t_L g615 ( .A(n_463), .B(n_616), .Y(n_615) );
AND2x2_ASAP7_75t_L g620 ( .A(n_463), .B(n_587), .Y(n_620) );
OR2x2_ASAP7_75t_L g628 ( .A(n_463), .B(n_629), .Y(n_628) );
AND2x2_ASAP7_75t_L g700 ( .A(n_463), .B(n_496), .Y(n_700) );
NAND2xp5_ASAP7_75t_L g714 ( .A(n_463), .B(n_649), .Y(n_714) );
INVx3_ASAP7_75t_SL g463 ( .A(n_464), .Y(n_463) );
AND2x2_ASAP7_75t_L g559 ( .A(n_464), .B(n_473), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_464), .B(n_496), .Y(n_560) );
AND2x4_ASAP7_75t_L g582 ( .A(n_464), .B(n_513), .Y(n_582) );
AND2x2_ASAP7_75t_L g612 ( .A(n_464), .B(n_484), .Y(n_612) );
AND2x2_ASAP7_75t_L g621 ( .A(n_464), .B(n_611), .Y(n_621) );
AND2x2_ASAP7_75t_L g637 ( .A(n_464), .B(n_497), .Y(n_637) );
OR2x2_ASAP7_75t_L g646 ( .A(n_464), .B(n_629), .Y(n_646) );
AND2x2_ASAP7_75t_L g652 ( .A(n_464), .B(n_587), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_464), .B(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g666 ( .A(n_464), .B(n_509), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_464), .B(n_555), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g705 ( .A(n_464), .B(n_616), .Y(n_705) );
OR2x6_ASAP7_75t_L g464 ( .A(n_465), .B(n_471), .Y(n_464) );
INVx2_ASAP7_75t_L g513 ( .A(n_473), .Y(n_513) );
AND2x2_ASAP7_75t_L g611 ( .A(n_473), .B(n_496), .Y(n_611) );
AND2x2_ASAP7_75t_L g616 ( .A(n_473), .B(n_497), .Y(n_616) );
INVx1_ASAP7_75t_L g672 ( .A(n_473), .Y(n_672) );
INVx1_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
AND2x2_ASAP7_75t_L g581 ( .A(n_483), .B(n_582), .Y(n_581) );
AND2x2_ASAP7_75t_L g483 ( .A(n_484), .B(n_496), .Y(n_483) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_484), .B(n_544), .Y(n_543) );
BUFx3_ASAP7_75t_L g558 ( .A(n_484), .Y(n_558) );
OR2x2_ASAP7_75t_L g629 ( .A(n_484), .B(n_496), .Y(n_629) );
OR2x2_ASAP7_75t_L g690 ( .A(n_484), .B(n_597), .Y(n_690) );
OA21x2_ASAP7_75t_L g484 ( .A1(n_485), .A2(n_488), .B(n_495), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AO21x2_ASAP7_75t_L g509 ( .A1(n_486), .A2(n_510), .B(n_511), .Y(n_509) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx1_ASAP7_75t_L g510 ( .A(n_488), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_495), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_496), .B(n_513), .Y(n_512) );
AND2x2_ASAP7_75t_L g649 ( .A(n_496), .B(n_509), .Y(n_649) );
INVx2_ASAP7_75t_SL g496 ( .A(n_497), .Y(n_496) );
BUFx2_ASAP7_75t_L g588 ( .A(n_497), .Y(n_588) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AOI221xp5_ASAP7_75t_L g693 ( .A1(n_508), .A2(n_694), .B1(n_698), .B2(n_701), .C(n_702), .Y(n_693) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_512), .Y(n_508) );
INVx1_ASAP7_75t_SL g556 ( .A(n_509), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_509), .B(n_672), .Y(n_671) );
AND2x2_ASAP7_75t_L g688 ( .A(n_509), .B(n_544), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g680 ( .A(n_512), .B(n_558), .Y(n_680) );
AND2x2_ASAP7_75t_L g587 ( .A(n_513), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_SL g591 ( .A(n_514), .Y(n_591) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_514), .B(n_597), .Y(n_627) );
AND2x2_ASAP7_75t_L g514 ( .A(n_515), .B(n_524), .Y(n_514) );
AND2x2_ASAP7_75t_L g552 ( .A(n_515), .B(n_525), .Y(n_552) );
INVx4_ASAP7_75t_L g564 ( .A(n_515), .Y(n_564) );
BUFx3_ASAP7_75t_L g607 ( .A(n_515), .Y(n_607) );
AND3x2_ASAP7_75t_L g622 ( .A(n_515), .B(n_623), .C(n_624), .Y(n_622) );
AND2x2_ASAP7_75t_L g704 ( .A(n_524), .B(n_618), .Y(n_704) );
AND2x2_ASAP7_75t_L g712 ( .A(n_524), .B(n_597), .Y(n_712) );
INVx1_ASAP7_75t_SL g717 ( .A(n_524), .Y(n_717) );
AND2x2_ASAP7_75t_L g524 ( .A(n_525), .B(n_534), .Y(n_524) );
INVx1_ASAP7_75t_SL g575 ( .A(n_525), .Y(n_575) );
AND2x2_ASAP7_75t_L g598 ( .A(n_525), .B(n_564), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g600 ( .A(n_525), .B(n_548), .Y(n_600) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_525), .Y(n_640) );
OR2x2_ASAP7_75t_L g645 ( .A(n_525), .B(n_564), .Y(n_645) );
INVx2_ASAP7_75t_L g550 ( .A(n_534), .Y(n_550) );
AND2x2_ASAP7_75t_L g585 ( .A(n_534), .B(n_565), .Y(n_585) );
OR2x2_ASAP7_75t_L g605 ( .A(n_534), .B(n_565), .Y(n_605) );
HB1xp67_ASAP7_75t_L g625 ( .A(n_534), .Y(n_625) );
INVx1_ASAP7_75t_SL g542 ( .A(n_543), .Y(n_542) );
AOI21xp33_ASAP7_75t_L g675 ( .A1(n_543), .A2(n_584), .B(n_676), .Y(n_675) );
AOI322xp5_ASAP7_75t_L g711 ( .A1(n_545), .A2(n_555), .A3(n_582), .B1(n_712), .B2(n_713), .C1(n_715), .C2(n_718), .Y(n_711) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
OR2x2_ASAP7_75t_L g546 ( .A(n_547), .B(n_551), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g654 ( .A(n_547), .B(n_655), .Y(n_654) );
INVx1_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_548), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
AND2x2_ASAP7_75t_L g574 ( .A(n_549), .B(n_575), .Y(n_574) );
INVx2_ASAP7_75t_L g549 ( .A(n_550), .Y(n_549) );
AND2x2_ASAP7_75t_L g642 ( .A(n_550), .B(n_564), .Y(n_642) );
AND2x2_ASAP7_75t_L g709 ( .A(n_550), .B(n_565), .Y(n_709) );
INVx1_ASAP7_75t_SL g551 ( .A(n_552), .Y(n_551) );
AND2x2_ASAP7_75t_L g650 ( .A(n_552), .B(n_604), .Y(n_650) );
AOI31xp33_ASAP7_75t_L g553 ( .A1(n_554), .A2(n_557), .A3(n_560), .B(n_561), .Y(n_553) );
AND2x2_ASAP7_75t_L g609 ( .A(n_555), .B(n_587), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_555), .B(n_579), .Y(n_691) );
AND2x2_ASAP7_75t_L g710 ( .A(n_555), .B(n_615), .Y(n_710) );
INVx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_558), .B(n_587), .Y(n_599) );
NAND2x1p5_ASAP7_75t_L g633 ( .A(n_558), .B(n_616), .Y(n_633) );
NAND2xp5_ASAP7_75t_SL g636 ( .A(n_558), .B(n_637), .Y(n_636) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_558), .B(n_700), .Y(n_699) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_559), .B(n_616), .Y(n_648) );
INVx1_ASAP7_75t_L g692 ( .A(n_559), .Y(n_692) );
INVx1_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_574), .Y(n_562) );
INVxp67_ASAP7_75t_L g644 ( .A(n_563), .Y(n_644) );
NOR2xp33_ASAP7_75t_L g563 ( .A(n_564), .B(n_565), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_564), .B(n_575), .Y(n_580) );
INVx1_ASAP7_75t_L g686 ( .A(n_564), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g697 ( .A(n_564), .B(n_663), .Y(n_697) );
BUFx3_ASAP7_75t_L g597 ( .A(n_565), .Y(n_597) );
AND2x2_ASAP7_75t_L g623 ( .A(n_565), .B(n_575), .Y(n_623) );
INVx2_ASAP7_75t_L g663 ( .A(n_565), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g695 ( .A(n_574), .B(n_696), .Y(n_695) );
AOI211xp5_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .B(n_583), .C(n_592), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
AOI21xp33_ASAP7_75t_L g626 ( .A1(n_578), .A2(n_627), .B(n_628), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_579), .B(n_585), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g617 ( .A(n_579), .B(n_618), .Y(n_617) );
INVx1_ASAP7_75t_L g579 ( .A(n_580), .Y(n_579) );
OR2x2_ASAP7_75t_L g659 ( .A(n_580), .B(n_605), .Y(n_659) );
INVx3_ASAP7_75t_L g590 ( .A(n_582), .Y(n_590) );
OAI22xp5_ASAP7_75t_SL g583 ( .A1(n_584), .A2(n_586), .B1(n_589), .B2(n_591), .Y(n_583) );
OAI21xp5_ASAP7_75t_SL g608 ( .A1(n_585), .A2(n_609), .B(n_610), .Y(n_608) );
AND2x2_ASAP7_75t_L g634 ( .A(n_585), .B(n_598), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_585), .B(n_686), .Y(n_685) );
INVxp67_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
OR2x2_ASAP7_75t_L g589 ( .A(n_588), .B(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g658 ( .A(n_588), .Y(n_658) );
OAI21xp5_ASAP7_75t_SL g602 ( .A1(n_589), .A2(n_603), .B(n_608), .Y(n_602) );
OAI22xp33_ASAP7_75t_SL g592 ( .A1(n_593), .A2(n_595), .B1(n_599), .B2(n_600), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
NOR2xp33_ASAP7_75t_L g669 ( .A(n_594), .B(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
AND2x2_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
INVx1_ASAP7_75t_L g618 ( .A(n_597), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_597), .B(n_640), .Y(n_639) );
NOR3xp33_ASAP7_75t_L g601 ( .A(n_602), .B(n_613), .C(n_626), .Y(n_601) );
OAI22xp5_ASAP7_75t_SL g668 ( .A1(n_603), .A2(n_669), .B1(n_673), .B2(n_674), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
OR2x2_ASAP7_75t_L g673 ( .A(n_605), .B(n_606), .Y(n_673) );
AND2x2_ASAP7_75t_L g681 ( .A(n_606), .B(n_662), .Y(n_681) );
CKINVDCx16_ASAP7_75t_R g606 ( .A(n_607), .Y(n_606) );
O2A1O1Ixp33_ASAP7_75t_SL g689 ( .A1(n_607), .A2(n_690), .B(n_691), .C(n_692), .Y(n_689) );
OR2x2_ASAP7_75t_L g716 ( .A(n_607), .B(n_717), .Y(n_716) );
AND2x2_ASAP7_75t_L g610 ( .A(n_611), .B(n_612), .Y(n_610) );
OAI21xp33_ASAP7_75t_L g613 ( .A1(n_614), .A2(n_617), .B(n_619), .Y(n_613) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
O2A1O1Ixp33_ASAP7_75t_L g651 ( .A1(n_615), .A2(n_652), .B(n_653), .C(n_656), .Y(n_651) );
OAI21xp33_ASAP7_75t_SL g619 ( .A1(n_620), .A2(n_621), .B(n_622), .Y(n_619) );
AND2x2_ASAP7_75t_L g684 ( .A(n_623), .B(n_642), .Y(n_684) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g662 ( .A(n_625), .B(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g667 ( .A(n_627), .Y(n_667) );
NAND3xp33_ASAP7_75t_SL g630 ( .A(n_631), .B(n_651), .C(n_664), .Y(n_630) );
AOI211xp5_ASAP7_75t_L g631 ( .A1(n_632), .A2(n_634), .B(n_635), .C(n_643), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_633), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
INVx1_ASAP7_75t_L g701 ( .A(n_638), .Y(n_701) );
OR2x2_ASAP7_75t_L g638 ( .A(n_639), .B(n_641), .Y(n_638) );
INVx1_ASAP7_75t_L g661 ( .A(n_640), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_640), .B(n_709), .Y(n_708) );
INVxp67_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
A2O1A1Ixp33_ASAP7_75t_L g643 ( .A1(n_644), .A2(n_645), .B(n_646), .C(n_647), .Y(n_643) );
INVx2_ASAP7_75t_SL g655 ( .A(n_645), .Y(n_655) );
OAI22xp5_ASAP7_75t_L g656 ( .A1(n_646), .A2(n_657), .B1(n_659), .B2(n_660), .Y(n_656) );
OAI21xp33_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_649), .B(n_650), .Y(n_647) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_661), .B(n_662), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g664 ( .A1(n_665), .A2(n_667), .B(n_668), .C(n_675), .Y(n_664) );
INVx1_ASAP7_75t_SL g665 ( .A(n_666), .Y(n_665) );
INVxp33_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g718 ( .A(n_672), .Y(n_718) );
NAND4xp25_ASAP7_75t_L g677 ( .A(n_678), .B(n_693), .C(n_706), .D(n_711), .Y(n_677) );
AOI211xp5_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_681), .B(n_682), .C(n_689), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI21xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_685), .B(n_687), .Y(n_682) );
AOI21xp33_ASAP7_75t_L g702 ( .A1(n_683), .A2(n_703), .B(n_705), .Y(n_702) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_690), .B(n_716), .Y(n_715) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_L g698 ( .A(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g706 ( .A(n_707), .B(n_710), .Y(n_706) );
INVxp67_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
INVx1_ASAP7_75t_L g726 ( .A(n_719), .Y(n_726) );
INVx2_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
INVx1_ASAP7_75t_SL g727 ( .A(n_728), .Y(n_727) );
endmodule