module real_jpeg_27267_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_28;
wire n_44;
wire n_62;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_118;
wire n_17;
wire n_116;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx11_ASAP7_75t_SL g39 ( 
.A(n_0),
.Y(n_39)
);

HB1xp67_ASAP7_75t_L g56 ( 
.A(n_1),
.Y(n_56)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_1),
.Y(n_72)
);

BUFx12_ASAP7_75t_L g69 ( 
.A(n_2),
.Y(n_69)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx8_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_5),
.A2(n_37),
.B1(n_38),
.B2(n_40),
.Y(n_36)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_5),
.A2(n_8),
.B(n_38),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g21 ( 
.A1(n_6),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_6),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_6),
.A2(n_18),
.B1(n_20),
.B2(n_24),
.Y(n_34)
);

AOI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_6),
.A2(n_24),
.B1(n_37),
.B2(n_38),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g17 ( 
.A1(n_7),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_17)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_7),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_8),
.A2(n_22),
.B1(n_23),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_8),
.A2(n_18),
.B1(n_20),
.B2(n_27),
.Y(n_42)
);

AOI21xp33_ASAP7_75t_SL g48 ( 
.A1(n_8),
.A2(n_18),
.B(n_30),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_8),
.A2(n_27),
.B1(n_37),
.B2(n_38),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_8),
.B(n_67),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_8),
.B(n_17),
.Y(n_93)
);

HAxp5_ASAP7_75t_SL g9 ( 
.A(n_10),
.B(n_85),
.CON(n_9),
.SN(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_84),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_58),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_13),
.B(n_58),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_32),
.C(n_46),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_14),
.A2(n_15),
.B1(n_32),
.B2(n_102),
.Y(n_117)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

OAI21xp5_ASAP7_75t_L g15 ( 
.A1(n_16),
.A2(n_21),
.B(n_25),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_16),
.A2(n_21),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_29),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g20 ( 
.A(n_18),
.Y(n_20)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_18),
.A2(n_20),
.B1(n_40),
.B2(n_45),
.Y(n_44)
);

A2O1A1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_18),
.A2(n_27),
.B(n_40),
.C(n_90),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_22),
.B1(n_23),
.B2(n_30),
.Y(n_29)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_22),
.A2(n_23),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

A2O1A1Ixp33_ASAP7_75t_L g47 ( 
.A1(n_23),
.A2(n_27),
.B(n_31),
.C(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

CKINVDCx14_ASAP7_75t_R g63 ( 
.A(n_26),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_27),
.B(n_107),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g110 ( 
.A(n_27),
.B(n_36),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g62 ( 
.A(n_28),
.Y(n_62)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_32),
.B(n_89),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_32),
.A2(n_89),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_32),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g32 ( 
.A1(n_33),
.A2(n_35),
.B(n_41),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_34),
.A2(n_36),
.B1(n_42),
.B2(n_43),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g105 ( 
.A(n_37),
.B(n_106),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_55),
.Y(n_54)
);

INVx11_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_43),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_46),
.B(n_117),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_49),
.B1(n_50),
.B2(n_57),
.Y(n_46)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_47),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_57),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_53),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_51),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_52),
.A2(n_54),
.B1(n_72),
.B2(n_73),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_54),
.Y(n_75)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_60),
.B1(n_78),
.B2(n_79),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g60 ( 
.A1(n_61),
.A2(n_64),
.B1(n_76),
.B2(n_77),
.Y(n_60)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_64),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_66),
.B1(n_70),
.B2(n_71),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_100),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_70),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_71),
.B(n_105),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_74),
.Y(n_71)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_80),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_81),
.A2(n_83),
.B1(n_93),
.B2(n_94),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_94),
.C(n_96),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_114),
.B(n_118),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_98),
.B(n_113),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_88),
.B(n_91),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_88),
.B(n_91),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_89),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_92),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_92),
.Y(n_97)
);

CKINVDCx16_ASAP7_75t_R g94 ( 
.A(n_93),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_96),
.B(n_110),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_96),
.B(n_110),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B(n_112),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_104),
.A2(n_109),
.B(n_111),
.Y(n_103)
);

INVx5_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_115),
.B(n_116),
.Y(n_118)
);


endmodule