module fake_jpeg_12385_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_137;
wire n_74;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_122;
wire n_75;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

INVx1_ASAP7_75t_SL g16 ( 
.A(n_13),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

BUFx12_ASAP7_75t_L g18 ( 
.A(n_2),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx5_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_3),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_3),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_4),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_9),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_25),
.B(n_14),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_40),
.B(n_41),
.Y(n_78)
);

AOI21xp33_ASAP7_75t_L g41 ( 
.A1(n_25),
.A2(n_14),
.B(n_12),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_42),
.B(n_44),
.Y(n_86)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_27),
.Y(n_43)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_32),
.B(n_12),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_45),
.Y(n_92)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_15),
.Y(n_46)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_46),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_34),
.B(n_16),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_47),
.B(n_51),
.Y(n_89)
);

BUFx16f_ASAP7_75t_L g48 ( 
.A(n_30),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g90 ( 
.A(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_16),
.A2(n_12),
.B1(n_10),
.B2(n_9),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_49),
.B(n_19),
.C(n_20),
.Y(n_95)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_30),
.Y(n_50)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_50),
.Y(n_80)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_34),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_18),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_52),
.B(n_54),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_22),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_53),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g54 ( 
.A(n_26),
.B(n_8),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx16f_ASAP7_75t_L g56 ( 
.A(n_30),
.Y(n_56)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_56),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_22),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

BUFx6f_ASAP7_75t_SL g58 ( 
.A(n_23),
.Y(n_58)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_58),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_22),
.Y(n_59)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_59),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_60),
.Y(n_74)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_61),
.B(n_62),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_18),
.Y(n_62)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_15),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g116 ( 
.A(n_63),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_64),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_18),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_65),
.B(n_24),
.Y(n_119)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_24),
.Y(n_66)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_15),
.Y(n_67)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_29),
.Y(n_68)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_68),
.Y(n_83)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_69),
.Y(n_96)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_72),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_53),
.A2(n_21),
.B1(n_38),
.B2(n_16),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_81),
.A2(n_100),
.B1(n_35),
.B2(n_18),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_49),
.A2(n_38),
.B1(n_21),
.B2(n_28),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_82),
.A2(n_85),
.B1(n_117),
.B2(n_80),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_30),
.Y(n_85)
);

AND2x2_ASAP7_75t_L g163 ( 
.A(n_85),
.B(n_95),
.Y(n_163)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_43),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_87),
.B(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_29),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_98),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_66),
.A2(n_21),
.B1(n_28),
.B2(n_19),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_91),
.A2(n_97),
.B1(n_101),
.B2(n_35),
.Y(n_139)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_58),
.A2(n_28),
.B1(n_19),
.B2(n_20),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_52),
.B(n_31),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_57),
.A2(n_64),
.B1(n_59),
.B2(n_38),
.Y(n_100)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_54),
.A2(n_20),
.B1(n_38),
.B2(n_36),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_62),
.B(n_33),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_102),
.B(n_108),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_45),
.A2(n_33),
.B1(n_31),
.B2(n_26),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_L g133 ( 
.A1(n_104),
.A2(n_17),
.B1(n_35),
.B2(n_18),
.Y(n_133)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_65),
.B(n_37),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g109 ( 
.A(n_48),
.Y(n_109)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_109),
.Y(n_167)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g137 ( 
.A(n_110),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_56),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_112),
.B(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_46),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_114),
.B(n_115),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_63),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_55),
.B(n_36),
.C(n_17),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_117),
.B(n_0),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_119),
.B(n_24),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_60),
.B(n_37),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_1),
.Y(n_150)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_60),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_121),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_88),
.B(n_40),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g185 ( 
.A(n_123),
.B(n_145),
.Y(n_185)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_108),
.Y(n_124)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_124),
.Y(n_174)
);

OR2x2_ASAP7_75t_SL g125 ( 
.A(n_78),
.B(n_60),
.Y(n_125)
);

OR2x2_ASAP7_75t_L g199 ( 
.A(n_125),
.B(n_159),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_100),
.A2(n_37),
.B1(n_36),
.B2(n_17),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_127),
.A2(n_152),
.B1(n_156),
.B2(n_162),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g128 ( 
.A(n_76),
.Y(n_128)
);

BUFx2_ASAP7_75t_L g175 ( 
.A(n_128),
.Y(n_175)
);

NAND3xp33_ASAP7_75t_L g181 ( 
.A(n_130),
.B(n_132),
.C(n_135),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_103),
.B(n_8),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_133),
.B(n_134),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_86),
.B(n_89),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_136),
.Y(n_179)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g198 ( 
.A(n_141),
.B(n_150),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_98),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_143),
.B(n_162),
.Y(n_186)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_83),
.Y(n_144)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_144),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_105),
.B(n_102),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_95),
.B(n_8),
.Y(n_146)
);

NAND3xp33_ASAP7_75t_L g192 ( 
.A(n_146),
.B(n_7),
.C(n_126),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_111),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_147),
.B(n_148),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_120),
.B(n_0),
.Y(n_148)
);

BUFx2_ASAP7_75t_SL g149 ( 
.A(n_90),
.Y(n_149)
);

BUFx24_ASAP7_75t_L g187 ( 
.A(n_149),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_73),
.Y(n_151)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_151),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_81),
.A2(n_35),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_153),
.A2(n_166),
.B1(n_168),
.B2(n_162),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g154 ( 
.A(n_90),
.Y(n_154)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_154),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_72),
.B(n_110),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_155),
.B(n_5),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_82),
.A2(n_118),
.B1(n_76),
.B2(n_106),
.Y(n_156)
);

INVx4_ASAP7_75t_SL g157 ( 
.A(n_84),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_157),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_73),
.B(n_1),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_158),
.B(n_164),
.Y(n_183)
);

OR2x2_ASAP7_75t_SL g159 ( 
.A(n_96),
.B(n_35),
.Y(n_159)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx2_ASAP7_75t_L g205 ( 
.A(n_161),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g162 ( 
.A(n_106),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_92),
.B(n_2),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_79),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_165),
.B(n_122),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_118),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_166)
);

OA21x2_ASAP7_75t_L g168 ( 
.A1(n_85),
.A2(n_5),
.B(n_6),
.Y(n_168)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_168),
.A2(n_129),
.B(n_137),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_156),
.A2(n_80),
.B1(n_71),
.B2(n_75),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_171),
.A2(n_195),
.B1(n_203),
.B2(n_169),
.Y(n_212)
);

AOI32xp33_ASAP7_75t_L g172 ( 
.A1(n_125),
.A2(n_80),
.A3(n_84),
.B1(n_71),
.B2(n_70),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_172),
.B(n_176),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_124),
.A2(n_75),
.B1(n_96),
.B2(n_99),
.Y(n_173)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_173),
.A2(n_180),
.B(n_182),
.Y(n_233)
);

XOR2xp5_ASAP7_75t_L g176 ( 
.A(n_163),
.B(n_116),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_176),
.B(n_178),
.C(n_199),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_163),
.B(n_94),
.C(n_107),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_153),
.A2(n_142),
.B1(n_143),
.B2(n_140),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_142),
.A2(n_94),
.B1(n_70),
.B2(n_74),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_140),
.A2(n_74),
.B(n_6),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g239 ( 
.A(n_184),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_188),
.B(n_191),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_163),
.A2(n_7),
.B(n_150),
.Y(n_189)
);

AND2x2_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_197),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_123),
.B(n_7),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_191),
.Y(n_227)
);

AOI32xp33_ASAP7_75t_L g193 ( 
.A1(n_158),
.A2(n_164),
.A3(n_159),
.B1(n_136),
.B2(n_144),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_193),
.B(n_207),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_127),
.A2(n_152),
.B1(n_141),
.B2(n_133),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_131),
.B(n_161),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_138),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_151),
.A2(n_128),
.B1(n_169),
.B2(n_138),
.Y(n_202)
);

OA21x2_ASAP7_75t_L g237 ( 
.A1(n_202),
.A2(n_205),
.B(n_200),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_204),
.B(n_177),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_168),
.A2(n_155),
.B1(n_122),
.B2(n_165),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_206),
.Y(n_240)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_179),
.Y(n_209)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_209),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_211),
.B(n_218),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_212),
.A2(n_217),
.B1(n_228),
.B2(n_229),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g214 ( 
.A(n_187),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_214),
.B(n_216),
.Y(n_253)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_215),
.B(n_232),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_187),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_203),
.A2(n_160),
.B1(n_154),
.B2(n_137),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_183),
.B(n_137),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_179),
.Y(n_219)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_219),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_183),
.B(n_160),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_220),
.B(n_221),
.Y(n_261)
);

AO22x1_ASAP7_75t_SL g221 ( 
.A1(n_174),
.A2(n_157),
.B1(n_167),
.B2(n_198),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_180),
.B(n_167),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_224),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_174),
.B(n_157),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_198),
.B(n_184),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_225),
.B(n_227),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_SL g226 ( 
.A1(n_190),
.A2(n_172),
.B1(n_187),
.B2(n_182),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_226),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_190),
.A2(n_199),
.B1(n_206),
.B2(n_198),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_207),
.B1(n_170),
.B2(n_189),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g246 ( 
.A1(n_230),
.A2(n_188),
.B(n_181),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_201),
.B(n_185),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_231),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_178),
.B(n_194),
.Y(n_232)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_194),
.Y(n_234)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_234),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_235),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_170),
.B(n_173),
.C(n_200),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_236),
.B(n_170),
.C(n_202),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_237),
.A2(n_187),
.B(n_196),
.Y(n_243)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_205),
.Y(n_238)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_238),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_246),
.C(n_257),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g269 ( 
.A1(n_243),
.A2(n_265),
.B(n_210),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_175),
.B1(n_208),
.B2(n_239),
.Y(n_247)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_247),
.Y(n_275)
);

AO21x1_ASAP7_75t_L g249 ( 
.A1(n_240),
.A2(n_222),
.B(n_229),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_249),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_225),
.A2(n_175),
.B1(n_208),
.B2(n_222),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_259),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_215),
.B(n_232),
.C(n_230),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g259 ( 
.A(n_238),
.Y(n_259)
);

OAI32xp33_ASAP7_75t_L g260 ( 
.A1(n_223),
.A2(n_220),
.A3(n_233),
.B1(n_218),
.B2(n_211),
.Y(n_260)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_260),
.Y(n_284)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_209),
.Y(n_263)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_228),
.A2(n_210),
.B(n_236),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_213),
.B(n_216),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g265 ( 
.A1(n_210),
.A2(n_233),
.B(n_221),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_219),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_266),
.B(n_248),
.Y(n_286)
);

OA21x2_ASAP7_75t_L g268 ( 
.A1(n_261),
.A2(n_265),
.B(n_262),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_268),
.A2(n_275),
.B1(n_277),
.B2(n_276),
.Y(n_305)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_269),
.B(n_288),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_257),
.B(n_233),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_271),
.B(n_276),
.C(n_278),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_248),
.A2(n_262),
.B1(n_242),
.B2(n_249),
.Y(n_272)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_217),
.B(n_214),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_SL g290 ( 
.A1(n_273),
.A2(n_281),
.B(n_247),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_258),
.B(n_233),
.C(n_221),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_258),
.B(n_221),
.C(n_224),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_264),
.B(n_234),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_279),
.B(n_280),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_251),
.A2(n_212),
.B1(n_213),
.B2(n_237),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_256),
.B(n_237),
.Y(n_282)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_254),
.Y(n_304)
);

NAND3xp33_ASAP7_75t_L g285 ( 
.A(n_256),
.B(n_237),
.C(n_246),
.Y(n_285)
);

OAI322xp33_ASAP7_75t_L g292 ( 
.A1(n_285),
.A2(n_245),
.A3(n_247),
.B1(n_241),
.B2(n_260),
.C1(n_266),
.C2(n_250),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_287),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g287 ( 
.A1(n_242),
.A2(n_249),
.B1(n_267),
.B2(n_261),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_267),
.A2(n_255),
.B(n_253),
.Y(n_288)
);

CKINVDCx16_ASAP7_75t_R g289 ( 
.A(n_253),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_254),
.Y(n_303)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_269),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g313 ( 
.A1(n_292),
.A2(n_273),
.B(n_275),
.Y(n_313)
);

MAJx2_ASAP7_75t_L g294 ( 
.A(n_270),
.B(n_245),
.C(n_244),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_294),
.B(n_278),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_L g295 ( 
.A(n_270),
.B(n_244),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_295),
.B(n_299),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_274),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_297),
.B(n_293),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_277),
.A2(n_250),
.B1(n_252),
.B2(n_263),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_298),
.A2(n_305),
.B1(n_284),
.B2(n_283),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g299 ( 
.A(n_271),
.B(n_252),
.Y(n_299)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_259),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_302),
.B(n_304),
.Y(n_315)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_303),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_306),
.B(n_291),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_307),
.B(n_311),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_280),
.C(n_282),
.Y(n_309)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_309),
.B(n_310),
.C(n_317),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_299),
.B(n_288),
.C(n_274),
.Y(n_310)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_301),
.A2(n_281),
.B(n_284),
.Y(n_312)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_312),
.A2(n_313),
.B(n_309),
.Y(n_325)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_314),
.A2(n_310),
.B1(n_308),
.B2(n_315),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_316),
.A2(n_298),
.B1(n_302),
.B2(n_291),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_296),
.B(n_268),
.C(n_283),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_296),
.B(n_268),
.C(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_300),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g319 ( 
.A1(n_306),
.A2(n_291),
.B1(n_305),
.B2(n_304),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_319),
.B(n_320),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_311),
.B(n_300),
.Y(n_320)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_321),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_322),
.B(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_325),
.C(n_326),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_317),
.C(n_318),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_331),
.B(n_327),
.C(n_323),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_334),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_331),
.A2(n_321),
.B(n_319),
.Y(n_334)
);

NAND3xp33_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_307),
.C(n_320),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_L g336 ( 
.A1(n_335),
.A2(n_329),
.B(n_330),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_329),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_337),
.B1(n_332),
.B2(n_315),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_332),
.Y(n_340)
);


endmodule