module fake_netlist_1_7958_n_716 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_716);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_420;
wire n_342;
wire n_423;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_597;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_406;
wire n_395;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_44), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_6), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_45), .Y(n_81) );
CKINVDCx20_ASAP7_75t_R g82 ( .A(n_38), .Y(n_82) );
CKINVDCx20_ASAP7_75t_R g83 ( .A(n_59), .Y(n_83) );
HB1xp67_ASAP7_75t_L g84 ( .A(n_62), .Y(n_84) );
BUFx3_ASAP7_75t_L g85 ( .A(n_5), .Y(n_85) );
INVx1_ASAP7_75t_SL g86 ( .A(n_6), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_3), .Y(n_87) );
CKINVDCx20_ASAP7_75t_R g88 ( .A(n_56), .Y(n_88) );
BUFx6f_ASAP7_75t_L g89 ( .A(n_41), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_37), .Y(n_90) );
BUFx3_ASAP7_75t_L g91 ( .A(n_35), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_25), .Y(n_92) );
CKINVDCx16_ASAP7_75t_R g93 ( .A(n_30), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_33), .Y(n_94) );
BUFx3_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_75), .Y(n_96) );
INVxp67_ASAP7_75t_L g97 ( .A(n_65), .Y(n_97) );
INVxp33_ASAP7_75t_SL g98 ( .A(n_0), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_42), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_77), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_46), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_47), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_36), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_68), .Y(n_104) );
HB1xp67_ASAP7_75t_L g105 ( .A(n_76), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_72), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_23), .Y(n_107) );
INVx2_ASAP7_75t_L g108 ( .A(n_28), .Y(n_108) );
CKINVDCx5p33_ASAP7_75t_R g109 ( .A(n_52), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_16), .Y(n_110) );
BUFx6f_ASAP7_75t_L g111 ( .A(n_19), .Y(n_111) );
BUFx6f_ASAP7_75t_L g112 ( .A(n_64), .Y(n_112) );
BUFx3_ASAP7_75t_L g113 ( .A(n_51), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_78), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_16), .Y(n_115) );
INVxp67_ASAP7_75t_L g116 ( .A(n_1), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_73), .Y(n_117) );
INVxp67_ASAP7_75t_SL g118 ( .A(n_61), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_53), .Y(n_119) );
CKINVDCx5p33_ASAP7_75t_R g120 ( .A(n_55), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_8), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_5), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_13), .Y(n_123) );
BUFx3_ASAP7_75t_L g124 ( .A(n_1), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_66), .Y(n_125) );
NOR2xp33_ASAP7_75t_L g126 ( .A(n_58), .B(n_71), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_43), .Y(n_127) );
INVx3_ASAP7_75t_L g128 ( .A(n_85), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_108), .Y(n_129) );
AND2x4_ASAP7_75t_L g130 ( .A(n_85), .B(n_0), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_93), .B(n_2), .Y(n_131) );
AND2x6_ASAP7_75t_L g132 ( .A(n_91), .B(n_113), .Y(n_132) );
CKINVDCx20_ASAP7_75t_R g133 ( .A(n_115), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_79), .Y(n_135) );
INVxp67_ASAP7_75t_L g136 ( .A(n_95), .Y(n_136) );
HB1xp67_ASAP7_75t_L g137 ( .A(n_115), .Y(n_137) );
NAND2xp5_ASAP7_75t_L g138 ( .A(n_84), .B(n_2), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_89), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_92), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_108), .Y(n_142) );
AND2x2_ASAP7_75t_L g143 ( .A(n_99), .B(n_3), .Y(n_143) );
AND2x2_ASAP7_75t_L g144 ( .A(n_105), .B(n_4), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_103), .Y(n_145) );
AND2x6_ASAP7_75t_L g146 ( .A(n_91), .B(n_27), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_103), .Y(n_147) );
INVx1_ASAP7_75t_L g148 ( .A(n_117), .Y(n_148) );
AND2x4_ASAP7_75t_L g149 ( .A(n_95), .B(n_4), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_124), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_116), .B(n_7), .Y(n_151) );
BUFx6f_ASAP7_75t_L g152 ( .A(n_89), .Y(n_152) );
AND2x2_ASAP7_75t_L g153 ( .A(n_124), .B(n_8), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_117), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_110), .Y(n_155) );
HB1xp67_ASAP7_75t_L g156 ( .A(n_110), .Y(n_156) );
BUFx6f_ASAP7_75t_L g157 ( .A(n_89), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_81), .Y(n_158) );
INVx3_ASAP7_75t_L g159 ( .A(n_80), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_94), .Y(n_160) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_89), .Y(n_161) );
XOR2xp5_ASAP7_75t_L g162 ( .A(n_98), .B(n_9), .Y(n_162) );
AND2x4_ASAP7_75t_L g163 ( .A(n_113), .B(n_9), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_100), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_101), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_102), .Y(n_166) );
AOI22xp5_ASAP7_75t_L g167 ( .A1(n_98), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_104), .Y(n_168) );
BUFx2_ASAP7_75t_L g169 ( .A(n_90), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_107), .Y(n_170) );
BUFx2_ASAP7_75t_L g171 ( .A(n_90), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_140), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_130), .Y(n_173) );
INVx1_ASAP7_75t_L g174 ( .A(n_130), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_169), .Y(n_175) );
INVx2_ASAP7_75t_L g176 ( .A(n_140), .Y(n_176) );
BUFx3_ASAP7_75t_L g177 ( .A(n_169), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g178 ( .A(n_171), .B(n_97), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_130), .Y(n_179) );
NAND2xp5_ASAP7_75t_SL g180 ( .A(n_171), .B(n_109), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_129), .Y(n_181) );
INVx1_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_140), .Y(n_183) );
NAND2xp5_ASAP7_75t_SL g184 ( .A(n_136), .B(n_109), .Y(n_184) );
INVx2_ASAP7_75t_L g185 ( .A(n_140), .Y(n_185) );
BUFx6f_ASAP7_75t_L g186 ( .A(n_140), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_158), .B(n_127), .Y(n_187) );
BUFx3_ASAP7_75t_L g188 ( .A(n_132), .Y(n_188) );
HB1xp67_ASAP7_75t_L g189 ( .A(n_137), .Y(n_189) );
AND2x4_ASAP7_75t_L g190 ( .A(n_163), .B(n_87), .Y(n_190) );
NOR2xp33_ASAP7_75t_L g191 ( .A(n_158), .B(n_125), .Y(n_191) );
INVx4_ASAP7_75t_SL g192 ( .A(n_146), .Y(n_192) );
AND2x4_ASAP7_75t_L g193 ( .A(n_163), .B(n_123), .Y(n_193) );
AND2x2_ASAP7_75t_L g194 ( .A(n_144), .B(n_127), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_134), .B(n_96), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_152), .Y(n_196) );
INVx4_ASAP7_75t_L g197 ( .A(n_146), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_163), .B(n_122), .Y(n_198) );
INVxp67_ASAP7_75t_L g199 ( .A(n_131), .Y(n_199) );
INVx2_ASAP7_75t_L g200 ( .A(n_152), .Y(n_200) );
OAI22xp5_ASAP7_75t_L g201 ( .A1(n_133), .A2(n_82), .B1(n_83), .B2(n_88), .Y(n_201) );
AND2x6_ASAP7_75t_L g202 ( .A(n_163), .B(n_112), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_152), .Y(n_203) );
OR2x2_ASAP7_75t_L g204 ( .A(n_156), .B(n_86), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_144), .A2(n_121), .B1(n_114), .B2(n_120), .Y(n_205) );
CKINVDCx11_ASAP7_75t_R g206 ( .A(n_149), .Y(n_206) );
NAND2xp5_ASAP7_75t_SL g207 ( .A(n_134), .B(n_135), .Y(n_207) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_160), .B(n_96), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_160), .B(n_114), .Y(n_209) );
BUFx3_ASAP7_75t_L g210 ( .A(n_132), .Y(n_210) );
CKINVDCx5p33_ASAP7_75t_R g211 ( .A(n_131), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_152), .Y(n_212) );
INVx2_ASAP7_75t_SL g213 ( .A(n_128), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_152), .Y(n_214) );
NOR2x1p5_ASAP7_75t_L g215 ( .A(n_159), .B(n_120), .Y(n_215) );
INVx1_ASAP7_75t_L g216 ( .A(n_129), .Y(n_216) );
INVx3_ASAP7_75t_L g217 ( .A(n_149), .Y(n_217) );
INVx1_ASAP7_75t_L g218 ( .A(n_142), .Y(n_218) );
INVx5_ASAP7_75t_L g219 ( .A(n_146), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_157), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_149), .Y(n_221) );
INVxp33_ASAP7_75t_SL g222 ( .A(n_143), .Y(n_222) );
INVx2_ASAP7_75t_L g223 ( .A(n_157), .Y(n_223) );
BUFx2_ASAP7_75t_L g224 ( .A(n_143), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_164), .B(n_119), .Y(n_225) );
NOR2xp33_ASAP7_75t_SL g226 ( .A(n_146), .B(n_119), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_149), .Y(n_227) );
BUFx3_ASAP7_75t_L g228 ( .A(n_132), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_164), .B(n_168), .Y(n_229) );
NOR2xp33_ASAP7_75t_L g230 ( .A(n_165), .B(n_106), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_153), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_153), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_165), .B(n_106), .Y(n_233) );
HB1xp67_ASAP7_75t_L g234 ( .A(n_162), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_128), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g236 ( .A(n_187), .B(n_139), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_213), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_178), .B(n_168), .Y(n_238) );
AND2x4_ASAP7_75t_SL g239 ( .A(n_175), .B(n_167), .Y(n_239) );
INVx5_ASAP7_75t_L g240 ( .A(n_202), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_208), .B(n_147), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_209), .B(n_147), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_235), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_233), .B(n_135), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_235), .Y(n_245) );
INVx4_ASAP7_75t_L g246 ( .A(n_206), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_213), .Y(n_247) );
OAI22xp5_ASAP7_75t_L g248 ( .A1(n_222), .A2(n_138), .B1(n_166), .B2(n_148), .Y(n_248) );
BUFx3_ASAP7_75t_L g249 ( .A(n_188), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_181), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_181), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_216), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_225), .B(n_230), .Y(n_253) );
BUFx3_ASAP7_75t_L g254 ( .A(n_188), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_231), .B(n_166), .Y(n_255) );
INVx4_ASAP7_75t_L g256 ( .A(n_206), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_194), .B(n_139), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g258 ( .A(n_194), .B(n_148), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g259 ( .A(n_229), .B(n_141), .Y(n_259) );
AND2x2_ASAP7_75t_L g260 ( .A(n_224), .B(n_151), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_232), .B(n_141), .Y(n_261) );
AOI22xp5_ASAP7_75t_L g262 ( .A1(n_222), .A2(n_132), .B1(n_170), .B2(n_146), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_195), .B(n_159), .Y(n_263) );
INVx3_ASAP7_75t_L g264 ( .A(n_217), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_190), .B(n_159), .Y(n_265) );
CKINVDCx20_ASAP7_75t_R g266 ( .A(n_201), .Y(n_266) );
INVx1_ASAP7_75t_L g267 ( .A(n_216), .Y(n_267) );
INVx2_ASAP7_75t_SL g268 ( .A(n_177), .Y(n_268) );
NAND2xp5_ASAP7_75t_SL g269 ( .A(n_197), .B(n_145), .Y(n_269) );
OAI22xp5_ASAP7_75t_SL g270 ( .A1(n_234), .A2(n_162), .B1(n_155), .B2(n_170), .Y(n_270) );
BUFx6f_ASAP7_75t_L g271 ( .A(n_197), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_218), .Y(n_272) );
AOI22xp33_ASAP7_75t_L g273 ( .A1(n_173), .A2(n_145), .B1(n_154), .B2(n_146), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_190), .B(n_150), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g275 ( .A(n_190), .B(n_150), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g276 ( .A1(n_199), .A2(n_128), .B1(n_150), .B2(n_154), .Y(n_276) );
AND2x4_ASAP7_75t_L g277 ( .A(n_215), .B(n_155), .Y(n_277) );
AND2x4_ASAP7_75t_L g278 ( .A(n_177), .B(n_146), .Y(n_278) );
INVx2_ASAP7_75t_SL g279 ( .A(n_204), .Y(n_279) );
HB1xp67_ASAP7_75t_L g280 ( .A(n_204), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_193), .B(n_132), .Y(n_281) );
A2O1A1Ixp33_ASAP7_75t_L g282 ( .A1(n_174), .A2(n_142), .B(n_118), .C(n_126), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_193), .B(n_132), .Y(n_283) );
AO22x1_ASAP7_75t_L g284 ( .A1(n_211), .A2(n_132), .B1(n_111), .B2(n_112), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_193), .B(n_112), .Y(n_285) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_198), .B(n_112), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_198), .B(n_112), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_198), .B(n_111), .Y(n_288) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_224), .B(n_111), .Y(n_289) );
BUFx6f_ASAP7_75t_L g290 ( .A(n_197), .Y(n_290) );
NAND2xp5_ASAP7_75t_L g291 ( .A(n_184), .B(n_111), .Y(n_291) );
OAI22xp5_ASAP7_75t_L g292 ( .A1(n_211), .A2(n_179), .B1(n_227), .B2(n_182), .Y(n_292) );
NAND2xp5_ASAP7_75t_SL g293 ( .A(n_219), .B(n_111), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_205), .B(n_89), .Y(n_294) );
A2O1A1Ixp33_ASAP7_75t_L g295 ( .A1(n_221), .A2(n_161), .B(n_157), .C(n_12), .Y(n_295) );
BUFx3_ASAP7_75t_L g296 ( .A(n_210), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_210), .Y(n_297) );
INVx1_ASAP7_75t_SL g298 ( .A(n_189), .Y(n_298) );
AOI22xp5_ASAP7_75t_L g299 ( .A1(n_180), .A2(n_157), .B1(n_161), .B2(n_13), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_191), .B(n_10), .Y(n_300) );
AND3x1_ASAP7_75t_L g301 ( .A(n_226), .B(n_11), .C(n_14), .Y(n_301) );
AOI22xp5_ASAP7_75t_L g302 ( .A1(n_217), .A2(n_161), .B1(n_157), .B2(n_14), .Y(n_302) );
AOI22xp5_ASAP7_75t_L g303 ( .A1(n_217), .A2(n_161), .B1(n_15), .B2(n_18), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_202), .B(n_161), .Y(n_304) );
NAND2xp5_ASAP7_75t_SL g305 ( .A(n_271), .B(n_219), .Y(n_305) );
INVx2_ASAP7_75t_L g306 ( .A(n_264), .Y(n_306) );
BUFx2_ASAP7_75t_L g307 ( .A(n_298), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_238), .B(n_207), .Y(n_308) );
AOI21xp5_ASAP7_75t_L g309 ( .A1(n_269), .A2(n_219), .B(n_228), .Y(n_309) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_279), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_280), .Y(n_311) );
NOR2x1_ASAP7_75t_L g312 ( .A(n_246), .B(n_218), .Y(n_312) );
OAI22xp5_ASAP7_75t_SL g313 ( .A1(n_266), .A2(n_219), .B1(n_15), .B2(n_228), .Y(n_313) );
AOI21x1_ASAP7_75t_SL g314 ( .A1(n_278), .A2(n_202), .B(n_192), .Y(n_314) );
INVxp67_ASAP7_75t_SL g315 ( .A(n_280), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_269), .A2(n_219), .B(n_192), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_246), .Y(n_317) );
OAI22xp5_ASAP7_75t_L g318 ( .A1(n_257), .A2(n_202), .B1(n_192), .B2(n_214), .Y(n_318) );
O2A1O1Ixp33_ASAP7_75t_SL g319 ( .A1(n_295), .A2(n_223), .B(n_214), .C(n_212), .Y(n_319) );
AND2x2_ASAP7_75t_L g320 ( .A(n_260), .B(n_202), .Y(n_320) );
O2A1O1Ixp33_ASAP7_75t_L g321 ( .A1(n_248), .A2(n_223), .B(n_212), .C(n_203), .Y(n_321) );
AO21x1_ASAP7_75t_L g322 ( .A1(n_285), .A2(n_203), .B(n_176), .Y(n_322) );
AOI21x1_ASAP7_75t_L g323 ( .A1(n_284), .A2(n_172), .B(n_185), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_274), .Y(n_324) );
INVx4_ASAP7_75t_L g325 ( .A(n_256), .Y(n_325) );
NOR2xp33_ASAP7_75t_L g326 ( .A(n_238), .B(n_202), .Y(n_326) );
NAND2xp5_ASAP7_75t_SL g327 ( .A(n_271), .B(n_192), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g328 ( .A1(n_258), .A2(n_185), .B1(n_200), .B2(n_196), .Y(n_328) );
OAI22xp5_ASAP7_75t_L g329 ( .A1(n_292), .A2(n_200), .B1(n_196), .B2(n_183), .Y(n_329) );
XNOR2xp5_ASAP7_75t_L g330 ( .A(n_270), .B(n_239), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_236), .B(n_17), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g332 ( .A1(n_277), .A2(n_183), .B1(n_176), .B2(n_172), .Y(n_332) );
AND2x4_ASAP7_75t_L g333 ( .A(n_256), .B(n_20), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_275), .Y(n_334) );
NAND3xp33_ASAP7_75t_SL g335 ( .A(n_282), .B(n_21), .C(n_22), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_241), .B(n_24), .Y(n_336) );
INVx3_ASAP7_75t_SL g337 ( .A(n_268), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_255), .B(n_26), .Y(n_338) );
O2A1O1Ixp33_ASAP7_75t_L g339 ( .A1(n_282), .A2(n_29), .B(n_31), .C(n_32), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_242), .A2(n_220), .B(n_186), .Y(n_340) );
AOI21xp5_ASAP7_75t_L g341 ( .A1(n_244), .A2(n_220), .B(n_186), .Y(n_341) );
AOI21xp33_ASAP7_75t_L g342 ( .A1(n_281), .A2(n_34), .B(n_39), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_265), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g344 ( .A(n_255), .B(n_40), .Y(n_344) );
NOR2xp33_ASAP7_75t_L g345 ( .A(n_243), .B(n_48), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_301), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_283), .A2(n_220), .B(n_186), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_259), .B(n_49), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_245), .B(n_50), .Y(n_349) );
INVx2_ASAP7_75t_L g350 ( .A(n_264), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_251), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_253), .B(n_54), .Y(n_352) );
BUFx2_ASAP7_75t_L g353 ( .A(n_278), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_277), .B(n_57), .Y(n_354) );
INVx2_ASAP7_75t_L g355 ( .A(n_272), .Y(n_355) );
A2O1A1Ixp33_ASAP7_75t_L g356 ( .A1(n_261), .A2(n_220), .B(n_186), .C(n_67), .Y(n_356) );
NAND2xp5_ASAP7_75t_SL g357 ( .A(n_271), .B(n_186), .Y(n_357) );
INVx2_ASAP7_75t_L g358 ( .A(n_351), .Y(n_358) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_307), .Y(n_359) );
AO31x2_ASAP7_75t_L g360 ( .A1(n_322), .A2(n_295), .A3(n_287), .B(n_286), .Y(n_360) );
OAI21xp5_ASAP7_75t_L g361 ( .A1(n_308), .A2(n_273), .B(n_262), .Y(n_361) );
AOI21xp5_ASAP7_75t_L g362 ( .A1(n_340), .A2(n_288), .B(n_273), .Y(n_362) );
AND2x2_ASAP7_75t_L g363 ( .A(n_315), .B(n_300), .Y(n_363) );
AO31x2_ASAP7_75t_L g364 ( .A1(n_356), .A2(n_276), .A3(n_294), .B(n_289), .Y(n_364) );
OR2x2_ASAP7_75t_L g365 ( .A(n_311), .B(n_252), .Y(n_365) );
O2A1O1Ixp33_ASAP7_75t_SL g366 ( .A1(n_352), .A2(n_291), .B(n_250), .C(n_267), .Y(n_366) );
NOR2xp33_ASAP7_75t_L g367 ( .A(n_310), .B(n_263), .Y(n_367) );
AO31x2_ASAP7_75t_L g368 ( .A1(n_356), .A2(n_263), .A3(n_304), .B(n_237), .Y(n_368) );
AO31x2_ASAP7_75t_L g369 ( .A1(n_329), .A2(n_247), .A3(n_303), .B(n_299), .Y(n_369) );
CKINVDCx9p33_ASAP7_75t_R g370 ( .A(n_326), .Y(n_370) );
NOR2xp33_ASAP7_75t_L g371 ( .A(n_330), .B(n_290), .Y(n_371) );
AO32x2_ASAP7_75t_L g372 ( .A1(n_313), .A2(n_302), .A3(n_293), .B1(n_240), .B2(n_220), .Y(n_372) );
NAND2xp5_ASAP7_75t_SL g373 ( .A(n_337), .B(n_240), .Y(n_373) );
OAI21x1_ASAP7_75t_L g374 ( .A1(n_341), .A2(n_293), .B(n_290), .Y(n_374) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_343), .B(n_290), .Y(n_375) );
AOI22xp5_ASAP7_75t_L g376 ( .A1(n_346), .A2(n_290), .B1(n_271), .B2(n_240), .Y(n_376) );
OAI21x1_ASAP7_75t_L g377 ( .A1(n_323), .A2(n_240), .B(n_297), .Y(n_377) );
NOR2xp33_ASAP7_75t_L g378 ( .A(n_325), .B(n_296), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_324), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_326), .A2(n_297), .B(n_296), .C(n_254), .Y(n_380) );
OAI21x1_ASAP7_75t_L g381 ( .A1(n_347), .A2(n_249), .B(n_254), .Y(n_381) );
INVx2_ASAP7_75t_L g382 ( .A(n_351), .Y(n_382) );
NAND2x1_ASAP7_75t_L g383 ( .A(n_355), .B(n_249), .Y(n_383) );
O2A1O1Ixp33_ASAP7_75t_SL g384 ( .A1(n_344), .A2(n_336), .B(n_331), .C(n_348), .Y(n_384) );
AO31x2_ASAP7_75t_L g385 ( .A1(n_345), .A2(n_60), .A3(n_63), .B(n_69), .Y(n_385) );
OAI21x1_ASAP7_75t_L g386 ( .A1(n_357), .A2(n_70), .B(n_74), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_334), .Y(n_387) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_355), .B(n_306), .Y(n_388) );
CKINVDCx6p67_ASAP7_75t_R g389 ( .A(n_325), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g390 ( .A(n_337), .B(n_353), .Y(n_390) );
OAI21x1_ASAP7_75t_L g391 ( .A1(n_374), .A2(n_357), .B(n_314), .Y(n_391) );
INVx1_ASAP7_75t_SL g392 ( .A(n_359), .Y(n_392) );
OAI21xp33_ASAP7_75t_L g393 ( .A1(n_363), .A2(n_338), .B(n_335), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_358), .Y(n_394) );
HB1xp67_ASAP7_75t_L g395 ( .A(n_359), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_379), .B(n_320), .Y(n_396) );
OR2x2_ASAP7_75t_L g397 ( .A(n_365), .B(n_333), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_382), .Y(n_398) );
OA21x2_ASAP7_75t_L g399 ( .A1(n_362), .A2(n_342), .B(n_349), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_381), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_367), .A2(n_387), .B1(n_390), .B2(n_361), .C(n_371), .Y(n_401) );
AO21x2_ASAP7_75t_L g402 ( .A1(n_362), .A2(n_319), .B(n_339), .Y(n_402) );
INVx1_ASAP7_75t_L g403 ( .A(n_375), .Y(n_403) );
AOI21xp5_ASAP7_75t_L g404 ( .A1(n_384), .A2(n_321), .B(n_319), .Y(n_404) );
AND2x2_ASAP7_75t_L g405 ( .A(n_375), .B(n_306), .Y(n_405) );
AOI22xp33_ASAP7_75t_SL g406 ( .A1(n_378), .A2(n_333), .B1(n_354), .B2(n_317), .Y(n_406) );
OA21x2_ASAP7_75t_L g407 ( .A1(n_386), .A2(n_328), .B(n_345), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_389), .B(n_354), .Y(n_408) );
O2A1O1Ixp33_ASAP7_75t_L g409 ( .A1(n_361), .A2(n_350), .B(n_312), .C(n_318), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_366), .A2(n_327), .B(n_305), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_388), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_360), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_360), .Y(n_413) );
AOI21xp5_ASAP7_75t_L g414 ( .A1(n_380), .A2(n_327), .B(n_305), .Y(n_414) );
OAI21x1_ASAP7_75t_L g415 ( .A1(n_377), .A2(n_316), .B(n_328), .Y(n_415) );
OAI21x1_ASAP7_75t_L g416 ( .A1(n_383), .A2(n_309), .B(n_350), .Y(n_416) );
OAI211xp5_ASAP7_75t_SL g417 ( .A1(n_373), .A2(n_332), .B(n_376), .C(n_372), .Y(n_417) );
INVx2_ASAP7_75t_L g418 ( .A(n_368), .Y(n_418) );
NAND3xp33_ASAP7_75t_L g419 ( .A(n_376), .B(n_372), .C(n_364), .Y(n_419) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_403), .B(n_364), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_400), .Y(n_421) );
AO21x2_ASAP7_75t_L g422 ( .A1(n_419), .A2(n_368), .B(n_364), .Y(n_422) );
OA21x2_ASAP7_75t_L g423 ( .A1(n_419), .A2(n_368), .B(n_360), .Y(n_423) );
BUFx3_ASAP7_75t_L g424 ( .A(n_405), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_403), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_394), .B(n_385), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_394), .B(n_385), .Y(n_427) );
INVx1_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_400), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_398), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_412), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_412), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g433 ( .A(n_405), .B(n_369), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_413), .Y(n_434) );
AND2x2_ASAP7_75t_L g435 ( .A(n_396), .B(n_385), .Y(n_435) );
BUFx3_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
AO21x2_ASAP7_75t_L g437 ( .A1(n_404), .A2(n_372), .B(n_369), .Y(n_437) );
BUFx2_ASAP7_75t_L g438 ( .A(n_400), .Y(n_438) );
AOI211xp5_ASAP7_75t_L g439 ( .A1(n_401), .A2(n_369), .B(n_370), .C(n_397), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_418), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_418), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_418), .Y(n_442) );
INVx3_ASAP7_75t_L g443 ( .A(n_391), .Y(n_443) );
INVx1_ASAP7_75t_L g444 ( .A(n_413), .Y(n_444) );
AOI21xp5_ASAP7_75t_L g445 ( .A1(n_393), .A2(n_370), .B(n_399), .Y(n_445) );
AND2x2_ASAP7_75t_L g446 ( .A(n_396), .B(n_411), .Y(n_446) );
AOI22xp5_ASAP7_75t_L g447 ( .A1(n_406), .A2(n_392), .B1(n_395), .B2(n_408), .Y(n_447) );
INVx1_ASAP7_75t_L g448 ( .A(n_411), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_393), .A2(n_409), .B1(n_417), .B2(n_414), .C(n_410), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_391), .B(n_415), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_415), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_416), .B(n_402), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_416), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_402), .A2(n_270), .B1(n_248), .B2(n_280), .C(n_401), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_402), .B(n_407), .Y(n_455) );
INVx4_ASAP7_75t_L g456 ( .A(n_424), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_425), .B(n_407), .Y(n_457) );
NOR2x1_ASAP7_75t_SL g458 ( .A(n_424), .B(n_407), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_425), .B(n_407), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g460 ( .A(n_446), .B(n_399), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_440), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_431), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_440), .Y(n_463) );
OAI221xp5_ASAP7_75t_L g464 ( .A1(n_454), .A2(n_399), .B1(n_447), .B2(n_439), .C(n_436), .Y(n_464) );
INVx2_ASAP7_75t_SL g465 ( .A(n_424), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_440), .Y(n_466) );
HB1xp67_ASAP7_75t_L g467 ( .A(n_438), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_431), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_435), .B(n_399), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_438), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_446), .B(n_435), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_432), .Y(n_472) );
AND2x2_ASAP7_75t_L g473 ( .A(n_446), .B(n_427), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_441), .Y(n_474) );
BUFx4f_ASAP7_75t_SL g475 ( .A(n_436), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_433), .B(n_444), .Y(n_476) );
AND2x4_ASAP7_75t_L g477 ( .A(n_432), .B(n_434), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_434), .Y(n_478) );
INVx3_ASAP7_75t_L g479 ( .A(n_452), .Y(n_479) );
HB1xp67_ASAP7_75t_L g480 ( .A(n_441), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_444), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_433), .B(n_420), .Y(n_482) );
BUFx6f_ASAP7_75t_L g483 ( .A(n_452), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_426), .B(n_427), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_441), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_442), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_442), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_448), .Y(n_488) );
INVx2_ASAP7_75t_L g489 ( .A(n_442), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_426), .B(n_428), .Y(n_490) );
AND2x2_ASAP7_75t_L g491 ( .A(n_428), .B(n_430), .Y(n_491) );
AND2x2_ASAP7_75t_L g492 ( .A(n_430), .B(n_448), .Y(n_492) );
BUFx3_ASAP7_75t_L g493 ( .A(n_436), .Y(n_493) );
OAI22xp5_ASAP7_75t_SL g494 ( .A1(n_447), .A2(n_439), .B1(n_420), .B2(n_423), .Y(n_494) );
INVx2_ASAP7_75t_L g495 ( .A(n_421), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_421), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_423), .B(n_422), .Y(n_497) );
INVx2_ASAP7_75t_L g498 ( .A(n_421), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_423), .B(n_422), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_429), .Y(n_500) );
NOR2x1_ASAP7_75t_SL g501 ( .A(n_429), .B(n_453), .Y(n_501) );
BUFx2_ASAP7_75t_L g502 ( .A(n_429), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_423), .B(n_422), .Y(n_503) );
AOI22xp33_ASAP7_75t_L g504 ( .A1(n_454), .A2(n_449), .B1(n_450), .B2(n_455), .Y(n_504) );
AND2x2_ASAP7_75t_L g505 ( .A(n_423), .B(n_422), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
INVx1_ASAP7_75t_L g507 ( .A(n_491), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_473), .B(n_455), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_475), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_491), .B(n_455), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g511 ( .A(n_492), .B(n_437), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_492), .B(n_437), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_473), .B(n_437), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_488), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_488), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_484), .B(n_437), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_484), .B(n_452), .Y(n_517) );
BUFx2_ASAP7_75t_L g518 ( .A(n_456), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_490), .B(n_449), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_462), .Y(n_521) );
OR2x2_ASAP7_75t_L g522 ( .A(n_471), .B(n_451), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_484), .B(n_452), .Y(n_523) );
INVx2_ASAP7_75t_SL g524 ( .A(n_456), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_462), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_479), .B(n_450), .Y(n_526) );
OA21x2_ASAP7_75t_SL g527 ( .A1(n_477), .A2(n_450), .B(n_445), .Y(n_527) );
INVx1_ASAP7_75t_L g528 ( .A(n_468), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_490), .B(n_451), .Y(n_529) );
AND2x4_ASAP7_75t_SL g530 ( .A(n_456), .B(n_450), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_471), .B(n_445), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_468), .Y(n_532) );
NAND2xp33_ASAP7_75t_R g533 ( .A(n_502), .B(n_443), .Y(n_533) );
INVx4_ASAP7_75t_L g534 ( .A(n_456), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_469), .B(n_443), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_469), .B(n_443), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_472), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_480), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_465), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_476), .B(n_443), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_472), .Y(n_541) );
NOR2xp33_ASAP7_75t_L g542 ( .A(n_475), .B(n_465), .Y(n_542) );
AND2x2_ASAP7_75t_L g543 ( .A(n_469), .B(n_477), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_477), .B(n_497), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_465), .Y(n_545) );
INVx2_ASAP7_75t_L g546 ( .A(n_487), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_477), .B(n_497), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_487), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_497), .B(n_505), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_495), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_503), .B(n_505), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_478), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_503), .B(n_482), .Y(n_553) );
INVx2_ASAP7_75t_L g554 ( .A(n_495), .Y(n_554) );
INVx2_ASAP7_75t_L g555 ( .A(n_495), .Y(n_555) );
NOR2xp67_ASAP7_75t_L g556 ( .A(n_464), .B(n_470), .Y(n_556) );
INVx6_ASAP7_75t_L g557 ( .A(n_493), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_478), .Y(n_558) );
INVx6_ASAP7_75t_L g559 ( .A(n_493), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_482), .B(n_476), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_460), .B(n_481), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_481), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_479), .B(n_483), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_460), .B(n_467), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_504), .B(n_502), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_549), .B(n_479), .Y(n_566) );
OR2x2_ASAP7_75t_L g567 ( .A(n_560), .B(n_470), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_507), .B(n_493), .Y(n_568) );
OAI221xp5_ASAP7_75t_SL g569 ( .A1(n_519), .A2(n_464), .B1(n_499), .B2(n_479), .C(n_467), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_549), .B(n_483), .Y(n_570) );
AND2x2_ASAP7_75t_L g571 ( .A(n_551), .B(n_483), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_553), .B(n_494), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_553), .B(n_494), .Y(n_573) );
INVx2_ASAP7_75t_L g574 ( .A(n_550), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_551), .B(n_483), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_560), .B(n_485), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_552), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_557), .Y(n_578) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_508), .B(n_485), .Y(n_579) );
INVxp67_ASAP7_75t_L g580 ( .A(n_518), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_543), .B(n_483), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_550), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_552), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_558), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_508), .B(n_485), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_543), .B(n_483), .Y(n_586) );
AND2x2_ASAP7_75t_L g587 ( .A(n_544), .B(n_501), .Y(n_587) );
OR2x2_ASAP7_75t_L g588 ( .A(n_510), .B(n_486), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_558), .Y(n_589) );
AND2x2_ASAP7_75t_L g590 ( .A(n_516), .B(n_499), .Y(n_590) );
HB1xp67_ASAP7_75t_L g591 ( .A(n_520), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_516), .B(n_458), .Y(n_592) );
NOR2xp33_ASAP7_75t_L g593 ( .A(n_561), .B(n_457), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_513), .B(n_486), .Y(n_594) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_556), .A2(n_457), .B1(n_459), .B2(n_506), .C(n_500), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_514), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_515), .Y(n_597) );
NOR2xp33_ASAP7_75t_L g598 ( .A(n_561), .B(n_459), .Y(n_598) );
OR2x6_ASAP7_75t_L g599 ( .A(n_534), .B(n_496), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_564), .B(n_489), .Y(n_600) );
INVx2_ASAP7_75t_L g601 ( .A(n_554), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_554), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_513), .B(n_489), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_521), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_564), .B(n_489), .Y(n_605) );
OR2x2_ASAP7_75t_L g606 ( .A(n_517), .B(n_523), .Y(n_606) );
OR2x2_ASAP7_75t_L g607 ( .A(n_517), .B(n_486), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_544), .B(n_458), .Y(n_608) );
INVxp67_ASAP7_75t_L g609 ( .A(n_518), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
AND2x4_ASAP7_75t_L g611 ( .A(n_547), .B(n_501), .Y(n_611) );
NAND2x1p5_ASAP7_75t_L g612 ( .A(n_534), .B(n_496), .Y(n_612) );
OR2x2_ASAP7_75t_L g613 ( .A(n_523), .B(n_461), .Y(n_613) );
AND2x2_ASAP7_75t_L g614 ( .A(n_547), .B(n_496), .Y(n_614) );
INVx2_ASAP7_75t_SL g615 ( .A(n_557), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_535), .B(n_506), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_528), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_532), .Y(n_618) );
OR2x2_ASAP7_75t_L g619 ( .A(n_579), .B(n_522), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_585), .B(n_522), .Y(n_620) );
OAI21xp5_ASAP7_75t_L g621 ( .A1(n_595), .A2(n_509), .B(n_542), .Y(n_621) );
OAI32xp33_ASAP7_75t_L g622 ( .A1(n_572), .A2(n_534), .A3(n_533), .B1(n_524), .B2(n_545), .Y(n_622) );
NAND4xp25_ASAP7_75t_L g623 ( .A(n_569), .B(n_527), .C(n_573), .D(n_565), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_593), .B(n_565), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_593), .B(n_512), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_590), .B(n_535), .Y(n_626) );
HB1xp67_ASAP7_75t_L g627 ( .A(n_591), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_598), .B(n_511), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_567), .Y(n_629) );
INVx1_ASAP7_75t_SL g630 ( .A(n_587), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_596), .Y(n_631) );
AND2x4_ASAP7_75t_L g632 ( .A(n_611), .B(n_563), .Y(n_632) );
OR2x2_ASAP7_75t_L g633 ( .A(n_590), .B(n_540), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_574), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_574), .Y(n_635) );
AND2x2_ASAP7_75t_L g636 ( .A(n_571), .B(n_536), .Y(n_636) );
AO21x1_ASAP7_75t_L g637 ( .A1(n_612), .A2(n_541), .B(n_562), .Y(n_637) );
AND2x2_ASAP7_75t_L g638 ( .A(n_571), .B(n_575), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_575), .B(n_536), .Y(n_639) );
INVx1_ASAP7_75t_SL g640 ( .A(n_600), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_570), .B(n_526), .Y(n_641) );
AOI22xp5_ASAP7_75t_L g642 ( .A1(n_592), .A2(n_531), .B1(n_559), .B2(n_557), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_578), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_597), .Y(n_644) );
OAI22xp33_ASAP7_75t_R g645 ( .A1(n_606), .A2(n_524), .B1(n_537), .B2(n_548), .Y(n_645) );
A2O1A1Ixp33_ASAP7_75t_L g646 ( .A1(n_611), .A2(n_530), .B(n_539), .C(n_526), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_582), .Y(n_647) );
AOI22xp5_ASAP7_75t_L g648 ( .A1(n_592), .A2(n_559), .B1(n_557), .B2(n_526), .Y(n_648) );
INVx1_ASAP7_75t_SL g649 ( .A(n_605), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g650 ( .A(n_598), .B(n_529), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_604), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_576), .B(n_520), .Y(n_652) );
NAND2xp33_ASAP7_75t_SL g653 ( .A(n_578), .B(n_548), .Y(n_653) );
INVx2_ASAP7_75t_L g654 ( .A(n_582), .Y(n_654) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_591), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_627), .Y(n_656) );
O2A1O1Ixp5_ASAP7_75t_L g657 ( .A1(n_637), .A2(n_611), .B(n_568), .C(n_618), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_623), .A2(n_570), .B1(n_566), .B2(n_599), .Y(n_658) );
INVxp67_ASAP7_75t_L g659 ( .A(n_655), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_630), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_645), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_622), .A2(n_615), .B(n_609), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_625), .B(n_616), .Y(n_663) );
O2A1O1Ixp33_ASAP7_75t_L g664 ( .A1(n_621), .A2(n_580), .B(n_599), .C(n_615), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_631), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_628), .A2(n_608), .B1(n_566), .B2(n_581), .Y(n_666) );
AND2x2_ASAP7_75t_L g667 ( .A(n_641), .B(n_586), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_624), .B(n_616), .Y(n_668) );
AOI222xp33_ASAP7_75t_L g669 ( .A1(n_629), .A2(n_608), .B1(n_610), .B2(n_617), .C1(n_603), .C2(n_594), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g670 ( .A(n_643), .B(n_577), .C(n_589), .D(n_584), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_640), .B(n_588), .Y(n_671) );
OAI21xp5_ASAP7_75t_L g672 ( .A1(n_646), .A2(n_612), .B(n_599), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_649), .B(n_613), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_644), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_651), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_650), .B(n_583), .Y(n_676) );
OAI322xp33_ASAP7_75t_L g677 ( .A1(n_619), .A2(n_607), .A3(n_586), .B1(n_581), .B2(n_614), .C1(n_601), .C2(n_602), .Y(n_677) );
AND2x4_ASAP7_75t_SL g678 ( .A(n_632), .B(n_614), .Y(n_678) );
XOR2xp5_ASAP7_75t_L g679 ( .A(n_658), .B(n_648), .Y(n_679) );
OAI22xp5_ASAP7_75t_L g680 ( .A1(n_658), .A2(n_646), .B1(n_642), .B2(n_632), .Y(n_680) );
OAI221xp5_ASAP7_75t_L g681 ( .A1(n_661), .A2(n_653), .B1(n_652), .B2(n_620), .C(n_633), .Y(n_681) );
NAND3xp33_ASAP7_75t_L g682 ( .A(n_657), .B(n_653), .C(n_647), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_L g683 ( .A1(n_657), .A2(n_637), .B(n_647), .C(n_634), .Y(n_683) );
OAI21xp5_ASAP7_75t_L g684 ( .A1(n_664), .A2(n_626), .B(n_641), .Y(n_684) );
NOR3xp33_ASAP7_75t_L g685 ( .A(n_662), .B(n_635), .C(n_634), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_672), .B(n_670), .Y(n_686) );
NOR2x1_ASAP7_75t_L g687 ( .A(n_677), .B(n_632), .Y(n_687) );
NOR2x1_ASAP7_75t_L g688 ( .A(n_660), .B(n_638), .Y(n_688) );
OAI211xp5_ASAP7_75t_L g689 ( .A1(n_669), .A2(n_626), .B(n_638), .C(n_639), .Y(n_689) );
INVx1_ASAP7_75t_L g690 ( .A(n_665), .Y(n_690) );
INVxp67_ASAP7_75t_L g691 ( .A(n_674), .Y(n_691) );
OAI21xp33_ASAP7_75t_SL g692 ( .A1(n_666), .A2(n_639), .B(n_636), .Y(n_692) );
O2A1O1Ixp33_ASAP7_75t_L g693 ( .A1(n_686), .A2(n_659), .B(n_656), .C(n_675), .Y(n_693) );
AOI221xp5_ASAP7_75t_L g694 ( .A1(n_681), .A2(n_676), .B1(n_659), .B2(n_671), .C(n_663), .Y(n_694) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_680), .A2(n_673), .B(n_668), .C(n_667), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g696 ( .A1(n_688), .A2(n_678), .B1(n_636), .B2(n_559), .Y(n_696) );
AOI22xp5_ASAP7_75t_L g697 ( .A1(n_687), .A2(n_678), .B1(n_559), .B2(n_635), .Y(n_697) );
O2A1O1Ixp33_ASAP7_75t_L g698 ( .A1(n_683), .A2(n_654), .B(n_602), .C(n_601), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_689), .A2(n_563), .B(n_654), .C(n_546), .Y(n_699) );
OAI211xp5_ASAP7_75t_L g700 ( .A1(n_679), .A2(n_546), .B(n_538), .C(n_506), .Y(n_700) );
NOR3xp33_ASAP7_75t_L g701 ( .A(n_693), .B(n_682), .C(n_692), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g702 ( .A1(n_697), .A2(n_684), .B(n_685), .C(n_691), .Y(n_702) );
OAI21xp33_ASAP7_75t_SL g703 ( .A1(n_696), .A2(n_690), .B(n_538), .Y(n_703) );
NAND3xp33_ASAP7_75t_L g704 ( .A(n_695), .B(n_563), .C(n_555), .Y(n_704) );
NAND3xp33_ASAP7_75t_SL g705 ( .A(n_699), .B(n_500), .C(n_555), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_701), .B(n_694), .Y(n_706) );
XNOR2xp5_ASAP7_75t_SL g707 ( .A(n_702), .B(n_700), .Y(n_707) );
NOR2x1_ASAP7_75t_L g708 ( .A(n_705), .B(n_698), .Y(n_708) );
OR2x2_ASAP7_75t_L g709 ( .A(n_706), .B(n_704), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_707), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_709), .Y(n_711) );
OAI22x1_ASAP7_75t_L g712 ( .A1(n_711), .A2(n_710), .B1(n_708), .B2(n_703), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g713 ( .A1(n_712), .A2(n_530), .B1(n_463), .B2(n_466), .C(n_474), .Y(n_713) );
AOI21xp33_ASAP7_75t_L g714 ( .A1(n_713), .A2(n_461), .B(n_463), .Y(n_714) );
AO21x2_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_461), .B(n_463), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_466), .B1(n_474), .B2(n_498), .Y(n_716) );
endmodule