module fake_jpeg_641_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

BUFx3_ASAP7_75t_L g10 ( 
.A(n_1),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

INVx2_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_3),
.B(n_2),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_5),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_14),
.B(n_0),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_17),
.B(n_8),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_18),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_SL g19 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_19)
);

OAI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_19),
.A2(n_24),
.B1(n_11),
.B2(n_13),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_6),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_20),
.B(n_22),
.Y(n_27)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_21),
.B(n_23),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_12),
.A2(n_7),
.B1(n_2),
.B2(n_3),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_30),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_22),
.B(n_12),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_29),
.B(n_32),
.C(n_18),
.Y(n_38)
);

AOI21xp33_ASAP7_75t_L g30 ( 
.A1(n_17),
.A2(n_20),
.B(n_23),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_31),
.A2(n_11),
.B1(n_19),
.B2(n_10),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_24),
.B(n_15),
.Y(n_32)
);

AND2x6_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_1),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_33),
.B(n_21),
.C(n_18),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g43 ( 
.A1(n_34),
.A2(n_35),
.B1(n_25),
.B2(n_28),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_32),
.A2(n_23),
.B1(n_13),
.B2(n_18),
.Y(n_35)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_38),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_39),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_40),
.B(n_41),
.C(n_38),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_18),
.C(n_21),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_27),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_46),
.C(n_33),
.Y(n_49)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_25),
.C(n_27),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_44),
.B(n_46),
.C(n_42),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_51),
.B(n_44),
.Y(n_54)
);

AOI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_46),
.B(n_42),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_52),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_L g56 ( 
.A1(n_54),
.A2(n_45),
.A3(n_47),
.B1(n_43),
.B2(n_48),
.C1(n_1),
.C2(n_4),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g57 ( 
.A1(n_56),
.A2(n_45),
.A3(n_53),
.B1(n_4),
.B2(n_5),
.C1(n_2),
.C2(n_3),
.Y(n_57)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_55),
.A3(n_45),
.B1(n_53),
.B2(n_4),
.C1(n_5),
.C2(n_3),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_55),
.C(n_5),
.Y(n_59)
);


endmodule