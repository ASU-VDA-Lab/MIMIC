module real_jpeg_25827_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx3_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_3),
.A2(n_42),
.B1(n_44),
.B2(n_49),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_3),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_3),
.A2(n_49),
.B1(n_52),
.B2(n_66),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_3),
.A2(n_22),
.B1(n_26),
.B2(n_49),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_3),
.A2(n_28),
.B1(n_29),
.B2(n_49),
.Y(n_131)
);

BUFx10_ASAP7_75t_L g59 ( 
.A(n_4),
.Y(n_59)
);

OAI22xp33_ASAP7_75t_SL g139 ( 
.A1(n_5),
.A2(n_53),
.B1(n_77),
.B2(n_140),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_5),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_5),
.A2(n_42),
.B1(n_44),
.B2(n_140),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_5),
.A2(n_22),
.B1(n_26),
.B2(n_140),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_5),
.A2(n_28),
.B1(n_29),
.B2(n_140),
.Y(n_255)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

INVx13_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_8),
.A2(n_52),
.B1(n_54),
.B2(n_55),
.Y(n_51)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_8),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_8),
.A2(n_42),
.B1(n_44),
.B2(n_54),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_54),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_8),
.A2(n_28),
.B1(n_29),
.B2(n_54),
.Y(n_165)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g32 ( 
.A1(n_10),
.A2(n_22),
.B1(n_26),
.B2(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_10),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g41 ( 
.A1(n_10),
.A2(n_33),
.B1(n_42),
.B2(n_44),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_10),
.A2(n_33),
.B1(n_53),
.B2(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_10),
.A2(n_28),
.B1(n_29),
.B2(n_33),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_10),
.A2(n_59),
.B(n_202),
.C(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_10),
.B(n_57),
.Y(n_215)
);

O2A1O1Ixp33_ASAP7_75t_L g225 ( 
.A1(n_10),
.A2(n_37),
.B(n_44),
.C(n_226),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_10),
.B(n_25),
.C(n_28),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_10),
.B(n_87),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_10),
.B(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_10),
.B(n_27),
.Y(n_272)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_11),
.Y(n_108)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_11),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_11),
.B(n_255),
.Y(n_260)
);

INVx6_ASAP7_75t_L g268 ( 
.A(n_11),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_80),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_78),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_73),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_73),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_67),
.C(n_68),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_16),
.A2(n_17),
.B1(n_316),
.B2(n_317),
.Y(n_315)
);

CKINVDCx14_ASAP7_75t_R g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_34),
.C(n_50),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_18),
.A2(n_97),
.B1(n_98),
.B2(n_101),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_18),
.A2(n_34),
.B1(n_101),
.B2(n_148),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_18),
.A2(n_101),
.B1(n_186),
.B2(n_211),
.Y(n_210)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_30),
.B(n_31),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_19),
.A2(n_112),
.B(n_113),
.Y(n_111)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_20),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_20),
.B(n_32),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_20),
.B(n_230),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx8_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g36 ( 
.A1(n_22),
.A2(n_26),
.B1(n_37),
.B2(n_39),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_22),
.B(n_243),
.Y(n_242)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g226 ( 
.A1(n_26),
.A2(n_33),
.B(n_39),
.Y(n_226)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_27),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_27),
.B(n_92),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_27),
.B(n_230),
.Y(n_240)
);

INVx1_ASAP7_75t_SL g29 ( 
.A(n_28),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_28),
.B(n_266),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_30),
.B(n_31),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g132 ( 
.A1(n_30),
.A2(n_91),
.B(n_112),
.Y(n_132)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_33),
.A2(n_44),
.B(n_58),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g148 ( 
.A(n_34),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_35),
.B(n_45),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_35),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_40),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g67 ( 
.A1(n_36),
.A2(n_40),
.B(n_46),
.Y(n_67)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_36),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_36),
.B(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_37),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_37),
.A2(n_39),
.B1(n_42),
.B2(n_44),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_41),
.B(n_99),
.Y(n_135)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_42),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g57 ( 
.A1(n_42),
.A2(n_44),
.B1(n_58),
.B2(n_59),
.Y(n_57)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_45),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_46),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_50),
.B(n_147),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_57),
.B(n_60),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_51),
.Y(n_71)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_53),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_53),
.A2(n_58),
.B1(n_59),
.B2(n_64),
.Y(n_63)
);

INVx8_ASAP7_75t_L g64 ( 
.A(n_53),
.Y(n_64)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_57),
.B(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_57),
.B(n_65),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_76),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_57),
.B(n_139),
.Y(n_172)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_60),
.B(n_74),
.Y(n_73)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_61),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_62),
.B(n_76),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_62),
.B(n_139),
.Y(n_138)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_64),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_67),
.B(n_162),
.C(n_171),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_67),
.A2(n_171),
.B1(n_301),
.B2(n_302),
.Y(n_300)
);

CKINVDCx14_ASAP7_75t_R g301 ( 
.A(n_67),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g316 ( 
.A1(n_67),
.A2(n_68),
.B1(n_69),
.B2(n_301),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_71),
.B(n_72),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_116),
.B(n_117),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_72),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_72),
.B(n_138),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_75),
.B(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_77),
.Y(n_203)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_314),
.B(n_319),
.Y(n_80)
);

OAI211xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_141),
.B(n_151),
.C(n_313),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_118),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_83),
.B(n_118),
.Y(n_152)
);

BUFx24_ASAP7_75t_SL g320 ( 
.A(n_83),
.Y(n_320)
);

FAx1_ASAP7_75t_SL g83 ( 
.A(n_84),
.B(n_93),
.CI(n_104),
.CON(n_83),
.SN(n_83)
);

OAI21xp5_ASAP7_75t_SL g123 ( 
.A1(n_84),
.A2(n_85),
.B(n_88),
.Y(n_123)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_84),
.B(n_93),
.C(n_104),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_87),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_89),
.B(n_228),
.Y(n_227)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_91),
.B(n_240),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_94),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_94),
.A2(n_102),
.B1(n_146),
.B2(n_149),
.Y(n_145)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_94),
.B(n_98),
.C(n_101),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_94),
.B(n_146),
.C(n_150),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_95),
.B(n_172),
.Y(n_185)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_100),
.B(n_195),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_184),
.C(n_186),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_110),
.B(n_114),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_105),
.B(n_111),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_105),
.A2(n_114),
.B1(n_115),
.B2(n_122),
.Y(n_121)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_105),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_111),
.B1(n_122),
.B2(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_105),
.B(n_225),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_105),
.A2(n_122),
.B1(n_225),
.B2(n_284),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_108),
.B(n_109),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g130 ( 
.A(n_106),
.B(n_131),
.Y(n_130)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_106),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_106),
.B(n_109),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_106),
.B(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_107),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_121),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_111),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_113),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_113),
.B(n_229),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_119),
.B(n_123),
.C(n_124),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_123),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_124),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_133),
.C(n_136),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_125),
.B(n_157),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_132),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_126),
.B(n_132),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_130),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_127),
.B(n_252),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_129),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_130),
.A2(n_165),
.B(n_168),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_130),
.B(n_260),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_131),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_133),
.A2(n_136),
.B1(n_137),
.B2(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_133),
.Y(n_158)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_135),
.B(n_188),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND3xp33_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_152),
.C(n_153),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_144),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_143),
.B(n_144),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_150),
.Y(n_144)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_146),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_176),
.B(n_312),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_173),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_155),
.B(n_173),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_159),
.C(n_161),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_156),
.B(n_159),
.Y(n_310)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_161),
.B(n_310),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_162),
.A2(n_163),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_169),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_169),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_167),
.B(n_217),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_167),
.B(n_253),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_170),
.B(n_240),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g302 ( 
.A(n_171),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_307),
.B(n_311),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_218),
.B(n_293),
.C(n_306),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_206),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_179),
.B(n_206),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_192),
.B2(n_205),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_191),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_182),
.B(n_191),
.C(n_205),
.Y(n_294)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_184),
.A2(n_185),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_192),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_194),
.B(n_199),
.C(n_200),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_204),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_201),
.B(n_204),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_212),
.C(n_213),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_207),
.A2(n_208),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g233 ( 
.A(n_212),
.B(n_213),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_215),
.C(n_216),
.Y(n_213)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_223),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_216),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_217),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_292),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_220),
.A2(n_234),
.B(n_291),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_231),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_221),
.B(n_231),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_222),
.B(n_224),
.C(n_227),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_222),
.B(n_289),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g289 ( 
.A(n_224),
.B(n_227),
.Y(n_289)
);

CKINVDCx14_ASAP7_75t_R g284 ( 
.A(n_225),
.Y(n_284)
);

INVxp33_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_286),
.B(n_290),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_236),
.A2(n_277),
.B(n_285),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_257),
.B(n_276),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_244),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_244),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_239),
.B(n_241),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_239),
.A2(n_241),
.B1(n_242),
.B2(n_262),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_239),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_256),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_247),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_247),
.B(n_250),
.C(n_256),
.Y(n_278)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_248),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_251),
.Y(n_256)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

INVxp33_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_258),
.A2(n_263),
.B(n_275),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_259),
.B(n_261),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_261),
.Y(n_275)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_260),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_271),
.B(n_274),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVx5_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_SL g274 ( 
.A(n_272),
.B(n_273),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_278),
.B(n_279),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_283),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_281),
.B(n_282),
.C(n_283),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g290 ( 
.A(n_287),
.B(n_288),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_295),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_294),
.B(n_295),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_305),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_303),
.B2(n_304),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_297),
.B(n_304),
.C(n_305),
.Y(n_308)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_300),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g303 ( 
.A(n_304),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_308),
.B(n_309),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_318),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g319 ( 
.A(n_315),
.B(n_318),
.Y(n_319)
);

CKINVDCx14_ASAP7_75t_R g317 ( 
.A(n_316),
.Y(n_317)
);


endmodule