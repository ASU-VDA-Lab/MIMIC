module fake_jpeg_21263_n_14 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_14);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_14;

wire n_13;
wire n_11;
wire n_10;
wire n_12;
wire n_8;
wire n_9;

NAND2xp33_ASAP7_75t_SL g8 ( 
.A(n_5),
.B(n_1),
.Y(n_8)
);

INVx6_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

AOI22xp5_ASAP7_75t_L g10 ( 
.A1(n_9),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_10)
);

AOI21xp5_ASAP7_75t_L g12 ( 
.A1(n_10),
.A2(n_11),
.B(n_0),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g11 ( 
.A(n_9),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_12),
.B(n_3),
.Y(n_13)
);

AOI322xp5_ASAP7_75t_L g14 ( 
.A1(n_13),
.A2(n_4),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.C1(n_9),
.C2(n_12),
.Y(n_14)
);


endmodule