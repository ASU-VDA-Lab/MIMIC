module real_jpeg_10248_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_332, n_7, n_331, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_332;
input n_7;
input n_331;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_176;
wire n_323;
wire n_166;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx24_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_24),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_1),
.A2(n_33),
.B1(n_58),
.B2(n_59),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_1),
.A2(n_33),
.B1(n_43),
.B2(n_45),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_1),
.A2(n_29),
.B1(n_30),
.B2(n_33),
.Y(n_279)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_3),
.A2(n_24),
.B1(n_32),
.B2(n_35),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g76 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_3),
.A2(n_35),
.B1(n_58),
.B2(n_59),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_3),
.A2(n_35),
.B1(n_43),
.B2(n_45),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g116 ( 
.A1(n_4),
.A2(n_45),
.B(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_4),
.B(n_45),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_4),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_4),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_4),
.B(n_89),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_4),
.A2(n_26),
.B(n_30),
.Y(n_203)
);

OAI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_4),
.A2(n_24),
.B1(n_32),
.B2(n_128),
.Y(n_221)
);

BUFx10_ASAP7_75t_L g109 ( 
.A(n_5),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_6),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g55 ( 
.A1(n_7),
.A2(n_45),
.B(n_56),
.C(n_57),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_7),
.B(n_45),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_7),
.A2(n_58),
.B1(n_59),
.B2(n_61),
.Y(n_57)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_7),
.Y(n_61)
);

BUFx6f_ASAP7_75t_SL g42 ( 
.A(n_8),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_10),
.A2(n_29),
.B1(n_30),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_10),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g63 ( 
.A1(n_10),
.A2(n_43),
.B1(n_45),
.B2(n_47),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_10),
.A2(n_47),
.B1(n_58),
.B2(n_59),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_10),
.A2(n_24),
.B1(n_32),
.B2(n_47),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_11),
.A2(n_29),
.B1(n_30),
.B2(n_53),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_11),
.Y(n_53)
);

OAI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_11),
.A2(n_24),
.B1(n_32),
.B2(n_53),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g167 ( 
.A1(n_11),
.A2(n_53),
.B1(n_58),
.B2(n_59),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_11),
.A2(n_43),
.B1(n_45),
.B2(n_53),
.Y(n_216)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_43),
.B1(n_45),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_13),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g130 ( 
.A1(n_13),
.A2(n_58),
.B1(n_59),
.B2(n_119),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_119),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g223 ( 
.A1(n_13),
.A2(n_24),
.B1(n_32),
.B2(n_119),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_14),
.A2(n_58),
.B1(n_59),
.B2(n_107),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g107 ( 
.A(n_14),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_14),
.A2(n_43),
.B1(n_45),
.B2(n_107),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_107),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_14),
.A2(n_24),
.B1(n_32),
.B2(n_107),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_15),
.A2(n_58),
.B1(n_59),
.B2(n_112),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_15),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_15),
.A2(n_43),
.B1(n_45),
.B2(n_112),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_112),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_15),
.A2(n_24),
.B1(n_32),
.B2(n_112),
.Y(n_251)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_95),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_SL g17 ( 
.A(n_18),
.B(n_93),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_80),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_19),
.B(n_80),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_67),
.C(n_71),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_20),
.A2(n_21),
.B1(n_67),
.B2(n_316),
.Y(n_322)
);

CKINVDCx14_ASAP7_75t_R g20 ( 
.A(n_21),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_36),
.B1(n_37),
.B2(n_66),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_22),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_SL g22 ( 
.A1(n_23),
.A2(n_28),
.B1(n_31),
.B2(n_34),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_23),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_23),
.A2(n_28),
.B1(n_223),
.B2(n_232),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_23),
.A2(n_28),
.B1(n_232),
.B2(n_251),
.Y(n_250)
);

OAI21xp5_ASAP7_75t_SL g275 ( 
.A1(n_23),
.A2(n_251),
.B(n_276),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g296 ( 
.A1(n_23),
.A2(n_88),
.B(n_297),
.Y(n_296)
);

A2O1A1Ixp33_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_24),
.B(n_25),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_24),
.Y(n_32)
);

A2O1A1Ixp33_ASAP7_75t_L g202 ( 
.A1(n_24),
.A2(n_25),
.B(n_128),
.C(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_25),
.A2(n_26),
.B1(n_29),
.B2(n_30),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g67 ( 
.A1(n_28),
.A2(n_31),
.B(n_68),
.Y(n_67)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_28),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_30),
.Y(n_29)
);

O2A1O1Ixp33_ASAP7_75t_L g49 ( 
.A1(n_30),
.A2(n_40),
.B(n_41),
.C(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_30),
.B(n_41),
.Y(n_50)
);

HAxp5_ASAP7_75t_SL g157 ( 
.A(n_30),
.B(n_128),
.CON(n_157),
.SN(n_157)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_34),
.Y(n_86)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g37 ( 
.A1(n_38),
.A2(n_54),
.B1(n_64),
.B2(n_65),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_48),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_39),
.A2(n_74),
.B(n_219),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_40),
.B(n_46),
.Y(n_39)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_40),
.Y(n_79)
);

OAI21xp5_ASAP7_75t_L g83 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_83)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_40),
.A2(n_49),
.B1(n_157),
.B2(n_158),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_40),
.A2(n_49),
.B1(n_76),
.B2(n_302),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_41),
.A2(n_42),
.B1(n_43),
.B2(n_45),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_41),
.B(n_45),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_42),
.Y(n_41)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_43),
.A2(n_50),
.B1(n_157),
.B2(n_163),
.Y(n_162)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_46),
.A2(n_49),
.B(n_78),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g278 ( 
.A1(n_48),
.A2(n_79),
.B(n_279),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_49),
.B(n_51),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g74 ( 
.A(n_49),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_52),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_52),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_54),
.B(n_64),
.C(n_66),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_54),
.A2(n_65),
.B1(n_72),
.B2(n_73),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_55),
.A2(n_57),
.B(n_62),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_55),
.A2(n_57),
.B1(n_116),
.B2(n_118),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_55),
.A2(n_57),
.B1(n_118),
.B2(n_145),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_55),
.A2(n_57),
.B1(n_145),
.B2(n_155),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_55),
.A2(n_155),
.B(n_191),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g214 ( 
.A(n_55),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g256 ( 
.A1(n_55),
.A2(n_57),
.B1(n_238),
.B2(n_257),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_SL g285 ( 
.A1(n_55),
.A2(n_257),
.B(n_286),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_56),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g127 ( 
.A(n_57),
.B(n_128),
.Y(n_127)
);

INVxp67_ASAP7_75t_L g192 ( 
.A(n_57),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_57),
.B(n_216),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_57),
.A2(n_238),
.B(n_239),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_58),
.B(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_58),
.B(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_58),
.B(n_136),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_59),
.A2(n_121),
.B1(n_122),
.B2(n_123),
.Y(n_120)
);

BUFx24_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_63),
.B(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_63),
.A2(n_214),
.B(n_215),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_65),
.B(n_67),
.C(n_72),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_67),
.A2(n_316),
.B1(n_317),
.B2(n_318),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_67),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_69),
.B(n_89),
.Y(n_88)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_70),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_70),
.A2(n_89),
.B1(n_221),
.B2(n_222),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g321 ( 
.A(n_71),
.B(n_322),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B(n_77),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_74),
.A2(n_79),
.B1(n_176),
.B2(n_177),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_74),
.A2(n_79),
.B1(n_177),
.B2(n_219),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_76),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_78),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_79),
.B(n_128),
.Y(n_143)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_82),
.A2(n_83),
.B1(n_84),
.B2(n_85),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_83),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_85),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_89),
.B(n_277),
.Y(n_276)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_91),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

OAI321xp33_ASAP7_75t_L g95 ( 
.A1(n_96),
.A2(n_313),
.A3(n_323),
.B1(n_328),
.B2(n_329),
.C(n_331),
.Y(n_95)
);

AOI321xp33_ASAP7_75t_L g96 ( 
.A1(n_97),
.A2(n_265),
.A3(n_289),
.B1(n_306),
.B2(n_312),
.C(n_332),
.Y(n_96)
);

NOR3xp33_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_225),
.C(n_261),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_196),
.B(n_224),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_170),
.B(n_195),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_150),
.B(n_169),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g101 ( 
.A1(n_102),
.A2(n_139),
.B(n_149),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_103),
.A2(n_125),
.B(n_138),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_113),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_104),
.B(n_113),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_108),
.B1(n_109),
.B2(n_110),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_106),
.A2(n_130),
.B1(n_131),
.B2(n_132),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_108),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_108),
.B(n_167),
.Y(n_182)
);

CKINVDCx16_ASAP7_75t_R g132 ( 
.A(n_109),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_109),
.B(n_148),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_109),
.B(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_111),
.Y(n_110)
);

OAI21xp5_ASAP7_75t_SL g146 ( 
.A1(n_111),
.A2(n_131),
.B(n_147),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_114),
.A2(n_115),
.B1(n_120),
.B2(n_124),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_114),
.B(n_124),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_115),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_117),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_120),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g125 ( 
.A1(n_126),
.A2(n_133),
.B(n_137),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_127),
.B(n_129),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_128),
.B(n_132),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_131),
.A2(n_165),
.B(n_166),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_131),
.A2(n_132),
.B1(n_181),
.B2(n_206),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_131),
.A2(n_166),
.B(n_206),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g284 ( 
.A1(n_131),
.A2(n_132),
.B(n_165),
.Y(n_284)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_132),
.A2(n_181),
.B(n_182),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_135),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_140),
.B(n_141),
.Y(n_149)
);

CKINVDCx5p33_ASAP7_75t_R g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_142),
.B(n_151),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g169 ( 
.A(n_142),
.B(n_151),
.Y(n_169)
);

FAx1_ASAP7_75t_SL g142 ( 
.A(n_143),
.B(n_144),
.CI(n_146),
.CON(n_142),
.SN(n_142)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_147),
.B(n_182),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_148),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_152),
.A2(n_153),
.B1(n_161),
.B2(n_168),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_153),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_154),
.A2(n_156),
.B1(n_159),
.B2(n_160),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_154),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_156),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_160),
.C(n_168),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_158),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_161),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_164),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_171),
.B(n_172),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_174),
.B1(n_187),
.B2(n_188),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_173),
.B(n_190),
.C(n_193),
.Y(n_197)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_178),
.B1(n_179),
.B2(n_186),
.Y(n_174)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_175),
.Y(n_186)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_183),
.B1(n_184),
.B2(n_185),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_180),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_184),
.C(n_186),
.Y(n_207)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_193),
.B2(n_194),
.Y(n_188)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_189),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_190),
.Y(n_194)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_191),
.B(n_239),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_198),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_197),
.B(n_198),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_210),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_207),
.B1(n_208),
.B2(n_209),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_200),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_200),
.B(n_209),
.C(n_210),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_204),
.B2(n_205),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_205),
.Y(n_228)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_207),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_220),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_213),
.B1(n_217),
.B2(n_218),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_213),
.B(n_217),
.C(n_220),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_214),
.B(n_240),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_215),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_216),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_218),
.Y(n_217)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_225),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_244),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_244),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_227),
.B(n_235),
.C(n_242),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_227),
.B(n_264),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_228),
.B(n_229),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_228),
.B(n_230),
.C(n_234),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_234),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_233),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_236),
.B1(n_242),
.B2(n_243),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_241),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_241),
.Y(n_247)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_244)
);

CKINVDCx14_ASAP7_75t_R g260 ( 
.A(n_245),
.Y(n_260)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_254),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_246),
.B(n_254),
.C(n_258),
.Y(n_267)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_248),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_247),
.B(n_249),
.C(n_253),
.Y(n_288)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_252),
.B2(n_253),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_256),
.Y(n_272)
);

CKINVDCx14_ASAP7_75t_R g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_262),
.B(n_263),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g309 ( 
.A(n_262),
.B(n_263),
.Y(n_309)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g306 ( 
.A1(n_266),
.A2(n_307),
.B(n_311),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_267),
.B(n_268),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_288),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g269 ( 
.A1(n_270),
.A2(n_271),
.B1(n_281),
.B2(n_282),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_282),
.C(n_288),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g270 ( 
.A(n_271),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_272),
.B(n_274),
.C(n_280),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B1(n_278),
.B2(n_280),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_275),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_277),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_278),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_279),
.Y(n_302)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_283),
.A2(n_284),
.B1(n_285),
.B2(n_287),
.Y(n_282)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_283),
.A2(n_284),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g320 ( 
.A1(n_283),
.A2(n_296),
.B(n_299),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_285),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g287 ( 
.A(n_285),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g312 ( 
.A(n_290),
.B(n_291),
.Y(n_312)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_291),
.Y(n_324)
);

FAx1_ASAP7_75t_SL g291 ( 
.A(n_292),
.B(n_300),
.CI(n_305),
.CON(n_291),
.SN(n_291)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_294),
.B1(n_298),
.B2(n_299),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g295 ( 
.A(n_296),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_298),
.Y(n_299)
);

OAI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_303),
.B(n_304),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_303),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_304),
.Y(n_319)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_304),
.A2(n_315),
.B1(n_319),
.B2(n_327),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_308),
.A2(n_309),
.B(n_310),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_321),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_314),
.B(n_321),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_315),
.B(n_319),
.C(n_320),
.Y(n_314)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_315),
.Y(n_327)
);

CKINVDCx16_ASAP7_75t_R g317 ( 
.A(n_318),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g325 ( 
.A(n_320),
.B(n_326),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_324),
.B(n_325),
.Y(n_328)
);


endmodule