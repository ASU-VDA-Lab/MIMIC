module fake_jpeg_1243_n_704 (n_13, n_1, n_10, n_6, n_14, n_19, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_704);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_704;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_696;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_657;
wire n_27;
wire n_664;
wire n_365;
wire n_179;
wire n_620;
wire n_686;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_678;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_699;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_635;
wire n_517;
wire n_629;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_643;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_647;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_641;
wire n_701;
wire n_48;
wire n_465;
wire n_638;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_623;
wire n_579;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_637;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_672;
wire n_309;
wire n_624;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_688;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_596;
wire n_569;
wire n_400;
wire n_646;
wire n_319;
wire n_689;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_663;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_634;
wire n_23;
wire n_69;
wire n_658;
wire n_698;
wire n_195;
wire n_450;
wire n_557;
wire n_681;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_666;
wire n_639;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_645;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_694;
wire n_692;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_622;
wire n_463;
wire n_667;
wire n_92;
wire n_332;
wire n_640;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_653;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_626;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_668;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_682;
wire n_305;
wire n_161;
wire n_441;
wire n_697;
wire n_555;
wire n_342;
wire n_642;
wire n_101;
wire n_226;
wire n_509;
wire n_644;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_656;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_649;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_679;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_691;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_615;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_662;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_676;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_648;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_670;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_683;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_631;
wire n_433;
wire n_636;
wire n_690;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_650;
wire n_218;
wire n_63;
wire n_652;
wire n_599;
wire n_239;
wire n_693;
wire n_674;
wire n_243;
wire n_481;
wire n_628;
wire n_619;
wire n_348;
wire n_587;
wire n_703;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_655;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_684;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_680;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_625;
wire n_147;
wire n_449;
wire n_627;
wire n_695;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_702;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_618;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_659;
wire n_125;
wire n_661;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_687;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_673;
wire n_58;
wire n_41;
wire n_613;
wire n_630;
wire n_266;
wire n_548;
wire n_665;
wire n_72;
wire n_512;
wire n_654;
wire n_445;
wire n_443;
wire n_677;
wire n_617;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_700;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_671;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_669;
wire n_524;
wire n_402;
wire n_563;
wire n_685;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_660;
wire n_373;
wire n_633;
wire n_112;
wire n_632;
wire n_616;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_651;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_675;
wire n_335;
wire n_120;
wire n_621;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_5),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_18),
.Y(n_32)
);

INVx11_ASAP7_75t_SL g33 ( 
.A(n_18),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_17),
.Y(n_34)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_6),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_12),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

INVx13_ASAP7_75t_L g42 ( 
.A(n_14),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_11),
.Y(n_48)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_8),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_15),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_9),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_2),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_13),
.Y(n_56)
);

INVxp67_ASAP7_75t_L g57 ( 
.A(n_7),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_19),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx11_ASAP7_75t_SL g60 ( 
.A(n_17),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_61),
.Y(n_142)
);

INVx6_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx4_ASAP7_75t_SL g205 ( 
.A(n_63),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_11),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_64),
.B(n_103),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_22),
.B(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_65),
.B(n_68),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_39),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_67),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_57),
.B(n_30),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_44),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_70),
.Y(n_195)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_SL g158 ( 
.A(n_71),
.Y(n_158)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_29),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g215 ( 
.A(n_72),
.Y(n_215)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_73),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_74),
.Y(n_147)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_75),
.Y(n_164)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_76),
.Y(n_136)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_77),
.Y(n_198)
);

INVx13_ASAP7_75t_L g78 ( 
.A(n_33),
.Y(n_78)
);

INVx13_ASAP7_75t_L g196 ( 
.A(n_78),
.Y(n_196)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g206 ( 
.A(n_79),
.Y(n_206)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_80),
.B(n_89),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_26),
.B(n_10),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_81),
.B(n_83),
.Y(n_151)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_20),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_26),
.B(n_10),
.Y(n_83)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_44),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g212 ( 
.A(n_84),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_85),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_38),
.Y(n_86)
);

INVx6_ASAP7_75t_L g144 ( 
.A(n_86),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_38),
.Y(n_87)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_87),
.Y(n_154)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_30),
.Y(n_88)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_88),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_60),
.Y(n_89)
);

INVx8_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_90),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_47),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_91),
.Y(n_188)
);

INVx6_ASAP7_75t_L g92 ( 
.A(n_38),
.Y(n_92)
);

INVx8_ASAP7_75t_L g146 ( 
.A(n_92),
.Y(n_146)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_93),
.Y(n_216)
);

BUFx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_94),
.Y(n_180)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_24),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_95),
.B(n_101),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_43),
.Y(n_97)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_97),
.Y(n_145)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx6_ASAP7_75t_L g193 ( 
.A(n_98),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_24),
.Y(n_99)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_20),
.Y(n_100)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_100),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_21),
.B(n_10),
.Y(n_101)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_29),
.Y(n_102)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_102),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_21),
.B(n_12),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_20),
.Y(n_104)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_104),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_23),
.Y(n_105)
);

INVx6_ASAP7_75t_L g221 ( 
.A(n_105),
.Y(n_221)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_106),
.Y(n_171)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx8_ASAP7_75t_L g169 ( 
.A(n_107),
.Y(n_169)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_108),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_23),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g189 ( 
.A(n_109),
.Y(n_189)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_43),
.Y(n_110)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_110),
.Y(n_156)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_111),
.Y(n_170)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_27),
.Y(n_112)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_27),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g225 ( 
.A(n_113),
.Y(n_225)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_41),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g173 ( 
.A(n_114),
.Y(n_173)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_49),
.Y(n_115)
);

INVx4_ASAP7_75t_L g200 ( 
.A(n_115),
.Y(n_200)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_46),
.Y(n_116)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_116),
.Y(n_191)
);

INVx13_ASAP7_75t_L g117 ( 
.A(n_42),
.Y(n_117)
);

BUFx24_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_27),
.Y(n_118)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_118),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_27),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g227 ( 
.A(n_119),
.Y(n_227)
);

BUFx16f_ASAP7_75t_L g120 ( 
.A(n_42),
.Y(n_120)
);

BUFx5_ASAP7_75t_L g137 ( 
.A(n_120),
.Y(n_137)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_50),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_121),
.B(n_131),
.Y(n_175)
);

BUFx24_ASAP7_75t_L g122 ( 
.A(n_42),
.Y(n_122)
);

INVx11_ASAP7_75t_L g222 ( 
.A(n_122),
.Y(n_222)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_41),
.Y(n_123)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_123),
.Y(n_192)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_27),
.Y(n_124)
);

INVx3_ASAP7_75t_L g229 ( 
.A(n_124),
.Y(n_229)
);

INVx11_ASAP7_75t_L g125 ( 
.A(n_35),
.Y(n_125)
);

INVx4_ASAP7_75t_L g211 ( 
.A(n_125),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_35),
.Y(n_126)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_126),
.Y(n_184)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_35),
.Y(n_127)
);

INVx5_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

INVx11_ASAP7_75t_L g128 ( 
.A(n_35),
.Y(n_128)
);

INVx4_ASAP7_75t_L g217 ( 
.A(n_128),
.Y(n_217)
);

INVx6_ASAP7_75t_L g129 ( 
.A(n_35),
.Y(n_129)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_58),
.B(n_12),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_130),
.B(n_19),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_50),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_52),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_132),
.B(n_37),
.Y(n_187)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_56),
.Y(n_133)
);

INVx2_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_71),
.B(n_75),
.C(n_108),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_134),
.B(n_122),
.C(n_78),
.Y(n_267)
);

BUFx5_ASAP7_75t_L g148 ( 
.A(n_120),
.Y(n_148)
);

INVx4_ASAP7_75t_L g238 ( 
.A(n_148),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_106),
.B(n_56),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_SL g244 ( 
.A(n_149),
.B(n_157),
.Y(n_244)
);

AOI22xp33_ASAP7_75t_SL g155 ( 
.A1(n_72),
.A2(n_32),
.B1(n_54),
.B2(n_58),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_155),
.A2(n_32),
.B1(n_45),
.B2(n_48),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g157 ( 
.A(n_94),
.Y(n_157)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_92),
.Y(n_160)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_160),
.Y(n_230)
);

OR2x2_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_54),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_161),
.B(n_182),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_129),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_163),
.B(n_194),
.Y(n_257)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_62),
.Y(n_167)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_167),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_168),
.B(n_178),
.Y(n_259)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_67),
.Y(n_176)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_118),
.B(n_55),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_84),
.Y(n_179)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_179),
.Y(n_254)
);

OR2x2_ASAP7_75t_L g182 ( 
.A(n_124),
.B(n_36),
.Y(n_182)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_98),
.Y(n_185)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_185),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_187),
.B(n_190),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_91),
.B(n_36),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_82),
.B(n_55),
.Y(n_194)
);

INVx5_ASAP7_75t_L g202 ( 
.A(n_123),
.Y(n_202)
);

INVx4_ASAP7_75t_L g278 ( 
.A(n_202),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_86),
.B(n_34),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_203),
.B(n_207),
.Y(n_289)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_204),
.B(n_224),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_87),
.B(n_34),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_96),
.B(n_31),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_208),
.B(n_213),
.Y(n_292)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_104),
.Y(n_210)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_210),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_61),
.B(n_31),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_66),
.A2(n_37),
.B1(n_28),
.B2(n_25),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_214),
.A2(n_53),
.B1(n_51),
.B2(n_49),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_70),
.A2(n_45),
.B1(n_28),
.B2(n_25),
.Y(n_218)
);

NAND2x1_ASAP7_75t_L g312 ( 
.A(n_218),
.B(n_7),
.Y(n_312)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_93),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g251 ( 
.A(n_219),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_105),
.Y(n_224)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_107),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_226),
.B(n_126),
.Y(n_241)
);

INVx4_ASAP7_75t_L g228 ( 
.A(n_125),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_228),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_231),
.Y(n_338)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_138),
.Y(n_232)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_232),
.Y(n_371)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_141),
.Y(n_233)
);

INVx2_ASAP7_75t_SL g339 ( 
.A(n_233),
.Y(n_339)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_215),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_234),
.Y(n_348)
);

BUFx6f_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

INVx5_ASAP7_75t_L g325 ( 
.A(n_235),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g236 ( 
.A1(n_200),
.A2(n_32),
.B1(n_123),
.B2(n_114),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g326 ( 
.A1(n_236),
.A2(n_237),
.B1(n_245),
.B2(n_264),
.Y(n_326)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_149),
.A2(n_128),
.B1(n_100),
.B2(n_90),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g239 ( 
.A(n_223),
.Y(n_239)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_239),
.Y(n_336)
);

NAND2x1p5_ASAP7_75t_L g240 ( 
.A(n_159),
.B(n_127),
.Y(n_240)
);

AO21x1_ASAP7_75t_L g340 ( 
.A1(n_240),
.A2(n_247),
.B(n_312),
.Y(n_340)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_241),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_139),
.B(n_48),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_242),
.B(n_246),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_173),
.A2(n_119),
.B1(n_113),
.B2(n_109),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_139),
.B(n_79),
.Y(n_246)
);

OR2x2_ASAP7_75t_SL g247 ( 
.A(n_151),
.B(n_117),
.Y(n_247)
);

CKINVDCx12_ASAP7_75t_R g248 ( 
.A(n_223),
.Y(n_248)
);

INVx13_ASAP7_75t_L g361 ( 
.A(n_248),
.Y(n_361)
);

INVx6_ASAP7_75t_L g250 ( 
.A(n_142),
.Y(n_250)
);

INVx3_ASAP7_75t_SL g318 ( 
.A(n_250),
.Y(n_318)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_145),
.Y(n_252)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_156),
.B(n_53),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_253),
.B(n_274),
.C(n_276),
.Y(n_323)
);

BUFx12f_ASAP7_75t_L g256 ( 
.A(n_137),
.Y(n_256)
);

INVx4_ASAP7_75t_L g337 ( 
.A(n_256),
.Y(n_337)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_165),
.Y(n_258)
);

INVx3_ASAP7_75t_SL g358 ( 
.A(n_258),
.Y(n_358)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_170),
.Y(n_260)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_260),
.Y(n_327)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_158),
.Y(n_262)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_262),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g264 ( 
.A1(n_153),
.A2(n_85),
.B1(n_29),
.B2(n_122),
.Y(n_264)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_150),
.Y(n_265)
);

INVx4_ASAP7_75t_L g347 ( 
.A(n_265),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g266 ( 
.A(n_165),
.Y(n_266)
);

INVx3_ASAP7_75t_L g335 ( 
.A(n_266),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_267),
.B(n_300),
.Y(n_328)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_158),
.Y(n_268)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g269 ( 
.A1(n_215),
.A2(n_53),
.B1(n_51),
.B2(n_49),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g353 ( 
.A1(n_269),
.A2(n_284),
.B1(n_299),
.B2(n_303),
.Y(n_353)
);

BUFx2_ASAP7_75t_L g270 ( 
.A(n_166),
.Y(n_270)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_270),
.Y(n_330)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_271),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_272),
.A2(n_269),
.B1(n_264),
.B2(n_155),
.Y(n_313)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_175),
.Y(n_273)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_273),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_151),
.B(n_51),
.Y(n_274)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_152),
.Y(n_275)
);

INVx2_ASAP7_75t_L g331 ( 
.A(n_275),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_172),
.B(n_175),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_172),
.B(n_9),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_279),
.B(n_285),
.Y(n_354)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_135),
.B(n_9),
.C(n_18),
.Y(n_281)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_281),
.B(n_166),
.Y(n_332)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_195),
.Y(n_282)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_282),
.Y(n_372)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_147),
.Y(n_283)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_283),
.Y(n_343)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_198),
.A2(n_194),
.B1(n_192),
.B2(n_164),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_187),
.B(n_13),
.Y(n_285)
);

INVx5_ASAP7_75t_L g286 ( 
.A(n_169),
.Y(n_286)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_286),
.Y(n_344)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_222),
.Y(n_287)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_287),
.Y(n_352)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_147),
.Y(n_288)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_288),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_177),
.B(n_13),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_290),
.B(n_298),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_180),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g359 ( 
.A(n_293),
.B(n_296),
.Y(n_359)
);

INVx6_ASAP7_75t_SL g294 ( 
.A(n_196),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_294),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_195),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_295),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_182),
.B(n_19),
.Y(n_296)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_174),
.Y(n_297)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_297),
.Y(n_367)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_161),
.B(n_8),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_206),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_201),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_171),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_306),
.Y(n_320)
);

INVx5_ASAP7_75t_L g302 ( 
.A(n_169),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g360 ( 
.A(n_302),
.B(n_305),
.Y(n_360)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_206),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_188),
.A2(n_8),
.B1(n_18),
.B2(n_2),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_SL g362 ( 
.A1(n_304),
.A2(n_217),
.B1(n_146),
.B2(n_227),
.Y(n_362)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_140),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_136),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_205),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_307),
.B(n_311),
.Y(n_345)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_183),
.Y(n_308)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_308),
.B(n_310),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_199),
.B(n_7),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_309),
.B(n_19),
.Y(n_363)
);

INVx2_ASAP7_75t_L g310 ( 
.A(n_220),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_205),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_L g413 ( 
.A1(n_313),
.A2(n_315),
.B1(n_303),
.B2(n_235),
.Y(n_413)
);

OAI22xp33_ASAP7_75t_SL g315 ( 
.A1(n_289),
.A2(n_162),
.B1(n_186),
.B2(n_212),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_292),
.A2(n_197),
.B1(n_193),
.B2(n_186),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_321),
.A2(n_357),
.B1(n_258),
.B2(n_287),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_253),
.A2(n_212),
.B1(n_162),
.B2(n_146),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_324),
.A2(n_368),
.B1(n_282),
.B2(n_250),
.Y(n_396)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_332),
.B(n_251),
.Y(n_409)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_240),
.A2(n_180),
.B(n_211),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g418 ( 
.A1(n_333),
.A2(n_251),
.B(n_266),
.Y(n_418)
);

OR2x4_ASAP7_75t_L g342 ( 
.A(n_247),
.B(n_196),
.Y(n_342)
);

AO21x1_ASAP7_75t_L g402 ( 
.A1(n_342),
.A2(n_263),
.B(n_239),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_240),
.B(n_274),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_346),
.B(n_349),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_276),
.B(n_229),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g355 ( 
.A1(n_291),
.A2(n_216),
.B1(n_188),
.B2(n_184),
.Y(n_355)
);

OAI22xp33_ASAP7_75t_SL g383 ( 
.A1(n_355),
.A2(n_237),
.B1(n_236),
.B2(n_245),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_257),
.B(n_221),
.Y(n_356)
);

NOR2xp33_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_294),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_231),
.A2(n_193),
.B1(n_197),
.B2(n_144),
.Y(n_357)
);

A2O1A1Ixp33_ASAP7_75t_SL g398 ( 
.A1(n_362),
.A2(n_239),
.B(n_304),
.C(n_256),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g392 ( 
.A(n_363),
.B(n_375),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_259),
.B(n_181),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_364),
.B(n_366),
.Y(n_408)
);

AOI22xp33_ASAP7_75t_SL g365 ( 
.A1(n_267),
.A2(n_227),
.B1(n_225),
.B2(n_189),
.Y(n_365)
);

INVxp67_ASAP7_75t_SL g416 ( 
.A(n_365),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_280),
.B(n_181),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_244),
.A2(n_144),
.B1(n_154),
.B2(n_143),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_281),
.B(n_154),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_369),
.B(n_373),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g373 ( 
.A(n_277),
.B(n_143),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_230),
.B(n_221),
.Y(n_375)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_370),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_376),
.B(n_399),
.Y(n_437)
);

INVx13_ASAP7_75t_L g377 ( 
.A(n_361),
.Y(n_377)
);

BUFx4f_ASAP7_75t_L g430 ( 
.A(n_377),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_378),
.B(n_387),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_323),
.B(n_284),
.C(n_301),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_379),
.B(n_380),
.C(n_424),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_323),
.B(n_254),
.C(n_243),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_339),
.Y(n_381)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_381),
.Y(n_439)
);

INVx2_ASAP7_75t_L g382 ( 
.A(n_339),
.Y(n_382)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_382),
.Y(n_433)
);

AOI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_383),
.A2(n_398),
.B1(n_401),
.B2(n_351),
.Y(n_466)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_333),
.B(n_312),
.Y(n_384)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

INVx6_ASAP7_75t_SL g385 ( 
.A(n_361),
.Y(n_385)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_385),
.Y(n_427)
);

INVx4_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_386),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_316),
.B(n_234),
.Y(n_387)
);

INVx3_ASAP7_75t_L g388 ( 
.A(n_347),
.Y(n_388)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_388),
.Y(n_449)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_345),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_389),
.B(n_390),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g390 ( 
.A(n_370),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_347),
.Y(n_391)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_391),
.Y(n_456)
);

INVx13_ASAP7_75t_L g393 ( 
.A(n_314),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_393),
.Y(n_431)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g458 ( 
.A(n_394),
.Y(n_458)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_342),
.B(n_265),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_395),
.B(n_397),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g453 ( 
.A1(n_396),
.A2(n_423),
.B1(n_321),
.B2(n_381),
.Y(n_453)
);

OR2x2_ASAP7_75t_L g397 ( 
.A(n_340),
.B(n_297),
.Y(n_397)
);

NOR2xp33_ASAP7_75t_L g399 ( 
.A(n_341),
.B(n_374),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_341),
.B(n_249),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_400),
.B(n_414),
.Y(n_441)
);

OAI22xp33_ASAP7_75t_SL g401 ( 
.A1(n_373),
.A2(n_300),
.B1(n_270),
.B2(n_299),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g450 ( 
.A1(n_402),
.A2(n_405),
.B(n_418),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_359),
.B(n_261),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_403),
.B(n_407),
.Y(n_447)
);

XNOR2xp5_ASAP7_75t_SL g404 ( 
.A(n_349),
.B(n_346),
.Y(n_404)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_404),
.B(n_409),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g405 ( 
.A(n_328),
.B(n_255),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g407 ( 
.A(n_366),
.B(n_278),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_354),
.B(n_278),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_411),
.B(n_422),
.Y(n_462)
);

INVx3_ASAP7_75t_L g412 ( 
.A(n_325),
.Y(n_412)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_412),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_413),
.A2(n_368),
.B1(n_358),
.B2(n_318),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_369),
.B(n_302),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_364),
.B(n_286),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_415),
.B(n_417),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_332),
.B(n_295),
.Y(n_417)
);

INVx4_ASAP7_75t_L g419 ( 
.A(n_344),
.Y(n_419)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_419),
.Y(n_459)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_339),
.Y(n_420)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_420),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_340),
.B(n_209),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_421),
.B(n_348),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g422 ( 
.A(n_371),
.B(n_238),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g424 ( 
.A(n_328),
.B(n_238),
.C(n_209),
.Y(n_424)
);

BUFx2_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_425),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g428 ( 
.A1(n_410),
.A2(n_324),
.B1(n_338),
.B2(n_328),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g500 ( 
.A1(n_428),
.A2(n_429),
.B1(n_451),
.B2(n_467),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_410),
.A2(n_338),
.B1(n_326),
.B2(n_353),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_397),
.A2(n_357),
.B(n_337),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g482 ( 
.A1(n_432),
.A2(n_450),
.B(n_461),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g436 ( 
.A(n_409),
.B(n_319),
.C(n_334),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_436),
.B(n_442),
.C(n_443),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_404),
.B(n_334),
.Y(n_442)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_406),
.B(n_319),
.Y(n_443)
);

OAI22xp5_ASAP7_75t_L g501 ( 
.A1(n_444),
.A2(n_453),
.B1(n_454),
.B2(n_466),
.Y(n_501)
);

MAJx2_ASAP7_75t_L g446 ( 
.A(n_406),
.B(n_327),
.C(n_317),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g488 ( 
.A(n_446),
.B(n_393),
.C(n_343),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_380),
.B(n_327),
.C(n_343),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_448),
.B(n_464),
.C(n_350),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_408),
.A2(n_414),
.B1(n_397),
.B2(n_421),
.Y(n_451)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_396),
.A2(n_372),
.B1(n_367),
.B2(n_318),
.Y(n_454)
);

INVxp67_ASAP7_75t_L g490 ( 
.A(n_455),
.Y(n_490)
);

OAI21xp5_ASAP7_75t_SL g461 ( 
.A1(n_395),
.A2(n_402),
.B(n_384),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g484 ( 
.A1(n_461),
.A2(n_420),
.B(n_385),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g464 ( 
.A(n_417),
.B(n_320),
.Y(n_464)
);

OAI22xp5_ASAP7_75t_SL g467 ( 
.A1(n_408),
.A2(n_372),
.B1(n_367),
.B2(n_335),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_433),
.Y(n_468)
);

INVx13_ASAP7_75t_L g528 ( 
.A(n_468),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g469 ( 
.A(n_431),
.B(n_402),
.Y(n_469)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_469),
.Y(n_521)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_439),
.Y(n_470)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_470),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_435),
.B(n_389),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g514 ( 
.A(n_471),
.B(n_475),
.Y(n_514)
);

AOI22xp5_ASAP7_75t_SL g472 ( 
.A1(n_429),
.A2(n_416),
.B1(n_384),
.B2(n_376),
.Y(n_472)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_472),
.A2(n_482),
.B(n_484),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_453),
.A2(n_415),
.B1(n_423),
.B2(n_395),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g510 ( 
.A1(n_473),
.A2(n_478),
.B1(n_434),
.B2(n_455),
.Y(n_510)
);

XOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_446),
.B(n_379),
.Y(n_474)
);

XNOR2x1_ASAP7_75t_L g533 ( 
.A(n_474),
.B(n_488),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_427),
.B(n_403),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_439),
.Y(n_476)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_476),
.Y(n_513)
);

NAND2x1p5_ASAP7_75t_L g477 ( 
.A(n_434),
.B(n_405),
.Y(n_477)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_477),
.A2(n_489),
.B(n_450),
.Y(n_507)
);

OAI22xp5_ASAP7_75t_SL g478 ( 
.A1(n_432),
.A2(n_405),
.B1(n_390),
.B2(n_418),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_441),
.B(n_424),
.Y(n_479)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_441),
.B(n_400),
.Y(n_480)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_480),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_SL g481 ( 
.A(n_437),
.B(n_392),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_481),
.B(n_491),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_452),
.B(n_382),
.Y(n_483)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_483),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g485 ( 
.A(n_433),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_485),
.B(n_487),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_452),
.B(n_392),
.Y(n_486)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_486),
.Y(n_534)
);

AND2x6_ASAP7_75t_L g487 ( 
.A(n_445),
.B(n_393),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g489 ( 
.A(n_431),
.B(n_419),
.Y(n_489)
);

CKINVDCx16_ASAP7_75t_R g491 ( 
.A(n_462),
.Y(n_491)
);

AND2x6_ASAP7_75t_L g492 ( 
.A(n_445),
.B(n_398),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_492),
.B(n_493),
.Y(n_518)
);

INVx1_ASAP7_75t_SL g493 ( 
.A(n_430),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g494 ( 
.A(n_438),
.B(n_350),
.Y(n_494)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_494),
.B(n_370),
.Y(n_523)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_427),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_495),
.B(n_502),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_506),
.Y(n_527)
);

NOR2xp33_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_386),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_L g539 ( 
.A(n_498),
.B(n_499),
.Y(n_539)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_447),
.B(n_329),
.Y(n_499)
);

AO22x1_ASAP7_75t_L g502 ( 
.A1(n_451),
.A2(n_360),
.B1(n_398),
.B2(n_388),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_448),
.B(n_464),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_503),
.B(n_348),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_428),
.A2(n_398),
.B1(n_412),
.B2(n_425),
.Y(n_504)
);

OAI22xp5_ASAP7_75t_SL g512 ( 
.A1(n_504),
.A2(n_463),
.B1(n_458),
.B2(n_440),
.Y(n_512)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_467),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_505),
.B(n_457),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_329),
.C(n_322),
.Y(n_506)
);

OR2x2_ASAP7_75t_L g552 ( 
.A(n_507),
.B(n_469),
.Y(n_552)
);

OAI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_510),
.A2(n_517),
.B1(n_520),
.B2(n_522),
.Y(n_550)
);

OAI22xp5_ASAP7_75t_L g511 ( 
.A1(n_500),
.A2(n_466),
.B1(n_454),
.B2(n_443),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_511),
.A2(n_512),
.B1(n_537),
.B2(n_544),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g517 ( 
.A1(n_501),
.A2(n_444),
.B1(n_426),
.B2(n_438),
.Y(n_517)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_500),
.A2(n_442),
.B1(n_436),
.B2(n_458),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g522 ( 
.A1(n_473),
.A2(n_440),
.B1(n_463),
.B2(n_457),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_523),
.B(n_496),
.C(n_497),
.Y(n_547)
);

AOI21xp5_ASAP7_75t_L g525 ( 
.A1(n_482),
.A2(n_430),
.B(n_398),
.Y(n_525)
);

AOI21xp5_ASAP7_75t_L g565 ( 
.A1(n_525),
.A2(n_484),
.B(n_492),
.Y(n_565)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_526),
.Y(n_554)
);

AOI22x1_ASAP7_75t_SL g530 ( 
.A1(n_478),
.A2(n_465),
.B1(n_456),
.B2(n_449),
.Y(n_530)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_SL g531 ( 
.A1(n_472),
.A2(n_456),
.B(n_449),
.Y(n_531)
);

CKINVDCx14_ASAP7_75t_R g560 ( 
.A(n_531),
.Y(n_560)
);

NAND2xp5_ASAP7_75t_L g535 ( 
.A(n_495),
.B(n_459),
.Y(n_535)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_535),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g536 ( 
.A(n_468),
.B(n_485),
.Y(n_536)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_536),
.Y(n_576)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_505),
.A2(n_465),
.B1(n_459),
.B2(n_430),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_483),
.Y(n_538)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_538),
.Y(n_569)
);

XNOR2x2_ASAP7_75t_L g540 ( 
.A(n_477),
.B(n_488),
.Y(n_540)
);

NAND2xp5_ASAP7_75t_L g574 ( 
.A(n_540),
.B(n_502),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_541),
.B(n_494),
.Y(n_549)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_470),
.Y(n_542)
);

INVx1_ASAP7_75t_SL g551 ( 
.A(n_542),
.Y(n_551)
);

NOR2xp33_ASAP7_75t_L g543 ( 
.A(n_481),
.B(n_391),
.Y(n_543)
);

CKINVDCx14_ASAP7_75t_R g563 ( 
.A(n_543),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_L g544 ( 
.A1(n_504),
.A2(n_430),
.B1(n_425),
.B2(n_335),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_511),
.A2(n_524),
.B1(n_509),
.B2(n_515),
.Y(n_546)
);

OAI22xp5_ASAP7_75t_SL g583 ( 
.A1(n_546),
.A2(n_575),
.B1(n_577),
.B2(n_522),
.Y(n_583)
);

XOR2xp5_ASAP7_75t_L g580 ( 
.A(n_547),
.B(n_558),
.Y(n_580)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_535),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g581 ( 
.A(n_548),
.B(n_549),
.Y(n_581)
);

INVxp67_ASAP7_75t_L g593 ( 
.A(n_552),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g553 ( 
.A(n_536),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_553),
.B(n_557),
.Y(n_592)
);

OAI21xp33_ASAP7_75t_L g557 ( 
.A1(n_515),
.A2(n_486),
.B(n_479),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_527),
.B(n_506),
.C(n_517),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g585 ( 
.A(n_558),
.B(n_564),
.C(n_568),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g559 ( 
.A(n_514),
.B(n_496),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_559),
.B(n_544),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_SL g561 ( 
.A1(n_510),
.A2(n_490),
.B1(n_469),
.B2(n_480),
.Y(n_561)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_561),
.Y(n_582)
);

NOR2xp33_ASAP7_75t_L g562 ( 
.A(n_516),
.B(n_490),
.Y(n_562)
);

CKINVDCx16_ASAP7_75t_R g584 ( 
.A(n_562),
.Y(n_584)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_527),
.B(n_474),
.C(n_477),
.Y(n_564)
);

OAI22xp5_ASAP7_75t_L g595 ( 
.A1(n_565),
.A2(n_530),
.B1(n_525),
.B2(n_518),
.Y(n_595)
);

AOI21xp5_ASAP7_75t_L g566 ( 
.A1(n_519),
.A2(n_487),
.B(n_489),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g599 ( 
.A(n_566),
.Y(n_599)
);

INVx3_ASAP7_75t_SL g567 ( 
.A(n_509),
.Y(n_567)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_567),
.Y(n_594)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_520),
.B(n_476),
.C(n_489),
.Y(n_568)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_507),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g589 ( 
.A(n_570),
.B(n_531),
.Y(n_589)
);

OAI22xp5_ASAP7_75t_SL g571 ( 
.A1(n_534),
.A2(n_524),
.B1(n_532),
.B2(n_538),
.Y(n_571)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_571),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g572 ( 
.A(n_523),
.B(n_344),
.C(n_322),
.Y(n_572)
);

MAJIxp5_ASAP7_75t_L g587 ( 
.A(n_572),
.B(n_573),
.C(n_578),
.Y(n_587)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_533),
.B(n_502),
.C(n_331),
.Y(n_573)
);

XNOR2xp5_ASAP7_75t_L g586 ( 
.A(n_574),
.B(n_540),
.Y(n_586)
);

AOI22xp5_ASAP7_75t_L g575 ( 
.A1(n_526),
.A2(n_521),
.B1(n_534),
.B2(n_512),
.Y(n_575)
);

AOI22xp5_ASAP7_75t_L g577 ( 
.A1(n_521),
.A2(n_532),
.B1(n_518),
.B2(n_529),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_533),
.B(n_331),
.C(n_360),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g579 ( 
.A(n_540),
.B(n_360),
.C(n_337),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g597 ( 
.A(n_579),
.B(n_537),
.C(n_542),
.Y(n_597)
);

XNOR2xp5_ASAP7_75t_L g624 ( 
.A(n_580),
.B(n_588),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_583),
.A2(n_576),
.B1(n_554),
.B2(n_556),
.Y(n_612)
);

INVxp67_ASAP7_75t_L g628 ( 
.A(n_586),
.Y(n_628)
);

XOR2xp5_ASAP7_75t_L g588 ( 
.A(n_550),
.B(n_519),
.Y(n_588)
);

INVx1_ASAP7_75t_L g608 ( 
.A(n_589),
.Y(n_608)
);

NAND2xp5_ASAP7_75t_L g590 ( 
.A(n_571),
.B(n_529),
.Y(n_590)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_590),
.Y(n_613)
);

CKINVDCx16_ASAP7_75t_R g591 ( 
.A(n_561),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_591),
.B(n_596),
.Y(n_617)
);

XNOR2xp5_ASAP7_75t_L g625 ( 
.A(n_595),
.B(n_597),
.Y(n_625)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_568),
.B(n_539),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g598 ( 
.A(n_563),
.B(n_550),
.Y(n_598)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_598),
.B(n_600),
.Y(n_626)
);

MAJIxp5_ASAP7_75t_L g600 ( 
.A(n_547),
.B(n_528),
.C(n_513),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_577),
.B(n_513),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_601),
.B(n_605),
.Y(n_614)
);

OAI22xp5_ASAP7_75t_L g603 ( 
.A1(n_546),
.A2(n_545),
.B1(n_567),
.B2(n_575),
.Y(n_603)
);

AOI22xp5_ASAP7_75t_L g622 ( 
.A1(n_603),
.A2(n_555),
.B1(n_551),
.B2(n_578),
.Y(n_622)
);

XNOR2xp5_ASAP7_75t_L g604 ( 
.A(n_564),
.B(n_528),
.Y(n_604)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_604),
.B(n_570),
.Y(n_615)
);

MAJIxp5_ASAP7_75t_L g605 ( 
.A(n_572),
.B(n_528),
.C(n_508),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_576),
.B(n_508),
.Y(n_606)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_606),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g627 ( 
.A(n_607),
.B(n_325),
.Y(n_627)
);

XNOR2xp5_ASAP7_75t_SL g609 ( 
.A(n_586),
.B(n_574),
.Y(n_609)
);

XNOR2xp5_ASAP7_75t_L g642 ( 
.A(n_609),
.B(n_597),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_594),
.Y(n_610)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_610),
.Y(n_650)
);

OAI22xp5_ASAP7_75t_L g636 ( 
.A1(n_612),
.A2(n_620),
.B1(n_622),
.B2(n_630),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_615),
.B(n_627),
.Y(n_640)
);

NOR3xp33_ASAP7_75t_L g616 ( 
.A(n_592),
.B(n_566),
.C(n_579),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g637 ( 
.A(n_616),
.B(n_599),
.Y(n_637)
);

AOI21xp5_ASAP7_75t_L g618 ( 
.A1(n_600),
.A2(n_560),
.B(n_565),
.Y(n_618)
);

OAI21x1_ASAP7_75t_L g643 ( 
.A1(n_618),
.A2(n_621),
.B(n_593),
.Y(n_643)
);

MAJIxp5_ASAP7_75t_L g619 ( 
.A(n_580),
.B(n_573),
.C(n_554),
.Y(n_619)
);

MAJIxp5_ASAP7_75t_L g634 ( 
.A(n_619),
.B(n_623),
.C(n_629),
.Y(n_634)
);

AOI22xp5_ASAP7_75t_L g620 ( 
.A1(n_603),
.A2(n_556),
.B1(n_545),
.B2(n_569),
.Y(n_620)
);

AOI21xp5_ASAP7_75t_L g621 ( 
.A1(n_604),
.A2(n_552),
.B(n_555),
.Y(n_621)
);

MAJIxp5_ASAP7_75t_L g623 ( 
.A(n_585),
.B(n_551),
.C(n_493),
.Y(n_623)
);

MAJIxp5_ASAP7_75t_L g629 ( 
.A(n_585),
.B(n_351),
.C(n_394),
.Y(n_629)
);

AOI22xp5_ASAP7_75t_L g630 ( 
.A1(n_584),
.A2(n_330),
.B1(n_352),
.B2(n_394),
.Y(n_630)
);

A2O1A1Ixp33_ASAP7_75t_SL g631 ( 
.A1(n_589),
.A2(n_377),
.B(n_352),
.C(n_330),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_631),
.B(n_594),
.Y(n_644)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_610),
.Y(n_632)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_632),
.Y(n_655)
);

NOR2xp33_ASAP7_75t_SL g633 ( 
.A(n_626),
.B(n_581),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_633),
.B(n_638),
.Y(n_654)
);

INVx1_ASAP7_75t_L g635 ( 
.A(n_612),
.Y(n_635)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_635),
.Y(n_660)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_637),
.Y(n_664)
);

MAJIxp5_ASAP7_75t_L g638 ( 
.A(n_623),
.B(n_605),
.C(n_591),
.Y(n_638)
);

MAJIxp5_ASAP7_75t_L g639 ( 
.A(n_619),
.B(n_588),
.C(n_587),
.Y(n_639)
);

XNOR2xp5_ASAP7_75t_L g652 ( 
.A(n_639),
.B(n_645),
.Y(n_652)
);

XOR2x1_ASAP7_75t_SL g641 ( 
.A(n_609),
.B(n_593),
.Y(n_641)
);

OAI21xp33_ASAP7_75t_L g665 ( 
.A1(n_641),
.A2(n_646),
.B(n_651),
.Y(n_665)
);

XOR2xp5_ASAP7_75t_L g662 ( 
.A(n_642),
.B(n_647),
.Y(n_662)
);

AND2x2_ASAP7_75t_L g659 ( 
.A(n_643),
.B(n_624),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_SL g657 ( 
.A1(n_644),
.A2(n_583),
.B1(n_636),
.B2(n_635),
.Y(n_657)
);

MAJIxp5_ASAP7_75t_L g645 ( 
.A(n_624),
.B(n_587),
.C(n_582),
.Y(n_645)
);

OAI21xp5_ASAP7_75t_SL g646 ( 
.A1(n_617),
.A2(n_599),
.B(n_595),
.Y(n_646)
);

OA21x2_ASAP7_75t_L g647 ( 
.A1(n_608),
.A2(n_582),
.B(n_602),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_SL g648 ( 
.A(n_614),
.B(n_590),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_SL g656 ( 
.A(n_648),
.B(n_625),
.Y(n_656)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_620),
.Y(n_649)
);

XNOR2xp5_ASAP7_75t_L g653 ( 
.A(n_649),
.B(n_625),
.Y(n_653)
);

OAI21xp5_ASAP7_75t_SL g651 ( 
.A1(n_611),
.A2(n_602),
.B(n_606),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_653),
.B(n_656),
.Y(n_678)
);

OAI22xp33_ASAP7_75t_SL g671 ( 
.A1(n_657),
.A2(n_667),
.B1(n_632),
.B2(n_650),
.Y(n_671)
);

XNOR2xp5_ASAP7_75t_L g658 ( 
.A(n_639),
.B(n_629),
.Y(n_658)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_658),
.B(n_661),
.Y(n_669)
);

AND2x2_ASAP7_75t_SL g673 ( 
.A(n_659),
.B(n_645),
.Y(n_673)
);

MAJIxp5_ASAP7_75t_L g661 ( 
.A(n_638),
.B(n_628),
.C(n_613),
.Y(n_661)
);

XNOR2xp5_ASAP7_75t_L g663 ( 
.A(n_634),
.B(n_628),
.Y(n_663)
);

MAJIxp5_ASAP7_75t_L g674 ( 
.A(n_663),
.B(n_666),
.C(n_642),
.Y(n_674)
);

MAJIxp5_ASAP7_75t_L g666 ( 
.A(n_634),
.B(n_631),
.C(n_377),
.Y(n_666)
);

AOI22xp5_ASAP7_75t_SL g667 ( 
.A1(n_649),
.A2(n_631),
.B1(n_256),
.B2(n_227),
.Y(n_667)
);

OAI22xp5_ASAP7_75t_SL g668 ( 
.A1(n_644),
.A2(n_631),
.B1(n_225),
.B2(n_189),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g676 ( 
.A(n_668),
.B(n_225),
.Y(n_676)
);

NAND2x1p5_ASAP7_75t_L g670 ( 
.A(n_660),
.B(n_651),
.Y(n_670)
);

AO21x1_ASAP7_75t_L g690 ( 
.A1(n_670),
.A2(n_679),
.B(n_680),
.Y(n_690)
);

XOR2xp5_ASAP7_75t_L g688 ( 
.A(n_671),
.B(n_6),
.Y(n_688)
);

CKINVDCx16_ASAP7_75t_R g672 ( 
.A(n_659),
.Y(n_672)
);

AOI22xp5_ASAP7_75t_L g689 ( 
.A1(n_672),
.A2(n_676),
.B1(n_677),
.B2(n_681),
.Y(n_689)
);

CKINVDCx20_ASAP7_75t_R g684 ( 
.A(n_673),
.Y(n_684)
);

OR2x2_ASAP7_75t_L g683 ( 
.A(n_674),
.B(n_675),
.Y(n_683)
);

MAJIxp5_ASAP7_75t_L g675 ( 
.A(n_652),
.B(n_646),
.C(n_640),
.Y(n_675)
);

INVxp67_ASAP7_75t_L g677 ( 
.A(n_654),
.Y(n_677)
);

OAI21xp5_ASAP7_75t_SL g679 ( 
.A1(n_664),
.A2(n_647),
.B(n_640),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_662),
.B(n_647),
.Y(n_680)
);

OAI21xp5_ASAP7_75t_L g681 ( 
.A1(n_665),
.A2(n_641),
.B(n_189),
.Y(n_681)
);

NOR2xp33_ASAP7_75t_L g682 ( 
.A(n_669),
.B(n_655),
.Y(n_682)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_682),
.Y(n_695)
);

NOR2xp33_ASAP7_75t_SL g685 ( 
.A(n_669),
.B(n_661),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_685),
.B(n_686),
.Y(n_692)
);

XNOR2xp5_ASAP7_75t_L g686 ( 
.A(n_673),
.B(n_662),
.Y(n_686)
);

AOI322xp5_ASAP7_75t_L g687 ( 
.A1(n_680),
.A2(n_665),
.A3(n_657),
.B1(n_667),
.B2(n_666),
.C1(n_6),
.C2(n_14),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_687),
.B(n_688),
.Y(n_694)
);

OAI21xp5_ASAP7_75t_SL g691 ( 
.A1(n_684),
.A2(n_678),
.B(n_670),
.Y(n_691)
);

NOR3xp33_ASAP7_75t_L g698 ( 
.A(n_691),
.B(n_2),
.C(n_5),
.Y(n_698)
);

MAJIxp5_ASAP7_75t_L g693 ( 
.A(n_683),
.B(n_17),
.C(n_2),
.Y(n_693)
);

NOR2xp33_ASAP7_75t_L g696 ( 
.A(n_693),
.B(n_0),
.Y(n_696)
);

OAI21xp5_ASAP7_75t_L g699 ( 
.A1(n_696),
.A2(n_697),
.B(n_698),
.Y(n_699)
);

AOI322xp5_ASAP7_75t_L g697 ( 
.A1(n_695),
.A2(n_690),
.A3(n_682),
.B1(n_689),
.B2(n_687),
.C1(n_15),
.C2(n_16),
.Y(n_697)
);

MAJIxp5_ASAP7_75t_L g700 ( 
.A(n_697),
.B(n_692),
.C(n_694),
.Y(n_700)
);

AOI322xp5_ASAP7_75t_L g701 ( 
.A1(n_700),
.A2(n_0),
.A3(n_1),
.B1(n_5),
.B2(n_15),
.C1(n_16),
.C2(n_699),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_701),
.Y(n_702)
);

AOI31xp33_ASAP7_75t_L g703 ( 
.A1(n_702),
.A2(n_5),
.A3(n_15),
.B(n_0),
.Y(n_703)
);

AOI21xp5_ASAP7_75t_L g704 ( 
.A1(n_703),
.A2(n_0),
.B(n_1),
.Y(n_704)
);


endmodule