module fake_jpeg_3421_n_194 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_194);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_194;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_16),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_23),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_5),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_47),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_33),
.Y(n_55)
);

BUFx4f_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_39),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx14_ASAP7_75t_R g59 ( 
.A(n_9),
.Y(n_59)
);

BUFx3_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_13),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_22),
.Y(n_62)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_8),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_19),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_9),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_22),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_29),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_57),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g79 ( 
.A(n_68),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx6_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx6_ASAP7_75t_SL g70 ( 
.A(n_57),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_73),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_75),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_51),
.Y(n_72)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_72),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_59),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_50),
.Y(n_74)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_74),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_56),
.B(n_45),
.Y(n_75)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_77),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g78 ( 
.A1(n_70),
.A2(n_51),
.B1(n_60),
.B2(n_63),
.Y(n_78)
);

O2A1O1Ixp33_ASAP7_75t_L g104 ( 
.A1(n_78),
.A2(n_77),
.B(n_87),
.C(n_62),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_69),
.A2(n_60),
.B1(n_63),
.B2(n_53),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_81),
.A2(n_69),
.B1(n_72),
.B2(n_62),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_66),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_82),
.B(n_84),
.Y(n_92)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_74),
.Y(n_83)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_75),
.A2(n_48),
.B1(n_61),
.B2(n_56),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_85),
.A2(n_64),
.B1(n_65),
.B2(n_49),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_72),
.B(n_54),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_58),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_84),
.A2(n_61),
.B1(n_48),
.B2(n_50),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_94),
.B1(n_105),
.B2(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_92),
.B(n_98),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_85),
.A2(n_72),
.B1(n_66),
.B2(n_53),
.Y(n_93)
);

AO22x2_ASAP7_75t_L g112 ( 
.A1(n_93),
.A2(n_101),
.B1(n_76),
.B2(n_1),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_95),
.Y(n_113)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_88),
.Y(n_96)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_96),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_78),
.A2(n_69),
.B1(n_64),
.B2(n_67),
.Y(n_97)
);

INVxp67_ASAP7_75t_L g117 ( 
.A(n_97),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_80),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_100),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_86),
.B(n_52),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_88),
.A2(n_67),
.B1(n_55),
.B2(n_52),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_83),
.Y(n_102)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_102),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_78),
.B(n_55),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_104),
.Y(n_123)
);

O2A1O1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_104),
.A2(n_0),
.B(n_3),
.C(n_4),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g105 ( 
.A1(n_78),
.A2(n_87),
.B1(n_76),
.B2(n_79),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_100),
.B(n_98),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_106),
.B(n_107),
.C(n_124),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_79),
.C(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_91),
.Y(n_110)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_110),
.Y(n_129)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_91),
.Y(n_111)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_116),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g114 ( 
.A1(n_94),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g141 ( 
.A1(n_114),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_141)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_102),
.Y(n_115)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_115),
.Y(n_145)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

A2O1A1Ixp33_ASAP7_75t_SL g133 ( 
.A1(n_118),
.A2(n_6),
.B(n_7),
.C(n_8),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_125),
.B1(n_10),
.B2(n_11),
.Y(n_135)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_89),
.Y(n_122)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_123),
.B(n_11),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_103),
.B(n_3),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_105),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_125)
);

XOR2xp5_ASAP7_75t_L g127 ( 
.A(n_108),
.B(n_93),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_127),
.B(n_130),
.C(n_134),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g130 ( 
.A(n_109),
.B(n_89),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_122),
.B(n_101),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_132),
.B(n_136),
.Y(n_151)
);

CKINVDCx14_ASAP7_75t_R g160 ( 
.A(n_133),
.Y(n_160)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_117),
.A2(n_7),
.B(n_10),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_135),
.A2(n_141),
.B1(n_142),
.B2(n_25),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_121),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_138),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_118),
.B(n_12),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_117),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_113),
.B1(n_112),
.B2(n_23),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_119),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_140),
.B(n_146),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_142)
);

AOI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_113),
.A2(n_17),
.B(n_19),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_144),
.B(n_133),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_112),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g169 ( 
.A(n_148),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_149),
.B(n_152),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_128),
.A2(n_112),
.B1(n_21),
.B2(n_20),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_155),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_32),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g153 ( 
.A(n_134),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_153),
.B(n_162),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_131),
.Y(n_154)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_154),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_127),
.B(n_31),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_126),
.B(n_34),
.C(n_40),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_27),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_139),
.A2(n_145),
.B1(n_143),
.B2(n_133),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_158),
.A2(n_141),
.B1(n_28),
.B2(n_30),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_126),
.B(n_20),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_140),
.B(n_21),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_164),
.Y(n_167)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_144),
.B(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g181 ( 
.A(n_171),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_172),
.A2(n_149),
.B1(n_158),
.B2(n_165),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g176 ( 
.A(n_173),
.B(n_157),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_166),
.B(n_159),
.Y(n_175)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_175),
.Y(n_183)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_176),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_168),
.B(n_156),
.C(n_152),
.Y(n_177)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_177),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_178),
.A2(n_179),
.B1(n_180),
.B2(n_174),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_173),
.B(n_156),
.C(n_155),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_171),
.A2(n_148),
.B(n_151),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_182),
.A2(n_181),
.B1(n_169),
.B2(n_174),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_186),
.A2(n_187),
.B1(n_181),
.B2(n_160),
.Y(n_188)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_183),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_188),
.B(n_182),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_189),
.B(n_185),
.C(n_184),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_190),
.B(n_177),
.Y(n_191)
);

AOI321xp33_ASAP7_75t_L g192 ( 
.A1(n_191),
.A2(n_167),
.A3(n_170),
.B1(n_38),
.B2(n_42),
.C(n_37),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g193 ( 
.A(n_192),
.B(n_172),
.C(n_36),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_193),
.B(n_150),
.Y(n_194)
);


endmodule