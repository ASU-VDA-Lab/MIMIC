module fake_jpeg_8981_n_284 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_284);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_284;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

INVx2_ASAP7_75t_L g13 ( 
.A(n_7),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

BUFx3_ASAP7_75t_L g15 ( 
.A(n_4),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_11),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_0),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_26),
.Y(n_28)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_28),
.Y(n_47)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_13),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_30),
.Y(n_51)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_34),
.Y(n_43)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx4_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_20),
.Y(n_37)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_38),
.B(n_40),
.Y(n_67)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g64 ( 
.A(n_41),
.B(n_49),
.Y(n_64)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_42),
.Y(n_60)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_45),
.Y(n_73)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_50),
.B(n_52),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_33),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_54),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_L g55 ( 
.A1(n_35),
.A2(n_13),
.B1(n_27),
.B2(n_16),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_55),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_56),
.Y(n_81)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_57),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_47),
.A2(n_13),
.B1(n_17),
.B2(n_18),
.Y(n_58)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_58),
.A2(n_59),
.B1(n_61),
.B2(n_72),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_47),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_61)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_49),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_62),
.B(n_63),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_65),
.A2(n_70),
.B1(n_60),
.B2(n_44),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

CKINVDCx14_ASAP7_75t_R g86 ( 
.A(n_66),
.Y(n_86)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_70),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_52),
.B(n_29),
.Y(n_71)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_71),
.A2(n_75),
.B(n_69),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_42),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_22),
.B1(n_20),
.B2(n_23),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_74),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_80)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_39),
.B(n_19),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_48),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_76),
.Y(n_94)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx11_ASAP7_75t_L g101 ( 
.A(n_77),
.Y(n_101)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_64),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_79),
.Y(n_100)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_80),
.A2(n_83),
.B1(n_65),
.B2(n_60),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_82),
.B(n_90),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

INVx3_ASAP7_75t_SL g102 ( 
.A(n_85),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_75),
.B(n_71),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_46),
.B1(n_16),
.B2(n_21),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_89),
.A2(n_73),
.B1(n_25),
.B2(n_24),
.Y(n_112)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_67),
.Y(n_90)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_67),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_93),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_69),
.A2(n_21),
.B1(n_16),
.B2(n_27),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_97),
.B1(n_21),
.B2(n_27),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_95),
.Y(n_104)
);

OAI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_63),
.A2(n_75),
.B1(n_60),
.B2(n_65),
.Y(n_97)
);

BUFx24_ASAP7_75t_SL g99 ( 
.A(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_99),
.B(n_116),
.Y(n_128)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_96),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_103),
.B(n_106),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_105),
.B(n_22),
.Y(n_143)
);

CKINVDCx16_ASAP7_75t_R g106 ( 
.A(n_96),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_107),
.A2(n_111),
.B1(n_119),
.B2(n_81),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_71),
.Y(n_108)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_108),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_91),
.B(n_68),
.Y(n_109)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

AOI32xp33_ASAP7_75t_L g110 ( 
.A1(n_84),
.A2(n_72),
.A3(n_30),
.B1(n_28),
.B2(n_15),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_110),
.A2(n_117),
.B1(n_106),
.B2(n_103),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_112),
.A2(n_98),
.B1(n_94),
.B2(n_81),
.Y(n_133)
);

NAND2xp33_ASAP7_75t_SL g115 ( 
.A(n_87),
.B(n_0),
.Y(n_115)
);

NAND2xp33_ASAP7_75t_SL g125 ( 
.A(n_115),
.B(n_0),
.Y(n_125)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_80),
.Y(n_116)
);

NAND3xp33_ASAP7_75t_L g117 ( 
.A(n_93),
.B(n_79),
.C(n_92),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_89),
.B(n_15),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_118),
.B(n_86),
.C(n_88),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_86),
.A2(n_73),
.B1(n_25),
.B2(n_24),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_82),
.B(n_56),
.Y(n_120)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_121),
.B(n_126),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_122),
.B(n_109),
.C(n_100),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_123),
.B(n_133),
.Y(n_146)
);

AND2x6_ASAP7_75t_L g124 ( 
.A(n_115),
.B(n_12),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_124),
.Y(n_164)
);

NAND3xp33_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_12),
.C(n_2),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_116),
.A2(n_107),
.B1(n_110),
.B2(n_108),
.Y(n_126)
);

OAI32xp33_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_88),
.A3(n_15),
.B1(n_23),
.B2(n_22),
.Y(n_127)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_127),
.Y(n_144)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_102),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_131),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_105),
.B(n_1),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_130),
.A2(n_140),
.B(n_114),
.Y(n_150)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_132),
.Y(n_159)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_101),
.Y(n_134)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_135),
.B(n_142),
.Y(n_153)
);

AND2x2_ASAP7_75t_L g140 ( 
.A(n_118),
.B(n_1),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_101),
.B(n_98),
.Y(n_141)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_141),
.Y(n_155)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_120),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g157 ( 
.A(n_143),
.B(n_30),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_145),
.B(n_129),
.C(n_85),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_123),
.A2(n_142),
.B1(n_138),
.B2(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_147),
.A2(n_148),
.B1(n_151),
.B2(n_152),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_138),
.A2(n_113),
.B1(n_114),
.B2(n_117),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_150),
.B(n_132),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_136),
.A2(n_113),
.B1(n_100),
.B2(n_112),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g152 ( 
.A1(n_137),
.A2(n_111),
.B1(n_81),
.B2(n_104),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_136),
.A2(n_119),
.B1(n_98),
.B2(n_104),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_154),
.A2(n_161),
.B1(n_168),
.B2(n_166),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g156 ( 
.A1(n_143),
.A2(n_102),
.A3(n_22),
.B1(n_23),
.B2(n_28),
.Y(n_156)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g186 ( 
.A(n_157),
.B(n_1),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_139),
.B(n_95),
.Y(n_158)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_158),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_122),
.A2(n_56),
.B1(n_76),
.B2(n_77),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_162),
.B(n_163),
.Y(n_170)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_133),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_140),
.B(n_23),
.Y(n_165)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_165),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_127),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_167),
.B(n_168),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_76),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_157),
.B(n_130),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_171),
.B(n_179),
.C(n_185),
.Y(n_198)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_159),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_172),
.B(n_173),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

AOI21xp5_ASAP7_75t_SL g174 ( 
.A1(n_164),
.A2(n_130),
.B(n_124),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_174),
.A2(n_188),
.B(n_150),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_163),
.A2(n_135),
.B1(n_128),
.B2(n_131),
.Y(n_175)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_175),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_153),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_176),
.B(n_181),
.Y(n_199)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_178),
.B(n_186),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_180),
.A2(n_161),
.B1(n_164),
.B2(n_156),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_158),
.Y(n_181)
);

INVxp33_ASAP7_75t_L g183 ( 
.A(n_160),
.Y(n_183)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_183),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_151),
.B(n_134),
.Y(n_184)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_184),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_145),
.B(n_85),
.C(n_2),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_147),
.B(n_1),
.C(n_2),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_187),
.B(n_3),
.Y(n_203)
);

XOR2x2_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_12),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_154),
.B(n_2),
.Y(n_190)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_190),
.Y(n_205)
);

OA21x2_ASAP7_75t_L g192 ( 
.A1(n_169),
.A2(n_167),
.B(n_144),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_193),
.B(n_196),
.Y(n_213)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_178),
.B(n_166),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_144),
.Y(n_201)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_201),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_172),
.Y(n_202)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_202),
.Y(n_218)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_203),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_204),
.A2(n_182),
.B1(n_146),
.B2(n_148),
.Y(n_212)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_184),
.Y(n_206)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_183),
.B(n_155),
.Y(n_207)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_207),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g208 ( 
.A(n_188),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_208),
.B(n_210),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_155),
.Y(n_210)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_179),
.C(n_185),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_217),
.C(n_219),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_194),
.B1(n_197),
.B2(n_195),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_200),
.A2(n_177),
.B1(n_191),
.B2(n_174),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_215),
.B1(n_194),
.B2(n_199),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_200),
.A2(n_177),
.B1(n_182),
.B2(n_159),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_171),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_186),
.C(n_149),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_209),
.B(n_187),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_221),
.B(n_226),
.C(n_205),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_170),
.B1(n_149),
.B2(n_165),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_222),
.A2(n_197),
.B1(n_201),
.B2(n_192),
.Y(n_235)
);

FAx1_ASAP7_75t_SL g224 ( 
.A(n_193),
.B(n_170),
.CI(n_152),
.CON(n_224),
.SN(n_224)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_224),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_206),
.B(n_3),
.C(n_4),
.Y(n_226)
);

XNOR2xp5_ASAP7_75t_SL g229 ( 
.A(n_213),
.B(n_196),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_229),
.B(n_233),
.Y(n_243)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_231),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_205),
.Y(n_232)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_232),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_SL g233 ( 
.A(n_214),
.B(n_196),
.Y(n_233)
);

CKINVDCx14_ASAP7_75t_R g253 ( 
.A(n_234),
.Y(n_253)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_217),
.B(n_221),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_237),
.C(n_11),
.Y(n_250)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_226),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g244 ( 
.A1(n_238),
.A2(n_241),
.B1(n_201),
.B2(n_192),
.Y(n_244)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_215),
.A2(n_220),
.B1(n_216),
.B2(n_224),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_239),
.A2(n_242),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_225),
.B(n_202),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g249 ( 
.A(n_240),
.Y(n_249)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_222),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_224),
.A2(n_227),
.B1(n_219),
.B2(n_211),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_244),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_233),
.B(n_218),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_245),
.B(n_250),
.C(n_254),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_246),
.B(n_248),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_228),
.A2(n_3),
.B(n_5),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_230),
.B(n_236),
.C(n_237),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_254),
.B(n_230),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_255),
.B(n_259),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_249),
.B(n_235),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_257),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_250),
.B(n_229),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_252),
.B(n_5),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_260),
.B(n_261),
.Y(n_268)
);

CKINVDCx16_ASAP7_75t_R g261 ( 
.A(n_248),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_6),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_263),
.B(n_253),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_243),
.B(n_6),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g267 ( 
.A(n_264),
.B(n_246),
.Y(n_267)
);

AOI21xp5_ASAP7_75t_SL g266 ( 
.A1(n_262),
.A2(n_251),
.B(n_247),
.Y(n_266)
);

AOI21x1_ASAP7_75t_SL g275 ( 
.A1(n_266),
.A2(n_264),
.B(n_7),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g272 ( 
.A(n_267),
.B(n_269),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_256),
.B(n_258),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_270),
.B(n_256),
.C(n_258),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_273),
.A2(n_275),
.B(n_268),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g274 ( 
.A1(n_265),
.A2(n_251),
.B(n_243),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_274),
.A2(n_271),
.B(n_268),
.Y(n_277)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_276),
.A2(n_277),
.B(n_272),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_278),
.B(n_6),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_L g280 ( 
.A1(n_279),
.A2(n_6),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C1(n_10),
.C2(n_11),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_280),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g282 ( 
.A1(n_281),
.A2(n_9),
.B(n_11),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_282),
.B(n_9),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_283),
.B(n_9),
.Y(n_284)
);


endmodule