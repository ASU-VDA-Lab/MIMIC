module fake_aes_2762_n_1037 (n_303, n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_300, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_292, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_297, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_304, n_127, n_291, n_170, n_294, n_40, n_111, n_157, n_296, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_295, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_298, n_283, n_299, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_293, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_305, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_301, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_302, n_145, n_270, n_246, n_153, n_61, n_259, n_290, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1037);
input n_303;
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_300;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_292;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_297;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_304;
input n_127;
input n_291;
input n_170;
input n_294;
input n_40;
input n_111;
input n_157;
input n_296;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_295;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_298;
input n_283;
input n_299;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_293;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_305;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_301;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_302;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_290;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1037;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_1034;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_1031;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_667;
wire n_496;
wire n_311;
wire n_801;
wire n_988;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_1032;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_917;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_1030;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_617;
wire n_384;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_599;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_975;
wire n_968;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_809;
wire n_567;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_455;
wire n_312;
wire n_529;
wire n_1025;
wire n_1011;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_624;
wire n_426;
wire n_769;
wire n_725;
wire n_818;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1033;
wire n_1014;
wire n_767;
wire n_828;
wire n_533;
wire n_506;
wire n_393;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_826;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_1028;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_935;
wire n_427;
wire n_910;
wire n_950;
wire n_460;
wire n_478;
wire n_415;
wire n_482;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_813;
wire n_938;
wire n_928;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_699;
wire n_338;
wire n_519;
wire n_729;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_1036;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_902;
wire n_905;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_1035;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_420;
wire n_621;
wire n_446;
wire n_342;
wire n_423;
wire n_666;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_937;
wire n_388;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_822;
wire n_823;
wire n_970;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_899;
wire n_654;
wire n_894;
wire n_495;
wire n_428;
wire n_364;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_1029;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_553;
wire n_440;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_498;
wire n_349;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_763;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_875;
wire n_620;
wire n_841;
wire n_947;
wire n_912;
wire n_924;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_1027;
wire n_859;
wire n_994;
wire n_930;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_991;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
INVxp33_ASAP7_75t_SL g306 ( .A(n_200), .Y(n_306) );
BUFx3_ASAP7_75t_L g307 ( .A(n_178), .Y(n_307) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_196), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_302), .Y(n_309) );
CKINVDCx20_ASAP7_75t_R g310 ( .A(n_141), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_209), .Y(n_311) );
INVxp67_ASAP7_75t_SL g312 ( .A(n_259), .Y(n_312) );
CKINVDCx16_ASAP7_75t_R g313 ( .A(n_222), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_86), .Y(n_314) );
INVxp33_ASAP7_75t_SL g315 ( .A(n_56), .Y(n_315) );
INVx3_ASAP7_75t_L g316 ( .A(n_130), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_176), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_229), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_91), .Y(n_319) );
INVx1_ASAP7_75t_L g320 ( .A(n_170), .Y(n_320) );
BUFx3_ASAP7_75t_L g321 ( .A(n_134), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_64), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_0), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_203), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_79), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_193), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_246), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_255), .Y(n_328) );
INVx1_ASAP7_75t_L g329 ( .A(n_301), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_160), .Y(n_330) );
BUFx2_ASAP7_75t_SL g331 ( .A(n_224), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_169), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_202), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_150), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_228), .Y(n_335) );
INVx1_ASAP7_75t_L g336 ( .A(n_295), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_281), .Y(n_337) );
BUFx2_ASAP7_75t_L g338 ( .A(n_101), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_193), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_305), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_115), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_292), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_136), .Y(n_343) );
BUFx2_ASAP7_75t_L g344 ( .A(n_100), .Y(n_344) );
CKINVDCx5p33_ASAP7_75t_R g345 ( .A(n_304), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_263), .Y(n_346) );
INVxp33_ASAP7_75t_L g347 ( .A(n_72), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_172), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_205), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_104), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_283), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_149), .B(n_236), .Y(n_352) );
INVxp67_ASAP7_75t_SL g353 ( .A(n_105), .Y(n_353) );
INVx1_ASAP7_75t_L g354 ( .A(n_221), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_248), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_210), .Y(n_356) );
INVxp67_ASAP7_75t_SL g357 ( .A(n_287), .Y(n_357) );
CKINVDCx20_ASAP7_75t_R g358 ( .A(n_294), .Y(n_358) );
INVxp67_ASAP7_75t_SL g359 ( .A(n_5), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_233), .Y(n_360) );
INVx2_ASAP7_75t_SL g361 ( .A(n_260), .Y(n_361) );
INVxp33_ASAP7_75t_SL g362 ( .A(n_93), .Y(n_362) );
CKINVDCx16_ASAP7_75t_R g363 ( .A(n_118), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_284), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_270), .Y(n_365) );
INVx2_ASAP7_75t_L g366 ( .A(n_219), .Y(n_366) );
INVxp33_ASAP7_75t_L g367 ( .A(n_290), .Y(n_367) );
INVxp67_ASAP7_75t_L g368 ( .A(n_217), .Y(n_368) );
INVxp33_ASAP7_75t_SL g369 ( .A(n_288), .Y(n_369) );
HB1xp67_ASAP7_75t_L g370 ( .A(n_182), .Y(n_370) );
INVxp33_ASAP7_75t_SL g371 ( .A(n_241), .Y(n_371) );
HB1xp67_ASAP7_75t_L g372 ( .A(n_5), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_195), .Y(n_373) );
CKINVDCx20_ASAP7_75t_R g374 ( .A(n_12), .Y(n_374) );
CKINVDCx16_ASAP7_75t_R g375 ( .A(n_277), .Y(n_375) );
CKINVDCx5p33_ASAP7_75t_R g376 ( .A(n_22), .Y(n_376) );
INVxp33_ASAP7_75t_SL g377 ( .A(n_253), .Y(n_377) );
INVxp67_ASAP7_75t_SL g378 ( .A(n_276), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_293), .Y(n_379) );
INVx1_ASAP7_75t_L g380 ( .A(n_98), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_63), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_92), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_190), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_289), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_266), .Y(n_385) );
INVx1_ASAP7_75t_L g386 ( .A(n_104), .Y(n_386) );
INVxp33_ASAP7_75t_L g387 ( .A(n_39), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_173), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_225), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_192), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_66), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_256), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_118), .Y(n_393) );
CKINVDCx5p33_ASAP7_75t_R g394 ( .A(n_102), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_156), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_88), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_52), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_66), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_1), .Y(n_399) );
INVxp33_ASAP7_75t_SL g400 ( .A(n_122), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_272), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_174), .Y(n_402) );
INVx2_ASAP7_75t_L g403 ( .A(n_142), .Y(n_403) );
INVx1_ASAP7_75t_L g404 ( .A(n_198), .Y(n_404) );
INVxp67_ASAP7_75t_SL g405 ( .A(n_3), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_123), .Y(n_406) );
CKINVDCx16_ASAP7_75t_R g407 ( .A(n_89), .Y(n_407) );
BUFx6f_ASAP7_75t_L g408 ( .A(n_131), .Y(n_408) );
INVx2_ASAP7_75t_L g409 ( .A(n_34), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_136), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_216), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_19), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_82), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_250), .Y(n_414) );
CKINVDCx14_ASAP7_75t_R g415 ( .A(n_291), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_286), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_258), .Y(n_417) );
BUFx3_ASAP7_75t_L g418 ( .A(n_189), .Y(n_418) );
INVx2_ASAP7_75t_L g419 ( .A(n_211), .Y(n_419) );
CKINVDCx5p33_ASAP7_75t_R g420 ( .A(n_273), .Y(n_420) );
INVx1_ASAP7_75t_L g421 ( .A(n_194), .Y(n_421) );
INVx1_ASAP7_75t_L g422 ( .A(n_23), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_303), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_129), .Y(n_424) );
CKINVDCx5p33_ASAP7_75t_R g425 ( .A(n_257), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_195), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_96), .Y(n_427) );
BUFx2_ASAP7_75t_SL g428 ( .A(n_101), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_252), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_127), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_70), .Y(n_431) );
INVx1_ASAP7_75t_L g432 ( .A(n_235), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_142), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_151), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_148), .Y(n_435) );
INVxp33_ASAP7_75t_L g436 ( .A(n_102), .Y(n_436) );
INVx2_ASAP7_75t_L g437 ( .A(n_285), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_208), .Y(n_438) );
INVx2_ASAP7_75t_SL g439 ( .A(n_59), .Y(n_439) );
BUFx6f_ASAP7_75t_L g440 ( .A(n_127), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_100), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_80), .Y(n_442) );
INVxp67_ASAP7_75t_SL g443 ( .A(n_230), .Y(n_443) );
INVxp67_ASAP7_75t_L g444 ( .A(n_215), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_140), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_71), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_162), .Y(n_447) );
CKINVDCx20_ASAP7_75t_R g448 ( .A(n_251), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_242), .Y(n_449) );
CKINVDCx5p33_ASAP7_75t_R g450 ( .A(n_358), .Y(n_450) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_318), .A2(n_1), .B(n_2), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_316), .Y(n_452) );
OA21x2_ASAP7_75t_L g453 ( .A1(n_318), .A2(n_2), .B(n_3), .Y(n_453) );
CKINVDCx20_ASAP7_75t_R g454 ( .A(n_363), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_338), .B(n_344), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_316), .Y(n_456) );
INVx3_ASAP7_75t_L g457 ( .A(n_316), .Y(n_457) );
CKINVDCx20_ASAP7_75t_R g458 ( .A(n_407), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_324), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_313), .Y(n_460) );
NAND2xp5_ASAP7_75t_SL g461 ( .A(n_361), .B(n_4), .Y(n_461) );
CKINVDCx16_ASAP7_75t_R g462 ( .A(n_375), .Y(n_462) );
NAND2xp33_ASAP7_75t_SL g463 ( .A(n_347), .B(n_4), .Y(n_463) );
AND2x4_ASAP7_75t_L g464 ( .A(n_361), .B(n_6), .Y(n_464) );
BUFx6f_ASAP7_75t_L g465 ( .A(n_335), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_335), .Y(n_466) );
OR2x6_ASAP7_75t_L g467 ( .A(n_331), .B(n_6), .Y(n_467) );
INVx1_ASAP7_75t_L g468 ( .A(n_324), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_344), .B(n_7), .Y(n_469) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_308), .Y(n_470) );
CKINVDCx5p33_ASAP7_75t_R g471 ( .A(n_448), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_335), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_335), .Y(n_473) );
INVx2_ASAP7_75t_L g474 ( .A(n_335), .Y(n_474) );
CKINVDCx5p33_ASAP7_75t_R g475 ( .A(n_309), .Y(n_475) );
CKINVDCx5p33_ASAP7_75t_R g476 ( .A(n_415), .Y(n_476) );
BUFx2_ASAP7_75t_L g477 ( .A(n_475), .Y(n_477) );
AND2x4_ASAP7_75t_L g478 ( .A(n_464), .B(n_439), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_455), .A2(n_315), .B1(n_362), .B2(n_306), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_457), .Y(n_480) );
INVx3_ASAP7_75t_L g481 ( .A(n_464), .Y(n_481) );
AND2x4_ASAP7_75t_L g482 ( .A(n_464), .B(n_439), .Y(n_482) );
OAI22xp5_ASAP7_75t_L g483 ( .A1(n_455), .A2(n_436), .B1(n_387), .B2(n_315), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_470), .B(n_350), .Y(n_484) );
AND2x6_ASAP7_75t_L g485 ( .A(n_464), .B(n_352), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g486 ( .A(n_462), .B(n_367), .Y(n_486) );
INVx2_ASAP7_75t_L g487 ( .A(n_457), .Y(n_487) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_465), .Y(n_488) );
AND2x6_ASAP7_75t_L g489 ( .A(n_464), .B(n_352), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_457), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_457), .B(n_314), .Y(n_491) );
BUFx6f_ASAP7_75t_L g492 ( .A(n_465), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_459), .B(n_314), .Y(n_493) );
NOR2xp33_ASAP7_75t_L g494 ( .A(n_476), .B(n_368), .Y(n_494) );
AND2x4_ASAP7_75t_L g495 ( .A(n_464), .B(n_307), .Y(n_495) );
BUFx3_ASAP7_75t_L g496 ( .A(n_452), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_452), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
AND2x4_ASAP7_75t_L g499 ( .A(n_456), .B(n_307), .Y(n_499) );
NOR2xp33_ASAP7_75t_L g500 ( .A(n_460), .B(n_444), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_451), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_451), .Y(n_502) );
BUFx6f_ASAP7_75t_L g503 ( .A(n_465), .Y(n_503) );
NOR2xp33_ASAP7_75t_R g504 ( .A(n_460), .B(n_309), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_487), .Y(n_505) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_496), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_491), .B(n_493), .Y(n_507) );
BUFx4f_ASAP7_75t_L g508 ( .A(n_485), .Y(n_508) );
NOR2xp33_ASAP7_75t_SL g509 ( .A(n_477), .B(n_467), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_485), .B(n_459), .Y(n_510) );
INVx5_ASAP7_75t_L g511 ( .A(n_485), .Y(n_511) );
INVx2_ASAP7_75t_L g512 ( .A(n_487), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g513 ( .A1(n_481), .A2(n_468), .B(n_461), .Y(n_513) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_485), .A2(n_467), .B1(n_451), .B2(n_453), .Y(n_514) );
CKINVDCx5p33_ASAP7_75t_R g515 ( .A(n_504), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_481), .Y(n_516) );
HB1xp67_ASAP7_75t_L g517 ( .A(n_484), .Y(n_517) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_482), .B(n_345), .Y(n_518) );
NOR2x1_ASAP7_75t_R g519 ( .A(n_478), .B(n_450), .Y(n_519) );
NAND2xp5_ASAP7_75t_L g520 ( .A(n_485), .B(n_468), .Y(n_520) );
BUFx3_ASAP7_75t_L g521 ( .A(n_485), .Y(n_521) );
BUFx12f_ASAP7_75t_L g522 ( .A(n_482), .Y(n_522) );
INVx2_ASAP7_75t_L g523 ( .A(n_480), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g524 ( .A1(n_489), .A2(n_467), .B1(n_451), .B2(n_453), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_480), .Y(n_525) );
AND2x4_ASAP7_75t_L g526 ( .A(n_478), .B(n_467), .Y(n_526) );
INVx1_ASAP7_75t_L g527 ( .A(n_490), .Y(n_527) );
INVx3_ASAP7_75t_L g528 ( .A(n_495), .Y(n_528) );
BUFx10_ASAP7_75t_L g529 ( .A(n_489), .Y(n_529) );
CKINVDCx11_ASAP7_75t_R g530 ( .A(n_483), .Y(n_530) );
AO22x1_ASAP7_75t_L g531 ( .A1(n_489), .A2(n_371), .B1(n_377), .B2(n_369), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_501), .A2(n_461), .B(n_467), .Y(n_532) );
AND2x4_ASAP7_75t_L g533 ( .A(n_478), .B(n_467), .Y(n_533) );
OR2x6_ASAP7_75t_L g534 ( .A(n_495), .B(n_469), .Y(n_534) );
INVx5_ASAP7_75t_L g535 ( .A(n_489), .Y(n_535) );
INVx1_ASAP7_75t_L g536 ( .A(n_490), .Y(n_536) );
BUFx2_ASAP7_75t_L g537 ( .A(n_489), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_501), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_495), .B(n_469), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_496), .B(n_420), .Y(n_540) );
OR2x4_ASAP7_75t_L g541 ( .A(n_486), .B(n_317), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_497), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_495), .B(n_420), .Y(n_543) );
BUFx3_ASAP7_75t_L g544 ( .A(n_502), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_499), .B(n_370), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_499), .B(n_425), .Y(n_546) );
INVx5_ASAP7_75t_L g547 ( .A(n_488), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_494), .B(n_425), .Y(n_548) );
INVx2_ASAP7_75t_L g549 ( .A(n_502), .Y(n_549) );
AOI22xp5_ASAP7_75t_L g550 ( .A1(n_479), .A2(n_463), .B1(n_499), .B2(n_498), .Y(n_550) );
AND2x4_ASAP7_75t_L g551 ( .A(n_498), .B(n_372), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_500), .B(n_451), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_503), .A2(n_453), .B1(n_451), .B2(n_463), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_488), .Y(n_554) );
BUFx8_ASAP7_75t_L g555 ( .A(n_488), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_488), .Y(n_556) );
BUFx6f_ASAP7_75t_L g557 ( .A(n_492), .Y(n_557) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_492), .B(n_369), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_492), .Y(n_559) );
BUFx3_ASAP7_75t_L g560 ( .A(n_555), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_538), .A2(n_453), .B(n_312), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_538), .A2(n_453), .B(n_357), .Y(n_562) );
AOI21xp5_ASAP7_75t_L g563 ( .A1(n_549), .A2(n_453), .B(n_378), .Y(n_563) );
AOI21xp5_ASAP7_75t_L g564 ( .A1(n_549), .A2(n_443), .B(n_311), .Y(n_564) );
NAND2x1p5_ASAP7_75t_L g565 ( .A(n_511), .B(n_321), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_528), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g567 ( .A1(n_509), .A2(n_471), .B1(n_310), .B2(n_374), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_541), .B(n_306), .Y(n_568) );
INVx4_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_517), .B(n_454), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_539), .B(n_322), .Y(n_571) );
AOI22xp5_ASAP7_75t_L g572 ( .A1(n_526), .A2(n_458), .B1(n_454), .B2(n_400), .Y(n_572) );
INVx1_ASAP7_75t_L g573 ( .A(n_528), .Y(n_573) );
INVx5_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
INVxp67_ASAP7_75t_L g575 ( .A(n_519), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_542), .Y(n_576) );
AO21x1_ASAP7_75t_L g577 ( .A1(n_532), .A2(n_328), .B(n_327), .Y(n_577) );
INVx4_ASAP7_75t_L g578 ( .A(n_511), .Y(n_578) );
INVx3_ASAP7_75t_L g579 ( .A(n_555), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g580 ( .A(n_541), .B(n_362), .Y(n_580) );
INVx3_ASAP7_75t_L g581 ( .A(n_555), .Y(n_581) );
AND2x2_ASAP7_75t_L g582 ( .A(n_551), .B(n_458), .Y(n_582) );
AOI22xp33_ASAP7_75t_L g583 ( .A1(n_526), .A2(n_400), .B1(n_371), .B2(n_377), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g584 ( .A(n_515), .Y(n_584) );
INVx2_ASAP7_75t_L g585 ( .A(n_544), .Y(n_585) );
OA22x2_ASAP7_75t_L g586 ( .A1(n_550), .A2(n_339), .B1(n_376), .B2(n_334), .Y(n_586) );
NOR2xp33_ASAP7_75t_SL g587 ( .A(n_508), .B(n_519), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_525), .Y(n_588) );
O2A1O1Ixp5_ASAP7_75t_L g589 ( .A1(n_518), .A2(n_349), .B(n_366), .C(n_337), .Y(n_589) );
BUFx6f_ASAP7_75t_L g590 ( .A(n_544), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g591 ( .A1(n_526), .A2(n_533), .B1(n_539), .B2(n_552), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_551), .B(n_545), .Y(n_592) );
INVx1_ASAP7_75t_SL g593 ( .A(n_551), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_544), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_516), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_507), .A2(n_328), .B(n_327), .Y(n_596) );
BUFx4_ASAP7_75t_SL g597 ( .A(n_534), .Y(n_597) );
OR2x6_ASAP7_75t_L g598 ( .A(n_521), .B(n_428), .Y(n_598) );
AND2x2_ASAP7_75t_SL g599 ( .A(n_508), .B(n_317), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_555), .Y(n_600) );
CKINVDCx6p67_ASAP7_75t_R g601 ( .A(n_511), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_526), .B(n_334), .Y(n_602) );
INVx6_ASAP7_75t_L g603 ( .A(n_522), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
AOI21xp5_ASAP7_75t_L g605 ( .A1(n_516), .A2(n_336), .B(n_329), .Y(n_605) );
INVx2_ASAP7_75t_SL g606 ( .A(n_511), .Y(n_606) );
INVx3_ASAP7_75t_L g607 ( .A(n_529), .Y(n_607) );
AOI21xp5_ASAP7_75t_L g608 ( .A1(n_527), .A2(n_336), .B(n_329), .Y(n_608) );
INVx3_ASAP7_75t_L g609 ( .A(n_529), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_536), .A2(n_342), .B(n_340), .Y(n_610) );
INVx1_ASAP7_75t_SL g611 ( .A(n_546), .Y(n_611) );
INVx2_ASAP7_75t_SL g612 ( .A(n_535), .Y(n_612) );
OR2x6_ASAP7_75t_L g613 ( .A(n_521), .B(n_331), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_533), .B(n_353), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_523), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_534), .Y(n_616) );
BUFx8_ASAP7_75t_SL g617 ( .A(n_508), .Y(n_617) );
INVx4_ASAP7_75t_L g618 ( .A(n_535), .Y(n_618) );
BUFx3_ASAP7_75t_L g619 ( .A(n_506), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_533), .B(n_394), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_550), .B(n_397), .Y(n_621) );
INVx1_ASAP7_75t_SL g622 ( .A(n_534), .Y(n_622) );
OR2x6_ASAP7_75t_L g623 ( .A(n_537), .B(n_319), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_537), .Y(n_624) );
BUFx12f_ASAP7_75t_L g625 ( .A(n_530), .Y(n_625) );
INVx6_ASAP7_75t_L g626 ( .A(n_506), .Y(n_626) );
AND2x4_ASAP7_75t_L g627 ( .A(n_535), .B(n_359), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_510), .Y(n_628) );
BUFx6f_ASAP7_75t_L g629 ( .A(n_506), .Y(n_629) );
A2O1A1Ixp33_ASAP7_75t_L g630 ( .A1(n_552), .A2(n_323), .B(n_326), .C(n_320), .Y(n_630) );
BUFx6f_ASAP7_75t_L g631 ( .A(n_506), .Y(n_631) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_520), .A2(n_342), .B(n_340), .Y(n_632) );
INVx3_ASAP7_75t_L g633 ( .A(n_529), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_531), .B(n_405), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_592), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_593), .B(n_531), .Y(n_636) );
OAI22xp5_ASAP7_75t_L g637 ( .A1(n_591), .A2(n_514), .B1(n_524), .B2(n_543), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g638 ( .A1(n_623), .A2(n_541), .B1(n_326), .B2(n_330), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_591), .A2(n_540), .B1(n_553), .B2(n_513), .Y(n_639) );
OAI22xp5_ASAP7_75t_L g640 ( .A1(n_623), .A2(n_512), .B1(n_505), .B2(n_558), .Y(n_640) );
AOI21xp33_ASAP7_75t_L g641 ( .A1(n_568), .A2(n_548), .B(n_512), .Y(n_641) );
AOI22xp33_ASAP7_75t_L g642 ( .A1(n_586), .A2(n_321), .B1(n_418), .B2(n_408), .Y(n_642) );
INVx4_ASAP7_75t_L g643 ( .A(n_560), .Y(n_643) );
BUFx6f_ASAP7_75t_L g644 ( .A(n_590), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_614), .B(n_373), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_586), .A2(n_418), .B1(n_408), .B2(n_333), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_615), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_561), .A2(n_556), .B(n_554), .Y(n_648) );
INVx4_ASAP7_75t_L g649 ( .A(n_600), .Y(n_649) );
BUFx2_ASAP7_75t_L g650 ( .A(n_623), .Y(n_650) );
CKINVDCx5p33_ASAP7_75t_R g651 ( .A(n_625), .Y(n_651) );
AOI22xp5_ASAP7_75t_L g652 ( .A1(n_582), .A2(n_570), .B1(n_567), .B2(n_572), .Y(n_652) );
AO21x2_ASAP7_75t_L g653 ( .A1(n_577), .A2(n_351), .B(n_346), .Y(n_653) );
AOI21xp5_ASAP7_75t_L g654 ( .A1(n_562), .A2(n_556), .B(n_554), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_603), .B(n_325), .Y(n_655) );
CKINVDCx5p33_ASAP7_75t_R g656 ( .A(n_584), .Y(n_656) );
HB1xp67_ASAP7_75t_L g657 ( .A(n_597), .Y(n_657) );
AOI22xp33_ASAP7_75t_L g658 ( .A1(n_621), .A2(n_440), .B1(n_333), .B2(n_381), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_581), .Y(n_659) );
A2O1A1Ixp33_ASAP7_75t_L g660 ( .A1(n_576), .A2(n_332), .B(n_343), .C(n_341), .Y(n_660) );
O2A1O1Ixp33_ASAP7_75t_L g661 ( .A1(n_630), .A2(n_382), .B(n_383), .C(n_380), .Y(n_661) );
AOI221xp5_ASAP7_75t_L g662 ( .A1(n_568), .A2(n_390), .B1(n_391), .B2(n_388), .C(n_386), .Y(n_662) );
AND2x4_ASAP7_75t_L g663 ( .A(n_581), .B(n_332), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_583), .B(n_393), .Y(n_664) );
AOI22xp33_ASAP7_75t_SL g665 ( .A1(n_599), .A2(n_341), .B1(n_348), .B2(n_343), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g666 ( .A1(n_580), .A2(n_395), .B1(n_402), .B2(n_399), .C(n_396), .Y(n_666) );
AOI22xp33_ASAP7_75t_L g667 ( .A1(n_580), .A2(n_440), .B1(n_404), .B2(n_410), .Y(n_667) );
BUFx6f_ASAP7_75t_L g668 ( .A(n_590), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_588), .Y(n_669) );
INVx3_ASAP7_75t_L g670 ( .A(n_579), .Y(n_670) );
INVx2_ASAP7_75t_L g671 ( .A(n_595), .Y(n_671) );
AO21x2_ASAP7_75t_L g672 ( .A1(n_563), .A2(n_354), .B(n_351), .Y(n_672) );
INVx3_ASAP7_75t_L g673 ( .A(n_569), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_604), .Y(n_674) );
AOI22xp33_ASAP7_75t_SL g675 ( .A1(n_587), .A2(n_431), .B1(n_433), .B2(n_430), .Y(n_675) );
O2A1O1Ixp5_ASAP7_75t_SL g676 ( .A1(n_575), .A2(n_356), .B(n_432), .C(n_355), .Y(n_676) );
AOI22xp33_ASAP7_75t_L g677 ( .A1(n_634), .A2(n_413), .B1(n_421), .B2(n_412), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_622), .A2(n_434), .B1(n_435), .B2(n_433), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_616), .B(n_434), .Y(n_679) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_571), .A2(n_424), .B1(n_426), .B2(n_422), .Y(n_680) );
AND2x4_ASAP7_75t_L g681 ( .A(n_611), .B(n_435), .Y(n_681) );
INVx4_ASAP7_75t_L g682 ( .A(n_574), .Y(n_682) );
INVx2_ASAP7_75t_L g683 ( .A(n_566), .Y(n_683) );
NOR2xp33_ASAP7_75t_L g684 ( .A(n_602), .B(n_427), .Y(n_684) );
AOI21xp5_ASAP7_75t_L g685 ( .A1(n_596), .A2(n_559), .B(n_557), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g686 ( .A1(n_627), .A2(n_442), .B1(n_445), .B2(n_441), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_573), .Y(n_687) );
A2O1A1Ixp33_ASAP7_75t_L g688 ( .A1(n_630), .A2(n_446), .B(n_447), .C(n_445), .Y(n_688) );
NAND2xp33_ASAP7_75t_SL g689 ( .A(n_624), .B(n_446), .Y(n_689) );
NAND2xp5_ASAP7_75t_SL g690 ( .A(n_585), .B(n_547), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_620), .B(n_447), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_627), .Y(n_692) );
CKINVDCx8_ASAP7_75t_R g693 ( .A(n_627), .Y(n_693) );
CKINVDCx5p33_ASAP7_75t_R g694 ( .A(n_617), .Y(n_694) );
OR2x2_ASAP7_75t_L g695 ( .A(n_598), .B(n_398), .Y(n_695) );
CKINVDCx16_ASAP7_75t_R g696 ( .A(n_613), .Y(n_696) );
CKINVDCx5p33_ASAP7_75t_R g697 ( .A(n_617), .Y(n_697) );
AND2x6_ASAP7_75t_L g698 ( .A(n_594), .B(n_438), .Y(n_698) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_628), .A2(n_403), .B1(n_406), .B2(n_398), .Y(n_699) );
OAI21x1_ASAP7_75t_L g700 ( .A1(n_565), .A2(n_559), .B(n_349), .Y(n_700) );
INVx6_ASAP7_75t_L g701 ( .A(n_574), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_613), .B(n_409), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_608), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_610), .Y(n_704) );
OR2x2_ASAP7_75t_L g705 ( .A(n_565), .B(n_8), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_601), .A2(n_360), .B1(n_365), .B2(n_364), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_647), .Y(n_707) );
OAI22xp33_ASAP7_75t_L g708 ( .A1(n_696), .A2(n_601), .B1(n_631), .B2(n_629), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_635), .B(n_564), .Y(n_709) );
OAI211xp5_ASAP7_75t_SL g710 ( .A1(n_652), .A2(n_589), .B(n_384), .C(n_385), .Y(n_710) );
AND2x2_ASAP7_75t_L g711 ( .A(n_681), .B(n_605), .Y(n_711) );
AOI332xp33_ASAP7_75t_L g712 ( .A1(n_677), .A2(n_417), .A3(n_379), .B1(n_392), .B2(n_401), .B3(n_449), .C1(n_411), .C2(n_429), .Y(n_712) );
OA21x2_ASAP7_75t_L g713 ( .A1(n_648), .A2(n_654), .B(n_685), .Y(n_713) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_662), .A2(n_632), .B1(n_423), .B2(n_416), .C(n_414), .Y(n_714) );
OAI22xp33_ASAP7_75t_L g715 ( .A1(n_650), .A2(n_631), .B1(n_629), .B2(n_578), .Y(n_715) );
AND2x2_ASAP7_75t_L g716 ( .A(n_681), .B(n_9), .Y(n_716) );
OAI22xp33_ASAP7_75t_L g717 ( .A1(n_655), .A2(n_631), .B1(n_629), .B2(n_578), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_665), .B(n_9), .Y(n_718) );
AOI221xp5_ASAP7_75t_SL g719 ( .A1(n_638), .A2(n_389), .B1(n_419), .B2(n_366), .C(n_337), .Y(n_719) );
AO221x2_ASAP7_75t_L g720 ( .A1(n_638), .A2(n_437), .B1(n_419), .B2(n_389), .C(n_12), .Y(n_720) );
OAI21x1_ASAP7_75t_L g721 ( .A1(n_654), .A2(n_607), .B(n_609), .Y(n_721) );
BUFx3_ASAP7_75t_L g722 ( .A(n_643), .Y(n_722) );
AOI22xp33_ASAP7_75t_L g723 ( .A1(n_665), .A2(n_619), .B1(n_626), .B2(n_606), .Y(n_723) );
OR2x6_ASAP7_75t_L g724 ( .A(n_657), .B(n_578), .Y(n_724) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_684), .A2(n_626), .B1(n_612), .B2(n_618), .Y(n_725) );
OA21x2_ASAP7_75t_L g726 ( .A1(n_685), .A2(n_472), .B(n_466), .Y(n_726) );
OAI22xp5_ASAP7_75t_L g727 ( .A1(n_693), .A2(n_626), .B1(n_631), .B2(n_629), .Y(n_727) );
AO31x2_ASAP7_75t_L g728 ( .A1(n_639), .A2(n_466), .A3(n_473), .B(n_472), .Y(n_728) );
INVx2_ASAP7_75t_L g729 ( .A(n_671), .Y(n_729) );
BUFx12f_ASAP7_75t_L g730 ( .A(n_651), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_684), .A2(n_618), .B1(n_607), .B2(n_609), .Y(n_731) );
OAI221xp5_ASAP7_75t_L g732 ( .A1(n_666), .A2(n_633), .B1(n_472), .B2(n_474), .C(n_473), .Y(n_732) );
OAI22xp5_ASAP7_75t_L g733 ( .A1(n_655), .A2(n_466), .B1(n_473), .B2(n_472), .Y(n_733) );
INVx1_ASAP7_75t_L g734 ( .A(n_669), .Y(n_734) );
NOR2xp33_ASAP7_75t_L g735 ( .A(n_664), .B(n_10), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_689), .A2(n_547), .B1(n_474), .B2(n_557), .Y(n_736) );
INVx3_ASAP7_75t_L g737 ( .A(n_682), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_642), .A2(n_465), .B1(n_557), .B2(n_547), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_658), .A2(n_547), .B1(n_557), .B2(n_13), .Y(n_739) );
OA21x2_ASAP7_75t_L g740 ( .A1(n_700), .A2(n_503), .B(n_492), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g741 ( .A1(n_658), .A2(n_15), .B1(n_11), .B2(n_14), .Y(n_741) );
AOI21x1_ASAP7_75t_L g742 ( .A1(n_640), .A2(n_503), .B(n_204), .Y(n_742) );
OAI221xp5_ASAP7_75t_L g743 ( .A1(n_680), .A2(n_642), .B1(n_675), .B2(n_646), .C(n_667), .Y(n_743) );
OAI22xp5_ASAP7_75t_L g744 ( .A1(n_686), .A2(n_18), .B1(n_16), .B2(n_17), .Y(n_744) );
INVx1_ASAP7_75t_L g745 ( .A(n_674), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_663), .Y(n_746) );
OAI211xp5_ASAP7_75t_L g747 ( .A1(n_646), .A2(n_503), .B(n_20), .C(n_18), .Y(n_747) );
OAI22xp33_ASAP7_75t_L g748 ( .A1(n_705), .A2(n_21), .B1(n_19), .B2(n_20), .Y(n_748) );
INVx3_ASAP7_75t_L g749 ( .A(n_682), .Y(n_749) );
OR2x6_ASAP7_75t_L g750 ( .A(n_649), .B(n_24), .Y(n_750) );
AOI221xp5_ASAP7_75t_L g751 ( .A1(n_661), .A2(n_26), .B1(n_24), .B2(n_25), .C(n_27), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_695), .Y(n_752) );
INVx1_ASAP7_75t_L g753 ( .A(n_645), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g754 ( .A(n_667), .B(n_28), .Y(n_754) );
AOI22xp33_ASAP7_75t_L g755 ( .A1(n_637), .A2(n_31), .B1(n_29), .B2(n_30), .Y(n_755) );
AOI22xp33_ASAP7_75t_L g756 ( .A1(n_703), .A2(n_34), .B1(n_32), .B2(n_33), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_644), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_644), .Y(n_758) );
INVx2_ASAP7_75t_L g759 ( .A(n_644), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_704), .A2(n_37), .B1(n_35), .B2(n_36), .Y(n_760) );
AO31x2_ASAP7_75t_L g761 ( .A1(n_688), .A2(n_38), .A3(n_36), .B(n_37), .Y(n_761) );
INVx2_ASAP7_75t_L g762 ( .A(n_668), .Y(n_762) );
AOI22xp33_ASAP7_75t_L g763 ( .A1(n_679), .A2(n_702), .B1(n_678), .B2(n_691), .Y(n_763) );
AOI221xp5_ASAP7_75t_L g764 ( .A1(n_661), .A2(n_40), .B1(n_38), .B2(n_39), .C(n_41), .Y(n_764) );
INVx1_ASAP7_75t_L g765 ( .A(n_687), .Y(n_765) );
OAI221xp5_ASAP7_75t_SL g766 ( .A1(n_688), .A2(n_42), .B1(n_40), .B2(n_41), .C(n_43), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g767 ( .A1(n_660), .A2(n_44), .B1(n_42), .B2(n_43), .C(n_45), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_692), .A2(n_46), .B1(n_44), .B2(n_45), .Y(n_768) );
OR3x1_ASAP7_75t_L g769 ( .A(n_641), .B(n_47), .C(n_48), .Y(n_769) );
OAI22xp33_ASAP7_75t_L g770 ( .A1(n_636), .A2(n_51), .B1(n_49), .B2(n_50), .Y(n_770) );
AOI22xp33_ASAP7_75t_L g771 ( .A1(n_699), .A2(n_53), .B1(n_51), .B2(n_52), .Y(n_771) );
AO21x2_ASAP7_75t_L g772 ( .A1(n_653), .A2(n_207), .B(n_206), .Y(n_772) );
OAI22xp33_ASAP7_75t_L g773 ( .A1(n_706), .A2(n_55), .B1(n_53), .B2(n_54), .Y(n_773) );
NAND3xp33_ASAP7_75t_SL g774 ( .A(n_656), .B(n_54), .C(n_55), .Y(n_774) );
INVx2_ASAP7_75t_L g775 ( .A(n_672), .Y(n_775) );
NOR2xp33_ASAP7_75t_SL g776 ( .A(n_694), .B(n_57), .Y(n_776) );
INVx2_ASAP7_75t_L g777 ( .A(n_707), .Y(n_777) );
INVx3_ASAP7_75t_L g778 ( .A(n_722), .Y(n_778) );
OAI33xp33_ASAP7_75t_L g779 ( .A1(n_748), .A2(n_683), .A3(n_690), .B1(n_676), .B2(n_697), .B3(n_653), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_707), .Y(n_780) );
NOR3xp33_ASAP7_75t_L g781 ( .A(n_774), .B(n_659), .C(n_670), .Y(n_781) );
OR2x2_ASAP7_75t_L g782 ( .A(n_752), .B(n_673), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g783 ( .A(n_743), .B(n_698), .Y(n_783) );
OAI33xp33_ASAP7_75t_L g784 ( .A1(n_773), .A2(n_698), .A3(n_60), .B1(n_62), .B2(n_57), .B3(n_58), .Y(n_784) );
OAI22xp5_ASAP7_75t_L g785 ( .A1(n_763), .A2(n_701), .B1(n_698), .B2(n_61), .Y(n_785) );
AOI21xp5_ASAP7_75t_L g786 ( .A1(n_717), .A2(n_708), .B(n_715), .Y(n_786) );
AND2x4_ASAP7_75t_L g787 ( .A(n_722), .B(n_65), .Y(n_787) );
OR2x6_ASAP7_75t_L g788 ( .A(n_750), .B(n_67), .Y(n_788) );
OAI211xp5_ASAP7_75t_L g789 ( .A1(n_712), .A2(n_71), .B(n_68), .C(n_69), .Y(n_789) );
NAND2xp5_ASAP7_75t_L g790 ( .A(n_753), .B(n_72), .Y(n_790) );
AOI22xp33_ASAP7_75t_SL g791 ( .A1(n_720), .A2(n_75), .B1(n_73), .B2(n_74), .Y(n_791) );
AND2x2_ASAP7_75t_L g792 ( .A(n_716), .B(n_76), .Y(n_792) );
INVx2_ASAP7_75t_L g793 ( .A(n_729), .Y(n_793) );
INVx2_ASAP7_75t_L g794 ( .A(n_729), .Y(n_794) );
INVx1_ASAP7_75t_L g795 ( .A(n_734), .Y(n_795) );
AND2x2_ASAP7_75t_L g796 ( .A(n_718), .B(n_77), .Y(n_796) );
NAND2xp33_ASAP7_75t_R g797 ( .A(n_740), .B(n_78), .Y(n_797) );
AND2x4_ASAP7_75t_L g798 ( .A(n_737), .B(n_81), .Y(n_798) );
INVx1_ASAP7_75t_L g799 ( .A(n_745), .Y(n_799) );
OAI22xp33_ASAP7_75t_SL g800 ( .A1(n_776), .A2(n_85), .B1(n_83), .B2(n_84), .Y(n_800) );
INVx2_ASAP7_75t_L g801 ( .A(n_765), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g802 ( .A1(n_720), .A2(n_89), .B1(n_87), .B2(n_88), .Y(n_802) );
AO21x2_ASAP7_75t_L g803 ( .A1(n_775), .A2(n_87), .B(n_90), .Y(n_803) );
INVx2_ASAP7_75t_L g804 ( .A(n_728), .Y(n_804) );
BUFx2_ASAP7_75t_L g805 ( .A(n_724), .Y(n_805) );
OAI321xp33_ASAP7_75t_L g806 ( .A1(n_766), .A2(n_94), .A3(n_95), .B1(n_96), .B2(n_97), .C(n_98), .Y(n_806) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_735), .A2(n_99), .B1(n_95), .B2(n_97), .Y(n_807) );
INVxp67_ASAP7_75t_SL g808 ( .A(n_717), .Y(n_808) );
INVx3_ASAP7_75t_L g809 ( .A(n_737), .Y(n_809) );
OR2x6_ASAP7_75t_L g810 ( .A(n_749), .B(n_103), .Y(n_810) );
INVx1_ASAP7_75t_L g811 ( .A(n_761), .Y(n_811) );
OAI33xp33_ASAP7_75t_L g812 ( .A1(n_770), .A2(n_106), .A3(n_107), .B1(n_108), .B2(n_109), .B3(n_110), .Y(n_812) );
INVx5_ASAP7_75t_SL g813 ( .A(n_730), .Y(n_813) );
AOI221xp5_ASAP7_75t_L g814 ( .A1(n_744), .A2(n_107), .B1(n_108), .B2(n_109), .C(n_111), .Y(n_814) );
OA21x2_ASAP7_75t_L g815 ( .A1(n_719), .A2(n_213), .B(n_212), .Y(n_815) );
AOI33xp33_ASAP7_75t_L g816 ( .A1(n_755), .A2(n_112), .A3(n_113), .B1(n_114), .B2(n_115), .B3(n_116), .Y(n_816) );
OAI22xp5_ASAP7_75t_L g817 ( .A1(n_723), .A2(n_117), .B1(n_114), .B2(n_116), .Y(n_817) );
NOR2x1_ASAP7_75t_L g818 ( .A(n_769), .B(n_117), .Y(n_818) );
INVx2_ASAP7_75t_L g819 ( .A(n_728), .Y(n_819) );
OA21x2_ASAP7_75t_L g820 ( .A1(n_721), .A2(n_218), .B(n_214), .Y(n_820) );
AO21x2_ASAP7_75t_L g821 ( .A1(n_742), .A2(n_119), .B(n_120), .Y(n_821) );
INVx1_ASAP7_75t_L g822 ( .A(n_761), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_711), .A2(n_122), .B1(n_120), .B2(n_121), .Y(n_823) );
OAI221xp5_ASAP7_75t_L g824 ( .A1(n_755), .A2(n_121), .B1(n_123), .B2(n_124), .C(n_125), .Y(n_824) );
INVxp67_ASAP7_75t_SL g825 ( .A(n_708), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g826 ( .A1(n_751), .A2(n_129), .B1(n_126), .B2(n_128), .Y(n_826) );
AO21x2_ASAP7_75t_L g827 ( .A1(n_715), .A2(n_126), .B(n_130), .Y(n_827) );
OAI22xp33_ASAP7_75t_L g828 ( .A1(n_767), .A2(n_134), .B1(n_132), .B2(n_133), .Y(n_828) );
AOI22xp33_ASAP7_75t_L g829 ( .A1(n_764), .A2(n_137), .B1(n_133), .B2(n_135), .Y(n_829) );
OAI22xp5_ASAP7_75t_L g830 ( .A1(n_725), .A2(n_140), .B1(n_138), .B2(n_139), .Y(n_830) );
NAND2xp5_ASAP7_75t_L g831 ( .A(n_746), .B(n_139), .Y(n_831) );
INVx5_ASAP7_75t_SL g832 ( .A(n_772), .Y(n_832) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_710), .A2(n_145), .B1(n_143), .B2(n_144), .Y(n_833) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_757), .Y(n_834) );
OAI221xp5_ASAP7_75t_L g835 ( .A1(n_771), .A2(n_145), .B1(n_146), .B2(n_147), .C(n_148), .Y(n_835) );
INVx2_ASAP7_75t_L g836 ( .A(n_728), .Y(n_836) );
INVx2_ASAP7_75t_L g837 ( .A(n_728), .Y(n_837) );
INVx1_ASAP7_75t_L g838 ( .A(n_761), .Y(n_838) );
AND2x2_ASAP7_75t_SL g839 ( .A(n_738), .B(n_152), .Y(n_839) );
INVx2_ASAP7_75t_L g840 ( .A(n_726), .Y(n_840) );
INVx2_ASAP7_75t_L g841 ( .A(n_726), .Y(n_841) );
AOI22xp33_ASAP7_75t_L g842 ( .A1(n_741), .A2(n_153), .B1(n_154), .B2(n_155), .Y(n_842) );
HB1xp67_ASAP7_75t_L g843 ( .A(n_757), .Y(n_843) );
OAI221xp5_ASAP7_75t_SL g844 ( .A1(n_802), .A2(n_756), .B1(n_760), .B2(n_768), .C(n_747), .Y(n_844) );
NAND3xp33_ASAP7_75t_L g845 ( .A(n_791), .B(n_714), .C(n_733), .Y(n_845) );
OAI33xp33_ASAP7_75t_L g846 ( .A1(n_800), .A2(n_754), .A3(n_709), .B1(n_739), .B2(n_727), .B3(n_157), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_792), .B(n_154), .Y(n_847) );
INVx5_ASAP7_75t_L g848 ( .A(n_788), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_795), .Y(n_849) );
OAI221xp5_ASAP7_75t_SL g850 ( .A1(n_802), .A2(n_731), .B1(n_736), .B2(n_732), .C(n_762), .Y(n_850) );
INVx2_ASAP7_75t_L g851 ( .A(n_777), .Y(n_851) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_799), .B(n_713), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_801), .Y(n_853) );
AND2x2_ASAP7_75t_L g854 ( .A(n_796), .B(n_158), .Y(n_854) );
INVx1_ASAP7_75t_SL g855 ( .A(n_778), .Y(n_855) );
NOR3xp33_ASAP7_75t_L g856 ( .A(n_789), .B(n_759), .C(n_758), .Y(n_856) );
INVxp67_ASAP7_75t_L g857 ( .A(n_797), .Y(n_857) );
AND2x4_ASAP7_75t_L g858 ( .A(n_778), .B(n_805), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_787), .B(n_159), .Y(n_859) );
HB1xp67_ASAP7_75t_L g860 ( .A(n_834), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_782), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_780), .Y(n_862) );
OAI33xp33_ASAP7_75t_L g863 ( .A1(n_828), .A2(n_161), .A3(n_162), .B1(n_163), .B2(n_164), .B3(n_165), .Y(n_863) );
INVxp67_ASAP7_75t_SL g864 ( .A(n_797), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_810), .Y(n_865) );
HB1xp67_ASAP7_75t_L g866 ( .A(n_834), .Y(n_866) );
INVx3_ASAP7_75t_L g867 ( .A(n_809), .Y(n_867) );
NAND2xp5_ASAP7_75t_L g868 ( .A(n_811), .B(n_740), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_798), .Y(n_869) );
OAI33xp33_ASAP7_75t_L g870 ( .A1(n_830), .A2(n_166), .A3(n_167), .B1(n_168), .B2(n_169), .B3(n_170), .Y(n_870) );
HB1xp67_ASAP7_75t_L g871 ( .A(n_843), .Y(n_871) );
INVxp67_ASAP7_75t_SL g872 ( .A(n_840), .Y(n_872) );
INVxp67_ASAP7_75t_SL g873 ( .A(n_841), .Y(n_873) );
OR2x6_ASAP7_75t_L g874 ( .A(n_786), .B(n_171), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g875 ( .A(n_822), .B(n_838), .Y(n_875) );
OR2x2_ASAP7_75t_L g876 ( .A(n_793), .B(n_794), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g877 ( .A(n_843), .B(n_175), .Y(n_877) );
BUFx2_ASAP7_75t_L g878 ( .A(n_809), .Y(n_878) );
AOI211xp5_ASAP7_75t_SL g879 ( .A1(n_806), .A2(n_177), .B(n_179), .C(n_180), .Y(n_879) );
OR2x6_ASAP7_75t_L g880 ( .A(n_785), .B(n_177), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_818), .B(n_181), .C(n_182), .Y(n_881) );
INVx4_ASAP7_75t_L g882 ( .A(n_839), .Y(n_882) );
INVx1_ASAP7_75t_L g883 ( .A(n_790), .Y(n_883) );
AND2x2_ASAP7_75t_L g884 ( .A(n_823), .B(n_183), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_825), .B(n_184), .Y(n_885) );
INVx1_ASAP7_75t_L g886 ( .A(n_803), .Y(n_886) );
BUFx6f_ASAP7_75t_L g887 ( .A(n_804), .Y(n_887) );
INVx2_ASAP7_75t_L g888 ( .A(n_819), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_816), .Y(n_889) );
INVx3_ASAP7_75t_L g890 ( .A(n_827), .Y(n_890) );
INVx1_ASAP7_75t_L g891 ( .A(n_816), .Y(n_891) );
OAI21xp5_ASAP7_75t_SL g892 ( .A1(n_807), .A2(n_185), .B(n_186), .Y(n_892) );
INVx2_ASAP7_75t_L g893 ( .A(n_836), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_823), .B(n_187), .Y(n_894) );
INVx1_ASAP7_75t_L g895 ( .A(n_827), .Y(n_895) );
INVx5_ASAP7_75t_L g896 ( .A(n_813), .Y(n_896) );
AO22x1_ASAP7_75t_L g897 ( .A1(n_825), .A2(n_188), .B1(n_189), .B2(n_190), .Y(n_897) );
AND2x4_ASAP7_75t_L g898 ( .A(n_808), .B(n_191), .Y(n_898) );
INVx1_ASAP7_75t_SL g899 ( .A(n_831), .Y(n_899) );
INVx2_ASAP7_75t_L g900 ( .A(n_837), .Y(n_900) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_783), .B(n_808), .Y(n_901) );
INVx2_ASAP7_75t_L g902 ( .A(n_821), .Y(n_902) );
INVx1_ASAP7_75t_L g903 ( .A(n_817), .Y(n_903) );
AND2x2_ASAP7_75t_L g904 ( .A(n_861), .B(n_197), .Y(n_904) );
INVx5_ASAP7_75t_L g905 ( .A(n_896), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_849), .Y(n_906) );
INVx2_ASAP7_75t_L g907 ( .A(n_876), .Y(n_907) );
INVx3_ASAP7_75t_L g908 ( .A(n_848), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_853), .B(n_199), .Y(n_909) );
AND2x2_ASAP7_75t_L g910 ( .A(n_855), .B(n_199), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_877), .Y(n_911) );
INVx1_ASAP7_75t_L g912 ( .A(n_877), .Y(n_912) );
NAND2xp5_ASAP7_75t_L g913 ( .A(n_852), .B(n_826), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_860), .B(n_201), .Y(n_914) );
INVx2_ASAP7_75t_SL g915 ( .A(n_896), .Y(n_915) );
NAND2xp5_ASAP7_75t_L g916 ( .A(n_889), .B(n_829), .Y(n_916) );
INVx2_ASAP7_75t_L g917 ( .A(n_851), .Y(n_917) );
INVx2_ASAP7_75t_L g918 ( .A(n_862), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_891), .B(n_866), .Y(n_919) );
AND2x2_ASAP7_75t_L g920 ( .A(n_847), .B(n_201), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g921 ( .A1(n_882), .A2(n_784), .B1(n_781), .B2(n_812), .Y(n_921) );
NAND2xp5_ASAP7_75t_L g922 ( .A(n_871), .B(n_829), .Y(n_922) );
A2O1A1Ixp33_ASAP7_75t_L g923 ( .A1(n_892), .A2(n_824), .B(n_835), .C(n_814), .Y(n_923) );
AND2x2_ASAP7_75t_L g924 ( .A(n_854), .B(n_842), .Y(n_924) );
OR2x2_ASAP7_75t_L g925 ( .A(n_871), .B(n_832), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_901), .B(n_832), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g927 ( .A(n_857), .B(n_833), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_865), .Y(n_928) );
NAND2xp5_ASAP7_75t_L g929 ( .A(n_857), .B(n_833), .Y(n_929) );
AND2x2_ASAP7_75t_L g930 ( .A(n_859), .B(n_815), .Y(n_930) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_864), .B(n_815), .Y(n_931) );
NAND2xp5_ASAP7_75t_L g932 ( .A(n_864), .B(n_815), .Y(n_932) );
HB1xp67_ASAP7_75t_L g933 ( .A(n_878), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_875), .B(n_820), .Y(n_934) );
BUFx2_ASAP7_75t_L g935 ( .A(n_858), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_875), .B(n_779), .Y(n_936) );
NOR2xp67_ASAP7_75t_SL g937 ( .A(n_848), .B(n_220), .Y(n_937) );
INVx1_ASAP7_75t_L g938 ( .A(n_885), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_885), .Y(n_939) );
AND2x2_ASAP7_75t_L g940 ( .A(n_869), .B(n_223), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_872), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g942 ( .A(n_895), .B(n_226), .Y(n_942) );
AND2x2_ASAP7_75t_L g943 ( .A(n_898), .B(n_227), .Y(n_943) );
NAND2xp5_ASAP7_75t_L g944 ( .A(n_903), .B(n_231), .Y(n_944) );
NOR2x1_ASAP7_75t_L g945 ( .A(n_874), .B(n_232), .Y(n_945) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_883), .B(n_234), .Y(n_946) );
AOI221xp5_ASAP7_75t_L g947 ( .A1(n_863), .A2(n_237), .B1(n_238), .B2(n_239), .C(n_240), .Y(n_947) );
INVx1_ASAP7_75t_L g948 ( .A(n_873), .Y(n_948) );
NAND2xp5_ASAP7_75t_L g949 ( .A(n_890), .B(n_243), .Y(n_949) );
NOR3xp33_ASAP7_75t_L g950 ( .A(n_881), .B(n_244), .C(n_245), .Y(n_950) );
AND2x2_ASAP7_75t_L g951 ( .A(n_899), .B(n_247), .Y(n_951) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_890), .B(n_249), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_867), .Y(n_953) );
AND2x4_ASAP7_75t_L g954 ( .A(n_935), .B(n_887), .Y(n_954) );
HB1xp67_ASAP7_75t_L g955 ( .A(n_933), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g956 ( .A(n_938), .B(n_886), .Y(n_956) );
INVx1_ASAP7_75t_L g957 ( .A(n_906), .Y(n_957) );
NAND2xp5_ASAP7_75t_L g958 ( .A(n_939), .B(n_902), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_919), .B(n_888), .Y(n_959) );
NAND2xp5_ASAP7_75t_L g960 ( .A(n_919), .B(n_893), .Y(n_960) );
AOI22xp5_ASAP7_75t_L g961 ( .A1(n_927), .A2(n_880), .B1(n_884), .B2(n_894), .Y(n_961) );
OR2x2_ASAP7_75t_L g962 ( .A(n_907), .B(n_900), .Y(n_962) );
INVxp67_ASAP7_75t_SL g963 ( .A(n_941), .Y(n_963) );
OAI21xp5_ASAP7_75t_L g964 ( .A1(n_945), .A2(n_879), .B(n_845), .Y(n_964) );
INVxp67_ASAP7_75t_L g965 ( .A(n_928), .Y(n_965) );
AOI221xp5_ASAP7_75t_L g966 ( .A1(n_911), .A2(n_870), .B1(n_846), .B2(n_897), .C(n_844), .Y(n_966) );
INVx1_ASAP7_75t_SL g967 ( .A(n_905), .Y(n_967) );
OAI22xp5_ASAP7_75t_L g968 ( .A1(n_921), .A2(n_844), .B1(n_850), .B2(n_856), .Y(n_968) );
OA211x2_ASAP7_75t_L g969 ( .A1(n_947), .A2(n_868), .B(n_850), .C(n_254), .Y(n_969) );
AND2x4_ASAP7_75t_L g970 ( .A(n_948), .B(n_868), .Y(n_970) );
HB1xp67_ASAP7_75t_L g971 ( .A(n_914), .Y(n_971) );
OAI21xp33_ASAP7_75t_L g972 ( .A1(n_936), .A2(n_261), .B(n_262), .Y(n_972) );
AOI21xp33_ASAP7_75t_L g973 ( .A1(n_929), .A2(n_264), .B(n_265), .Y(n_973) );
AOI221xp5_ASAP7_75t_L g974 ( .A1(n_912), .A2(n_267), .B1(n_268), .B2(n_269), .C(n_271), .Y(n_974) );
INVx2_ASAP7_75t_L g975 ( .A(n_917), .Y(n_975) );
INVx2_ASAP7_75t_SL g976 ( .A(n_915), .Y(n_976) );
AND2x2_ASAP7_75t_L g977 ( .A(n_918), .B(n_274), .Y(n_977) );
AOI21xp33_ASAP7_75t_L g978 ( .A1(n_916), .A2(n_275), .B(n_278), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g979 ( .A1(n_924), .A2(n_279), .B1(n_280), .B2(n_282), .Y(n_979) );
INVxp67_ASAP7_75t_L g980 ( .A(n_920), .Y(n_980) );
INVx2_ASAP7_75t_L g981 ( .A(n_970), .Y(n_981) );
INVx1_ASAP7_75t_L g982 ( .A(n_957), .Y(n_982) );
INVx2_ASAP7_75t_L g983 ( .A(n_970), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g984 ( .A(n_971), .B(n_922), .Y(n_984) );
OR2x2_ASAP7_75t_L g985 ( .A(n_955), .B(n_926), .Y(n_985) );
INVx2_ASAP7_75t_L g986 ( .A(n_975), .Y(n_986) );
INVx2_ASAP7_75t_L g987 ( .A(n_958), .Y(n_987) );
INVx1_ASAP7_75t_L g988 ( .A(n_965), .Y(n_988) );
NAND2x1p5_ASAP7_75t_L g989 ( .A(n_967), .B(n_908), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g990 ( .A1(n_968), .A2(n_904), .B1(n_910), .B2(n_923), .C(n_909), .Y(n_990) );
NAND2xp5_ASAP7_75t_L g991 ( .A(n_956), .B(n_913), .Y(n_991) );
BUFx2_ASAP7_75t_L g992 ( .A(n_963), .Y(n_992) );
INVxp67_ASAP7_75t_SL g993 ( .A(n_962), .Y(n_993) );
INVx1_ASAP7_75t_L g994 ( .A(n_958), .Y(n_994) );
INVx2_ASAP7_75t_SL g995 ( .A(n_976), .Y(n_995) );
NOR3xp33_ASAP7_75t_L g996 ( .A(n_964), .B(n_950), .C(n_951), .Y(n_996) );
XNOR2x1_ASAP7_75t_L g997 ( .A(n_961), .B(n_943), .Y(n_997) );
INVx1_ASAP7_75t_L g998 ( .A(n_992), .Y(n_998) );
AO22x2_ASAP7_75t_L g999 ( .A1(n_988), .A2(n_980), .B1(n_960), .B2(n_959), .Y(n_999) );
INVx1_ASAP7_75t_L g1000 ( .A(n_994), .Y(n_1000) );
HB1xp67_ASAP7_75t_L g1001 ( .A(n_993), .Y(n_1001) );
OAI22xp5_ASAP7_75t_L g1002 ( .A1(n_997), .A2(n_969), .B1(n_966), .B2(n_954), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_991), .B(n_959), .Y(n_1003) );
INVx2_ASAP7_75t_L g1004 ( .A(n_989), .Y(n_1004) );
OAI211xp5_ASAP7_75t_L g1005 ( .A1(n_990), .A2(n_972), .B(n_973), .C(n_978), .Y(n_1005) );
NAND3xp33_ASAP7_75t_L g1006 ( .A(n_996), .B(n_974), .C(n_953), .Y(n_1006) );
XOR2x2_ASAP7_75t_L g1007 ( .A(n_997), .B(n_979), .Y(n_1007) );
INVx1_ASAP7_75t_L g1008 ( .A(n_982), .Y(n_1008) );
NOR2xp33_ASAP7_75t_SL g1009 ( .A(n_995), .B(n_937), .Y(n_1009) );
OR2x2_ASAP7_75t_L g1010 ( .A(n_1001), .B(n_984), .Y(n_1010) );
INVx2_ASAP7_75t_L g1011 ( .A(n_998), .Y(n_1011) );
INVxp33_ASAP7_75t_SL g1012 ( .A(n_1002), .Y(n_1012) );
XNOR2x1_ASAP7_75t_L g1013 ( .A(n_1007), .B(n_985), .Y(n_1013) );
INVx1_ASAP7_75t_L g1014 ( .A(n_1000), .Y(n_1014) );
AO22x2_ASAP7_75t_L g1015 ( .A1(n_1004), .A2(n_981), .B1(n_983), .B2(n_987), .Y(n_1015) );
NOR2x1p5_ASAP7_75t_L g1016 ( .A(n_1006), .B(n_986), .Y(n_1016) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_999), .B(n_986), .Y(n_1017) );
NOR3xp33_ASAP7_75t_L g1018 ( .A(n_1005), .B(n_944), .C(n_946), .Y(n_1018) );
AND2x2_ASAP7_75t_L g1019 ( .A(n_999), .B(n_930), .Y(n_1019) );
OAI211xp5_ASAP7_75t_SL g1020 ( .A1(n_1003), .A2(n_932), .B(n_931), .C(n_925), .Y(n_1020) );
OAI321xp33_ASAP7_75t_L g1021 ( .A1(n_1008), .A2(n_952), .A3(n_949), .B1(n_942), .B2(n_934), .C(n_977), .Y(n_1021) );
AOI21xp5_ASAP7_75t_L g1022 ( .A1(n_1009), .A2(n_952), .B(n_934), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_999), .B(n_940), .Y(n_1023) );
CKINVDCx5p33_ASAP7_75t_R g1024 ( .A(n_1012), .Y(n_1024) );
INVx2_ASAP7_75t_L g1025 ( .A(n_1015), .Y(n_1025) );
NOR4xp75_ASAP7_75t_L g1026 ( .A(n_1023), .B(n_1017), .C(n_1013), .D(n_1019), .Y(n_1026) );
CKINVDCx5p33_ASAP7_75t_R g1027 ( .A(n_1016), .Y(n_1027) );
INVx1_ASAP7_75t_L g1028 ( .A(n_1010), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1029 ( .A(n_1014), .Y(n_1029) );
AO22x2_ASAP7_75t_L g1030 ( .A1(n_1025), .A2(n_1011), .B1(n_1018), .B2(n_1022), .Y(n_1030) );
NOR3xp33_ASAP7_75t_L g1031 ( .A(n_1024), .B(n_1021), .C(n_1020), .Y(n_1031) );
AOI22xp33_ASAP7_75t_SL g1032 ( .A1(n_1030), .A2(n_1027), .B1(n_1026), .B2(n_1028), .Y(n_1032) );
AND2x4_ASAP7_75t_L g1033 ( .A(n_1031), .B(n_1029), .Y(n_1033) );
INVx4_ASAP7_75t_L g1034 ( .A(n_1033), .Y(n_1034) );
INVxp33_ASAP7_75t_L g1035 ( .A(n_1032), .Y(n_1035) );
OAI21xp5_ASAP7_75t_L g1036 ( .A1(n_1035), .A2(n_296), .B(n_297), .Y(n_1036) );
AOI221x1_ASAP7_75t_L g1037 ( .A1(n_1036), .A2(n_1034), .B1(n_298), .B2(n_299), .C(n_300), .Y(n_1037) );
endmodule