module real_jpeg_3772_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVx1_ASAP7_75t_L g43 ( 
.A(n_0),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_0),
.A2(n_43),
.B1(n_125),
.B2(n_242),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_0),
.B(n_253),
.C(n_254),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_0),
.B(n_73),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_0),
.B(n_284),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_0),
.B(n_99),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_0),
.B(n_321),
.Y(n_320)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_1),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_2),
.A2(n_91),
.B1(n_94),
.B2(n_95),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_2),
.Y(n_94)
);

OAI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_2),
.A2(n_94),
.B1(n_163),
.B2(n_258),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_SL g314 ( 
.A1(n_2),
.A2(n_94),
.B1(n_127),
.B2(n_204),
.Y(n_314)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_3),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g109 ( 
.A(n_3),
.Y(n_109)
);

INVx2_ASAP7_75t_L g176 ( 
.A(n_3),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_4),
.A2(n_161),
.B1(n_162),
.B2(n_166),
.Y(n_160)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_4),
.Y(n_166)
);

OAI22xp33_ASAP7_75t_SL g202 ( 
.A1(n_4),
.A2(n_118),
.B1(n_166),
.B2(n_203),
.Y(n_202)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx8_ASAP7_75t_L g156 ( 
.A(n_6),
.Y(n_156)
);

INVx2_ASAP7_75t_L g261 ( 
.A(n_6),
.Y(n_261)
);

BUFx6f_ASAP7_75t_L g284 ( 
.A(n_6),
.Y(n_284)
);

BUFx5_ASAP7_75t_L g327 ( 
.A(n_6),
.Y(n_327)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g51 ( 
.A1(n_8),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_8),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_8),
.A2(n_52),
.B1(n_124),
.B2(n_127),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_8),
.A2(n_52),
.B1(n_84),
.B2(n_185),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g262 ( 
.A1(n_8),
.A2(n_52),
.B1(n_263),
.B2(n_265),
.Y(n_262)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_10),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_10),
.Y(n_53)
);

BUFx5_ASAP7_75t_L g144 ( 
.A(n_10),
.Y(n_144)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_10),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_11),
.A2(n_115),
.B1(n_118),
.B2(n_121),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_11),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g188 ( 
.A1(n_11),
.A2(n_121),
.B1(n_189),
.B2(n_192),
.Y(n_188)
);

AOI22xp33_ASAP7_75t_L g171 ( 
.A1(n_12),
.A2(n_172),
.B1(n_177),
.B2(n_178),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_12),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_13),
.A2(n_83),
.B1(n_87),
.B2(n_88),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_13),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_13),
.A2(n_88),
.B1(n_143),
.B2(n_225),
.Y(n_224)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_13),
.A2(n_88),
.B1(n_203),
.B2(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_13),
.A2(n_88),
.B1(n_263),
.B2(n_289),
.Y(n_288)
);

BUFx3_ASAP7_75t_L g103 ( 
.A(n_14),
.Y(n_103)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_14),
.Y(n_113)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_14),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_14),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_SL g209 ( 
.A1(n_15),
.A2(n_210),
.B1(n_213),
.B2(n_214),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_15),
.Y(n_213)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_233),
.B1(n_234),
.B2(n_355),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g355 ( 
.A(n_18),
.Y(n_355)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_19),
.B(n_232),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_196),
.Y(n_19)
);

OR2x2_ASAP7_75t_L g232 ( 
.A(n_20),
.B(n_196),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_138),
.C(n_180),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_21),
.B(n_352),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_23),
.B1(n_58),
.B2(n_137),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_22),
.B(n_59),
.C(n_97),
.Y(n_216)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

AOI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_41),
.B(n_49),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_24),
.B(n_51),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_30),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_25)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_26),
.Y(n_29)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_26),
.Y(n_146)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_34),
.B1(n_37),
.B2(n_39),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_33),
.Y(n_40)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_33),
.Y(n_148)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_36),
.Y(n_323)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_38),
.Y(n_96)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

OAI21xp33_ASAP7_75t_SL g41 ( 
.A1(n_42),
.A2(n_43),
.B(n_44),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_43),
.B(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_43),
.B(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g285 ( 
.A1(n_43),
.A2(n_153),
.B(n_260),
.Y(n_285)
);

OAI21xp33_ASAP7_75t_SL g317 ( 
.A1(n_43),
.A2(n_318),
.B(n_319),
.Y(n_317)
);

OAI32xp33_ASAP7_75t_L g141 ( 
.A1(n_44),
.A2(n_142),
.A3(n_143),
.B1(n_145),
.B2(n_147),
.Y(n_141)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_48),
.Y(n_56)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_57),
.Y(n_50)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_57),
.Y(n_195)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

XNOR2xp5_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_97),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_82),
.B1(n_89),
.B2(n_90),
.Y(n_59)
);

INVx2_ASAP7_75t_SL g186 ( 
.A(n_60),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_73),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_62),
.A2(n_64),
.B1(n_68),
.B2(n_71),
.Y(n_61)
);

INVx6_ASAP7_75t_L g336 ( 
.A(n_62),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_64),
.Y(n_185)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx3_ASAP7_75t_L g142 ( 
.A(n_67),
.Y(n_142)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_67),
.Y(n_318)
);

AO22x2_ASAP7_75t_L g73 ( 
.A1(n_68),
.A2(n_74),
.B1(n_78),
.B2(n_80),
.Y(n_73)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g333 ( 
.A(n_70),
.Y(n_333)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_73),
.Y(n_89)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_77),
.Y(n_79)
);

INVx11_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx3_ASAP7_75t_L g120 ( 
.A(n_77),
.Y(n_120)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_77),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_77),
.Y(n_127)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_77),
.Y(n_136)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_82),
.A2(n_89),
.B(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_89),
.B(n_184),
.Y(n_231)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_90),
.Y(n_230)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g150 ( 
.A(n_93),
.Y(n_150)
);

AOI32xp33_ASAP7_75t_L g328 ( 
.A1(n_95),
.A2(n_320),
.A3(n_329),
.B1(n_332),
.B2(n_334),
.Y(n_328)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_96),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_114),
.B(n_122),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_98),
.A2(n_114),
.B1(n_200),
.B2(n_201),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g313 ( 
.A1(n_98),
.A2(n_200),
.B1(n_269),
.B2(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_99),
.B(n_123),
.Y(n_245)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g128 ( 
.A(n_100),
.B(n_129),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g268 ( 
.A1(n_100),
.A2(n_122),
.B(n_269),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_104),
.B1(n_108),
.B2(n_110),
.Y(n_100)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g134 ( 
.A(n_103),
.Y(n_134)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g158 ( 
.A(n_107),
.Y(n_158)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_107),
.Y(n_161)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_107),
.Y(n_193)
);

BUFx8_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_109),
.Y(n_165)
);

BUFx3_ASAP7_75t_L g291 ( 
.A(n_109),
.Y(n_291)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_117),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_117),
.Y(n_244)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_117),
.Y(n_251)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_117),
.Y(n_272)
);

INVx4_ASAP7_75t_SL g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g129 ( 
.A1(n_119),
.A2(n_130),
.B1(n_133),
.B2(n_135),
.Y(n_129)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.Y(n_122)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_SL g200 ( 
.A(n_128),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_132),
.Y(n_131)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

BUFx3_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_136),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_138),
.A2(n_139),
.B1(n_180),
.B2(n_353),
.Y(n_352)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_140),
.A2(n_141),
.B1(n_151),
.B2(n_152),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_141),
.B(n_151),
.Y(n_220)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_SL g145 ( 
.A(n_146),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_149),
.Y(n_147)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_159),
.B1(n_167),
.B2(n_170),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_153),
.A2(n_257),
.B(n_260),
.Y(n_256)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_154),
.A2(n_160),
.B1(n_168),
.B2(n_188),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_154),
.A2(n_168),
.B1(n_171),
.B2(n_208),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g294 ( 
.A(n_154),
.B(n_262),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_154),
.A2(n_299),
.B1(n_300),
.B2(n_301),
.Y(n_298)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_157),
.Y(n_154)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_155),
.Y(n_293)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_156),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_156),
.Y(n_303)
);

INVx3_ASAP7_75t_L g265 ( 
.A(n_157),
.Y(n_265)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_174),
.Y(n_215)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

BUFx6f_ASAP7_75t_L g179 ( 
.A(n_176),
.Y(n_179)
);

BUFx3_ASAP7_75t_L g191 ( 
.A(n_176),
.Y(n_191)
);

INVx4_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

INVx8_ASAP7_75t_L g264 ( 
.A(n_179),
.Y(n_264)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_180),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.C(n_194),
.Y(n_180)
);

XNOR2xp5_ASAP7_75t_SL g345 ( 
.A(n_181),
.B(n_346),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_186),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_186),
.A2(n_230),
.B(n_231),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_186),
.A2(n_231),
.B(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_187),
.B(n_194),
.Y(n_346)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_188),
.Y(n_326)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_191),
.Y(n_282)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_224),
.B(n_227),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_219),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_198),
.A2(n_216),
.B1(n_217),
.B2(n_218),
.Y(n_197)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_207),
.Y(n_198)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_200),
.A2(n_241),
.B(n_245),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_SL g343 ( 
.A1(n_200),
.A2(n_245),
.B(n_314),
.Y(n_343)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx3_ASAP7_75t_L g204 ( 
.A(n_205),
.Y(n_204)
);

INVx5_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_SL g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_214),
.Y(n_254)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_216),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_223),
.B1(n_228),
.B2(n_229),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

AOI21x1_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_349),
.B(n_354),
.Y(n_234)
);

AO21x1_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_338),
.B(n_348),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g236 ( 
.A1(n_237),
.A2(n_308),
.B(n_337),
.Y(n_236)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_275),
.B(n_307),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_255),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_255),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_240),
.A2(n_246),
.B1(n_247),
.B2(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_240),
.Y(n_305)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx4_ASAP7_75t_L g243 ( 
.A(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_252),
.Y(n_247)
);

INVx2_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx2_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx6_ASAP7_75t_L g335 ( 
.A(n_251),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_266),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_256),
.B(n_267),
.C(n_274),
.Y(n_309)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_257),
.Y(n_300)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

AOI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_267),
.A2(n_268),
.B1(n_273),
.B2(n_274),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx11_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

OAI21xp5_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_297),
.B(n_306),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_277),
.A2(n_286),
.B(n_296),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_285),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_283),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

INVx6_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_295),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_287),
.B(n_295),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_288),
.A2(n_292),
.B(n_294),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_288),
.Y(n_299)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx5_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_294),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_304),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_304),
.Y(n_306)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx8_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_310),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_309),
.B(n_310),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_324),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_312),
.A2(n_313),
.B1(n_315),
.B2(n_316),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_313),
.B(n_315),
.C(n_324),
.Y(n_339)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVxp33_ASAP7_75t_L g319 ( 
.A(n_320),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_322),
.Y(n_321)
);

INVx6_ASAP7_75t_SL g322 ( 
.A(n_323),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g324 ( 
.A(n_325),
.B(n_328),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_325),
.B(n_328),
.Y(n_344)
);

INVx5_ASAP7_75t_SL g329 ( 
.A(n_330),
.Y(n_329)
);

INVx4_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVx5_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

NAND2xp33_ASAP7_75t_SL g334 ( 
.A(n_335),
.B(n_336),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_339),
.B(n_340),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_SL g348 ( 
.A(n_339),
.B(n_340),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_341),
.A2(n_342),
.B1(n_345),
.B2(n_347),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_342),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_343),
.B(n_344),
.C(n_347),
.Y(n_350)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_345),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g354 ( 
.A(n_350),
.B(n_351),
.Y(n_354)
);


endmodule