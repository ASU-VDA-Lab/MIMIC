module fake_netlist_1_1133_n_29 (n_1, n_2, n_6, n_4, n_3, n_5, n_7, n_8, n_0, n_29);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_5;
input n_7;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx1_ASAP7_75t_L g9 ( .A(n_2), .Y(n_9) );
HB1xp67_ASAP7_75t_L g10 ( .A(n_0), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
NAND2xp5_ASAP7_75t_L g12 ( .A(n_6), .B(n_0), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_3), .Y(n_13) );
INVx2_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx8_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
INVx4_ASAP7_75t_L g16 ( .A(n_13), .Y(n_16) );
OR2x2_ASAP7_75t_SL g17 ( .A(n_10), .B(n_1), .Y(n_17) );
NAND2xp5_ASAP7_75t_SL g18 ( .A(n_11), .B(n_2), .Y(n_18) );
BUFx3_ASAP7_75t_L g19 ( .A(n_14), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_19), .Y(n_20) );
AND2x4_ASAP7_75t_L g21 ( .A(n_16), .B(n_14), .Y(n_21) );
HB1xp67_ASAP7_75t_L g22 ( .A(n_15), .Y(n_22) );
BUFx6f_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
AND2x2_ASAP7_75t_L g24 ( .A(n_23), .B(n_22), .Y(n_24) );
NOR4xp25_ASAP7_75t_SL g25 ( .A(n_24), .B(n_18), .C(n_17), .D(n_20), .Y(n_25) );
INVx1_ASAP7_75t_SL g26 ( .A(n_25), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_26), .Y(n_27) );
INVxp67_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
AOI322xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_9), .A3(n_12), .B1(n_17), .B2(n_4), .C1(n_5), .C2(n_7), .Y(n_29) );
endmodule