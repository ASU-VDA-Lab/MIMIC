module fake_jpeg_14889_n_268 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_268);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_268;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_252;
wire n_251;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_264;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx3_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g19 ( 
.A(n_3),
.B(n_8),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx16f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

INVx11_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_32),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_19),
.B(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_36),
.Y(n_47)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

INVx5_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_31),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_37),
.Y(n_53)
);

OR2x2_ASAP7_75t_L g38 ( 
.A(n_16),
.B(n_0),
.Y(n_38)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_38),
.B(n_40),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_22),
.Y(n_40)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_41),
.A2(n_18),
.B1(n_23),
.B2(n_26),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_42),
.A2(n_44),
.B1(n_45),
.B2(n_46),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_23),
.B1(n_18),
.B2(n_22),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_21),
.B1(n_16),
.B2(n_30),
.Y(n_45)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_32),
.A2(n_21),
.B1(n_40),
.B2(n_30),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_37),
.A2(n_39),
.B1(n_40),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_57),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_37),
.A2(n_24),
.B1(n_15),
.B2(n_25),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_32),
.A2(n_30),
.B1(n_19),
.B2(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_29),
.Y(n_54)
);

OAI21xp33_ASAP7_75t_L g78 ( 
.A1(n_54),
.A2(n_59),
.B(n_60),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_24),
.B1(n_15),
.B2(n_27),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_38),
.B(n_29),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_20),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_61),
.B(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_34),
.B(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_35),
.Y(n_64)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_63),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_65),
.B(n_75),
.Y(n_108)
);

OR2x2_ASAP7_75t_SL g66 ( 
.A(n_52),
.B(n_32),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g97 ( 
.A(n_66),
.B(n_47),
.C(n_35),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_50),
.A2(n_39),
.B1(n_25),
.B2(n_20),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_67),
.A2(n_57),
.B1(n_59),
.B2(n_39),
.Y(n_92)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_62),
.Y(n_72)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_58),
.Y(n_74)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_74),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_61),
.Y(n_75)
);

CKINVDCx9p33_ASAP7_75t_R g76 ( 
.A(n_46),
.Y(n_76)
);

INVx11_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

BUFx8_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_77),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_53),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_SL g107 ( 
.A(n_79),
.B(n_83),
.Y(n_107)
);

INVx2_ASAP7_75t_SL g80 ( 
.A(n_64),
.Y(n_80)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_43),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g102 ( 
.A(n_82),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_53),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_55),
.Y(n_84)
);

OR2x2_ASAP7_75t_L g89 ( 
.A(n_84),
.B(n_85),
.Y(n_89)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_55),
.Y(n_85)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_65),
.B(n_54),
.C(n_60),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_87),
.B(n_36),
.C(n_77),
.Y(n_129)
);

AND2x6_ASAP7_75t_L g88 ( 
.A(n_78),
.B(n_52),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_88),
.A2(n_106),
.B(n_34),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_43),
.B1(n_62),
.B2(n_70),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_90),
.A2(n_99),
.B1(n_100),
.B2(n_77),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_92),
.A2(n_86),
.B1(n_79),
.B2(n_83),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_52),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_98),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_66),
.A2(n_47),
.B(n_48),
.C(n_42),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_95),
.B(n_109),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_28),
.B(n_17),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_68),
.B(n_34),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g99 ( 
.A1(n_81),
.A2(n_35),
.B1(n_62),
.B2(n_56),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_56),
.B1(n_35),
.B2(n_2),
.Y(n_100)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_73),
.A2(n_34),
.B(n_36),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_20),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_85),
.Y(n_110)
);

CKINVDCx14_ASAP7_75t_R g142 ( 
.A(n_110),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_111),
.A2(n_113),
.B1(n_114),
.B2(n_118),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_106),
.A2(n_74),
.B1(n_71),
.B2(n_69),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_108),
.A2(n_71),
.B1(n_69),
.B2(n_80),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_34),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_115),
.A2(n_124),
.B(n_126),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_80),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_116),
.B(n_117),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_82),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_95),
.A2(n_56),
.B1(n_1),
.B2(n_2),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_87),
.B(n_72),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_119),
.B(n_120),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_72),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_72),
.Y(n_121)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_121),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_92),
.Y(n_143)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_107),
.Y(n_123)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_123),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_0),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_125),
.B(n_132),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_109),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_128),
.B(n_101),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g128 ( 
.A1(n_88),
.A2(n_77),
.B(n_49),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_101),
.C(n_103),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_88),
.B(n_49),
.Y(n_130)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_130),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_96),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_134),
.B(n_136),
.C(n_129),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_119),
.B(n_96),
.C(n_103),
.Y(n_136)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_121),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_141),
.B(n_151),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_143),
.B(n_129),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_123),
.B(n_105),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_148),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_145),
.A2(n_128),
.B1(n_118),
.B2(n_127),
.Y(n_169)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_114),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_113),
.B(n_93),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_149),
.A2(n_152),
.B(n_142),
.Y(n_164)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_120),
.Y(n_150)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_150),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_117),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_126),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_153),
.B(n_155),
.Y(n_168)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_110),
.Y(n_154)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_154),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g155 ( 
.A(n_112),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_156),
.B(n_136),
.C(n_139),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_SL g160 ( 
.A(n_134),
.B(n_130),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_SL g185 ( 
.A(n_160),
.B(n_169),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_137),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_163),
.B(n_165),
.Y(n_183)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_164),
.A2(n_172),
.B(n_174),
.Y(n_195)
);

INVxp33_ASAP7_75t_L g165 ( 
.A(n_138),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_147),
.Y(n_166)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_166),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_155),
.B(n_112),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_167),
.B(n_170),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_137),
.Y(n_170)
);

NAND3xp33_ASAP7_75t_L g171 ( 
.A(n_153),
.B(n_132),
.C(n_128),
.Y(n_171)
);

NOR2xp67_ASAP7_75t_R g182 ( 
.A(n_171),
.B(n_145),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_122),
.B(n_131),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_152),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_173),
.A2(n_175),
.B1(n_176),
.B2(n_140),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_133),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_150),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_154),
.B(n_115),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_177),
.B(n_115),
.Y(n_189)
);

XOR2xp5_ASAP7_75t_L g188 ( 
.A(n_178),
.B(n_140),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_186),
.C(n_187),
.Y(n_200)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_162),
.A2(n_149),
.B1(n_146),
.B2(n_148),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_180),
.B(n_181),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_162),
.A2(n_146),
.B1(n_124),
.B2(n_125),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g206 ( 
.A(n_182),
.B(n_164),
.Y(n_206)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_184),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_156),
.B(n_143),
.C(n_135),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_178),
.B(n_135),
.C(n_131),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_188),
.B(n_185),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_189),
.B(n_198),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_159),
.A2(n_104),
.B1(n_111),
.B2(n_124),
.Y(n_190)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_190),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_160),
.B(n_49),
.C(n_36),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_191),
.B(n_194),
.C(n_176),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_124),
.B1(n_104),
.B2(n_105),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_175),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_158),
.B(n_102),
.C(n_93),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_173),
.A2(n_104),
.B1(n_93),
.B2(n_91),
.Y(n_197)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_197),
.B(n_177),
.Y(n_201)
);

INVx3_ASAP7_75t_SL g198 ( 
.A(n_161),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_201),
.A2(n_157),
.B1(n_91),
.B2(n_0),
.Y(n_227)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_203),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_205),
.C(n_207),
.Y(n_216)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_185),
.B(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_206),
.B(n_187),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_188),
.B(n_169),
.Y(n_207)
);

BUFx24_ASAP7_75t_SL g209 ( 
.A(n_195),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_209),
.B(n_212),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_168),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_210),
.B(n_214),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_198),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_183),
.B(n_102),
.Y(n_213)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_213),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_167),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_194),
.C(n_186),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_200),
.C(n_207),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_218),
.B(n_225),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_192),
.B1(n_196),
.B2(n_158),
.Y(n_220)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_220),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_166),
.Y(n_221)
);

AND2x2_ASAP7_75t_L g230 ( 
.A(n_221),
.B(n_227),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_208),
.A2(n_157),
.B1(n_197),
.B2(n_189),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_226),
.B(n_228),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_202),
.B(n_3),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_229),
.B(n_5),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_232),
.B(n_240),
.C(n_17),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_L g233 ( 
.A1(n_217),
.A2(n_205),
.B(n_204),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_233),
.B(n_235),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_216),
.B(n_4),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_234),
.B(n_7),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_227),
.B(n_5),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_236),
.B(n_239),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_219),
.B(n_6),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_224),
.B(n_28),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_231),
.B(n_223),
.Y(n_242)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_242),
.Y(n_251)
);

OAI21x1_ASAP7_75t_L g244 ( 
.A1(n_237),
.A2(n_224),
.B(n_222),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_244),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_238),
.B(n_229),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_245),
.B(n_246),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_230),
.A2(n_221),
.B(n_216),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_247),
.B(n_249),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_240),
.B(n_8),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_248),
.B(n_234),
.Y(n_252)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_241),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_252),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_243),
.B(n_232),
.Y(n_254)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_254),
.B(n_241),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_259),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g259 ( 
.A1(n_250),
.A2(n_230),
.B(n_9),
.Y(n_259)
);

AOI322xp5_ASAP7_75t_L g260 ( 
.A1(n_251),
.A2(n_256),
.A3(n_255),
.B1(n_253),
.B2(n_11),
.C1(n_12),
.C2(n_8),
.Y(n_260)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_260),
.A2(n_11),
.B(n_12),
.Y(n_263)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_250),
.A2(n_9),
.B(n_10),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_261),
.B(n_9),
.C(n_10),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_262),
.B(n_263),
.C(n_258),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_265),
.B(n_266),
.Y(n_267)
);

MAJx2_ASAP7_75t_L g266 ( 
.A(n_264),
.B(n_13),
.C(n_14),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_267),
.B(n_13),
.Y(n_268)
);


endmodule