module fake_jpeg_1462_n_229 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_229);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_229;

wire n_159;
wire n_117;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_10),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_35),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_52),
.Y(n_59)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_21),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_20),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_34),
.Y(n_64)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_11),
.Y(n_65)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_37),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_21),
.Y(n_69)
);

INVx2_ASAP7_75t_SL g70 ( 
.A(n_10),
.Y(n_70)
);

BUFx10_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_3),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_0),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_8),
.Y(n_75)
);

INVx11_ASAP7_75t_SL g76 ( 
.A(n_49),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_70),
.B(n_51),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_78),
.B(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_79),
.Y(n_87)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_66),
.Y(n_80)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_80),
.Y(n_88)
);

INVx11_ASAP7_75t_L g81 ( 
.A(n_66),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_81),
.A2(n_56),
.B1(n_66),
.B2(n_55),
.Y(n_89)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_84),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_76),
.Y(n_84)
);

BUFx12_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_85),
.A2(n_56),
.B1(n_55),
.B2(n_59),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g86 ( 
.A1(n_83),
.A2(n_72),
.B1(n_54),
.B2(n_75),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_86),
.A2(n_90),
.B1(n_92),
.B2(n_96),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g101 ( 
.A(n_89),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_79),
.A2(n_75),
.B1(n_54),
.B2(n_72),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_83),
.A2(n_79),
.B1(n_81),
.B2(n_80),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.C(n_53),
.Y(n_94)
);

FAx1_ASAP7_75t_SL g103 ( 
.A(n_94),
.B(n_56),
.CI(n_71),
.CON(n_103),
.SN(n_103)
);

BUFx3_ASAP7_75t_L g112 ( 
.A(n_95),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_82),
.A2(n_53),
.B1(n_68),
.B2(n_73),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_83),
.A2(n_69),
.B1(n_74),
.B2(n_62),
.Y(n_97)
);

OAI22xp33_ASAP7_75t_SL g105 ( 
.A1(n_97),
.A2(n_84),
.B1(n_57),
.B2(n_81),
.Y(n_105)
);

OAI22xp33_ASAP7_75t_SL g98 ( 
.A1(n_81),
.A2(n_82),
.B1(n_84),
.B2(n_68),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_L g116 ( 
.A1(n_98),
.A2(n_71),
.B1(n_65),
.B2(n_85),
.Y(n_116)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_88),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g128 ( 
.A(n_99),
.Y(n_128)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_88),
.Y(n_100)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_98),
.Y(n_102)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_103),
.B(n_96),
.C(n_71),
.Y(n_122)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_104),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_105),
.A2(n_117),
.B1(n_87),
.B2(n_92),
.Y(n_124)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_87),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_106),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_61),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_107),
.B(n_111),
.Y(n_125)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_109),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_94),
.B(n_63),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_110),
.B(n_65),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_94),
.B(n_64),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_91),
.B(n_67),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_115),
.Y(n_127)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_93),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_114),
.B(n_40),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_97),
.B(n_77),
.Y(n_115)
);

OR2x2_ASAP7_75t_L g131 ( 
.A(n_116),
.B(n_85),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_86),
.A2(n_82),
.B1(n_71),
.B2(n_65),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_L g118 ( 
.A1(n_101),
.A2(n_112),
.B(n_103),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_SL g157 ( 
.A1(n_118),
.A2(n_38),
.B(n_36),
.Y(n_157)
);

BUFx12_ASAP7_75t_L g121 ( 
.A(n_99),
.Y(n_121)
);

CKINVDCx14_ASAP7_75t_R g150 ( 
.A(n_121),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_122),
.B(n_133),
.C(n_60),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_106),
.B(n_87),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g147 ( 
.A(n_123),
.B(n_129),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_124),
.A2(n_138),
.B1(n_31),
.B2(n_29),
.Y(n_161)
);

NOR2x1_ASAP7_75t_L g126 ( 
.A(n_102),
.B(n_95),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_126),
.B(n_139),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_103),
.B(n_0),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_130),
.B(n_134),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_131),
.Y(n_142)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_100),
.B(n_85),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_104),
.B(n_1),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_137),
.B(n_39),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_108),
.A2(n_65),
.B1(n_60),
.B2(n_85),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_112),
.B(n_1),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_118),
.A2(n_101),
.B(n_85),
.Y(n_140)
);

INVxp67_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_136),
.Y(n_141)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_141),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_143),
.B(n_126),
.Y(n_164)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_132),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_144),
.B(n_146),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_135),
.A2(n_50),
.B1(n_48),
.B2(n_47),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_153),
.B1(n_124),
.B2(n_138),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_133),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_127),
.B(n_2),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_151),
.B(n_152),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_2),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_46),
.B1(n_44),
.B2(n_43),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_120),
.B(n_42),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_154),
.B(n_160),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_4),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_155),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g184 ( 
.A(n_156),
.B(n_159),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_157),
.A2(n_163),
.B(n_128),
.Y(n_165)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_132),
.Y(n_158)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_158),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_119),
.B(n_4),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_122),
.B(n_32),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_161),
.A2(n_8),
.B1(n_9),
.B2(n_11),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_133),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_162),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_121),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_170),
.C(n_158),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_165),
.B(n_174),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_166),
.B(n_168),
.Y(n_192)
);

OAI22x1_ASAP7_75t_L g167 ( 
.A1(n_148),
.A2(n_131),
.B1(n_121),
.B2(n_28),
.Y(n_167)
);

AOI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_167),
.A2(n_176),
.B1(n_154),
.B2(n_147),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g169 ( 
.A1(n_142),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_175),
.B1(n_179),
.B2(n_145),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_5),
.C(n_6),
.Y(n_170)
);

NOR2x1_ASAP7_75t_L g174 ( 
.A(n_142),
.B(n_7),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_140),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_141),
.Y(n_180)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_180),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g182 ( 
.A1(n_160),
.A2(n_15),
.B(n_16),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g186 ( 
.A(n_182),
.B(n_15),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_186),
.B(n_191),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_187),
.B(n_193),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_189),
.A2(n_192),
.B1(n_183),
.B2(n_181),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g190 ( 
.A1(n_172),
.A2(n_157),
.B(n_150),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_190),
.A2(n_170),
.B(n_171),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g191 ( 
.A(n_177),
.B(n_153),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g193 ( 
.A(n_173),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g203 ( 
.A(n_194),
.B(n_196),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_164),
.B(n_144),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_195),
.B(n_184),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_171),
.B(n_16),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_183),
.B(n_22),
.Y(n_197)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_197),
.Y(n_208)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_198),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_199),
.A2(n_195),
.B1(n_188),
.B2(n_194),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_190),
.A2(n_167),
.B1(n_174),
.B2(n_172),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_201),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g210 ( 
.A(n_204),
.B(n_205),
.Y(n_210)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_185),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_207),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g209 ( 
.A(n_200),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_209),
.B(n_212),
.Y(n_219)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_203),
.B(n_189),
.C(n_184),
.Y(n_213)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_213),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_193),
.C(n_18),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

NAND2x1_ASAP7_75t_L g217 ( 
.A(n_215),
.B(n_202),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_217),
.A2(n_214),
.B1(n_204),
.B2(n_209),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g222 ( 
.A(n_220),
.B(n_216),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_219),
.A2(n_210),
.B1(n_211),
.B2(n_208),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_221),
.A2(n_218),
.B1(n_210),
.B2(n_206),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g224 ( 
.A(n_222),
.B(n_223),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_224),
.B(n_217),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_225),
.A2(n_221),
.B(n_19),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_22),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_227),
.B(n_17),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_20),
.Y(n_229)
);


endmodule