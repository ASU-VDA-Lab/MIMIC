module fake_ariane_1316_n_768 (n_83, n_8, n_56, n_60, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_142, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_127, n_35, n_54, n_25, n_768);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_142;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_127;
input n_35;
input n_54;
input n_25;

output n_768;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_698;
wire n_695;
wire n_160;
wire n_180;
wire n_730;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_646;
wire n_197;
wire n_640;
wire n_463;
wire n_176;
wire n_691;
wire n_404;
wire n_172;
wire n_678;
wire n_651;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_726;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_610;
wire n_205;
wire n_752;
wire n_341;
wire n_245;
wire n_421;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_760;
wire n_690;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_713;
wire n_649;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_244;
wire n_679;
wire n_643;
wire n_226;
wire n_220;
wire n_261;
wire n_682;
wire n_663;
wire n_370;
wire n_706;
wire n_189;
wire n_717;
wire n_286;
wire n_443;
wire n_586;
wire n_686;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_524;
wire n_349;
wire n_391;
wire n_634;
wire n_466;
wire n_756;
wire n_346;
wire n_214;
wire n_764;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_670;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_162;
wire n_765;
wire n_264;
wire n_737;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_637;
wire n_327;
wire n_766;
wire n_372;
wire n_377;
wire n_396;
wire n_631;
wire n_399;
wire n_554;
wire n_520;
wire n_714;
wire n_279;
wire n_702;
wire n_207;
wire n_363;
wire n_720;
wire n_354;
wire n_725;
wire n_419;
wire n_230;
wire n_270;
wire n_194;
wire n_633;
wire n_154;
wire n_338;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_193;
wire n_733;
wire n_761;
wire n_500;
wire n_731;
wire n_336;
wire n_665;
wire n_754;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_668;
wire n_339;
wire n_738;
wire n_758;
wire n_672;
wire n_487;
wire n_740;
wire n_167;
wire n_422;
wire n_153;
wire n_648;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_446;
wire n_553;
wire n_753;
wire n_566;
wire n_578;
wire n_701;
wire n_625;
wire n_405;
wire n_557;
wire n_169;
wire n_173;
wire n_242;
wire n_645;
wire n_309;
wire n_331;
wire n_320;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_647;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_721;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_759;
wire n_247;
wire n_569;
wire n_567;
wire n_732;
wire n_240;
wire n_369;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_677;
wire n_222;
wire n_478;
wire n_703;
wire n_748;
wire n_510;
wire n_256;
wire n_326;
wire n_681;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_635;
wire n_707;
wire n_330;
wire n_400;
wire n_694;
wire n_689;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_699;
wire n_727;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_644;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_688;
wire n_636;
wire n_427;
wire n_587;
wire n_497;
wire n_693;
wire n_303;
wire n_671;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_654;
wire n_588;
wire n_638;
wire n_334;
wire n_192;
wire n_729;
wire n_661;
wire n_488;
wire n_667;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_390;
wire n_498;
wire n_501;
wire n_438;
wire n_314;
wire n_684;
wire n_440;
wire n_627;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_728;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_715;
wire n_579;
wire n_459;
wire n_685;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_711;
wire n_453;
wire n_734;
wire n_491;
wire n_181;
wire n_723;
wire n_617;
wire n_616;
wire n_705;
wire n_630;
wire n_658;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_709;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_281;
wire n_628;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_743;
wire n_225;
wire n_235;
wire n_660;
wire n_464;
wire n_735;
wire n_575;
wire n_546;
wire n_297;
wire n_662;
wire n_641;
wire n_503;
wire n_700;
wire n_290;
wire n_527;
wire n_741;
wire n_747;
wire n_371;
wire n_199;
wire n_639;
wire n_217;
wire n_452;
wire n_673;
wire n_676;
wire n_178;
wire n_551;
wire n_308;
wire n_708;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_680;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_284;
wire n_448;
wire n_593;
wire n_755;
wire n_710;
wire n_249;
wire n_534;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_652;
wire n_451;
wire n_613;
wire n_745;
wire n_475;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_716;
wire n_742;
wire n_182;
wire n_696;
wire n_674;
wire n_482;
wire n_316;
wire n_196;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_744;
wire n_762;
wire n_656;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_252;
wire n_215;
wire n_629;
wire n_664;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_763;
wire n_655;
wire n_540;
wire n_216;
wire n_544;
wire n_692;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_750;
wire n_389;
wire n_657;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_304;
wire n_659;
wire n_509;
wire n_583;
wire n_724;
wire n_306;
wire n_666;
wire n_313;
wire n_430;
wire n_626;
wire n_493;
wire n_722;
wire n_203;
wire n_378;
wire n_436;
wire n_757;
wire n_375;
wire n_324;
wire n_585;
wire n_669;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_622;
wire n_697;
wire n_472;
wire n_296;
wire n_265;
wire n_746;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_704;
wire n_204;
wire n_751;
wire n_615;
wire n_521;
wire n_496;
wire n_739;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_580;
wire n_608;
wire n_494;
wire n_719;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_317;
wire n_243;
wire n_329;
wire n_718;
wire n_185;
wire n_340;
wire n_749;
wire n_289;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_632;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_650;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_618;
wire n_411;
wire n_484;
wire n_712;
wire n_353;
wire n_736;
wire n_767;
wire n_241;
wire n_357;
wire n_412;
wire n_687;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_642;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_653;
wire n_359;
wire n_155;
wire n_573;
wire n_531;
wire n_675;

INVx2_ASAP7_75t_L g153 ( 
.A(n_141),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_28),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_60),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_5),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_78),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_49),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_45),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_20),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_115),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_31),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_25),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_135),
.Y(n_165)
);

BUFx2_ASAP7_75t_L g166 ( 
.A(n_17),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_26),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_34),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_11),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_5),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_144),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_139),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_130),
.Y(n_174)
);

CKINVDCx6p67_ASAP7_75t_R g175 ( 
.A(n_147),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_110),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_101),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_40),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_10),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_133),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_63),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_136),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_68),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_38),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_109),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_124),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_21),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_1),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_39),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_104),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_119),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_9),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_143),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_13),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_7),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_151),
.Y(n_198)
);

NOR2xp67_ASAP7_75t_L g199 ( 
.A(n_55),
.B(n_36),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_33),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_54),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_97),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g203 ( 
.A(n_82),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_67),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_150),
.Y(n_205)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_4),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_84),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_118),
.Y(n_209)
);

BUFx8_ASAP7_75t_SL g210 ( 
.A(n_206),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_166),
.B(n_0),
.Y(n_211)
);

OAI21x1_ASAP7_75t_L g212 ( 
.A1(n_153),
.A2(n_73),
.B(n_146),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_161),
.Y(n_213)
);

INVx4_ASAP7_75t_L g214 ( 
.A(n_186),
.Y(n_214)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

BUFx8_ASAP7_75t_L g216 ( 
.A(n_153),
.Y(n_216)
);

INVx3_ASAP7_75t_L g217 ( 
.A(n_156),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_193),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_155),
.B(n_0),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_196),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_163),
.Y(n_221)
);

INVx4_ASAP7_75t_L g222 ( 
.A(n_186),
.Y(n_222)
);

INVxp67_ASAP7_75t_L g223 ( 
.A(n_169),
.Y(n_223)
);

BUFx6f_ASAP7_75t_L g224 ( 
.A(n_186),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_175),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_165),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g227 ( 
.A(n_154),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_171),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_174),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_180),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_159),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_181),
.Y(n_232)
);

BUFx8_ASAP7_75t_SL g233 ( 
.A(n_159),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_154),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_184),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_178),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

BUFx8_ASAP7_75t_SL g238 ( 
.A(n_172),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_208),
.B(n_2),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_168),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_170),
.Y(n_244)
);

BUFx8_ASAP7_75t_SL g245 ( 
.A(n_179),
.Y(n_245)
);

AND2x4_ASAP7_75t_L g246 ( 
.A(n_185),
.B(n_3),
.Y(n_246)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_189),
.Y(n_247)
);

AOI22x1_ASAP7_75t_SL g248 ( 
.A1(n_197),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_248)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_203),
.B(n_207),
.Y(n_249)
);

INVx5_ASAP7_75t_L g250 ( 
.A(n_202),
.Y(n_250)
);

AND2x4_ASAP7_75t_L g251 ( 
.A(n_202),
.B(n_8),
.Y(n_251)
);

INVx4_ASAP7_75t_L g252 ( 
.A(n_157),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_158),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_242),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_218),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_244),
.B(n_160),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_224),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g258 ( 
.A(n_245),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_241),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g260 ( 
.A(n_241),
.B(n_162),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_220),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_214),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_233),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_227),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_238),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_227),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_227),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_R g270 ( 
.A(n_225),
.B(n_164),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_245),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_201),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_210),
.Y(n_273)
);

OAI22xp5_ASAP7_75t_L g274 ( 
.A1(n_219),
.A2(n_209),
.B1(n_205),
.B2(n_204),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_210),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_253),
.Y(n_276)
);

NAND2xp33_ASAP7_75t_L g277 ( 
.A(n_249),
.B(n_167),
.Y(n_277)
);

NOR2xp67_ASAP7_75t_L g278 ( 
.A(n_223),
.B(n_252),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_253),
.Y(n_279)
);

INVx2_ASAP7_75t_L g280 ( 
.A(n_224),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_R g281 ( 
.A(n_253),
.B(n_173),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_253),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_247),
.Y(n_283)
);

INVx3_ASAP7_75t_L g284 ( 
.A(n_214),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_216),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_216),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g287 ( 
.A(n_223),
.Y(n_287)
);

INVx2_ASAP7_75t_L g288 ( 
.A(n_222),
.Y(n_288)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_224),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_R g290 ( 
.A(n_221),
.B(n_176),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_222),
.Y(n_291)
);

OA21x2_ASAP7_75t_L g292 ( 
.A1(n_239),
.A2(n_199),
.B(n_200),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_227),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_226),
.Y(n_294)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_224),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_234),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_234),
.Y(n_297)
);

INVx2_ASAP7_75t_SL g298 ( 
.A(n_229),
.Y(n_298)
);

HB1xp67_ASAP7_75t_L g299 ( 
.A(n_213),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_232),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_234),
.Y(n_301)
);

INVxp33_ASAP7_75t_L g302 ( 
.A(n_260),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_299),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_284),
.B(n_246),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_294),
.A2(n_211),
.B1(n_251),
.B2(n_246),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_284),
.B(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_255),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_296),
.Y(n_308)
);

NAND3xp33_ASAP7_75t_L g309 ( 
.A(n_300),
.B(n_231),
.C(n_251),
.Y(n_309)
);

AND2x4_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_213),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_263),
.B(n_250),
.Y(n_311)
);

NOR2xp67_ASAP7_75t_L g312 ( 
.A(n_285),
.B(n_250),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_262),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_254),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_272),
.B(n_228),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_290),
.B(n_228),
.Y(n_316)
);

NOR2xp67_ASAP7_75t_L g317 ( 
.A(n_286),
.B(n_250),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_288),
.Y(n_318)
);

NOR3xp33_ASAP7_75t_L g319 ( 
.A(n_274),
.B(n_217),
.C(n_230),
.Y(n_319)
);

NOR2xp67_ASAP7_75t_L g320 ( 
.A(n_258),
.B(n_250),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_290),
.B(n_230),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_276),
.B(n_235),
.Y(n_322)
);

INVx2_ASAP7_75t_SL g323 ( 
.A(n_287),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_297),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_265),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_279),
.B(n_237),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_282),
.B(n_217),
.Y(n_327)
);

INVxp67_ASAP7_75t_L g328 ( 
.A(n_256),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_268),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_291),
.B(n_234),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_277),
.B(n_236),
.Y(n_331)
);

INVx2_ASAP7_75t_SL g332 ( 
.A(n_283),
.Y(n_332)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_271),
.B(n_248),
.C(n_212),
.Y(n_333)
);

INVxp33_ASAP7_75t_L g334 ( 
.A(n_270),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_269),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_293),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g337 ( 
.A(n_278),
.B(n_236),
.Y(n_337)
);

NAND3xp33_ASAP7_75t_L g338 ( 
.A(n_292),
.B(n_243),
.C(n_240),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_292),
.A2(n_243),
.B1(n_236),
.B2(n_240),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_301),
.B(n_236),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_257),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_292),
.B(n_240),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_257),
.B(n_240),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_SL g344 ( 
.A(n_270),
.B(n_177),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_295),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_280),
.B(n_243),
.Y(n_346)
);

INVx2_ASAP7_75t_SL g347 ( 
.A(n_281),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_280),
.B(n_243),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_289),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_289),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_281),
.B(n_182),
.Y(n_351)
);

NAND2xp5_ASAP7_75t_SL g352 ( 
.A(n_295),
.B(n_183),
.Y(n_352)
);

NOR2xp67_ASAP7_75t_L g353 ( 
.A(n_273),
.B(n_215),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_295),
.Y(n_354)
);

NOR3xp33_ASAP7_75t_L g355 ( 
.A(n_261),
.B(n_188),
.C(n_190),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_275),
.B(n_215),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_295),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_264),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_266),
.B(n_215),
.Y(n_359)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_259),
.Y(n_360)
);

HB1xp67_ASAP7_75t_L g361 ( 
.A(n_267),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_284),
.B(n_215),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_284),
.B(n_191),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_284),
.B(n_192),
.Y(n_364)
);

NAND3xp33_ASAP7_75t_L g365 ( 
.A(n_294),
.B(n_198),
.C(n_195),
.Y(n_365)
);

OR2x2_ASAP7_75t_SL g366 ( 
.A(n_309),
.B(n_8),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_336),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_328),
.A2(n_194),
.B1(n_10),
.B2(n_11),
.Y(n_368)
);

NAND2x1p5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_353),
.Y(n_369)
);

INVx5_ASAP7_75t_L g370 ( 
.A(n_310),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_318),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_315),
.B(n_9),
.Y(n_372)
);

INVx2_ASAP7_75t_L g373 ( 
.A(n_308),
.Y(n_373)
);

INVx2_ASAP7_75t_SL g374 ( 
.A(n_323),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_345),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_307),
.Y(n_376)
);

NOR2x1_ASAP7_75t_L g377 ( 
.A(n_356),
.B(n_16),
.Y(n_377)
);

INVx3_ASAP7_75t_L g378 ( 
.A(n_345),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_313),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_332),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_322),
.B(n_12),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_326),
.B(n_13),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_L g383 ( 
.A1(n_305),
.A2(n_14),
.B1(n_15),
.B2(n_18),
.Y(n_383)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_334),
.B(n_14),
.Y(n_384)
);

NOR2x1p5_ASAP7_75t_L g385 ( 
.A(n_314),
.B(n_15),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_358),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_350),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_310),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_342),
.B(n_331),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_327),
.Y(n_390)
);

INVx3_ASAP7_75t_L g391 ( 
.A(n_345),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_304),
.B(n_148),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_365),
.B(n_19),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_324),
.Y(n_394)
);

AND2x6_ASAP7_75t_SL g395 ( 
.A(n_359),
.B(n_22),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g396 ( 
.A(n_304),
.B(n_23),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_319),
.B(n_24),
.Y(n_397)
);

INVx5_ASAP7_75t_L g398 ( 
.A(n_358),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_341),
.Y(n_399)
);

BUFx6f_ASAP7_75t_L g400 ( 
.A(n_357),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_306),
.B(n_27),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_325),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_343),
.Y(n_403)
);

INVx2_ASAP7_75t_SL g404 ( 
.A(n_360),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_306),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_405)
);

AND2x2_ASAP7_75t_SL g406 ( 
.A(n_358),
.B(n_35),
.Y(n_406)
);

AND2x4_ASAP7_75t_L g407 ( 
.A(n_320),
.B(n_37),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_363),
.B(n_41),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_302),
.A2(n_42),
.B1(n_43),
.B2(n_44),
.Y(n_409)
);

INVx5_ASAP7_75t_L g410 ( 
.A(n_349),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_361),
.Y(n_411)
);

BUFx3_ASAP7_75t_L g412 ( 
.A(n_303),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_329),
.Y(n_413)
);

A2O1A1Ixp33_ASAP7_75t_L g414 ( 
.A1(n_337),
.A2(n_46),
.B(n_47),
.C(n_48),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_316),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_415)
);

NOR2x1p5_ASAP7_75t_L g416 ( 
.A(n_355),
.B(n_53),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_330),
.B(n_321),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_363),
.B(n_145),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_364),
.B(n_56),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_344),
.B(n_142),
.Y(n_420)
);

NOR3xp33_ASAP7_75t_SL g421 ( 
.A(n_352),
.B(n_57),
.C(n_58),
.Y(n_421)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_312),
.Y(n_422)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_335),
.Y(n_423)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_317),
.Y(n_424)
);

INVx2_ASAP7_75t_SL g425 ( 
.A(n_340),
.Y(n_425)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_364),
.B(n_59),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_340),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_343),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_346),
.Y(n_429)
);

BUFx3_ASAP7_75t_L g430 ( 
.A(n_354),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_351),
.B(n_140),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g432 ( 
.A(n_348),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_392),
.A2(n_362),
.B(n_338),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_390),
.B(n_333),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_379),
.Y(n_437)
);

O2A1O1Ixp33_ASAP7_75t_L g438 ( 
.A1(n_372),
.A2(n_362),
.B(n_311),
.C(n_339),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_380),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_371),
.Y(n_440)
);

OR2x2_ASAP7_75t_L g441 ( 
.A(n_412),
.B(n_61),
.Y(n_441)
);

BUFx2_ASAP7_75t_L g442 ( 
.A(n_411),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g443 ( 
.A(n_370),
.B(n_62),
.Y(n_443)
);

OAI22xp33_ASAP7_75t_L g444 ( 
.A1(n_381),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_386),
.Y(n_445)
);

NAND2xp33_ASAP7_75t_L g446 ( 
.A(n_418),
.B(n_69),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_399),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_370),
.B(n_70),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_370),
.B(n_425),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_373),
.Y(n_450)
);

AOI22xp33_ASAP7_75t_L g451 ( 
.A1(n_388),
.A2(n_71),
.B1(n_72),
.B2(n_74),
.Y(n_451)
);

INVx6_ASAP7_75t_L g452 ( 
.A(n_398),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_387),
.Y(n_453)
);

O2A1O1Ixp33_ASAP7_75t_L g454 ( 
.A1(n_382),
.A2(n_75),
.B(n_76),
.C(n_77),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_427),
.B(n_79),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_394),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_387),
.Y(n_457)
);

AOI21xp5_ASAP7_75t_L g458 ( 
.A1(n_396),
.A2(n_80),
.B(n_81),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_402),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g460 ( 
.A1(n_401),
.A2(n_83),
.B(n_85),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_403),
.B(n_86),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_398),
.B(n_87),
.Y(n_462)
);

INVx1_ASAP7_75t_SL g463 ( 
.A(n_374),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_413),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_404),
.B(n_138),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_398),
.Y(n_466)
);

NAND2xp5_ASAP7_75t_SL g467 ( 
.A(n_406),
.B(n_88),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_384),
.B(n_89),
.Y(n_468)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_417),
.B(n_90),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_395),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_423),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_428),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_432),
.B(n_137),
.Y(n_473)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_419),
.A2(n_426),
.B(n_397),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_385),
.B(n_91),
.Y(n_475)
);

INVx1_ASAP7_75t_SL g476 ( 
.A(n_366),
.Y(n_476)
);

A2O1A1Ixp33_ASAP7_75t_L g477 ( 
.A1(n_383),
.A2(n_92),
.B(n_93),
.C(n_94),
.Y(n_477)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_408),
.A2(n_95),
.B(n_96),
.Y(n_478)
);

OR2x6_ASAP7_75t_L g479 ( 
.A(n_369),
.B(n_98),
.Y(n_479)
);

AOI22xp33_ASAP7_75t_L g480 ( 
.A1(n_403),
.A2(n_99),
.B1(n_100),
.B2(n_102),
.Y(n_480)
);

O2A1O1Ixp33_ASAP7_75t_SL g481 ( 
.A1(n_393),
.A2(n_103),
.B(n_105),
.C(n_106),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_422),
.B(n_108),
.Y(n_482)
);

OAI221xp5_ASAP7_75t_L g483 ( 
.A1(n_368),
.A2(n_111),
.B1(n_112),
.B2(n_114),
.C(n_116),
.Y(n_483)
);

A2O1A1Ixp33_ASAP7_75t_L g484 ( 
.A1(n_431),
.A2(n_117),
.B(n_120),
.C(n_121),
.Y(n_484)
);

AND2x2_ASAP7_75t_L g485 ( 
.A(n_424),
.B(n_122),
.Y(n_485)
);

BUFx6f_ASAP7_75t_L g486 ( 
.A(n_452),
.Y(n_486)
);

OAI21x1_ASAP7_75t_L g487 ( 
.A1(n_433),
.A2(n_377),
.B(n_405),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_434),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_453),
.Y(n_489)
);

AO21x2_ASAP7_75t_L g490 ( 
.A1(n_474),
.A2(n_429),
.B(n_415),
.Y(n_490)
);

INVx4_ASAP7_75t_L g491 ( 
.A(n_452),
.Y(n_491)
);

INVx2_ASAP7_75t_SL g492 ( 
.A(n_452),
.Y(n_492)
);

AO21x2_ASAP7_75t_L g493 ( 
.A1(n_474),
.A2(n_421),
.B(n_414),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_457),
.Y(n_494)
);

BUFx6f_ASAP7_75t_L g495 ( 
.A(n_436),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_437),
.Y(n_496)
);

BUFx2_ASAP7_75t_R g497 ( 
.A(n_445),
.Y(n_497)
);

OAI21xp5_ASAP7_75t_L g498 ( 
.A1(n_472),
.A2(n_420),
.B(n_389),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_459),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g500 ( 
.A(n_435),
.B(n_430),
.Y(n_500)
);

AO21x2_ASAP7_75t_L g501 ( 
.A1(n_433),
.A2(n_407),
.B(n_389),
.Y(n_501)
);

AOI22x1_ASAP7_75t_L g502 ( 
.A1(n_478),
.A2(n_416),
.B1(n_375),
.B2(n_378),
.Y(n_502)
);

OAI21xp5_ASAP7_75t_L g503 ( 
.A1(n_473),
.A2(n_389),
.B(n_375),
.Y(n_503)
);

INVx3_ASAP7_75t_L g504 ( 
.A(n_479),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_464),
.Y(n_505)
);

INVx1_ASAP7_75t_SL g506 ( 
.A(n_439),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_442),
.Y(n_507)
);

INVxp67_ASAP7_75t_SL g508 ( 
.A(n_441),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_471),
.Y(n_509)
);

OAI21xp5_ASAP7_75t_L g510 ( 
.A1(n_438),
.A2(n_389),
.B(n_391),
.Y(n_510)
);

BUFx2_ASAP7_75t_L g511 ( 
.A(n_466),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_461),
.A2(n_391),
.B(n_378),
.Y(n_512)
);

AND2x4_ASAP7_75t_L g513 ( 
.A(n_440),
.B(n_410),
.Y(n_513)
);

INVx1_ASAP7_75t_SL g514 ( 
.A(n_463),
.Y(n_514)
);

INVx3_ASAP7_75t_L g515 ( 
.A(n_479),
.Y(n_515)
);

HB1xp67_ASAP7_75t_L g516 ( 
.A(n_476),
.Y(n_516)
);

INVx3_ASAP7_75t_L g517 ( 
.A(n_479),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_447),
.Y(n_518)
);

OAI21x1_ASAP7_75t_L g519 ( 
.A1(n_458),
.A2(n_460),
.B(n_478),
.Y(n_519)
);

INVx3_ASAP7_75t_L g520 ( 
.A(n_450),
.Y(n_520)
);

AO21x2_ASAP7_75t_L g521 ( 
.A1(n_468),
.A2(n_407),
.B(n_400),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_456),
.Y(n_522)
);

OAI21x1_ASAP7_75t_L g523 ( 
.A1(n_458),
.A2(n_400),
.B(n_410),
.Y(n_523)
);

AND2x2_ASAP7_75t_L g524 ( 
.A(n_467),
.B(n_410),
.Y(n_524)
);

OAI21x1_ASAP7_75t_L g525 ( 
.A1(n_460),
.A2(n_400),
.B(n_409),
.Y(n_525)
);

BUFx6f_ASAP7_75t_L g526 ( 
.A(n_462),
.Y(n_526)
);

OAI21x1_ASAP7_75t_L g527 ( 
.A1(n_454),
.A2(n_123),
.B(n_125),
.Y(n_527)
);

OR2x6_ASAP7_75t_L g528 ( 
.A(n_485),
.B(n_126),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_449),
.B(n_127),
.Y(n_529)
);

AOI22x1_ASAP7_75t_L g530 ( 
.A1(n_475),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_530)
);

BUFx8_ASAP7_75t_SL g531 ( 
.A(n_511),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_489),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_489),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_494),
.Y(n_534)
);

INVx11_ASAP7_75t_L g535 ( 
.A(n_497),
.Y(n_535)
);

AOI22xp33_ASAP7_75t_L g536 ( 
.A1(n_508),
.A2(n_483),
.B1(n_465),
.B2(n_455),
.Y(n_536)
);

OAI22xp5_ASAP7_75t_L g537 ( 
.A1(n_500),
.A2(n_469),
.B1(n_477),
.B2(n_470),
.Y(n_537)
);

INVx2_ASAP7_75t_L g538 ( 
.A(n_494),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_518),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_488),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_486),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g542 ( 
.A(n_511),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_496),
.B(n_482),
.Y(n_543)
);

OAI22x1_ASAP7_75t_L g544 ( 
.A1(n_504),
.A2(n_448),
.B1(n_443),
.B2(n_444),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_499),
.Y(n_545)
);

CKINVDCx11_ASAP7_75t_R g546 ( 
.A(n_514),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_522),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g548 ( 
.A1(n_519),
.A2(n_446),
.B(n_481),
.Y(n_548)
);

AND2x4_ASAP7_75t_SL g549 ( 
.A(n_491),
.B(n_451),
.Y(n_549)
);

BUFx2_ASAP7_75t_L g550 ( 
.A(n_510),
.Y(n_550)
);

AND2x4_ASAP7_75t_L g551 ( 
.A(n_504),
.B(n_484),
.Y(n_551)
);

OA21x2_ASAP7_75t_L g552 ( 
.A1(n_512),
.A2(n_480),
.B(n_132),
.Y(n_552)
);

OAI21xp33_ASAP7_75t_SL g553 ( 
.A1(n_528),
.A2(n_134),
.B(n_503),
.Y(n_553)
);

BUFx2_ASAP7_75t_R g554 ( 
.A(n_504),
.Y(n_554)
);

AO21x2_ASAP7_75t_L g555 ( 
.A1(n_501),
.A2(n_498),
.B(n_519),
.Y(n_555)
);

BUFx3_ASAP7_75t_L g556 ( 
.A(n_486),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_506),
.B(n_516),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_505),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_491),
.Y(n_559)
);

BUFx12f_ASAP7_75t_L g560 ( 
.A(n_486),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_486),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_509),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_507),
.Y(n_563)
);

INVx3_ASAP7_75t_L g564 ( 
.A(n_491),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_520),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_520),
.Y(n_566)
);

AOI22xp33_ASAP7_75t_L g567 ( 
.A1(n_528),
.A2(n_517),
.B1(n_515),
.B2(n_520),
.Y(n_567)
);

AO21x1_ASAP7_75t_L g568 ( 
.A1(n_525),
.A2(n_487),
.B(n_527),
.Y(n_568)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_486),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_L g570 ( 
.A1(n_528),
.A2(n_502),
.B1(n_517),
.B2(n_515),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_517),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_539),
.Y(n_572)
);

NAND3xp33_ASAP7_75t_SL g573 ( 
.A(n_537),
.B(n_524),
.C(n_528),
.Y(n_573)
);

OAI22xp5_ASAP7_75t_L g574 ( 
.A1(n_536),
.A2(n_515),
.B1(n_502),
.B2(n_524),
.Y(n_574)
);

HB1xp67_ASAP7_75t_L g575 ( 
.A(n_569),
.Y(n_575)
);

AND2x4_ASAP7_75t_L g576 ( 
.A(n_541),
.B(n_513),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_R g577 ( 
.A(n_546),
.B(n_492),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_539),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_560),
.B(n_492),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_547),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_543),
.B(n_513),
.Y(n_581)
);

OR2x2_ASAP7_75t_L g582 ( 
.A(n_540),
.B(n_495),
.Y(n_582)
);

AND2x4_ASAP7_75t_L g583 ( 
.A(n_541),
.B(n_513),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_547),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_R g585 ( 
.A(n_542),
.B(n_526),
.Y(n_585)
);

INVx8_ASAP7_75t_L g586 ( 
.A(n_560),
.Y(n_586)
);

OAI22xp5_ASAP7_75t_SL g587 ( 
.A1(n_567),
.A2(n_529),
.B1(n_526),
.B2(n_525),
.Y(n_587)
);

NOR2x1_ASAP7_75t_L g588 ( 
.A(n_556),
.B(n_529),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_540),
.Y(n_589)
);

OR2x2_ASAP7_75t_L g590 ( 
.A(n_545),
.B(n_495),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_541),
.B(n_529),
.Y(n_591)
);

AND2x2_ASAP7_75t_L g592 ( 
.A(n_543),
.B(n_495),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_557),
.B(n_495),
.Y(n_593)
);

OAI21xp5_ASAP7_75t_L g594 ( 
.A1(n_553),
.A2(n_487),
.B(n_527),
.Y(n_594)
);

OR2x2_ASAP7_75t_L g595 ( 
.A(n_545),
.B(n_495),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_535),
.Y(n_596)
);

AOI22xp33_ASAP7_75t_L g597 ( 
.A1(n_550),
.A2(n_521),
.B1(n_501),
.B2(n_530),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_533),
.B(n_521),
.Y(n_598)
);

INVx4_ASAP7_75t_L g599 ( 
.A(n_535),
.Y(n_599)
);

AND2x2_ASAP7_75t_L g600 ( 
.A(n_554),
.B(n_501),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_558),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_561),
.B(n_526),
.Y(n_602)
);

CKINVDCx11_ASAP7_75t_R g603 ( 
.A(n_556),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_558),
.Y(n_604)
);

NOR3xp33_ASAP7_75t_SL g605 ( 
.A(n_553),
.B(n_493),
.C(n_530),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_533),
.Y(n_607)
);

AND2x4_ASAP7_75t_L g608 ( 
.A(n_561),
.B(n_526),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_531),
.Y(n_609)
);

NAND2x1p5_ASAP7_75t_L g610 ( 
.A(n_561),
.B(n_523),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_562),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_559),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_562),
.B(n_490),
.Y(n_613)
);

INVx1_ASAP7_75t_L g614 ( 
.A(n_534),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_R g615 ( 
.A(n_559),
.B(n_564),
.Y(n_615)
);

NAND2xp33_ASAP7_75t_R g616 ( 
.A(n_551),
.B(n_523),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_607),
.Y(n_617)
);

INVx2_ASAP7_75t_SL g618 ( 
.A(n_575),
.Y(n_618)
);

NOR2x1_ASAP7_75t_SL g619 ( 
.A(n_573),
.B(n_570),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_607),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_592),
.B(n_555),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_L g622 ( 
.A(n_581),
.B(n_593),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_601),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_604),
.Y(n_624)
);

AND2x4_ASAP7_75t_L g625 ( 
.A(n_608),
.B(n_534),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_571),
.B(n_538),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_608),
.B(n_589),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_611),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_587),
.A2(n_551),
.B1(n_549),
.B2(n_544),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_614),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_612),
.B(n_538),
.Y(n_631)
);

AND2x4_ASAP7_75t_L g632 ( 
.A(n_591),
.B(n_551),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_613),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_572),
.Y(n_634)
);

HB1xp67_ASAP7_75t_L g635 ( 
.A(n_582),
.Y(n_635)
);

INVx2_ASAP7_75t_SL g636 ( 
.A(n_590),
.Y(n_636)
);

AOI22xp33_ASAP7_75t_L g637 ( 
.A1(n_600),
.A2(n_551),
.B1(n_544),
.B2(n_566),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_578),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_576),
.B(n_566),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_595),
.B(n_555),
.Y(n_640)
);

AND2x2_ASAP7_75t_L g641 ( 
.A(n_580),
.B(n_555),
.Y(n_641)
);

HB1xp67_ASAP7_75t_L g642 ( 
.A(n_585),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_584),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_606),
.Y(n_644)
);

OR2x2_ASAP7_75t_L g645 ( 
.A(n_598),
.B(n_565),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_610),
.Y(n_646)
);

INVx4_ASAP7_75t_L g647 ( 
.A(n_603),
.Y(n_647)
);

HB1xp67_ASAP7_75t_L g648 ( 
.A(n_602),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_602),
.Y(n_649)
);

NAND3xp33_ASAP7_75t_L g650 ( 
.A(n_637),
.B(n_605),
.C(n_594),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_617),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_623),
.Y(n_652)
);

INVx2_ASAP7_75t_SL g653 ( 
.A(n_618),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_617),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_621),
.B(n_597),
.Y(n_655)
);

AND2x2_ASAP7_75t_L g656 ( 
.A(n_621),
.B(n_568),
.Y(n_656)
);

AND2x4_ASAP7_75t_L g657 ( 
.A(n_627),
.B(n_591),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_627),
.B(n_576),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_624),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_618),
.Y(n_660)
);

OR2x2_ASAP7_75t_L g661 ( 
.A(n_633),
.B(n_568),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_628),
.Y(n_662)
);

INVx2_ASAP7_75t_L g663 ( 
.A(n_620),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_640),
.B(n_583),
.Y(n_664)
);

AND2x2_ASAP7_75t_L g665 ( 
.A(n_640),
.B(n_583),
.Y(n_665)
);

AND2x2_ASAP7_75t_L g666 ( 
.A(n_633),
.B(n_574),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_630),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_L g668 ( 
.A(n_635),
.B(n_615),
.Y(n_668)
);

BUFx2_ASAP7_75t_L g669 ( 
.A(n_627),
.Y(n_669)
);

AND2x2_ASAP7_75t_SL g670 ( 
.A(n_632),
.B(n_629),
.Y(n_670)
);

NOR2x1p5_ASAP7_75t_L g671 ( 
.A(n_647),
.B(n_599),
.Y(n_671)
);

AND2x2_ASAP7_75t_L g672 ( 
.A(n_620),
.B(n_552),
.Y(n_672)
);

OR2x2_ASAP7_75t_L g673 ( 
.A(n_636),
.B(n_645),
.Y(n_673)
);

BUFx2_ASAP7_75t_L g674 ( 
.A(n_647),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_667),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_652),
.Y(n_676)
);

AND2x2_ASAP7_75t_L g677 ( 
.A(n_669),
.B(n_636),
.Y(n_677)
);

AND2x2_ASAP7_75t_L g678 ( 
.A(n_669),
.B(n_632),
.Y(n_678)
);

AND2x2_ASAP7_75t_L g679 ( 
.A(n_660),
.B(n_647),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_653),
.B(n_622),
.Y(n_680)
);

AND2x2_ASAP7_75t_L g681 ( 
.A(n_656),
.B(n_632),
.Y(n_681)
);

INVx2_ASAP7_75t_L g682 ( 
.A(n_651),
.Y(n_682)
);

INVx2_ASAP7_75t_SL g683 ( 
.A(n_653),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_657),
.B(n_646),
.Y(n_684)
);

OAI221xp5_ASAP7_75t_L g685 ( 
.A1(n_650),
.A2(n_631),
.B1(n_626),
.B2(n_588),
.C(n_639),
.Y(n_685)
);

OR2x2_ASAP7_75t_L g686 ( 
.A(n_673),
.B(n_645),
.Y(n_686)
);

AND2x2_ASAP7_75t_L g687 ( 
.A(n_656),
.B(n_641),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_657),
.B(n_630),
.Y(n_688)
);

AND2x4_ASAP7_75t_L g689 ( 
.A(n_657),
.B(n_641),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_675),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_682),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_676),
.Y(n_692)
);

OR2x2_ASAP7_75t_L g693 ( 
.A(n_686),
.B(n_673),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_682),
.Y(n_694)
);

HB1xp67_ASAP7_75t_L g695 ( 
.A(n_677),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_687),
.B(n_666),
.Y(n_696)
);

OAI22xp5_ASAP7_75t_L g697 ( 
.A1(n_685),
.A2(n_670),
.B1(n_668),
.B2(n_674),
.Y(n_697)
);

INVx2_ASAP7_75t_L g698 ( 
.A(n_688),
.Y(n_698)
);

OR2x2_ASAP7_75t_L g699 ( 
.A(n_687),
.B(n_661),
.Y(n_699)
);

XOR2x2_ASAP7_75t_L g700 ( 
.A(n_697),
.B(n_670),
.Y(n_700)
);

INVxp67_ASAP7_75t_L g701 ( 
.A(n_692),
.Y(n_701)
);

XNOR2x1_ASAP7_75t_L g702 ( 
.A(n_693),
.B(n_679),
.Y(n_702)
);

OR2x2_ASAP7_75t_L g703 ( 
.A(n_696),
.B(n_680),
.Y(n_703)
);

INVx1_ASAP7_75t_L g704 ( 
.A(n_701),
.Y(n_704)
);

NOR2xp33_ASAP7_75t_L g705 ( 
.A(n_702),
.B(n_609),
.Y(n_705)
);

INVx1_ASAP7_75t_L g706 ( 
.A(n_703),
.Y(n_706)
);

INVx2_ASAP7_75t_SL g707 ( 
.A(n_700),
.Y(n_707)
);

NOR3xp33_ASAP7_75t_SL g708 ( 
.A(n_700),
.B(n_596),
.C(n_671),
.Y(n_708)
);

INVx1_ASAP7_75t_SL g709 ( 
.A(n_705),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_704),
.B(n_599),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_706),
.Y(n_711)
);

AOI21xp5_ASAP7_75t_L g712 ( 
.A1(n_707),
.A2(n_690),
.B(n_683),
.Y(n_712)
);

AOI211xp5_ASAP7_75t_L g713 ( 
.A1(n_712),
.A2(n_577),
.B(n_708),
.C(n_690),
.Y(n_713)
);

AOI22xp5_ASAP7_75t_L g714 ( 
.A1(n_709),
.A2(n_655),
.B1(n_666),
.B2(n_659),
.Y(n_714)
);

AOI211xp5_ASAP7_75t_L g715 ( 
.A1(n_711),
.A2(n_699),
.B(n_662),
.C(n_642),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_714),
.B(n_710),
.Y(n_716)
);

AOI211xp5_ASAP7_75t_L g717 ( 
.A1(n_713),
.A2(n_695),
.B(n_661),
.C(n_655),
.Y(n_717)
);

INVxp67_ASAP7_75t_L g718 ( 
.A(n_715),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_SL g719 ( 
.A1(n_718),
.A2(n_564),
.B(n_559),
.C(n_677),
.Y(n_719)
);

NOR2x1_ASAP7_75t_L g720 ( 
.A(n_716),
.B(n_579),
.Y(n_720)
);

NOR2x1_ASAP7_75t_L g721 ( 
.A(n_717),
.B(n_579),
.Y(n_721)
);

AOI22xp5_ASAP7_75t_L g722 ( 
.A1(n_718),
.A2(n_684),
.B1(n_616),
.B2(n_694),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_716),
.Y(n_723)
);

NOR2xp33_ASAP7_75t_L g724 ( 
.A(n_718),
.B(n_683),
.Y(n_724)
);

AND2x2_ASAP7_75t_SL g725 ( 
.A(n_723),
.B(n_724),
.Y(n_725)
);

NAND4xp25_ASAP7_75t_L g726 ( 
.A(n_719),
.B(n_678),
.C(n_681),
.D(n_684),
.Y(n_726)
);

AND2x2_ASAP7_75t_L g727 ( 
.A(n_720),
.B(n_681),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_721),
.Y(n_728)
);

AOI221xp5_ASAP7_75t_L g729 ( 
.A1(n_722),
.A2(n_672),
.B1(n_691),
.B2(n_493),
.C(n_634),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_723),
.B(n_678),
.Y(n_730)
);

NAND3x1_ASAP7_75t_L g731 ( 
.A(n_723),
.B(n_586),
.C(n_564),
.Y(n_731)
);

INVx2_ASAP7_75t_SL g732 ( 
.A(n_730),
.Y(n_732)
);

INVx2_ASAP7_75t_SL g733 ( 
.A(n_725),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_728),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_727),
.Y(n_735)
);

NOR2xp33_ASAP7_75t_R g736 ( 
.A(n_731),
.B(n_586),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_726),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_729),
.B(n_698),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_730),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_725),
.B(n_684),
.Y(n_740)
);

AOI22xp5_ASAP7_75t_L g741 ( 
.A1(n_735),
.A2(n_688),
.B1(n_689),
.B2(n_625),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_733),
.B(n_732),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_739),
.Y(n_743)
);

AOI22x1_ASAP7_75t_L g744 ( 
.A1(n_734),
.A2(n_689),
.B1(n_688),
.B2(n_658),
.Y(n_744)
);

HB1xp67_ASAP7_75t_L g745 ( 
.A(n_737),
.Y(n_745)
);

AND3x1_ASAP7_75t_L g746 ( 
.A(n_740),
.B(n_665),
.C(n_664),
.Y(n_746)
);

OAI22x1_ASAP7_75t_L g747 ( 
.A1(n_738),
.A2(n_689),
.B1(n_658),
.B2(n_648),
.Y(n_747)
);

NOR2xp33_ASAP7_75t_R g748 ( 
.A(n_736),
.B(n_548),
.Y(n_748)
);

AO22x2_ASAP7_75t_L g749 ( 
.A1(n_736),
.A2(n_638),
.B1(n_643),
.B2(n_649),
.Y(n_749)
);

XOR2xp5_ASAP7_75t_L g750 ( 
.A(n_735),
.B(n_619),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_742),
.Y(n_751)
);

HB1xp67_ASAP7_75t_L g752 ( 
.A(n_743),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_745),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_746),
.Y(n_754)
);

INVx5_ASAP7_75t_L g755 ( 
.A(n_750),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_741),
.B(n_658),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_752),
.Y(n_757)
);

OAI22xp5_ASAP7_75t_SL g758 ( 
.A1(n_753),
.A2(n_747),
.B1(n_744),
.B2(n_748),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_751),
.B(n_749),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_754),
.Y(n_760)
);

AOI22xp5_ASAP7_75t_SL g761 ( 
.A1(n_755),
.A2(n_749),
.B1(n_552),
.B2(n_672),
.Y(n_761)
);

BUFx2_ASAP7_75t_L g762 ( 
.A(n_757),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_SL g763 ( 
.A1(n_760),
.A2(n_755),
.B1(n_756),
.B2(n_552),
.Y(n_763)
);

AOI22x1_ASAP7_75t_L g764 ( 
.A1(n_761),
.A2(n_651),
.B1(n_654),
.B2(n_663),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_762),
.B(n_759),
.Y(n_765)
);

AOI22xp5_ASAP7_75t_L g766 ( 
.A1(n_765),
.A2(n_758),
.B1(n_763),
.B2(n_764),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_766),
.A2(n_490),
.B1(n_663),
.B2(n_654),
.Y(n_767)
);

AOI22xp33_ASAP7_75t_L g768 ( 
.A1(n_767),
.A2(n_490),
.B1(n_644),
.B2(n_549),
.Y(n_768)
);


endmodule