module fake_jpeg_3185_n_62 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_62);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_62;

wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_19;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;

INVx6_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

BUFx4f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_22),
.Y(n_25)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_27),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_26),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx4_ASAP7_75t_SL g28 ( 
.A(n_24),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_28),
.B(n_29),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_29),
.A2(n_24),
.B1(n_23),
.B2(n_19),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_30),
.B(n_33),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_SL g33 ( 
.A(n_28),
.B(n_24),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_28),
.A2(n_19),
.B1(n_1),
.B2(n_3),
.Y(n_34)
);

INVxp33_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_31),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g42 ( 
.A(n_37),
.B(n_40),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_32),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_0),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g49 ( 
.A(n_44),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_34),
.Y(n_45)
);

XNOR2xp5_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_1),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_38),
.B(n_10),
.C(n_16),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_38),
.B1(n_4),
.B2(n_5),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_43),
.Y(n_53)
);

AO21x2_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_9),
.B(n_13),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_8),
.Y(n_54)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_54),
.B(n_55),
.C(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_6),
.C(n_11),
.Y(n_55)
);

MAJx2_ASAP7_75t_L g56 ( 
.A(n_48),
.B(n_12),
.C(n_18),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_52),
.B(n_49),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g60 ( 
.A1(n_59),
.A2(n_57),
.B(n_4),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_3),
.Y(n_62)
);


endmodule