module fake_jpeg_11510_n_56 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_56);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_56;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_25;
wire n_31;
wire n_17;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

AOI21xp33_ASAP7_75t_L g8 ( 
.A1(n_7),
.A2(n_4),
.B(n_3),
.Y(n_8)
);

INVxp67_ASAP7_75t_L g9 ( 
.A(n_5),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_3),
.Y(n_11)
);

INVx3_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_7),
.B(n_5),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_2),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g18 ( 
.A(n_14),
.B(n_0),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_18),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g19 ( 
.A(n_14),
.B(n_0),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_19),
.B(n_22),
.Y(n_30)
);

CKINVDCx9p33_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

INVx5_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_15),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_23),
.A2(n_9),
.B1(n_16),
.B2(n_13),
.Y(n_31)
);

INVx4_ASAP7_75t_SL g24 ( 
.A(n_10),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx3_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_25),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_26),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_8),
.B1(n_15),
.B2(n_10),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_18),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_31),
.B(n_25),
.Y(n_43)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_21),
.A2(n_15),
.B1(n_10),
.B2(n_11),
.Y(n_33)
);

OAI21xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_20),
.B(n_22),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g35 ( 
.A(n_23),
.B(n_17),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_17),
.C(n_16),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_43),
.B(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_26),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_36),
.B(n_34),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_41),
.B(n_42),
.C(n_35),
.Y(n_45)
);

MAJIxp5_ASAP7_75t_L g42 ( 
.A(n_28),
.B(n_19),
.C(n_10),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_45),
.B(n_46),
.Y(n_50)
);

BUFx24_ASAP7_75t_SL g47 ( 
.A(n_43),
.Y(n_47)
);

OAI211xp5_ASAP7_75t_L g51 ( 
.A1(n_47),
.A2(n_48),
.B(n_36),
.C(n_31),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_44),
.B(n_30),
.C(n_33),
.Y(n_49)
);

MAJx2_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_51),
.C(n_50),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_47),
.A2(n_11),
.B1(n_25),
.B2(n_32),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_52),
.A2(n_32),
.B1(n_24),
.B2(n_4),
.Y(n_53)
);

AOI322xp5_ASAP7_75t_L g55 ( 
.A1(n_53),
.A2(n_54),
.A3(n_49),
.B1(n_2),
.B2(n_6),
.C1(n_1),
.C2(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_55),
.B(n_1),
.Y(n_56)
);


endmodule