module fake_netlist_1_143_n_18 (n_3, n_1, n_2, n_0, n_18);
input n_3;
input n_1;
input n_2;
input n_0;
output n_18;
wire n_11;
wire n_13;
wire n_16;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_17;
wire n_5;
wire n_14;
wire n_8;
wire n_15;
wire n_10;
wire n_7;
INVx4_ASAP7_75t_L g4 ( .A(n_1), .Y(n_4) );
INVx2_ASAP7_75t_L g5 ( .A(n_1), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_3), .B(n_2), .Y(n_6) );
BUFx4f_ASAP7_75t_L g7 ( .A(n_2), .Y(n_7) );
AND2x2_ASAP7_75t_L g8 ( .A(n_4), .B(n_0), .Y(n_8) );
INVx1_ASAP7_75t_L g9 ( .A(n_5), .Y(n_9) );
O2A1O1Ixp33_ASAP7_75t_SL g10 ( .A1(n_6), .A2(n_0), .B(n_3), .C(n_4), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AOI22xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_8), .B1(n_10), .B2(n_7), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_12), .B(n_9), .Y(n_14) );
AOI211xp5_ASAP7_75t_L g15 ( .A1(n_13), .A2(n_12), .B(n_7), .C(n_0), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
AND2x4_ASAP7_75t_L g17 ( .A(n_16), .B(n_15), .Y(n_17) );
AOI21xp5_ASAP7_75t_L g18 ( .A1(n_17), .A2(n_11), .B(n_16), .Y(n_18) );
endmodule