module real_aes_8374_n_98 (n_17, n_28, n_76, n_56, n_34, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_98);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_98;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_211;
wire n_693;
wire n_496;
wire n_281;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_363;
wire n_417;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_691;
wire n_481;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_456;
wire n_156;
wire n_359;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_99;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g420 ( .A(n_0), .Y(n_420) );
A2O1A1Ixp33_ASAP7_75t_L g432 ( .A1(n_1), .A2(n_118), .B(n_130), .C(n_433), .Y(n_432) );
INVx1_ASAP7_75t_L g237 ( .A(n_2), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_3), .A2(n_145), .B(n_472), .Y(n_471) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_4), .B(n_141), .Y(n_477) );
AOI21xp33_ASAP7_75t_L g144 ( .A1(n_5), .A2(n_145), .B(n_146), .Y(n_144) );
AND2x6_ASAP7_75t_L g118 ( .A(n_6), .B(n_119), .Y(n_118) );
AOI21xp5_ASAP7_75t_L g212 ( .A1(n_7), .A2(n_213), .B(n_214), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g421 ( .A(n_8), .B(n_39), .Y(n_421) );
INVx1_ASAP7_75t_L g448 ( .A(n_9), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g436 ( .A(n_10), .B(n_151), .Y(n_436) );
INVx1_ASAP7_75t_L g153 ( .A(n_11), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_12), .B(n_205), .Y(n_204) );
INVx1_ASAP7_75t_L g115 ( .A(n_13), .Y(n_115) );
INVx1_ASAP7_75t_L g219 ( .A(n_14), .Y(n_219) );
A2O1A1Ixp33_ASAP7_75t_L g456 ( .A1(n_15), .A2(n_154), .B(n_220), .C(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_16), .B(n_141), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_17), .B(n_164), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g173 ( .A(n_18), .B(n_145), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_19), .B(n_490), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_20), .A2(n_121), .B(n_205), .C(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g167 ( .A(n_21), .B(n_141), .Y(n_167) );
NAND2xp5_ASAP7_75t_SL g511 ( .A(n_22), .B(n_151), .Y(n_511) );
A2O1A1Ixp33_ASAP7_75t_L g216 ( .A1(n_23), .A2(n_217), .B(n_218), .C(n_220), .Y(n_216) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_24), .B(n_151), .Y(n_498) );
CKINVDCx16_ASAP7_75t_R g507 ( .A(n_25), .Y(n_507) );
INVx1_ASAP7_75t_L g497 ( .A(n_26), .Y(n_497) );
BUFx6f_ASAP7_75t_L g126 ( .A(n_27), .Y(n_126) );
CKINVDCx20_ASAP7_75t_R g431 ( .A(n_28), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g238 ( .A(n_29), .B(n_151), .Y(n_238) );
INVx1_ASAP7_75t_L g486 ( .A(n_30), .Y(n_486) );
INVx1_ASAP7_75t_L g129 ( .A(n_31), .Y(n_129) );
INVx2_ASAP7_75t_L g123 ( .A(n_32), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g438 ( .A(n_33), .Y(n_438) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_34), .A2(n_155), .B(n_205), .C(n_475), .Y(n_474) );
INVxp67_ASAP7_75t_L g487 ( .A(n_35), .Y(n_487) );
A2O1A1Ixp33_ASAP7_75t_L g174 ( .A1(n_36), .A2(n_118), .B(n_130), .C(n_175), .Y(n_174) );
CKINVDCx14_ASAP7_75t_R g473 ( .A(n_37), .Y(n_473) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_38), .A2(n_130), .B(n_496), .C(n_500), .Y(n_495) );
INVx1_ASAP7_75t_L g127 ( .A(n_40), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g446 ( .A1(n_41), .A2(n_150), .B(n_180), .C(n_447), .Y(n_446) );
NAND2xp5_ASAP7_75t_SL g190 ( .A(n_42), .B(n_151), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g502 ( .A(n_43), .Y(n_502) );
CKINVDCx20_ASAP7_75t_R g483 ( .A(n_44), .Y(n_483) );
INVx1_ASAP7_75t_L g463 ( .A(n_45), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g715 ( .A(n_46), .Y(n_715) );
CKINVDCx16_ASAP7_75t_R g133 ( .A(n_47), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_48), .B(n_145), .Y(n_207) );
AOI222xp33_ASAP7_75t_SL g100 ( .A1(n_49), .A2(n_58), .B1(n_101), .B2(n_690), .C1(n_691), .C2(n_695), .Y(n_100) );
AOI22xp5_ASAP7_75t_L g120 ( .A1(n_50), .A2(n_121), .B1(n_124), .B2(n_130), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g184 ( .A(n_51), .Y(n_184) );
CKINVDCx16_ASAP7_75t_R g234 ( .A(n_52), .Y(n_234) );
A2O1A1Ixp33_ASAP7_75t_L g149 ( .A1(n_53), .A2(n_150), .B(n_152), .C(n_155), .Y(n_149) );
CKINVDCx14_ASAP7_75t_R g445 ( .A(n_54), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_55), .Y(n_194) );
INVx1_ASAP7_75t_L g147 ( .A(n_56), .Y(n_147) );
INVx1_ASAP7_75t_L g119 ( .A(n_57), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_58), .Y(n_690) );
INVx1_ASAP7_75t_L g114 ( .A(n_59), .Y(n_114) );
INVx1_ASAP7_75t_SL g476 ( .A(n_60), .Y(n_476) );
CKINVDCx20_ASAP7_75t_R g704 ( .A(n_61), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_62), .B(n_141), .Y(n_467) );
AOI222xp33_ASAP7_75t_L g98 ( .A1(n_63), .A2(n_99), .B1(n_699), .B2(n_708), .C1(n_716), .C2(n_722), .Y(n_98) );
OAI22xp5_ASAP7_75t_SL g710 ( .A1(n_63), .A2(n_422), .B1(n_692), .B2(n_711), .Y(n_710) );
CKINVDCx20_ASAP7_75t_R g711 ( .A(n_63), .Y(n_711) );
INVx1_ASAP7_75t_L g510 ( .A(n_64), .Y(n_510) );
A2O1A1Ixp33_ASAP7_75t_SL g163 ( .A1(n_65), .A2(n_155), .B(n_164), .C(n_165), .Y(n_163) );
INVxp67_ASAP7_75t_L g166 ( .A(n_66), .Y(n_166) );
INVx1_ASAP7_75t_L g703 ( .A(n_67), .Y(n_703) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_68), .A2(n_145), .B(n_444), .Y(n_443) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_69), .Y(n_514) );
CKINVDCx20_ASAP7_75t_R g138 ( .A(n_70), .Y(n_138) );
AOI21xp5_ASAP7_75t_L g453 ( .A1(n_71), .A2(n_145), .B(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g187 ( .A(n_72), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g481 ( .A1(n_73), .A2(n_213), .B(n_482), .Y(n_481) );
INVx1_ASAP7_75t_L g455 ( .A(n_74), .Y(n_455) );
CKINVDCx16_ASAP7_75t_R g494 ( .A(n_75), .Y(n_494) );
A2O1A1Ixp33_ASAP7_75t_L g188 ( .A1(n_76), .A2(n_118), .B(n_130), .C(n_189), .Y(n_188) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_77), .A2(n_145), .B(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g458 ( .A(n_78), .Y(n_458) );
NAND2xp5_ASAP7_75t_SL g176 ( .A(n_79), .B(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g112 ( .A(n_80), .Y(n_112) );
INVx1_ASAP7_75t_L g434 ( .A(n_81), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g178 ( .A(n_82), .B(n_164), .Y(n_178) );
A2O1A1Ixp33_ASAP7_75t_L g235 ( .A1(n_83), .A2(n_118), .B(n_130), .C(n_236), .Y(n_235) );
INVx2_ASAP7_75t_L g418 ( .A(n_84), .Y(n_418) );
OR2x2_ASAP7_75t_L g689 ( .A(n_84), .B(n_419), .Y(n_689) );
OR2x2_ASAP7_75t_L g707 ( .A(n_84), .B(n_698), .Y(n_707) );
A2O1A1Ixp33_ASAP7_75t_L g508 ( .A1(n_85), .A2(n_130), .B(n_509), .C(n_512), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g157 ( .A(n_86), .B(n_158), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g241 ( .A(n_87), .Y(n_241) );
A2O1A1Ixp33_ASAP7_75t_L g201 ( .A1(n_88), .A2(n_118), .B(n_130), .C(n_202), .Y(n_201) );
CKINVDCx20_ASAP7_75t_R g209 ( .A(n_89), .Y(n_209) );
INVx1_ASAP7_75t_L g162 ( .A(n_90), .Y(n_162) );
CKINVDCx16_ASAP7_75t_R g215 ( .A(n_91), .Y(n_215) );
NAND2xp5_ASAP7_75t_SL g203 ( .A(n_92), .B(n_177), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_93), .B(n_143), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_94), .B(n_143), .Y(n_221) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_95), .A2(n_145), .B(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g466 ( .A(n_96), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_97), .B(n_703), .Y(n_702) );
INVxp67_ASAP7_75t_L g99 ( .A(n_100), .Y(n_99) );
OAI22xp5_ASAP7_75t_SL g101 ( .A1(n_102), .A2(n_415), .B1(n_422), .B2(n_689), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_103), .Y(n_102) );
OAI22xp5_ASAP7_75t_SL g691 ( .A1(n_103), .A2(n_415), .B1(n_692), .B2(n_693), .Y(n_691) );
AND3x1_ASAP7_75t_L g103 ( .A(n_104), .B(n_340), .C(n_389), .Y(n_103) );
NOR3xp33_ASAP7_75t_SL g104 ( .A(n_105), .B(n_247), .C(n_285), .Y(n_104) );
OAI222xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_168), .B1(n_222), .B2(n_228), .C1(n_242), .C2(n_245), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_139), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_107), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_107), .B(n_290), .Y(n_381) );
BUFx2_ASAP7_75t_L g107 ( .A(n_108), .Y(n_107) );
OR2x2_ASAP7_75t_L g258 ( .A(n_108), .B(n_159), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_108), .B(n_140), .Y(n_266) );
AND2x2_ASAP7_75t_L g301 ( .A(n_108), .B(n_278), .Y(n_301) );
OR2x2_ASAP7_75t_L g325 ( .A(n_108), .B(n_140), .Y(n_325) );
OR2x2_ASAP7_75t_L g333 ( .A(n_108), .B(n_232), .Y(n_333) );
AND2x2_ASAP7_75t_L g336 ( .A(n_108), .B(n_159), .Y(n_336) );
INVx3_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
OR2x2_ASAP7_75t_L g230 ( .A(n_109), .B(n_231), .Y(n_230) );
AND2x2_ASAP7_75t_L g244 ( .A(n_109), .B(n_159), .Y(n_244) );
AND2x2_ASAP7_75t_L g294 ( .A(n_109), .B(n_232), .Y(n_294) );
AND2x2_ASAP7_75t_L g307 ( .A(n_109), .B(n_140), .Y(n_307) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_109), .B(n_393), .Y(n_414) );
AO21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_116), .B(n_137), .Y(n_109) );
NOR2xp33_ASAP7_75t_L g137 ( .A(n_110), .B(n_138), .Y(n_137) );
INVx2_ASAP7_75t_L g182 ( .A(n_110), .Y(n_182) );
AO21x2_ASAP7_75t_L g232 ( .A1(n_110), .A2(n_233), .B(n_240), .Y(n_232) );
INVx1_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_111), .Y(n_143) );
AND2x2_ASAP7_75t_L g111 ( .A(n_112), .B(n_113), .Y(n_111) );
AND2x2_ASAP7_75t_SL g158 ( .A(n_112), .B(n_113), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g113 ( .A(n_114), .B(n_115), .Y(n_113) );
OAI22xp33_ASAP7_75t_L g116 ( .A1(n_117), .A2(n_120), .B1(n_133), .B2(n_134), .Y(n_116) );
O2A1O1Ixp33_ASAP7_75t_L g146 ( .A1(n_117), .A2(n_147), .B(n_148), .C(n_149), .Y(n_146) );
O2A1O1Ixp33_ASAP7_75t_L g161 ( .A1(n_117), .A2(n_148), .B(n_162), .C(n_163), .Y(n_161) );
O2A1O1Ixp33_ASAP7_75t_L g214 ( .A1(n_117), .A2(n_148), .B(n_215), .C(n_216), .Y(n_214) );
O2A1O1Ixp33_ASAP7_75t_SL g444 ( .A1(n_117), .A2(n_148), .B(n_445), .C(n_446), .Y(n_444) );
O2A1O1Ixp33_ASAP7_75t_SL g454 ( .A1(n_117), .A2(n_148), .B(n_455), .C(n_456), .Y(n_454) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_117), .A2(n_148), .B(n_463), .C(n_464), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_L g472 ( .A1(n_117), .A2(n_148), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g482 ( .A1(n_117), .A2(n_148), .B(n_483), .C(n_484), .Y(n_482) );
INVx1_ASAP7_75t_L g512 ( .A(n_117), .Y(n_512) );
INVx4_ASAP7_75t_SL g117 ( .A(n_118), .Y(n_117) );
NAND2x1p5_ASAP7_75t_L g134 ( .A(n_118), .B(n_135), .Y(n_134) );
AND2x4_ASAP7_75t_L g145 ( .A(n_118), .B(n_135), .Y(n_145) );
BUFx3_ASAP7_75t_L g500 ( .A(n_118), .Y(n_500) );
INVx2_ASAP7_75t_L g239 ( .A(n_121), .Y(n_239) );
INVx3_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
INVx2_ASAP7_75t_L g131 ( .A(n_123), .Y(n_131) );
INVx1_ASAP7_75t_L g136 ( .A(n_123), .Y(n_136) );
OAI22xp5_ASAP7_75t_SL g124 ( .A1(n_125), .A2(n_127), .B1(n_128), .B2(n_129), .Y(n_124) );
INVx2_ASAP7_75t_L g128 ( .A(n_125), .Y(n_128) );
INVx4_ASAP7_75t_L g217 ( .A(n_125), .Y(n_217) );
BUFx6f_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
INVx1_ASAP7_75t_L g132 ( .A(n_126), .Y(n_132) );
AND2x2_ASAP7_75t_L g135 ( .A(n_126), .B(n_136), .Y(n_135) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_126), .Y(n_151) );
INVx3_ASAP7_75t_L g154 ( .A(n_126), .Y(n_154) );
INVx1_ASAP7_75t_L g164 ( .A(n_126), .Y(n_164) );
INVx2_ASAP7_75t_L g435 ( .A(n_128), .Y(n_435) );
INVx5_ASAP7_75t_L g148 ( .A(n_130), .Y(n_148) );
AND2x6_ASAP7_75t_L g130 ( .A(n_131), .B(n_132), .Y(n_130) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_131), .Y(n_156) );
BUFx3_ASAP7_75t_L g181 ( .A(n_131), .Y(n_181) );
OAI21xp5_ASAP7_75t_L g186 ( .A1(n_134), .A2(n_187), .B(n_188), .Y(n_186) );
OAI21xp5_ASAP7_75t_L g233 ( .A1(n_134), .A2(n_234), .B(n_235), .Y(n_233) );
OAI21xp5_ASAP7_75t_L g430 ( .A1(n_134), .A2(n_431), .B(n_432), .Y(n_430) );
O2A1O1Ixp33_ASAP7_75t_L g493 ( .A1(n_134), .A2(n_158), .B(n_494), .C(n_495), .Y(n_493) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_134), .A2(n_507), .B(n_508), .Y(n_506) );
INVx1_ASAP7_75t_L g488 ( .A(n_136), .Y(n_488) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_139), .A2(n_333), .B(n_334), .C(n_337), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g361 ( .A(n_139), .B(n_362), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_139), .B(n_277), .Y(n_399) );
AND2x2_ASAP7_75t_L g139 ( .A(n_140), .B(n_159), .Y(n_139) );
AND2x2_ASAP7_75t_SL g243 ( .A(n_140), .B(n_244), .Y(n_243) );
INVx2_ASAP7_75t_L g257 ( .A(n_140), .Y(n_257) );
AND2x2_ASAP7_75t_L g284 ( .A(n_140), .B(n_278), .Y(n_284) );
INVx1_ASAP7_75t_SL g292 ( .A(n_140), .Y(n_292) );
AND2x2_ASAP7_75t_L g315 ( .A(n_140), .B(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g393 ( .A(n_140), .Y(n_393) );
OA21x2_ASAP7_75t_L g140 ( .A1(n_141), .A2(n_144), .B(n_157), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_142), .Y(n_141) );
NOR2xp33_ASAP7_75t_SL g183 ( .A(n_142), .B(n_184), .Y(n_183) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_142), .B(n_438), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g501 ( .A(n_142), .B(n_502), .Y(n_501) );
AO21x2_ASAP7_75t_L g505 ( .A1(n_142), .A2(n_506), .B(n_513), .Y(n_505) );
INVx4_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
OA21x2_ASAP7_75t_L g159 ( .A1(n_143), .A2(n_160), .B(n_167), .Y(n_159) );
HB1xp67_ASAP7_75t_L g452 ( .A(n_143), .Y(n_452) );
BUFx2_ASAP7_75t_L g213 ( .A(n_145), .Y(n_213) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx4_ASAP7_75t_L g205 ( .A(n_151), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_153), .B(n_154), .Y(n_152) );
NOR2xp33_ASAP7_75t_L g165 ( .A(n_154), .B(n_166), .Y(n_165) );
INVx5_ASAP7_75t_L g177 ( .A(n_154), .Y(n_177) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_154), .B(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
HB1xp67_ASAP7_75t_L g206 ( .A(n_156), .Y(n_206) );
INVx1_ASAP7_75t_L g195 ( .A(n_158), .Y(n_195) );
INVx2_ASAP7_75t_L g199 ( .A(n_158), .Y(n_199) );
OA21x2_ASAP7_75t_L g211 ( .A1(n_158), .A2(n_212), .B(n_221), .Y(n_211) );
OA21x2_ASAP7_75t_L g442 ( .A1(n_158), .A2(n_443), .B(n_449), .Y(n_442) );
BUFx2_ASAP7_75t_L g229 ( .A(n_159), .Y(n_229) );
INVx1_ASAP7_75t_L g291 ( .A(n_159), .Y(n_291) );
INVx3_ASAP7_75t_L g316 ( .A(n_159), .Y(n_316) );
NAND2xp5_ASAP7_75t_SL g249 ( .A(n_168), .B(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g168 ( .A(n_169), .B(n_196), .Y(n_168) );
INVx1_ASAP7_75t_L g312 ( .A(n_169), .Y(n_312) );
OAI32xp33_ASAP7_75t_L g318 ( .A1(n_169), .A2(n_257), .A3(n_319), .B1(n_320), .B2(n_321), .Y(n_318) );
OAI22xp5_ASAP7_75t_L g322 ( .A1(n_169), .A2(n_323), .B1(n_326), .B2(n_331), .Y(n_322) );
INVx4_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
AND2x2_ASAP7_75t_L g260 ( .A(n_170), .B(n_261), .Y(n_260) );
AND2x2_ASAP7_75t_L g338 ( .A(n_170), .B(n_339), .Y(n_338) );
AND2x2_ASAP7_75t_L g408 ( .A(n_170), .B(n_354), .Y(n_408) );
AND2x2_ASAP7_75t_L g170 ( .A(n_171), .B(n_185), .Y(n_170) );
AND2x2_ASAP7_75t_L g223 ( .A(n_171), .B(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g253 ( .A(n_171), .Y(n_253) );
INVx1_ASAP7_75t_L g272 ( .A(n_171), .Y(n_272) );
OR2x2_ASAP7_75t_L g280 ( .A(n_171), .B(n_281), .Y(n_280) );
AND2x2_ASAP7_75t_L g287 ( .A(n_171), .B(n_261), .Y(n_287) );
NOR2xp33_ASAP7_75t_L g295 ( .A(n_171), .B(n_296), .Y(n_295) );
AND2x2_ASAP7_75t_L g308 ( .A(n_171), .B(n_226), .Y(n_308) );
INVx3_ASAP7_75t_L g330 ( .A(n_171), .Y(n_330) );
AND2x2_ASAP7_75t_L g355 ( .A(n_171), .B(n_227), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_171), .B(n_320), .Y(n_403) );
OR2x6_ASAP7_75t_L g171 ( .A(n_172), .B(n_183), .Y(n_171) );
AOI21xp5_ASAP7_75t_SL g172 ( .A1(n_173), .A2(n_174), .B(n_182), .Y(n_172) );
AOI21xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_178), .B(n_179), .Y(n_175) );
O2A1O1Ixp33_ASAP7_75t_L g236 ( .A1(n_177), .A2(n_237), .B(n_238), .C(n_239), .Y(n_236) );
OAI22xp33_ASAP7_75t_L g485 ( .A1(n_177), .A2(n_217), .B1(n_486), .B2(n_487), .Y(n_485) );
O2A1O1Ixp33_ASAP7_75t_L g496 ( .A1(n_177), .A2(n_497), .B(n_498), .C(n_499), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g189 ( .A1(n_179), .A2(n_190), .B(n_191), .Y(n_189) );
O2A1O1Ixp5_ASAP7_75t_L g433 ( .A1(n_179), .A2(n_434), .B(n_435), .C(n_436), .Y(n_433) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_179), .A2(n_435), .B(n_510), .C(n_511), .Y(n_509) );
INVx2_ASAP7_75t_L g179 ( .A(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
INVx1_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
INVx1_ASAP7_75t_L g192 ( .A(n_182), .Y(n_192) );
INVx2_ASAP7_75t_L g227 ( .A(n_185), .Y(n_227) );
AND2x2_ASAP7_75t_L g359 ( .A(n_185), .B(n_197), .Y(n_359) );
AO21x2_ASAP7_75t_L g185 ( .A1(n_186), .A2(n_192), .B(n_193), .Y(n_185) );
INVx1_ASAP7_75t_L g480 ( .A(n_192), .Y(n_480) );
AO21x2_ASAP7_75t_L g532 ( .A1(n_192), .A2(n_533), .B(n_534), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_195), .B(n_209), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_195), .B(n_241), .Y(n_240) );
AO21x2_ASAP7_75t_L g429 ( .A1(n_195), .A2(n_430), .B(n_437), .Y(n_429) );
INVx2_ASAP7_75t_L g401 ( .A(n_196), .Y(n_401) );
OR2x2_ASAP7_75t_L g196 ( .A(n_197), .B(n_210), .Y(n_196) );
INVx1_ASAP7_75t_L g246 ( .A(n_197), .Y(n_246) );
AND2x2_ASAP7_75t_L g273 ( .A(n_197), .B(n_274), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_197), .B(n_227), .Y(n_281) );
AND2x2_ASAP7_75t_L g339 ( .A(n_197), .B(n_262), .Y(n_339) );
INVx2_ASAP7_75t_L g197 ( .A(n_198), .Y(n_197) );
INVx1_ASAP7_75t_L g225 ( .A(n_198), .Y(n_225) );
AND2x2_ASAP7_75t_L g252 ( .A(n_198), .B(n_253), .Y(n_252) );
AND2x2_ASAP7_75t_L g261 ( .A(n_198), .B(n_262), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_198), .B(n_227), .Y(n_327) );
AO21x2_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_208), .Y(n_198) );
INVx1_ASAP7_75t_L g490 ( .A(n_199), .Y(n_490) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_199), .B(n_514), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_201), .B(n_207), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_206), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_205), .B(n_476), .Y(n_475) );
NAND2xp5_ASAP7_75t_L g254 ( .A(n_210), .B(n_255), .Y(n_254) );
INVx2_ASAP7_75t_L g274 ( .A(n_210), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g320 ( .A(n_210), .B(n_227), .Y(n_320) );
AND2x2_ASAP7_75t_L g329 ( .A(n_210), .B(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g354 ( .A(n_210), .Y(n_354) );
INVx2_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
AND2x2_ASAP7_75t_L g226 ( .A(n_211), .B(n_227), .Y(n_226) );
INVx1_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_217), .B(n_219), .Y(n_218) );
NOR2xp33_ASAP7_75t_L g457 ( .A(n_217), .B(n_458), .Y(n_457) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_217), .B(n_466), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g390 ( .A1(n_222), .A2(n_232), .B1(n_391), .B2(n_394), .Y(n_390) );
INVx1_ASAP7_75t_SL g222 ( .A(n_223), .Y(n_222) );
OAI21xp5_ASAP7_75t_SL g413 ( .A1(n_224), .A2(n_335), .B(n_414), .Y(n_413) );
AND2x2_ASAP7_75t_L g224 ( .A(n_225), .B(n_226), .Y(n_224) );
NOR2xp33_ASAP7_75t_L g347 ( .A(n_225), .B(n_330), .Y(n_347) );
INVx1_ASAP7_75t_L g372 ( .A(n_225), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_226), .B(n_246), .Y(n_245) );
AND2x2_ASAP7_75t_L g299 ( .A(n_226), .B(n_252), .Y(n_299) );
INVx2_ASAP7_75t_L g255 ( .A(n_227), .Y(n_255) );
INVx1_ASAP7_75t_L g305 ( .A(n_227), .Y(n_305) );
OAI221xp5_ASAP7_75t_L g396 ( .A1(n_228), .A2(n_380), .B1(n_397), .B2(n_400), .C(n_402), .Y(n_396) );
OR2x2_ASAP7_75t_L g228 ( .A(n_229), .B(n_230), .Y(n_228) );
INVx1_ASAP7_75t_L g267 ( .A(n_229), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_229), .B(n_278), .Y(n_319) );
NOR2xp33_ASAP7_75t_L g288 ( .A(n_230), .B(n_289), .Y(n_288) );
OR2x2_ASAP7_75t_L g321 ( .A(n_230), .B(n_267), .Y(n_321) );
INVx3_ASAP7_75t_SL g362 ( .A(n_230), .Y(n_362) );
AND2x2_ASAP7_75t_L g306 ( .A(n_231), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g335 ( .A(n_231), .B(n_336), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g350 ( .A(n_231), .B(n_244), .Y(n_350) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_231), .B(n_290), .Y(n_376) );
INVx3_ASAP7_75t_L g231 ( .A(n_232), .Y(n_231) );
INVx3_ASAP7_75t_L g278 ( .A(n_232), .Y(n_278) );
OAI322xp33_ASAP7_75t_L g373 ( .A1(n_232), .A2(n_304), .A3(n_326), .B1(n_374), .B2(n_376), .C1(n_377), .C2(n_378), .Y(n_373) );
INVx1_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
AOI21xp33_ASAP7_75t_L g397 ( .A1(n_243), .A2(n_246), .B(n_398), .Y(n_397) );
NOR2xp33_ASAP7_75t_SL g323 ( .A(n_244), .B(n_324), .Y(n_323) );
AND2x2_ASAP7_75t_L g345 ( .A(n_244), .B(n_257), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_244), .B(n_284), .Y(n_360) );
INVxp67_ASAP7_75t_L g311 ( .A(n_246), .Y(n_311) );
AOI211xp5_ASAP7_75t_L g317 ( .A1(n_246), .A2(n_318), .B(n_322), .C(n_332), .Y(n_317) );
OAI221xp5_ASAP7_75t_SL g247 ( .A1(n_248), .A2(n_256), .B1(n_259), .B2(n_263), .C(n_268), .Y(n_247) );
INVxp67_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_254), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g271 ( .A(n_255), .B(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g388 ( .A(n_255), .Y(n_388) );
OAI221xp5_ASAP7_75t_L g404 ( .A1(n_256), .A2(n_405), .B1(n_410), .B2(n_411), .C(n_413), .Y(n_404) );
OR2x2_ASAP7_75t_L g256 ( .A(n_257), .B(n_258), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_257), .B(n_301), .Y(n_300) );
INVx1_ASAP7_75t_SL g304 ( .A(n_257), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_257), .B(n_335), .Y(n_342) );
AND2x2_ASAP7_75t_L g384 ( .A(n_257), .B(n_362), .Y(n_384) );
NOR2xp33_ASAP7_75t_L g282 ( .A(n_258), .B(n_283), .Y(n_282) );
OAI22xp33_ASAP7_75t_L g379 ( .A1(n_258), .A2(n_270), .B1(n_380), .B2(n_381), .Y(n_379) );
OR2x2_ASAP7_75t_L g410 ( .A(n_258), .B(n_278), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g259 ( .A(n_260), .Y(n_259) );
INVx1_ASAP7_75t_L g387 ( .A(n_261), .Y(n_387) );
AND2x2_ASAP7_75t_L g412 ( .A(n_261), .B(n_355), .Y(n_412) );
INVxp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NOR2xp33_ASAP7_75t_SL g264 ( .A(n_265), .B(n_267), .Y(n_264) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
OR2x2_ASAP7_75t_L g276 ( .A(n_266), .B(n_277), .Y(n_276) );
AOI22xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_275), .B1(n_279), .B2(n_282), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_271), .B(n_273), .Y(n_270) );
INVx1_ASAP7_75t_L g343 ( .A(n_271), .Y(n_343) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_271), .B(n_311), .Y(n_378) );
AOI322xp5_ASAP7_75t_L g302 ( .A1(n_273), .A2(n_303), .A3(n_305), .B1(n_306), .B2(n_308), .C1(n_309), .C2(n_313), .Y(n_302) );
INVxp67_ASAP7_75t_L g296 ( .A(n_274), .Y(n_296) );
INVx1_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
OAI22xp5_ASAP7_75t_L g297 ( .A1(n_276), .A2(n_281), .B1(n_298), .B2(n_300), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g377 ( .A(n_277), .B(n_290), .Y(n_377) );
INVx1_ASAP7_75t_SL g277 ( .A(n_278), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g386 ( .A(n_278), .B(n_316), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g392 ( .A(n_278), .B(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
OR2x2_ASAP7_75t_L g374 ( .A(n_280), .B(n_375), .Y(n_374) );
INVx1_ASAP7_75t_SL g283 ( .A(n_284), .Y(n_283) );
NAND3xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_302), .C(n_317), .Y(n_285) );
AOI221xp5_ASAP7_75t_L g286 ( .A1(n_287), .A2(n_288), .B1(n_293), .B2(n_295), .C(n_297), .Y(n_286) );
AND2x2_ASAP7_75t_L g293 ( .A(n_289), .B(n_294), .Y(n_293) );
INVx3_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
AND2x4_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
AND2x2_ASAP7_75t_L g303 ( .A(n_294), .B(n_304), .Y(n_303) );
HB1xp67_ASAP7_75t_L g375 ( .A(n_296), .Y(n_375) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_301), .B(n_315), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g368 ( .A(n_304), .B(n_362), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_305), .B(n_365), .Y(n_364) );
INVx1_ASAP7_75t_SL g380 ( .A(n_308), .Y(n_380) );
AND2x2_ASAP7_75t_L g395 ( .A(n_308), .B(n_372), .Y(n_395) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_311), .B(n_312), .Y(n_310) );
INVx1_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
AOI211xp5_ASAP7_75t_L g389 ( .A1(n_319), .A2(n_390), .B(n_396), .C(n_404), .Y(n_389) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
OR2x2_ASAP7_75t_L g326 ( .A(n_327), .B(n_328), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g358 ( .A(n_329), .B(n_359), .Y(n_358) );
NAND2x1_ASAP7_75t_SL g400 ( .A(n_330), .B(n_401), .Y(n_400) );
CKINVDCx16_ASAP7_75t_R g370 ( .A(n_333), .Y(n_370) );
INVx1_ASAP7_75t_SL g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g365 ( .A(n_339), .Y(n_365) );
AND2x2_ASAP7_75t_L g369 ( .A(n_339), .B(n_355), .Y(n_369) );
NOR5xp2_ASAP7_75t_L g340 ( .A(n_341), .B(n_356), .C(n_373), .D(n_379), .E(n_382), .Y(n_340) );
OAI221xp5_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B1(n_344), .B2(n_346), .C(n_348), .Y(n_341) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_345), .B(n_403), .Y(n_402) );
INVxp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_349), .B(n_351), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_353), .B(n_355), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_354), .Y(n_353) );
AND2x2_ASAP7_75t_L g371 ( .A(n_355), .B(n_372), .Y(n_371) );
OAI221xp5_ASAP7_75t_SL g356 ( .A1(n_357), .A2(n_360), .B1(n_361), .B2(n_363), .C(n_366), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_367), .A2(n_369), .B1(n_370), .B2(n_371), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx1_ASAP7_75t_L g409 ( .A(n_369), .Y(n_409) );
AOI211xp5_ASAP7_75t_SL g382 ( .A1(n_383), .A2(n_385), .B(n_387), .C(n_388), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVxp67_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_409), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
CKINVDCx14_ASAP7_75t_R g411 ( .A(n_412), .Y(n_411) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
NOR2x2_ASAP7_75t_L g697 ( .A(n_418), .B(n_698), .Y(n_697) );
INVx2_ASAP7_75t_L g698 ( .A(n_419), .Y(n_698) );
AND2x2_ASAP7_75t_L g419 ( .A(n_420), .B(n_421), .Y(n_419) );
INVx2_ASAP7_75t_L g692 ( .A(n_422), .Y(n_692) );
OR2x2_ASAP7_75t_SL g422 ( .A(n_423), .B(n_644), .Y(n_422) );
NAND5xp2_ASAP7_75t_L g423 ( .A(n_424), .B(n_556), .C(n_594), .D(n_615), .E(n_632), .Y(n_423) );
NOR3xp33_ASAP7_75t_L g424 ( .A(n_425), .B(n_528), .C(n_549), .Y(n_424) );
OAI221xp5_ASAP7_75t_SL g425 ( .A1(n_426), .A2(n_468), .B1(n_491), .B2(n_515), .C(n_519), .Y(n_425) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_427), .B(n_439), .Y(n_426) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_428), .B(n_517), .Y(n_536) );
OR2x2_ASAP7_75t_L g563 ( .A(n_428), .B(n_451), .Y(n_563) );
AND2x2_ASAP7_75t_L g577 ( .A(n_428), .B(n_451), .Y(n_577) );
NOR2xp33_ASAP7_75t_L g591 ( .A(n_428), .B(n_442), .Y(n_591) );
AND2x2_ASAP7_75t_L g629 ( .A(n_428), .B(n_593), .Y(n_629) );
AND2x2_ASAP7_75t_L g658 ( .A(n_428), .B(n_568), .Y(n_658) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_428), .B(n_540), .Y(n_675) );
INVx4_ASAP7_75t_L g428 ( .A(n_429), .Y(n_428) );
AND2x2_ASAP7_75t_L g555 ( .A(n_429), .B(n_450), .Y(n_555) );
BUFx3_ASAP7_75t_L g580 ( .A(n_429), .Y(n_580) );
AND2x2_ASAP7_75t_L g609 ( .A(n_429), .B(n_451), .Y(n_609) );
AND3x2_ASAP7_75t_L g622 ( .A(n_429), .B(n_623), .C(n_624), .Y(n_622) );
INVx1_ASAP7_75t_L g545 ( .A(n_439), .Y(n_545) );
AND2x2_ASAP7_75t_L g439 ( .A(n_440), .B(n_450), .Y(n_439) );
AOI32xp33_ASAP7_75t_L g600 ( .A1(n_440), .A2(n_552), .A3(n_601), .B1(n_604), .B2(n_605), .Y(n_600) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
AND2x2_ASAP7_75t_L g527 ( .A(n_441), .B(n_450), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g598 ( .A(n_441), .B(n_555), .Y(n_598) );
AND2x2_ASAP7_75t_L g605 ( .A(n_441), .B(n_577), .Y(n_605) );
OR2x2_ASAP7_75t_L g611 ( .A(n_441), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g636 ( .A(n_441), .B(n_566), .Y(n_636) );
OR2x2_ASAP7_75t_L g654 ( .A(n_441), .B(n_479), .Y(n_654) );
BUFx3_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
AND2x2_ASAP7_75t_L g518 ( .A(n_442), .B(n_460), .Y(n_518) );
INVx2_ASAP7_75t_L g540 ( .A(n_442), .Y(n_540) );
OR2x2_ASAP7_75t_L g562 ( .A(n_442), .B(n_460), .Y(n_562) );
AND2x2_ASAP7_75t_L g567 ( .A(n_442), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_442), .B(n_619), .Y(n_618) );
AND2x2_ASAP7_75t_L g623 ( .A(n_442), .B(n_517), .Y(n_623) );
INVx1_ASAP7_75t_SL g674 ( .A(n_450), .Y(n_674) );
AND2x2_ASAP7_75t_L g450 ( .A(n_451), .B(n_460), .Y(n_450) );
INVx1_ASAP7_75t_SL g517 ( .A(n_451), .Y(n_517) );
HB1xp67_ASAP7_75t_L g566 ( .A(n_451), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_451), .B(n_603), .Y(n_602) );
NAND3xp33_ASAP7_75t_L g669 ( .A(n_451), .B(n_540), .C(n_658), .Y(n_669) );
OA21x2_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_453), .B(n_459), .Y(n_451) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_452), .A2(n_461), .B(n_467), .Y(n_460) );
OA21x2_ASAP7_75t_L g470 ( .A1(n_452), .A2(n_471), .B(n_477), .Y(n_470) );
INVx2_ASAP7_75t_L g568 ( .A(n_460), .Y(n_568) );
HB1xp67_ASAP7_75t_L g582 ( .A(n_460), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_469), .B(n_478), .Y(n_468) );
INVx1_ASAP7_75t_L g604 ( .A(n_469), .Y(n_604) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
AND2x2_ASAP7_75t_L g522 ( .A(n_470), .B(n_504), .Y(n_522) );
INVx2_ASAP7_75t_L g539 ( .A(n_470), .Y(n_539) );
AND2x2_ASAP7_75t_L g544 ( .A(n_470), .B(n_505), .Y(n_544) );
AND2x2_ASAP7_75t_L g559 ( .A(n_470), .B(n_492), .Y(n_559) );
AND2x2_ASAP7_75t_L g571 ( .A(n_470), .B(n_543), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_478), .B(n_587), .Y(n_586) );
NAND2x1p5_ASAP7_75t_L g643 ( .A(n_478), .B(n_544), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_478), .B(n_663), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_478), .B(n_538), .Y(n_666) );
BUFx3_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
OR2x2_ASAP7_75t_L g503 ( .A(n_479), .B(n_504), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_479), .B(n_522), .Y(n_521) );
AND2x2_ASAP7_75t_L g548 ( .A(n_479), .B(n_492), .Y(n_548) );
AND2x2_ASAP7_75t_L g574 ( .A(n_479), .B(n_504), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_479), .B(n_614), .Y(n_613) );
OA21x2_ASAP7_75t_L g479 ( .A1(n_480), .A2(n_481), .B(n_489), .Y(n_479) );
INVx1_ASAP7_75t_L g533 ( .A(n_481), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_485), .B(n_488), .Y(n_484) );
INVx2_ASAP7_75t_L g499 ( .A(n_488), .Y(n_499) );
INVx1_ASAP7_75t_L g534 ( .A(n_489), .Y(n_534) );
OR2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_503), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_492), .B(n_525), .Y(n_524) );
AND2x4_ASAP7_75t_L g538 ( .A(n_492), .B(n_539), .Y(n_538) );
INVx3_ASAP7_75t_SL g543 ( .A(n_492), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_492), .B(n_530), .Y(n_596) );
OR2x2_ASAP7_75t_L g606 ( .A(n_492), .B(n_532), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_492), .B(n_574), .Y(n_634) );
OR2x2_ASAP7_75t_L g664 ( .A(n_492), .B(n_504), .Y(n_664) );
AND2x2_ASAP7_75t_L g668 ( .A(n_492), .B(n_505), .Y(n_668) );
NAND2xp5_ASAP7_75t_SL g681 ( .A(n_492), .B(n_544), .Y(n_681) );
AND2x2_ASAP7_75t_L g688 ( .A(n_492), .B(n_570), .Y(n_688) );
OR2x6_ASAP7_75t_L g492 ( .A(n_493), .B(n_501), .Y(n_492) );
INVx1_ASAP7_75t_SL g631 ( .A(n_503), .Y(n_631) );
AND2x2_ASAP7_75t_L g570 ( .A(n_504), .B(n_532), .Y(n_570) );
AND2x2_ASAP7_75t_L g584 ( .A(n_504), .B(n_539), .Y(n_584) );
AND2x2_ASAP7_75t_L g587 ( .A(n_504), .B(n_543), .Y(n_587) );
INVx1_ASAP7_75t_L g614 ( .A(n_504), .Y(n_614) );
INVx2_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
BUFx2_ASAP7_75t_L g526 ( .A(n_505), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_516), .B(n_518), .Y(n_515) );
A2O1A1Ixp33_ASAP7_75t_L g685 ( .A1(n_516), .A2(n_562), .B(n_686), .C(n_687), .Y(n_685) );
HB1xp67_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
AND2x2_ASAP7_75t_L g592 ( .A(n_517), .B(n_593), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_518), .B(n_535), .Y(n_550) );
AND2x2_ASAP7_75t_L g576 ( .A(n_518), .B(n_577), .Y(n_576) );
OAI21xp5_ASAP7_75t_SL g519 ( .A1(n_520), .A2(n_523), .B(n_527), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_521), .B(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g547 ( .A(n_522), .B(n_548), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_522), .B(n_543), .Y(n_588) );
AND2x2_ASAP7_75t_L g679 ( .A(n_522), .B(n_530), .Y(n_679) );
INVxp67_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx1_ASAP7_75t_L g525 ( .A(n_526), .Y(n_525) );
AND2x2_ASAP7_75t_L g552 ( .A(n_526), .B(n_539), .Y(n_552) );
OR2x2_ASAP7_75t_L g553 ( .A(n_526), .B(n_537), .Y(n_553) );
OAI322xp33_ASAP7_75t_L g528 ( .A1(n_529), .A2(n_536), .A3(n_537), .B1(n_540), .B2(n_541), .C1(n_545), .C2(n_546), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_530), .B(n_535), .Y(n_529) );
AND2x2_ASAP7_75t_L g640 ( .A(n_530), .B(n_552), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g686 ( .A(n_530), .B(n_604), .Y(n_686) );
INVx2_ASAP7_75t_L g530 ( .A(n_531), .Y(n_530) );
INVx1_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g583 ( .A(n_532), .B(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g535 ( .A(n_536), .Y(n_535) );
OR2x2_ASAP7_75t_L g649 ( .A(n_536), .B(n_562), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_537), .B(n_631), .Y(n_630) );
INVx3_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_538), .B(n_570), .Y(n_627) );
AND2x2_ASAP7_75t_L g573 ( .A(n_539), .B(n_543), .Y(n_573) );
AND2x2_ASAP7_75t_L g581 ( .A(n_540), .B(n_582), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g678 ( .A1(n_540), .A2(n_619), .B(n_679), .C(n_680), .Y(n_678) );
AOI21xp33_ASAP7_75t_L g651 ( .A1(n_541), .A2(n_554), .B(n_652), .Y(n_651) );
INVx1_ASAP7_75t_SL g541 ( .A(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_543), .B(n_570), .Y(n_610) );
AND2x2_ASAP7_75t_L g616 ( .A(n_543), .B(n_584), .Y(n_616) );
AND2x2_ASAP7_75t_L g650 ( .A(n_543), .B(n_552), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g558 ( .A(n_544), .B(n_559), .Y(n_558) );
INVx2_ASAP7_75t_SL g660 ( .A(n_544), .Y(n_660) );
INVx1_ASAP7_75t_L g546 ( .A(n_547), .Y(n_546) );
AOI22xp5_ASAP7_75t_L g575 ( .A1(n_548), .A2(n_576), .B1(n_578), .B2(n_583), .Y(n_575) );
OAI22xp5_ASAP7_75t_SL g549 ( .A1(n_550), .A2(n_551), .B1(n_553), .B2(n_554), .Y(n_549) );
OAI22xp33_ASAP7_75t_L g585 ( .A1(n_550), .A2(n_586), .B1(n_588), .B2(n_589), .Y(n_585) );
INVxp67_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
INVx1_ASAP7_75t_SL g554 ( .A(n_555), .Y(n_554) );
AOI221xp5_ASAP7_75t_L g656 ( .A1(n_555), .A2(n_657), .B1(n_659), .B2(n_661), .C(n_665), .Y(n_656) );
AOI211xp5_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_560), .B(n_564), .C(n_585), .Y(n_556) );
INVxp67_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_562), .B(n_563), .Y(n_561) );
OR2x2_ASAP7_75t_L g626 ( .A(n_562), .B(n_579), .Y(n_626) );
INVx1_ASAP7_75t_L g677 ( .A(n_562), .Y(n_677) );
OAI221xp5_ASAP7_75t_L g564 ( .A1(n_563), .A2(n_565), .B1(n_569), .B2(n_572), .C(n_575), .Y(n_564) );
INVx2_ASAP7_75t_SL g619 ( .A(n_563), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
INVx1_ASAP7_75t_L g684 ( .A(n_566), .Y(n_684) );
AND2x2_ASAP7_75t_L g608 ( .A(n_567), .B(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g593 ( .A(n_568), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_570), .B(n_571), .Y(n_569) );
INVx1_ASAP7_75t_L g655 ( .A(n_571), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
AND2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .Y(n_578) );
NOR2xp33_ASAP7_75t_L g680 ( .A(n_579), .B(n_681), .Y(n_680) );
CKINVDCx16_ASAP7_75t_R g579 ( .A(n_580), .Y(n_579) );
INVxp67_ASAP7_75t_L g624 ( .A(n_582), .Y(n_624) );
O2A1O1Ixp33_ASAP7_75t_L g594 ( .A1(n_583), .A2(n_595), .B(n_597), .C(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g672 ( .A(n_586), .Y(n_672) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_590), .B(n_648), .Y(n_647) );
AND2x2_ASAP7_75t_L g590 ( .A(n_591), .B(n_592), .Y(n_590) );
INVx2_ASAP7_75t_L g603 ( .A(n_593), .Y(n_603) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx1_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
OAI222xp33_ASAP7_75t_L g599 ( .A1(n_600), .A2(n_606), .B1(n_607), .B2(n_610), .C1(n_611), .C2(n_613), .Y(n_599) );
INVx1_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
INVx1_ASAP7_75t_SL g639 ( .A(n_603), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g659 ( .A(n_606), .B(n_660), .Y(n_659) );
NAND2xp33_ASAP7_75t_SL g637 ( .A(n_607), .B(n_638), .Y(n_637) );
INVx1_ASAP7_75t_SL g607 ( .A(n_608), .Y(n_607) );
INVx1_ASAP7_75t_SL g612 ( .A(n_609), .Y(n_612) );
AND2x2_ASAP7_75t_L g676 ( .A(n_609), .B(n_677), .Y(n_676) );
OR2x2_ASAP7_75t_L g642 ( .A(n_612), .B(n_639), .Y(n_642) );
INVx1_ASAP7_75t_L g671 ( .A(n_613), .Y(n_671) );
AOI211xp5_ASAP7_75t_L g615 ( .A1(n_616), .A2(n_617), .B(n_620), .C(n_625), .Y(n_615) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_619), .B(n_639), .Y(n_638) );
INVx2_ASAP7_75t_SL g621 ( .A(n_622), .Y(n_621) );
AOI322xp5_ASAP7_75t_L g670 ( .A1(n_622), .A2(n_650), .A3(n_655), .B1(n_671), .B2(n_672), .C1(n_673), .C2(n_676), .Y(n_670) );
AND2x2_ASAP7_75t_L g657 ( .A(n_623), .B(n_658), .Y(n_657) );
OAI22xp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B1(n_628), .B2(n_630), .Y(n_625) );
INVxp33_ASAP7_75t_L g628 ( .A(n_629), .Y(n_628) );
AOI221xp5_ASAP7_75t_L g632 ( .A1(n_633), .A2(n_635), .B1(n_637), .B2(n_640), .C(n_641), .Y(n_632) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g641 ( .A(n_642), .B(n_643), .Y(n_641) );
NAND5xp2_ASAP7_75t_L g644 ( .A(n_645), .B(n_656), .C(n_670), .D(n_678), .E(n_682), .Y(n_644) );
AOI21xp5_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B(n_651), .Y(n_645) );
INVxp67_ASAP7_75t_L g646 ( .A(n_647), .Y(n_646) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVxp33_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_655), .Y(n_653) );
A2O1A1Ixp33_ASAP7_75t_L g682 ( .A1(n_658), .A2(n_683), .B(n_684), .C(n_685), .Y(n_682) );
AOI31xp33_ASAP7_75t_L g665 ( .A1(n_660), .A2(n_666), .A3(n_667), .B(n_669), .Y(n_665) );
INVx1_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
INVx1_ASAP7_75t_L g663 ( .A(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g667 ( .A(n_668), .Y(n_667) );
NOR2xp33_ASAP7_75t_L g673 ( .A(n_674), .B(n_675), .Y(n_673) );
INVx1_ASAP7_75t_L g683 ( .A(n_681), .Y(n_683) );
INVx1_ASAP7_75t_L g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g694 ( .A(n_689), .Y(n_694) );
INVx2_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
INVx2_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
NAND2xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_705), .Y(n_700) );
NOR2xp33_ASAP7_75t_SL g701 ( .A(n_702), .B(n_704), .Y(n_701) );
INVx1_ASAP7_75t_SL g721 ( .A(n_702), .Y(n_721) );
INVx1_ASAP7_75t_L g720 ( .A(n_704), .Y(n_720) );
OA21x2_ASAP7_75t_L g723 ( .A1(n_704), .A2(n_721), .B(n_724), .Y(n_723) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_705), .A2(n_710), .B(n_712), .Y(n_709) );
INVx1_ASAP7_75t_SL g705 ( .A(n_706), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_707), .Y(n_706) );
INVx1_ASAP7_75t_SL g714 ( .A(n_707), .Y(n_714) );
BUFx2_ASAP7_75t_L g724 ( .A(n_707), .Y(n_724) );
INVxp67_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
NOR2xp33_ASAP7_75t_SL g712 ( .A(n_713), .B(n_715), .Y(n_712) );
INVx1_ASAP7_75t_SL g713 ( .A(n_714), .Y(n_713) );
CKINVDCx20_ASAP7_75t_R g716 ( .A(n_717), .Y(n_716) );
CKINVDCx6p67_ASAP7_75t_R g717 ( .A(n_718), .Y(n_717) );
AND2x2_ASAP7_75t_L g718 ( .A(n_719), .B(n_721), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
CKINVDCx20_ASAP7_75t_R g722 ( .A(n_723), .Y(n_722) );
endmodule