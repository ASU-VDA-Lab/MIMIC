module fake_jpeg_26464_n_106 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_106);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_106;

wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_24),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_8),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_26),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_22),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx5_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_48),
.Y(n_66)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_49),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_0),
.B(n_1),
.Y(n_50)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_37),
.C(n_38),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

INVx3_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

INVx6_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

INVx5_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g56 ( 
.A1(n_53),
.A2(n_40),
.B1(n_42),
.B2(n_12),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_56),
.B(n_60),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_61),
.Y(n_70)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_45),
.B1(n_38),
.B2(n_37),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_62),
.A2(n_64),
.B1(n_41),
.B2(n_36),
.Y(n_75)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_67),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_53),
.A2(n_45),
.B1(n_46),
.B2(n_44),
.Y(n_64)
);

INVx13_ASAP7_75t_L g67 ( 
.A(n_49),
.Y(n_67)
);

INVx4_ASAP7_75t_SL g68 ( 
.A(n_67),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_69),
.Y(n_91)
);

CKINVDCx14_ASAP7_75t_R g69 ( 
.A(n_66),
.Y(n_69)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_66),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_71),
.B(n_72),
.Y(n_88)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_82),
.C(n_3),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_89)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_57),
.Y(n_76)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_76),
.A2(n_79),
.B(n_80),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_65),
.B(n_15),
.C(n_33),
.Y(n_78)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_78),
.B(n_18),
.C(n_28),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_59),
.B(n_0),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_1),
.Y(n_80)
);

OAI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_81),
.A2(n_73),
.B1(n_70),
.B2(n_68),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_60),
.B(n_2),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_2),
.B(n_3),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_84),
.B(n_86),
.C(n_90),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_85),
.B(n_89),
.Y(n_94)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_75),
.A2(n_81),
.B1(n_78),
.B2(n_19),
.Y(n_90)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_88),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_92),
.B(n_91),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_92),
.B(n_95),
.C(n_94),
.Y(n_96)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_96),
.A2(n_98),
.B1(n_91),
.B2(n_83),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g97 ( 
.A(n_93),
.Y(n_97)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_97),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_86),
.Y(n_101)
);

FAx1_ASAP7_75t_SL g102 ( 
.A(n_101),
.B(n_99),
.CI(n_21),
.CON(n_102),
.SN(n_102)
);

BUFx24_ASAP7_75t_SL g103 ( 
.A(n_102),
.Y(n_103)
);

AOI322xp5_ASAP7_75t_L g104 ( 
.A1(n_103),
.A2(n_102),
.A3(n_13),
.B1(n_23),
.B2(n_9),
.C1(n_10),
.C2(n_34),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_25),
.B(n_27),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_SL g106 ( 
.A(n_105),
.B(n_5),
.Y(n_106)
);


endmodule