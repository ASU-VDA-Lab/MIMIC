module fake_netlist_5_170_n_1933 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1933);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1933;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_343;
wire n_1449;
wire n_308;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_182;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1883;
wire n_1906;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_434;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1571;
wire n_187;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_368;
wire n_433;
wire n_314;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_204;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_185;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_239;
wire n_630;
wire n_1902;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_174;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1768;
wire n_321;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_212;
wire n_385;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_814;
wire n_192;
wire n_1549;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_178;
wire n_1814;
wire n_1035;
wire n_287;
wire n_783;
wire n_555;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_990;
wire n_836;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_917;
wire n_601;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1059;
wire n_1345;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_177;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_179;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1184;
wire n_1011;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1530;
wire n_1497;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_186;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_428;
wire n_379;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_273;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_180;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_437;
wire n_1642;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_175;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_1089;
wire n_927;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_35),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_125),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_4),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_91),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_97),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx10_ASAP7_75t_L g179 ( 
.A(n_88),
.Y(n_179)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_157),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_76),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_55),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_22),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_78),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_69),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_152),
.Y(n_186)
);

BUFx10_ASAP7_75t_L g187 ( 
.A(n_143),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_59),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_165),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_16),
.Y(n_190)
);

BUFx5_ASAP7_75t_L g191 ( 
.A(n_60),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_132),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_160),
.Y(n_194)
);

BUFx10_ASAP7_75t_L g195 ( 
.A(n_109),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_32),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_87),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_158),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_93),
.Y(n_199)
);

BUFx10_ASAP7_75t_L g200 ( 
.A(n_35),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_101),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_130),
.Y(n_202)
);

BUFx3_ASAP7_75t_L g203 ( 
.A(n_73),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_21),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_139),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_124),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_46),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_129),
.Y(n_209)
);

INVx2_ASAP7_75t_SL g210 ( 
.A(n_162),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_172),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_136),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_45),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_89),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_40),
.Y(n_215)
);

BUFx2_ASAP7_75t_L g216 ( 
.A(n_84),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_33),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_123),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_42),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_127),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_153),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g222 ( 
.A(n_71),
.Y(n_222)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_167),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_114),
.Y(n_224)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_6),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_140),
.Y(n_226)
);

BUFx3_ASAP7_75t_L g227 ( 
.A(n_67),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_112),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_29),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_58),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_61),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_18),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_135),
.Y(n_234)
);

BUFx3_ASAP7_75t_L g235 ( 
.A(n_142),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_66),
.Y(n_236)
);

INVx1_ASAP7_75t_SL g237 ( 
.A(n_24),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_147),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_42),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_20),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_0),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_83),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_19),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_126),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_96),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_3),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_154),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_15),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_169),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_6),
.Y(n_250)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_111),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_45),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_95),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_44),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_141),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_39),
.Y(n_256)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_11),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_77),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_155),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_55),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_108),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_52),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_102),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_62),
.Y(n_265)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_104),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_105),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_103),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_34),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_47),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_9),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_119),
.Y(n_272)
);

BUFx3_ASAP7_75t_L g273 ( 
.A(n_47),
.Y(n_273)
);

BUFx3_ASAP7_75t_L g274 ( 
.A(n_23),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_100),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_117),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_70),
.Y(n_277)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_22),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_9),
.Y(n_279)
);

BUFx3_ASAP7_75t_L g280 ( 
.A(n_74),
.Y(n_280)
);

INVx1_ASAP7_75t_SL g281 ( 
.A(n_56),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_2),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_43),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_18),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_121),
.Y(n_285)
);

BUFx10_ASAP7_75t_L g286 ( 
.A(n_51),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_29),
.Y(n_287)
);

BUFx5_ASAP7_75t_L g288 ( 
.A(n_0),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_53),
.Y(n_289)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_85),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_37),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_38),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_128),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_90),
.Y(n_294)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_38),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_113),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_156),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_23),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_159),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_80),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_64),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_19),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_65),
.Y(n_303)
);

CKINVDCx5p33_ASAP7_75t_R g304 ( 
.A(n_41),
.Y(n_304)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_59),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_31),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_137),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_32),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_118),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_170),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_115),
.Y(n_311)
);

INVx1_ASAP7_75t_SL g312 ( 
.A(n_50),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_53),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_148),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_138),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_122),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_13),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_120),
.Y(n_318)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_163),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_50),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_133),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_49),
.Y(n_322)
);

BUFx6f_ASAP7_75t_L g323 ( 
.A(n_54),
.Y(n_323)
);

BUFx6f_ASAP7_75t_L g324 ( 
.A(n_82),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_8),
.Y(n_325)
);

CKINVDCx16_ASAP7_75t_R g326 ( 
.A(n_46),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_33),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_51),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_72),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_39),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_3),
.Y(n_331)
);

BUFx2_ASAP7_75t_R g332 ( 
.A(n_106),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_7),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_4),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_43),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_26),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_60),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_86),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_28),
.Y(n_339)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_161),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_61),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_81),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_166),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_92),
.Y(n_344)
);

CKINVDCx16_ASAP7_75t_R g345 ( 
.A(n_305),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_177),
.Y(n_346)
);

BUFx2_ASAP7_75t_L g347 ( 
.A(n_295),
.Y(n_347)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_257),
.Y(n_348)
);

NOR2xp67_ASAP7_75t_L g349 ( 
.A(n_225),
.B(n_1),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_191),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_175),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_206),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_191),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_191),
.Y(n_354)
);

INVxp67_ASAP7_75t_SL g355 ( 
.A(n_216),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_207),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_201),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_191),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_339),
.B(n_1),
.Y(n_359)
);

NOR2xp33_ASAP7_75t_L g360 ( 
.A(n_210),
.B(n_2),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_209),
.Y(n_361)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_249),
.Y(n_362)
);

CKINVDCx20_ASAP7_75t_R g363 ( 
.A(n_258),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_211),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_212),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_191),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_191),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_214),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_220),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_191),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_210),
.B(n_223),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_262),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_191),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_288),
.Y(n_375)
);

HB1xp67_ASAP7_75t_L g376 ( 
.A(n_326),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_288),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_288),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_273),
.B(n_5),
.Y(n_379)
);

INVxp33_ASAP7_75t_L g380 ( 
.A(n_182),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_288),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_221),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_224),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_288),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_288),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_228),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_288),
.Y(n_387)
);

BUFx2_ASAP7_75t_L g388 ( 
.A(n_273),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_288),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_233),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_233),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_233),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_234),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_236),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_233),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_233),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_323),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_173),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_275),
.Y(n_399)
);

BUFx10_ASAP7_75t_L g400 ( 
.A(n_251),
.Y(n_400)
);

CKINVDCx16_ASAP7_75t_R g401 ( 
.A(n_180),
.Y(n_401)
);

AND2x2_ASAP7_75t_L g402 ( 
.A(n_274),
.B(n_5),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_238),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_323),
.Y(n_404)
);

CKINVDCx16_ASAP7_75t_R g405 ( 
.A(n_222),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_323),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_242),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_247),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g409 ( 
.A(n_179),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g410 ( 
.A(n_188),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_255),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g412 ( 
.A(n_259),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_261),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_264),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_267),
.Y(n_415)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_272),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_277),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_223),
.B(n_7),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_323),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_285),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_293),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_294),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_297),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_323),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g425 ( 
.A(n_173),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_299),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g427 ( 
.A(n_183),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_251),
.Y(n_428)
);

INVxp67_ASAP7_75t_L g429 ( 
.A(n_229),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_303),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_428),
.Y(n_431)
);

BUFx10_ASAP7_75t_L g432 ( 
.A(n_352),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_404),
.B(n_203),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g434 ( 
.A(n_346),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_404),
.B(n_372),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g436 ( 
.A(n_345),
.Y(n_436)
);

HB1xp67_ASAP7_75t_L g437 ( 
.A(n_376),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_390),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_390),
.Y(n_439)
);

NOR2xp67_ASAP7_75t_L g440 ( 
.A(n_350),
.B(n_176),
.Y(n_440)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_428),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g442 ( 
.A(n_345),
.B(n_179),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_356),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_391),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_357),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_362),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_391),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

INVx2_ASAP7_75t_L g449 ( 
.A(n_381),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_361),
.Y(n_450)
);

AND2x4_ASAP7_75t_L g451 ( 
.A(n_379),
.B(n_203),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g452 ( 
.A(n_359),
.B(n_179),
.Y(n_452)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_360),
.B(n_290),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_392),
.Y(n_454)
);

BUFx3_ASAP7_75t_L g455 ( 
.A(n_400),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_409),
.B(n_185),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_392),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_381),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_395),
.Y(n_459)
);

BUFx2_ASAP7_75t_L g460 ( 
.A(n_388),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_363),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g462 ( 
.A(n_355),
.B(n_290),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_364),
.Y(n_463)
);

BUFx2_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_365),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_368),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_369),
.Y(n_468)
);

INVx2_ASAP7_75t_L g469 ( 
.A(n_381),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

INVx4_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_396),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_396),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_379),
.B(n_227),
.Y(n_474)
);

CKINVDCx5p33_ASAP7_75t_R g475 ( 
.A(n_370),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_397),
.Y(n_476)
);

AND2x4_ASAP7_75t_L g477 ( 
.A(n_402),
.B(n_227),
.Y(n_477)
);

BUFx2_ASAP7_75t_L g478 ( 
.A(n_398),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_384),
.Y(n_479)
);

BUFx2_ASAP7_75t_L g480 ( 
.A(n_425),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_382),
.Y(n_481)
);

BUFx2_ASAP7_75t_L g482 ( 
.A(n_427),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_397),
.Y(n_483)
);

INVx2_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

BUFx6f_ASAP7_75t_L g485 ( 
.A(n_350),
.Y(n_485)
);

HB1xp67_ASAP7_75t_L g486 ( 
.A(n_347),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_383),
.Y(n_487)
);

BUFx6f_ASAP7_75t_L g488 ( 
.A(n_353),
.Y(n_488)
);

OA21x2_ASAP7_75t_L g489 ( 
.A1(n_353),
.A2(n_240),
.B(n_225),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_386),
.Y(n_490)
);

INVx3_ASAP7_75t_L g491 ( 
.A(n_354),
.Y(n_491)
);

INVx2_ASAP7_75t_L g492 ( 
.A(n_354),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_406),
.Y(n_493)
);

INVx3_ASAP7_75t_L g494 ( 
.A(n_358),
.Y(n_494)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_348),
.B(n_319),
.Y(n_495)
);

BUFx3_ASAP7_75t_L g496 ( 
.A(n_400),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_406),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_419),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_419),
.B(n_174),
.Y(n_499)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_373),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_399),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_358),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_366),
.Y(n_503)
);

INVxp67_ASAP7_75t_L g504 ( 
.A(n_347),
.Y(n_504)
);

BUFx6f_ASAP7_75t_L g505 ( 
.A(n_366),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_402),
.B(n_235),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_393),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_489),
.Y(n_508)
);

INVx3_ASAP7_75t_L g509 ( 
.A(n_479),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_449),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_435),
.B(n_394),
.Y(n_511)
);

AND2x2_ASAP7_75t_L g512 ( 
.A(n_506),
.B(n_424),
.Y(n_512)
);

AOI22xp33_ASAP7_75t_L g513 ( 
.A1(n_453),
.A2(n_418),
.B1(n_349),
.B2(n_348),
.Y(n_513)
);

BUFx6f_ASAP7_75t_L g514 ( 
.A(n_479),
.Y(n_514)
);

BUFx3_ASAP7_75t_L g515 ( 
.A(n_433),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_434),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_452),
.B(n_403),
.Y(n_517)
);

OR2x6_ASAP7_75t_L g518 ( 
.A(n_456),
.B(n_351),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_479),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_452),
.B(n_411),
.Y(n_520)
);

INVxp67_ASAP7_75t_SL g521 ( 
.A(n_479),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_489),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_479),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_432),
.B(n_401),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_489),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_489),
.Y(n_526)
);

INVx2_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

BUFx6f_ASAP7_75t_L g528 ( 
.A(n_479),
.Y(n_528)
);

NAND3xp33_ASAP7_75t_L g529 ( 
.A(n_453),
.B(n_414),
.C(n_413),
.Y(n_529)
);

NOR2x1p5_ASAP7_75t_L g530 ( 
.A(n_443),
.B(n_274),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_489),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_435),
.B(n_415),
.Y(n_532)
);

AOI22xp33_ASAP7_75t_L g533 ( 
.A1(n_462),
.A2(n_349),
.B1(n_240),
.B2(n_336),
.Y(n_533)
);

BUFx2_ASAP7_75t_L g534 ( 
.A(n_460),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_491),
.Y(n_535)
);

BUFx6f_ASAP7_75t_L g536 ( 
.A(n_479),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_492),
.Y(n_537)
);

AND2x2_ASAP7_75t_L g538 ( 
.A(n_506),
.B(n_424),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_492),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_492),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_460),
.Y(n_541)
);

NOR2xp33_ASAP7_75t_L g542 ( 
.A(n_450),
.B(n_420),
.Y(n_542)
);

AND2x2_ASAP7_75t_L g543 ( 
.A(n_506),
.B(n_380),
.Y(n_543)
);

AOI22xp33_ASAP7_75t_L g544 ( 
.A1(n_462),
.A2(n_278),
.B1(n_336),
.B2(n_291),
.Y(n_544)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_486),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_485),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_503),
.Y(n_547)
);

INVx3_ASAP7_75t_L g548 ( 
.A(n_485),
.Y(n_548)
);

INVx3_ASAP7_75t_L g549 ( 
.A(n_485),
.Y(n_549)
);

INVx4_ASAP7_75t_SL g550 ( 
.A(n_485),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_449),
.Y(n_551)
);

INVx2_ASAP7_75t_L g552 ( 
.A(n_458),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g553 ( 
.A1(n_456),
.A2(n_416),
.B1(n_407),
.B2(n_408),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_503),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_485),
.Y(n_555)
);

AOI22xp33_ASAP7_75t_L g556 ( 
.A1(n_433),
.A2(n_278),
.B1(n_270),
.B2(n_263),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_442),
.A2(n_417),
.B1(n_412),
.B2(n_401),
.Y(n_557)
);

INVx1_ASAP7_75t_L g558 ( 
.A(n_503),
.Y(n_558)
);

BUFx4f_ASAP7_75t_L g559 ( 
.A(n_485),
.Y(n_559)
);

BUFx3_ASAP7_75t_L g560 ( 
.A(n_433),
.Y(n_560)
);

AO21x2_ASAP7_75t_L g561 ( 
.A1(n_440),
.A2(n_193),
.B(n_186),
.Y(n_561)
);

NAND3xp33_ASAP7_75t_L g562 ( 
.A(n_495),
.B(n_422),
.C(n_421),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_458),
.Y(n_563)
);

OR2x6_ASAP7_75t_L g564 ( 
.A(n_464),
.B(n_351),
.Y(n_564)
);

INVx1_ASAP7_75t_SL g565 ( 
.A(n_464),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_433),
.B(n_423),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_463),
.B(n_426),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_491),
.Y(n_568)
);

NOR2xp67_ASAP7_75t_L g569 ( 
.A(n_471),
.B(n_430),
.Y(n_569)
);

INVx2_ASAP7_75t_L g570 ( 
.A(n_458),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_485),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_469),
.Y(n_573)
);

CKINVDCx5p33_ASAP7_75t_R g574 ( 
.A(n_445),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_466),
.B(n_405),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_432),
.B(n_405),
.Y(n_576)
);

INVx5_ASAP7_75t_L g577 ( 
.A(n_488),
.Y(n_577)
);

INVxp67_ASAP7_75t_SL g578 ( 
.A(n_491),
.Y(n_578)
);

OR2x6_ASAP7_75t_L g579 ( 
.A(n_478),
.B(n_410),
.Y(n_579)
);

INVx6_ASAP7_75t_L g580 ( 
.A(n_471),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_494),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_433),
.Y(n_582)
);

BUFx6f_ASAP7_75t_L g583 ( 
.A(n_488),
.Y(n_583)
);

AND2x4_ASAP7_75t_L g584 ( 
.A(n_451),
.B(n_474),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_494),
.Y(n_585)
);

AND2x2_ASAP7_75t_L g586 ( 
.A(n_451),
.B(n_410),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_469),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_471),
.B(n_235),
.Y(n_588)
);

INVx3_ASAP7_75t_R g589 ( 
.A(n_478),
.Y(n_589)
);

INVx4_ASAP7_75t_SL g590 ( 
.A(n_488),
.Y(n_590)
);

BUFx2_ASAP7_75t_L g591 ( 
.A(n_437),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_494),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_494),
.Y(n_593)
);

INVx3_ASAP7_75t_L g594 ( 
.A(n_488),
.Y(n_594)
);

BUFx2_ASAP7_75t_L g595 ( 
.A(n_437),
.Y(n_595)
);

BUFx3_ASAP7_75t_L g596 ( 
.A(n_455),
.Y(n_596)
);

INVx4_ASAP7_75t_L g597 ( 
.A(n_488),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_469),
.Y(n_598)
);

INVx3_ASAP7_75t_L g599 ( 
.A(n_488),
.Y(n_599)
);

AND2x4_ASAP7_75t_L g600 ( 
.A(n_451),
.B(n_266),
.Y(n_600)
);

INVx4_ASAP7_75t_L g601 ( 
.A(n_488),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_451),
.B(n_367),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_451),
.B(n_367),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_438),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_436),
.Y(n_605)
);

AO21x2_ASAP7_75t_L g606 ( 
.A1(n_440),
.A2(n_204),
.B(n_202),
.Y(n_606)
);

NAND2xp5_ASAP7_75t_SL g607 ( 
.A(n_432),
.B(n_409),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

INVx4_ASAP7_75t_L g609 ( 
.A(n_502),
.Y(n_609)
);

BUFx6f_ASAP7_75t_L g610 ( 
.A(n_502),
.Y(n_610)
);

AND2x2_ASAP7_75t_SL g611 ( 
.A(n_474),
.B(n_319),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_SL g612 ( 
.A(n_432),
.B(n_185),
.Y(n_612)
);

NOR2xp33_ASAP7_75t_L g613 ( 
.A(n_467),
.B(n_429),
.Y(n_613)
);

NAND2xp33_ASAP7_75t_R g614 ( 
.A(n_480),
.B(n_482),
.Y(n_614)
);

INVx1_ASAP7_75t_L g615 ( 
.A(n_438),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_432),
.B(n_468),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_470),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_475),
.B(n_185),
.Y(n_618)
);

INVx2_ASAP7_75t_L g619 ( 
.A(n_470),
.Y(n_619)
);

HB1xp67_ASAP7_75t_L g620 ( 
.A(n_486),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_474),
.B(n_371),
.Y(n_621)
);

AND2x4_ASAP7_75t_SL g622 ( 
.A(n_446),
.B(n_187),
.Y(n_622)
);

AND2x2_ASAP7_75t_L g623 ( 
.A(n_474),
.B(n_429),
.Y(n_623)
);

AND2x2_ASAP7_75t_L g624 ( 
.A(n_474),
.B(n_371),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_439),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_477),
.Y(n_626)
);

INVx1_ASAP7_75t_L g627 ( 
.A(n_439),
.Y(n_627)
);

INVx4_ASAP7_75t_L g628 ( 
.A(n_502),
.Y(n_628)
);

OAI22xp33_ASAP7_75t_SL g629 ( 
.A1(n_499),
.A2(n_280),
.B1(n_266),
.B2(n_301),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_481),
.B(n_174),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_444),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_455),
.Y(n_632)
);

INVx4_ASAP7_75t_L g633 ( 
.A(n_502),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_470),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_484),
.Y(n_635)
);

NOR2xp33_ASAP7_75t_L g636 ( 
.A(n_487),
.B(n_178),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_490),
.B(n_187),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_477),
.B(n_374),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_484),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_444),
.Y(n_640)
);

BUFx6f_ASAP7_75t_L g641 ( 
.A(n_502),
.Y(n_641)
);

INVx1_ASAP7_75t_SL g642 ( 
.A(n_461),
.Y(n_642)
);

AND2x6_ASAP7_75t_L g643 ( 
.A(n_477),
.B(n_251),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_SL g644 ( 
.A(n_507),
.B(n_187),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_484),
.Y(n_645)
);

BUFx6f_ASAP7_75t_L g646 ( 
.A(n_502),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_447),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_447),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_500),
.Y(n_649)
);

AND2x4_ASAP7_75t_L g650 ( 
.A(n_477),
.B(n_280),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_505),
.Y(n_651)
);

INVxp67_ASAP7_75t_SL g652 ( 
.A(n_505),
.Y(n_652)
);

INVx3_ASAP7_75t_L g653 ( 
.A(n_505),
.Y(n_653)
);

INVx2_ASAP7_75t_L g654 ( 
.A(n_454),
.Y(n_654)
);

INVx3_ASAP7_75t_L g655 ( 
.A(n_505),
.Y(n_655)
);

BUFx3_ASAP7_75t_L g656 ( 
.A(n_455),
.Y(n_656)
);

INVx4_ASAP7_75t_L g657 ( 
.A(n_505),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_454),
.Y(n_658)
);

AND2x4_ASAP7_75t_L g659 ( 
.A(n_477),
.B(n_301),
.Y(n_659)
);

BUFx4f_ASAP7_75t_L g660 ( 
.A(n_505),
.Y(n_660)
);

AOI21xp5_ASAP7_75t_L g661 ( 
.A1(n_582),
.A2(n_603),
.B(n_602),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_532),
.B(n_471),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_611),
.A2(n_508),
.B1(n_525),
.B2(n_522),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_511),
.B(n_496),
.Y(n_664)
);

INVx2_ASAP7_75t_SL g665 ( 
.A(n_543),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_582),
.B(n_496),
.Y(n_666)
);

NAND2x1_ASAP7_75t_L g667 ( 
.A(n_580),
.B(n_584),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_510),
.Y(n_668)
);

NOR2xp33_ASAP7_75t_L g669 ( 
.A(n_529),
.B(n_504),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_588),
.B(n_307),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_611),
.B(n_496),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_515),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_515),
.B(n_499),
.Y(n_673)
);

NOR2xp33_ASAP7_75t_L g674 ( 
.A(n_517),
.B(n_504),
.Y(n_674)
);

NOR2xp33_ASAP7_75t_L g675 ( 
.A(n_520),
.B(n_613),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_510),
.Y(n_676)
);

NOR2x1p5_ASAP7_75t_L g677 ( 
.A(n_562),
.B(n_183),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_566),
.B(n_480),
.Y(n_678)
);

INVx2_ASAP7_75t_L g679 ( 
.A(n_527),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_560),
.B(n_624),
.Y(n_680)
);

NAND2xp5_ASAP7_75t_SL g681 ( 
.A(n_584),
.B(n_436),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_560),
.B(n_505),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_584),
.B(n_251),
.Y(n_683)
);

NAND2x1_ASAP7_75t_L g684 ( 
.A(n_580),
.B(n_457),
.Y(n_684)
);

NOR2xp33_ASAP7_75t_L g685 ( 
.A(n_630),
.B(n_482),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_527),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_L g687 ( 
.A(n_636),
.B(n_495),
.Y(n_687)
);

A2O1A1Ixp33_ASAP7_75t_L g688 ( 
.A1(n_624),
.A2(n_374),
.B(n_375),
.C(n_377),
.Y(n_688)
);

INVx2_ASAP7_75t_SL g689 ( 
.A(n_543),
.Y(n_689)
);

INVx2_ASAP7_75t_L g690 ( 
.A(n_551),
.Y(n_690)
);

INVx2_ASAP7_75t_L g691 ( 
.A(n_551),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_626),
.B(n_457),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_552),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_626),
.Y(n_694)
);

INVx2_ASAP7_75t_L g695 ( 
.A(n_552),
.Y(n_695)
);

AOI21xp5_ASAP7_75t_L g696 ( 
.A1(n_621),
.A2(n_465),
.B(n_459),
.Y(n_696)
);

AOI22xp33_ASAP7_75t_L g697 ( 
.A1(n_508),
.A2(n_241),
.B1(n_306),
.B2(n_243),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_512),
.B(n_459),
.Y(n_698)
);

BUFx6f_ASAP7_75t_L g699 ( 
.A(n_600),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_512),
.Y(n_700)
);

CKINVDCx5p33_ASAP7_75t_R g701 ( 
.A(n_516),
.Y(n_701)
);

AOI22xp5_ASAP7_75t_L g702 ( 
.A1(n_586),
.A2(n_316),
.B1(n_184),
.B2(n_181),
.Y(n_702)
);

OAI22xp5_ASAP7_75t_L g703 ( 
.A1(n_580),
.A2(n_245),
.B1(n_310),
.B2(n_314),
.Y(n_703)
);

INVx8_ASAP7_75t_L g704 ( 
.A(n_564),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_538),
.B(n_465),
.Y(n_705)
);

AND2x6_ASAP7_75t_SL g706 ( 
.A(n_575),
.B(n_232),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_538),
.B(n_472),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_580),
.B(n_472),
.Y(n_708)
);

INVxp67_ASAP7_75t_L g709 ( 
.A(n_614),
.Y(n_709)
);

BUFx3_ASAP7_75t_L g710 ( 
.A(n_596),
.Y(n_710)
);

INVx1_ASAP7_75t_L g711 ( 
.A(n_638),
.Y(n_711)
);

AOI22xp5_ASAP7_75t_L g712 ( 
.A1(n_586),
.A2(n_178),
.B1(n_181),
.B2(n_184),
.Y(n_712)
);

INVxp67_ASAP7_75t_L g713 ( 
.A(n_534),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_578),
.B(n_473),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_623),
.B(n_473),
.Y(n_715)
);

INVx2_ASAP7_75t_L g716 ( 
.A(n_563),
.Y(n_716)
);

NAND2xp33_ASAP7_75t_L g717 ( 
.A(n_588),
.B(n_251),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_623),
.B(n_476),
.Y(n_718)
);

AND2x4_ASAP7_75t_L g719 ( 
.A(n_600),
.B(n_226),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_SL g720 ( 
.A(n_588),
.B(n_300),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_563),
.Y(n_721)
);

O2A1O1Ixp33_ASAP7_75t_L g722 ( 
.A1(n_522),
.A2(n_254),
.B(n_282),
.C(n_284),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_525),
.B(n_476),
.Y(n_723)
);

NAND2xp5_ASAP7_75t_SL g724 ( 
.A(n_569),
.B(n_300),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_564),
.B(n_237),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_534),
.Y(n_726)
);

NAND2xp33_ASAP7_75t_L g727 ( 
.A(n_643),
.B(n_300),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_604),
.Y(n_728)
);

NOR2xp33_ASAP7_75t_L g729 ( 
.A(n_564),
.B(n_281),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_604),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_600),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_526),
.B(n_300),
.Y(n_732)
);

AOI22xp5_ASAP7_75t_L g733 ( 
.A1(n_518),
.A2(n_318),
.B1(n_192),
.B2(n_194),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_526),
.B(n_300),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_531),
.B(n_483),
.Y(n_735)
);

INVx3_ASAP7_75t_L g736 ( 
.A(n_650),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_570),
.Y(n_737)
);

OAI22xp5_ASAP7_75t_L g738 ( 
.A1(n_513),
.A2(n_244),
.B1(n_253),
.B2(n_276),
.Y(n_738)
);

INVx8_ASAP7_75t_L g739 ( 
.A(n_564),
.Y(n_739)
);

INVx2_ASAP7_75t_L g740 ( 
.A(n_570),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_612),
.B(n_312),
.Y(n_741)
);

AOI22xp5_ASAP7_75t_L g742 ( 
.A1(n_518),
.A2(n_321),
.B1(n_192),
.B2(n_194),
.Y(n_742)
);

AOI22xp33_ASAP7_75t_L g743 ( 
.A1(n_531),
.A2(n_544),
.B1(n_606),
.B2(n_561),
.Y(n_743)
);

BUFx3_ASAP7_75t_L g744 ( 
.A(n_596),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_650),
.B(n_483),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_650),
.B(n_493),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_573),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_SL g748 ( 
.A(n_568),
.B(n_324),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_659),
.B(n_493),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_556),
.B(n_208),
.C(n_205),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_659),
.B(n_497),
.Y(n_751)
);

AND2x4_ASAP7_75t_L g752 ( 
.A(n_659),
.B(n_268),
.Y(n_752)
);

INVx2_ASAP7_75t_L g753 ( 
.A(n_573),
.Y(n_753)
);

AOI22xp33_ASAP7_75t_L g754 ( 
.A1(n_561),
.A2(n_313),
.B1(n_246),
.B2(n_327),
.Y(n_754)
);

OR2x2_ASAP7_75t_L g755 ( 
.A(n_565),
.B(n_335),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_615),
.Y(n_756)
);

NOR2xp33_ASAP7_75t_L g757 ( 
.A(n_518),
.B(n_189),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_587),
.Y(n_758)
);

HB1xp67_ASAP7_75t_L g759 ( 
.A(n_620),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_625),
.Y(n_760)
);

NOR2x1_ASAP7_75t_L g761 ( 
.A(n_542),
.B(n_315),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_SL g762 ( 
.A(n_568),
.B(n_324),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_561),
.A2(n_317),
.B1(n_298),
.B2(n_387),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_625),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_627),
.B(n_497),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_627),
.B(n_498),
.Y(n_766)
);

BUFx5_ASAP7_75t_L g767 ( 
.A(n_572),
.Y(n_767)
);

NAND2xp5_ASAP7_75t_L g768 ( 
.A(n_631),
.B(n_498),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_572),
.B(n_324),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_606),
.A2(n_385),
.B1(n_375),
.B2(n_377),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_631),
.Y(n_771)
);

A2O1A1Ixp33_ASAP7_75t_L g772 ( 
.A1(n_581),
.A2(n_378),
.B(n_385),
.C(n_387),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_640),
.B(n_338),
.Y(n_773)
);

INVx2_ASAP7_75t_SL g774 ( 
.A(n_541),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_518),
.B(n_189),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_640),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_647),
.B(n_378),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_579),
.B(n_332),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_L g779 ( 
.A(n_647),
.B(n_389),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_648),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_648),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_587),
.Y(n_782)
);

INVxp67_ASAP7_75t_L g783 ( 
.A(n_541),
.Y(n_783)
);

AOI22xp33_ASAP7_75t_L g784 ( 
.A1(n_606),
.A2(n_389),
.B1(n_320),
.B2(n_217),
.Y(n_784)
);

INVx1_ASAP7_75t_L g785 ( 
.A(n_658),
.Y(n_785)
);

INVx8_ASAP7_75t_L g786 ( 
.A(n_579),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_598),
.Y(n_787)
);

NOR2xp67_ASAP7_75t_L g788 ( 
.A(n_567),
.B(n_197),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_632),
.A2(n_197),
.B1(n_344),
.B2(n_343),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_658),
.Y(n_790)
);

NAND2x1p5_ASAP7_75t_L g791 ( 
.A(n_632),
.B(n_324),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_581),
.B(n_431),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_592),
.B(n_431),
.Y(n_793)
);

INVx2_ASAP7_75t_SL g794 ( 
.A(n_591),
.Y(n_794)
);

INVx4_ASAP7_75t_L g795 ( 
.A(n_546),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_598),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_654),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_592),
.B(n_431),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_593),
.B(n_441),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_593),
.B(n_441),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_516),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_533),
.A2(n_196),
.B1(n_289),
.B2(n_302),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_SL g803 ( 
.A(n_535),
.B(n_324),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_SL g804 ( 
.A(n_585),
.B(n_340),
.Y(n_804)
);

AOI22xp5_ASAP7_75t_L g805 ( 
.A1(n_530),
.A2(n_318),
.B1(n_344),
.B2(n_343),
.Y(n_805)
);

BUFx2_ASAP7_75t_L g806 ( 
.A(n_579),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_629),
.B(n_340),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_643),
.A2(n_340),
.B1(n_337),
.B2(n_334),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_521),
.B(n_441),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_654),
.B(n_340),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_SL g811 ( 
.A(n_514),
.B(n_340),
.Y(n_811)
);

OR2x2_ASAP7_75t_L g812 ( 
.A(n_591),
.B(n_190),
.Y(n_812)
);

A2O1A1Ixp33_ASAP7_75t_L g813 ( 
.A1(n_537),
.A2(n_190),
.B(n_308),
.C(n_322),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_579),
.B(n_200),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_SL g815 ( 
.A(n_514),
.B(n_198),
.Y(n_815)
);

BUFx6f_ASAP7_75t_SL g816 ( 
.A(n_589),
.Y(n_816)
);

AOI22xp5_ASAP7_75t_L g817 ( 
.A1(n_618),
.A2(n_637),
.B1(n_644),
.B2(n_607),
.Y(n_817)
);

BUFx3_ASAP7_75t_L g818 ( 
.A(n_656),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_514),
.B(n_198),
.Y(n_819)
);

INVxp67_ASAP7_75t_L g820 ( 
.A(n_595),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_652),
.B(n_448),
.Y(n_821)
);

INVx2_ASAP7_75t_SL g822 ( 
.A(n_595),
.Y(n_822)
);

BUFx6f_ASAP7_75t_L g823 ( 
.A(n_656),
.Y(n_823)
);

OR2x2_ASAP7_75t_L g824 ( 
.A(n_545),
.B(n_308),
.Y(n_824)
);

INVx3_ASAP7_75t_L g825 ( 
.A(n_617),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_514),
.B(n_199),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_524),
.B(n_199),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_509),
.B(n_448),
.Y(n_828)
);

NOR2xp67_ASAP7_75t_L g829 ( 
.A(n_553),
.B(n_309),
.Y(n_829)
);

AOI22xp5_ASAP7_75t_L g830 ( 
.A1(n_576),
.A2(n_311),
.B1(n_321),
.B2(n_309),
.Y(n_830)
);

AND2x4_ASAP7_75t_L g831 ( 
.A(n_550),
.B(n_311),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_509),
.B(n_448),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_675),
.B(n_537),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_797),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_728),
.Y(n_835)
);

NOR3xp33_ASAP7_75t_SL g836 ( 
.A(n_675),
.B(n_325),
.C(n_322),
.Y(n_836)
);

HB1xp67_ASAP7_75t_L g837 ( 
.A(n_794),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_730),
.Y(n_838)
);

NOR2x1_ASAP7_75t_L g839 ( 
.A(n_710),
.B(n_616),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_687),
.B(n_539),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_756),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_822),
.Y(n_842)
);

INVx3_ASAP7_75t_L g843 ( 
.A(n_699),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_699),
.Y(n_844)
);

INVx1_ASAP7_75t_SL g845 ( 
.A(n_774),
.Y(n_845)
);

INVx3_ASAP7_75t_L g846 ( 
.A(n_699),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_699),
.Y(n_847)
);

BUFx3_ASAP7_75t_L g848 ( 
.A(n_710),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_687),
.B(n_539),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_SL g850 ( 
.A(n_663),
.B(n_731),
.Y(n_850)
);

HB1xp67_ASAP7_75t_L g851 ( 
.A(n_759),
.Y(n_851)
);

NAND2xp33_ASAP7_75t_SL g852 ( 
.A(n_663),
.B(n_589),
.Y(n_852)
);

HB1xp67_ASAP7_75t_L g853 ( 
.A(n_759),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_731),
.B(n_557),
.Y(n_854)
);

INVx2_ASAP7_75t_L g855 ( 
.A(n_825),
.Y(n_855)
);

AND2x4_ASAP7_75t_L g856 ( 
.A(n_744),
.B(n_642),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_L g857 ( 
.A(n_674),
.B(n_622),
.Y(n_857)
);

BUFx2_ASAP7_75t_L g858 ( 
.A(n_713),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_760),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_744),
.Y(n_860)
);

NAND2x1p5_ASAP7_75t_L g861 ( 
.A(n_667),
.B(n_731),
.Y(n_861)
);

BUFx3_ASAP7_75t_L g862 ( 
.A(n_818),
.Y(n_862)
);

BUFx6f_ASAP7_75t_L g863 ( 
.A(n_731),
.Y(n_863)
);

INVx2_ASAP7_75t_L g864 ( 
.A(n_825),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_764),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_771),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_776),
.Y(n_867)
);

INVx2_ASAP7_75t_L g868 ( 
.A(n_668),
.Y(n_868)
);

INVx1_ASAP7_75t_SL g869 ( 
.A(n_755),
.Y(n_869)
);

NOR3xp33_ASAP7_75t_SL g870 ( 
.A(n_685),
.B(n_328),
.C(n_325),
.Y(n_870)
);

OR2x6_ASAP7_75t_L g871 ( 
.A(n_704),
.B(n_501),
.Y(n_871)
);

BUFx10_ASAP7_75t_L g872 ( 
.A(n_816),
.Y(n_872)
);

CKINVDCx20_ASAP7_75t_R g873 ( 
.A(n_701),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_780),
.Y(n_874)
);

AND2x2_ASAP7_75t_L g875 ( 
.A(n_674),
.B(n_622),
.Y(n_875)
);

INVx5_ASAP7_75t_L g876 ( 
.A(n_736),
.Y(n_876)
);

OR2x6_ASAP7_75t_L g877 ( 
.A(n_704),
.B(n_574),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_709),
.B(n_605),
.Y(n_878)
);

AOI22xp5_ASAP7_75t_L g879 ( 
.A1(n_669),
.A2(n_643),
.B1(n_605),
.B2(n_519),
.Y(n_879)
);

BUFx6f_ASAP7_75t_L g880 ( 
.A(n_823),
.Y(n_880)
);

INVx4_ASAP7_75t_L g881 ( 
.A(n_823),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_676),
.Y(n_882)
);

INVx8_ASAP7_75t_L g883 ( 
.A(n_786),
.Y(n_883)
);

INVx2_ASAP7_75t_SL g884 ( 
.A(n_824),
.Y(n_884)
);

BUFx12f_ASAP7_75t_L g885 ( 
.A(n_801),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_781),
.Y(n_886)
);

INVx2_ASAP7_75t_L g887 ( 
.A(n_679),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_662),
.B(n_540),
.Y(n_888)
);

NOR2x1_ASAP7_75t_L g889 ( 
.A(n_818),
.B(n_548),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_711),
.B(n_540),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_686),
.Y(n_891)
);

NOR2x1p5_ASAP7_75t_L g892 ( 
.A(n_778),
.B(n_574),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_785),
.Y(n_893)
);

BUFx2_ASAP7_75t_L g894 ( 
.A(n_726),
.Y(n_894)
);

AOI22xp5_ASAP7_75t_L g895 ( 
.A1(n_669),
.A2(n_643),
.B1(n_519),
.B2(n_509),
.Y(n_895)
);

NAND2xp33_ASAP7_75t_SL g896 ( 
.A(n_816),
.B(n_649),
.Y(n_896)
);

INVx3_ASAP7_75t_L g897 ( 
.A(n_736),
.Y(n_897)
);

INVx2_ASAP7_75t_SL g898 ( 
.A(n_812),
.Y(n_898)
);

INVx1_ASAP7_75t_L g899 ( 
.A(n_790),
.Y(n_899)
);

AOI22x1_ASAP7_75t_L g900 ( 
.A1(n_661),
.A2(n_519),
.B1(n_599),
.B2(n_655),
.Y(n_900)
);

INVxp67_ASAP7_75t_L g901 ( 
.A(n_725),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_690),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_694),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_664),
.B(n_547),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_672),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_745),
.Y(n_906)
);

INVx1_ASAP7_75t_SL g907 ( 
.A(n_814),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_691),
.Y(n_908)
);

NOR3xp33_ASAP7_75t_L g909 ( 
.A(n_741),
.B(n_649),
.C(n_329),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_693),
.Y(n_910)
);

NOR3xp33_ASAP7_75t_SL g911 ( 
.A(n_685),
.B(n_328),
.C(n_330),
.Y(n_911)
);

AND2x4_ASAP7_75t_L g912 ( 
.A(n_665),
.B(n_548),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_695),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_SL g914 ( 
.A(n_671),
.B(n_680),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_673),
.B(n_547),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_783),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_746),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_689),
.Y(n_918)
);

NOR2xp33_ASAP7_75t_R g919 ( 
.A(n_786),
.B(n_316),
.Y(n_919)
);

AND2x2_ASAP7_75t_L g920 ( 
.A(n_678),
.B(n_200),
.Y(n_920)
);

INVx2_ASAP7_75t_SL g921 ( 
.A(n_677),
.Y(n_921)
);

INVxp67_ASAP7_75t_SL g922 ( 
.A(n_823),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_715),
.B(n_554),
.Y(n_923)
);

BUFx2_ASAP7_75t_L g924 ( 
.A(n_820),
.Y(n_924)
);

HB1xp67_ASAP7_75t_L g925 ( 
.A(n_700),
.Y(n_925)
);

AND3x1_ASAP7_75t_L g926 ( 
.A(n_802),
.B(n_286),
.C(n_200),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_716),
.Y(n_927)
);

BUFx6f_ASAP7_75t_L g928 ( 
.A(n_823),
.Y(n_928)
);

NAND3xp33_ASAP7_75t_SL g929 ( 
.A(n_802),
.B(n_741),
.C(n_733),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_SL g930 ( 
.A(n_767),
.B(n_514),
.Y(n_930)
);

AND2x4_ASAP7_75t_SL g931 ( 
.A(n_719),
.B(n_195),
.Y(n_931)
);

NAND3xp33_ASAP7_75t_L g932 ( 
.A(n_678),
.B(n_256),
.C(n_269),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_749),
.Y(n_933)
);

INVx2_ASAP7_75t_L g934 ( 
.A(n_721),
.Y(n_934)
);

BUFx8_ASAP7_75t_SL g935 ( 
.A(n_806),
.Y(n_935)
);

BUFx2_ASAP7_75t_L g936 ( 
.A(n_786),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_718),
.B(n_554),
.Y(n_937)
);

INVx1_ASAP7_75t_SL g938 ( 
.A(n_725),
.Y(n_938)
);

HB1xp67_ASAP7_75t_L g939 ( 
.A(n_719),
.Y(n_939)
);

AND2x2_ASAP7_75t_L g940 ( 
.A(n_729),
.B(n_286),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_698),
.B(n_558),
.Y(n_941)
);

CKINVDCx20_ASAP7_75t_R g942 ( 
.A(n_704),
.Y(n_942)
);

INVx1_ASAP7_75t_SL g943 ( 
.A(n_729),
.Y(n_943)
);

BUFx6f_ASAP7_75t_L g944 ( 
.A(n_795),
.Y(n_944)
);

BUFx4f_ASAP7_75t_L g945 ( 
.A(n_739),
.Y(n_945)
);

INVx1_ASAP7_75t_L g946 ( 
.A(n_751),
.Y(n_946)
);

BUFx6f_ASAP7_75t_L g947 ( 
.A(n_795),
.Y(n_947)
);

AND2x2_ASAP7_75t_L g948 ( 
.A(n_757),
.B(n_286),
.Y(n_948)
);

AND2x6_ASAP7_75t_SL g949 ( 
.A(n_757),
.B(n_330),
.Y(n_949)
);

AND2x4_ASAP7_75t_L g950 ( 
.A(n_752),
.B(n_548),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_739),
.Y(n_951)
);

NOR2xp33_ASAP7_75t_L g952 ( 
.A(n_775),
.B(n_549),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_765),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_766),
.Y(n_954)
);

INVx4_ASAP7_75t_L g955 ( 
.A(n_739),
.Y(n_955)
);

BUFx3_ASAP7_75t_L g956 ( 
.A(n_752),
.Y(n_956)
);

INVx1_ASAP7_75t_L g957 ( 
.A(n_768),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_L g958 ( 
.A(n_705),
.B(n_707),
.Y(n_958)
);

HB1xp67_ASAP7_75t_L g959 ( 
.A(n_681),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_L g960 ( 
.A(n_697),
.B(n_558),
.Y(n_960)
);

AND3x1_ASAP7_75t_SL g961 ( 
.A(n_706),
.B(n_331),
.C(n_341),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_767),
.B(n_523),
.Y(n_962)
);

INVx3_ASAP7_75t_L g963 ( 
.A(n_767),
.Y(n_963)
);

INVx2_ASAP7_75t_L g964 ( 
.A(n_737),
.Y(n_964)
);

NOR2xp33_ASAP7_75t_R g965 ( 
.A(n_670),
.B(n_329),
.Y(n_965)
);

INVx2_ASAP7_75t_L g966 ( 
.A(n_740),
.Y(n_966)
);

NOR2xp33_ASAP7_75t_R g967 ( 
.A(n_775),
.B(n_827),
.Y(n_967)
);

BUFx8_ASAP7_75t_SL g968 ( 
.A(n_831),
.Y(n_968)
);

AND2x4_ASAP7_75t_L g969 ( 
.A(n_681),
.B(n_549),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_692),
.Y(n_970)
);

BUFx4f_ASAP7_75t_L g971 ( 
.A(n_831),
.Y(n_971)
);

NAND2x1_ASAP7_75t_L g972 ( 
.A(n_747),
.B(n_549),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_684),
.Y(n_973)
);

INVx1_ASAP7_75t_L g974 ( 
.A(n_753),
.Y(n_974)
);

CKINVDCx5p33_ASAP7_75t_R g975 ( 
.A(n_817),
.Y(n_975)
);

AND3x1_ASAP7_75t_SL g976 ( 
.A(n_784),
.B(n_331),
.C(n_341),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_758),
.Y(n_977)
);

INVx1_ASAP7_75t_L g978 ( 
.A(n_782),
.Y(n_978)
);

NOR2xp33_ASAP7_75t_L g979 ( 
.A(n_827),
.B(n_594),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_787),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_697),
.B(n_594),
.Y(n_981)
);

AND2x4_ASAP7_75t_L g982 ( 
.A(n_682),
.B(n_594),
.Y(n_982)
);

OAI22xp33_ASAP7_75t_L g983 ( 
.A1(n_742),
.A2(n_333),
.B1(n_334),
.B2(n_337),
.Y(n_983)
);

NAND2xp5_ASAP7_75t_L g984 ( 
.A(n_788),
.B(n_599),
.Y(n_984)
);

NOR2xp33_ASAP7_75t_R g985 ( 
.A(n_717),
.B(n_666),
.Y(n_985)
);

AOI22xp5_ASAP7_75t_SL g986 ( 
.A1(n_738),
.A2(n_333),
.B1(n_265),
.B2(n_260),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_683),
.A2(n_643),
.B1(n_599),
.B2(n_655),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_796),
.Y(n_988)
);

INVx2_ASAP7_75t_SL g989 ( 
.A(n_761),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_714),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_777),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_767),
.B(n_773),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_789),
.Y(n_993)
);

INVx3_ASAP7_75t_L g994 ( 
.A(n_767),
.Y(n_994)
);

INVx4_ASAP7_75t_L g995 ( 
.A(n_767),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_807),
.Y(n_996)
);

AOI221xp5_ASAP7_75t_L g997 ( 
.A1(n_784),
.A2(n_213),
.B1(n_292),
.B2(n_287),
.C(n_304),
.Y(n_997)
);

NOR3xp33_ASAP7_75t_SL g998 ( 
.A(n_813),
.B(n_250),
.C(n_215),
.Y(n_998)
);

INVxp67_ASAP7_75t_SL g999 ( 
.A(n_723),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_779),
.Y(n_1000)
);

NOR2xp33_ASAP7_75t_L g1001 ( 
.A(n_702),
.B(n_651),
.Y(n_1001)
);

INVx1_ASAP7_75t_L g1002 ( 
.A(n_792),
.Y(n_1002)
);

INVx2_ASAP7_75t_L g1003 ( 
.A(n_793),
.Y(n_1003)
);

NAND2xp33_ASAP7_75t_SL g1004 ( 
.A(n_808),
.B(n_546),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_SL g1005 ( 
.A(n_743),
.B(n_523),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_798),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_799),
.Y(n_1007)
);

NAND2xp33_ASAP7_75t_L g1008 ( 
.A(n_808),
.B(n_643),
.Y(n_1008)
);

INVx2_ASAP7_75t_SL g1009 ( 
.A(n_807),
.Y(n_1009)
);

BUFx3_ASAP7_75t_L g1010 ( 
.A(n_791),
.Y(n_1010)
);

BUFx6f_ASAP7_75t_L g1011 ( 
.A(n_791),
.Y(n_1011)
);

BUFx4f_ASAP7_75t_L g1012 ( 
.A(n_829),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_683),
.B(n_651),
.Y(n_1013)
);

CKINVDCx5p33_ASAP7_75t_R g1014 ( 
.A(n_805),
.Y(n_1014)
);

A2O1A1Ixp33_ASAP7_75t_L g1015 ( 
.A1(n_722),
.A2(n_231),
.B(n_279),
.C(n_271),
.Y(n_1015)
);

INVx2_ASAP7_75t_SL g1016 ( 
.A(n_815),
.Y(n_1016)
);

INVx4_ASAP7_75t_L g1017 ( 
.A(n_688),
.Y(n_1017)
);

AOI22xp33_ASAP7_75t_L g1018 ( 
.A1(n_754),
.A2(n_643),
.B1(n_639),
.B2(n_617),
.Y(n_1018)
);

BUFx6f_ASAP7_75t_L g1019 ( 
.A(n_735),
.Y(n_1019)
);

BUFx2_ASAP7_75t_L g1020 ( 
.A(n_813),
.Y(n_1020)
);

CKINVDCx5p33_ASAP7_75t_R g1021 ( 
.A(n_830),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_763),
.B(n_651),
.Y(n_1022)
);

AND2x4_ASAP7_75t_L g1023 ( 
.A(n_750),
.B(n_653),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_800),
.Y(n_1024)
);

AND2x2_ASAP7_75t_L g1025 ( 
.A(n_920),
.B(n_712),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_995),
.Y(n_1026)
);

NAND2xp33_ASAP7_75t_L g1027 ( 
.A(n_975),
.B(n_743),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_929),
.B(n_815),
.Y(n_1028)
);

OAI22xp5_ASAP7_75t_L g1029 ( 
.A1(n_999),
.A2(n_734),
.B1(n_732),
.B2(n_708),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_869),
.B(n_754),
.Y(n_1030)
);

AOI211x1_ASAP7_75t_L g1031 ( 
.A1(n_983),
.A2(n_734),
.B(n_732),
.C(n_826),
.Y(n_1031)
);

OAI21x1_ASAP7_75t_L g1032 ( 
.A1(n_900),
.A2(n_696),
.B(n_828),
.Y(n_1032)
);

INVx2_ASAP7_75t_L g1033 ( 
.A(n_868),
.Y(n_1033)
);

INVx3_ASAP7_75t_L g1034 ( 
.A(n_995),
.Y(n_1034)
);

AND2x4_ASAP7_75t_L g1035 ( 
.A(n_955),
.B(n_819),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_990),
.B(n_958),
.Y(n_1036)
);

INVx1_ASAP7_75t_L g1037 ( 
.A(n_925),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_SL g1038 ( 
.A1(n_1005),
.A2(n_720),
.B(n_944),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_953),
.B(n_763),
.Y(n_1039)
);

AND2x4_ASAP7_75t_L g1040 ( 
.A(n_955),
.B(n_819),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_1005),
.A2(n_832),
.B(n_809),
.Y(n_1041)
);

BUFx3_ASAP7_75t_L g1042 ( 
.A(n_885),
.Y(n_1042)
);

OAI21x1_ASAP7_75t_L g1043 ( 
.A1(n_930),
.A2(n_962),
.B(n_963),
.Y(n_1043)
);

AND2x2_ASAP7_75t_L g1044 ( 
.A(n_938),
.B(n_770),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_954),
.B(n_770),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_957),
.B(n_826),
.Y(n_1046)
);

NAND2xp5_ASAP7_75t_L g1047 ( 
.A(n_970),
.B(n_720),
.Y(n_1047)
);

BUFx2_ASAP7_75t_L g1048 ( 
.A(n_851),
.Y(n_1048)
);

OR2x2_ASAP7_75t_L g1049 ( 
.A(n_943),
.B(n_724),
.Y(n_1049)
);

OAI21x1_ASAP7_75t_L g1050 ( 
.A1(n_930),
.A2(n_821),
.B(n_811),
.Y(n_1050)
);

NAND2xp5_ASAP7_75t_L g1051 ( 
.A(n_833),
.B(n_724),
.Y(n_1051)
);

AO31x2_ASAP7_75t_L g1052 ( 
.A1(n_1020),
.A2(n_703),
.A3(n_772),
.B(n_635),
.Y(n_1052)
);

AOI21xp5_ASAP7_75t_L g1053 ( 
.A1(n_992),
.A2(n_559),
.B(n_660),
.Y(n_1053)
);

INVx1_ASAP7_75t_L g1054 ( 
.A(n_925),
.Y(n_1054)
);

AND2x4_ASAP7_75t_L g1055 ( 
.A(n_848),
.B(n_653),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_840),
.B(n_619),
.Y(n_1056)
);

OAI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_914),
.A2(n_769),
.B(n_762),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_849),
.B(n_906),
.Y(n_1058)
);

NAND2xp5_ASAP7_75t_L g1059 ( 
.A(n_917),
.B(n_619),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_967),
.B(n_523),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_933),
.B(n_634),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_946),
.B(n_634),
.Y(n_1062)
);

OAI21xp5_ASAP7_75t_L g1063 ( 
.A1(n_914),
.A2(n_762),
.B(n_748),
.Y(n_1063)
);

AOI21xp5_ASAP7_75t_L g1064 ( 
.A1(n_963),
.A2(n_559),
.B(n_660),
.Y(n_1064)
);

OAI21x1_ASAP7_75t_L g1065 ( 
.A1(n_962),
.A2(n_994),
.B(n_850),
.Y(n_1065)
);

OAI21x1_ASAP7_75t_L g1066 ( 
.A1(n_994),
.A2(n_811),
.B(n_655),
.Y(n_1066)
);

HB1xp67_ASAP7_75t_L g1067 ( 
.A(n_851),
.Y(n_1067)
);

OAI21x1_ASAP7_75t_L g1068 ( 
.A1(n_850),
.A2(n_653),
.B(n_769),
.Y(n_1068)
);

NOR2x1_ASAP7_75t_L g1069 ( 
.A(n_873),
.B(n_748),
.Y(n_1069)
);

BUFx2_ASAP7_75t_R g1070 ( 
.A(n_968),
.Y(n_1070)
);

AOI21xp5_ASAP7_75t_L g1071 ( 
.A1(n_1008),
.A2(n_559),
.B(n_660),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_868),
.Y(n_1072)
);

NAND2xp5_ASAP7_75t_L g1073 ( 
.A(n_991),
.B(n_635),
.Y(n_1073)
);

OAI21x1_ASAP7_75t_L g1074 ( 
.A1(n_984),
.A2(n_804),
.B(n_803),
.Y(n_1074)
);

NAND2xp5_ASAP7_75t_SL g1075 ( 
.A(n_967),
.B(n_523),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_835),
.Y(n_1076)
);

OAI21x1_ASAP7_75t_L g1077 ( 
.A1(n_889),
.A2(n_1022),
.B(n_981),
.Y(n_1077)
);

OAI21x1_ASAP7_75t_L g1078 ( 
.A1(n_861),
.A2(n_804),
.B(n_803),
.Y(n_1078)
);

AOI221x1_ASAP7_75t_L g1079 ( 
.A1(n_1004),
.A2(n_1015),
.B1(n_852),
.B2(n_952),
.C(n_979),
.Y(n_1079)
);

OAI21xp33_ASAP7_75t_SL g1080 ( 
.A1(n_1018),
.A2(n_810),
.B(n_628),
.Y(n_1080)
);

NAND3xp33_ASAP7_75t_L g1081 ( 
.A(n_997),
.B(n_239),
.C(n_219),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_SL g1082 ( 
.A(n_1019),
.B(n_523),
.Y(n_1082)
);

OAI21x1_ASAP7_75t_L g1083 ( 
.A1(n_861),
.A2(n_810),
.B(n_639),
.Y(n_1083)
);

OAI21xp5_ASAP7_75t_L g1084 ( 
.A1(n_979),
.A2(n_645),
.B(n_727),
.Y(n_1084)
);

AND2x4_ASAP7_75t_L g1085 ( 
.A(n_848),
.B(n_550),
.Y(n_1085)
);

NAND2x1_ASAP7_75t_L g1086 ( 
.A(n_944),
.B(n_947),
.Y(n_1086)
);

AND2x2_ASAP7_75t_L g1087 ( 
.A(n_901),
.B(n_230),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_1000),
.B(n_645),
.Y(n_1088)
);

AOI221x1_ASAP7_75t_L g1089 ( 
.A1(n_1004),
.A2(n_583),
.B1(n_646),
.B2(n_641),
.C(n_571),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_888),
.A2(n_550),
.B(n_590),
.Y(n_1090)
);

INVx2_ASAP7_75t_SL g1091 ( 
.A(n_853),
.Y(n_1091)
);

BUFx12f_ASAP7_75t_L g1092 ( 
.A(n_872),
.Y(n_1092)
);

OAI21xp5_ASAP7_75t_L g1093 ( 
.A1(n_952),
.A2(n_657),
.B(n_597),
.Y(n_1093)
);

OAI22xp5_ASAP7_75t_L g1094 ( 
.A1(n_996),
.A2(n_528),
.B1(n_536),
.B2(n_342),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_838),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_993),
.A2(n_248),
.B(n_252),
.C(n_283),
.Y(n_1096)
);

BUFx2_ASAP7_75t_L g1097 ( 
.A(n_853),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_1002),
.B(n_528),
.Y(n_1098)
);

A2O1A1Ixp33_ASAP7_75t_L g1099 ( 
.A1(n_857),
.A2(n_342),
.B(n_536),
.C(n_528),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_972),
.A2(n_550),
.B(n_590),
.Y(n_1100)
);

O2A1O1Ixp5_ASAP7_75t_SL g1101 ( 
.A1(n_854),
.A2(n_195),
.B(n_296),
.C(n_11),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_1006),
.B(n_528),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_915),
.A2(n_597),
.B(n_601),
.Y(n_1103)
);

AOI21xp33_ASAP7_75t_L g1104 ( 
.A1(n_948),
.A2(n_8),
.B(n_10),
.Y(n_1104)
);

NAND2xp5_ASAP7_75t_L g1105 ( 
.A(n_1007),
.B(n_528),
.Y(n_1105)
);

NAND2xp5_ASAP7_75t_L g1106 ( 
.A(n_1019),
.B(n_536),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_959),
.A2(n_597),
.B1(n_633),
.B2(n_628),
.Y(n_1107)
);

INVx2_ASAP7_75t_L g1108 ( 
.A(n_882),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1019),
.B(n_536),
.Y(n_1109)
);

NOR4xp25_ASAP7_75t_L g1110 ( 
.A(n_983),
.B(n_195),
.C(n_296),
.D(n_13),
.Y(n_1110)
);

NAND2xp33_ASAP7_75t_L g1111 ( 
.A(n_844),
.B(n_536),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1019),
.B(n_657),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_1003),
.B(n_657),
.Y(n_1113)
);

BUFx12f_ASAP7_75t_L g1114 ( 
.A(n_872),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_890),
.A2(n_590),
.B(n_601),
.Y(n_1115)
);

AO31x2_ASAP7_75t_L g1116 ( 
.A1(n_1015),
.A2(n_601),
.A3(n_609),
.B(n_628),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_SL g1117 ( 
.A1(n_1009),
.A2(n_1017),
.B(n_1016),
.Y(n_1117)
);

AO31x2_ASAP7_75t_L g1118 ( 
.A1(n_1017),
.A2(n_1001),
.A3(n_904),
.B(n_960),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_SL g1119 ( 
.A(n_876),
.B(n_646),
.Y(n_1119)
);

AND2x2_ASAP7_75t_L g1120 ( 
.A(n_875),
.B(n_296),
.Y(n_1120)
);

BUFx2_ASAP7_75t_L g1121 ( 
.A(n_856),
.Y(n_1121)
);

OAI21x1_ASAP7_75t_L g1122 ( 
.A1(n_923),
.A2(n_590),
.B(n_609),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1003),
.B(n_609),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_937),
.A2(n_633),
.B(n_641),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_857),
.A2(n_633),
.B1(n_641),
.B2(n_646),
.Y(n_1125)
);

NAND2xp5_ASAP7_75t_L g1126 ( 
.A(n_1024),
.B(n_841),
.Y(n_1126)
);

AND2x4_ASAP7_75t_L g1127 ( 
.A(n_860),
.B(n_646),
.Y(n_1127)
);

HB1xp67_ASAP7_75t_L g1128 ( 
.A(n_837),
.Y(n_1128)
);

AOI21xp5_ASAP7_75t_L g1129 ( 
.A1(n_941),
.A2(n_646),
.B(n_641),
.Y(n_1129)
);

OAI21x1_ASAP7_75t_SL g1130 ( 
.A1(n_879),
.A2(n_168),
.B(n_151),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_L g1131 ( 
.A(n_1024),
.B(n_641),
.Y(n_1131)
);

OAI21x1_ASAP7_75t_L g1132 ( 
.A1(n_897),
.A2(n_610),
.B(n_608),
.Y(n_1132)
);

HB1xp67_ASAP7_75t_L g1133 ( 
.A(n_837),
.Y(n_1133)
);

AOI21xp5_ASAP7_75t_L g1134 ( 
.A1(n_944),
.A2(n_610),
.B(n_608),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_859),
.B(n_610),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_897),
.A2(n_610),
.B(n_608),
.Y(n_1136)
);

INVx1_ASAP7_75t_L g1137 ( 
.A(n_865),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_866),
.B(n_610),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_SL g1139 ( 
.A(n_876),
.B(n_608),
.Y(n_1139)
);

OR2x6_ASAP7_75t_L g1140 ( 
.A(n_883),
.B(n_608),
.Y(n_1140)
);

OAI21x1_ASAP7_75t_L g1141 ( 
.A1(n_855),
.A2(n_583),
.B(n_571),
.Y(n_1141)
);

OAI21x1_ASAP7_75t_L g1142 ( 
.A1(n_855),
.A2(n_583),
.B(n_571),
.Y(n_1142)
);

INVxp67_ASAP7_75t_SL g1143 ( 
.A(n_844),
.Y(n_1143)
);

OAI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1001),
.A2(n_577),
.B(n_583),
.Y(n_1144)
);

AOI21xp5_ASAP7_75t_L g1145 ( 
.A1(n_944),
.A2(n_583),
.B(n_571),
.Y(n_1145)
);

OAI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_1018),
.A2(n_577),
.B(n_571),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_867),
.B(n_555),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_SL g1148 ( 
.A(n_909),
.B(n_10),
.C(n_12),
.Y(n_1148)
);

NOR2xp33_ASAP7_75t_L g1149 ( 
.A(n_959),
.B(n_12),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_874),
.B(n_555),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_864),
.A2(n_555),
.B(n_546),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_886),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_882),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_856),
.Y(n_1154)
);

AO31x2_ASAP7_75t_L g1155 ( 
.A1(n_834),
.A2(n_14),
.A3(n_15),
.B(n_16),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_947),
.A2(n_555),
.B(n_546),
.Y(n_1156)
);

OAI21x1_ASAP7_75t_L g1157 ( 
.A1(n_864),
.A2(n_555),
.B(n_546),
.Y(n_1157)
);

OAI21x1_ASAP7_75t_SL g1158 ( 
.A1(n_895),
.A2(n_150),
.B(n_149),
.Y(n_1158)
);

NAND3xp33_ASAP7_75t_L g1159 ( 
.A(n_926),
.B(n_577),
.C(n_17),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_893),
.B(n_577),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_887),
.A2(n_577),
.B(n_110),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_899),
.B(n_14),
.Y(n_1162)
);

AOI21x1_ASAP7_75t_L g1163 ( 
.A1(n_982),
.A2(n_400),
.B(n_145),
.Y(n_1163)
);

AND2x2_ASAP7_75t_L g1164 ( 
.A(n_940),
.B(n_17),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_903),
.B(n_20),
.Y(n_1165)
);

AOI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_947),
.A2(n_144),
.B(n_134),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_918),
.B(n_21),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_887),
.A2(n_131),
.B(n_116),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_918),
.B(n_24),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_876),
.B(n_107),
.Y(n_1170)
);

INVx3_ASAP7_75t_L g1171 ( 
.A(n_947),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_905),
.B(n_25),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_SL g1173 ( 
.A1(n_839),
.A2(n_99),
.B(n_98),
.Y(n_1173)
);

INVx2_ASAP7_75t_L g1174 ( 
.A(n_891),
.Y(n_1174)
);

AOI31xp67_ASAP7_75t_L g1175 ( 
.A1(n_854),
.A2(n_902),
.A3(n_891),
.B(n_980),
.Y(n_1175)
);

AO21x2_ASAP7_75t_L g1176 ( 
.A1(n_985),
.A2(n_987),
.B(n_965),
.Y(n_1176)
);

OAI21xp5_ASAP7_75t_L g1177 ( 
.A1(n_1013),
.A2(n_94),
.B(n_75),
.Y(n_1177)
);

OAI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1013),
.A2(n_68),
.B(n_26),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_852),
.A2(n_25),
.B(n_27),
.C(n_28),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_902),
.A2(n_27),
.B(n_30),
.Y(n_1180)
);

INVx4_ASAP7_75t_L g1181 ( 
.A(n_844),
.Y(n_1181)
);

OAI21xp33_ASAP7_75t_L g1182 ( 
.A1(n_1021),
.A2(n_30),
.B(n_31),
.Y(n_1182)
);

HB1xp67_ASAP7_75t_L g1183 ( 
.A(n_842),
.Y(n_1183)
);

INVx2_ASAP7_75t_SL g1184 ( 
.A(n_842),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_912),
.B(n_36),
.Y(n_1185)
);

AND2x2_ASAP7_75t_L g1186 ( 
.A(n_1030),
.B(n_878),
.Y(n_1186)
);

AOI21x1_ASAP7_75t_L g1187 ( 
.A1(n_1089),
.A2(n_974),
.B(n_988),
.Y(n_1187)
);

OAI21xp5_ASAP7_75t_L g1188 ( 
.A1(n_1028),
.A2(n_932),
.B(n_1023),
.Y(n_1188)
);

OAI21x1_ASAP7_75t_L g1189 ( 
.A1(n_1124),
.A2(n_908),
.B(n_910),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1076),
.Y(n_1190)
);

OAI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_1028),
.A2(n_1023),
.B(n_982),
.Y(n_1191)
);

OAI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1036),
.A2(n_969),
.B(n_912),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_1095),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_1092),
.Y(n_1194)
);

INVxp67_ASAP7_75t_L g1195 ( 
.A(n_1048),
.Y(n_1195)
);

NAND2xp5_ASAP7_75t_L g1196 ( 
.A(n_1058),
.B(n_989),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_SL g1197 ( 
.A1(n_1173),
.A2(n_921),
.B(n_881),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1137),
.Y(n_1198)
);

OA21x2_ASAP7_75t_L g1199 ( 
.A1(n_1079),
.A2(n_910),
.B(n_927),
.Y(n_1199)
);

BUFx8_ASAP7_75t_L g1200 ( 
.A(n_1092),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_1124),
.A2(n_908),
.B(n_934),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1115),
.A2(n_966),
.B(n_934),
.Y(n_1202)
);

NAND2xp5_ASAP7_75t_L g1203 ( 
.A(n_1044),
.B(n_907),
.Y(n_1203)
);

OAI21x1_ASAP7_75t_L g1204 ( 
.A1(n_1115),
.A2(n_927),
.B(n_966),
.Y(n_1204)
);

OA21x2_ASAP7_75t_L g1205 ( 
.A1(n_1077),
.A2(n_980),
.B(n_964),
.Y(n_1205)
);

AND2x2_ASAP7_75t_L g1206 ( 
.A(n_1025),
.B(n_1045),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1152),
.Y(n_1207)
);

OR2x2_ASAP7_75t_L g1208 ( 
.A(n_1121),
.B(n_878),
.Y(n_1208)
);

OAI21x1_ASAP7_75t_L g1209 ( 
.A1(n_1141),
.A2(n_913),
.B(n_964),
.Y(n_1209)
);

AOI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1027),
.A2(n_1014),
.B1(n_884),
.B2(n_856),
.Y(n_1210)
);

INVx5_ASAP7_75t_L g1211 ( 
.A(n_1140),
.Y(n_1211)
);

INVx4_ASAP7_75t_L g1212 ( 
.A(n_1181),
.Y(n_1212)
);

AOI22xp33_ASAP7_75t_L g1213 ( 
.A1(n_1027),
.A2(n_1104),
.B1(n_1182),
.B2(n_1148),
.Y(n_1213)
);

AND2x4_ASAP7_75t_L g1214 ( 
.A(n_1055),
.B(n_860),
.Y(n_1214)
);

OAI22xp5_ASAP7_75t_L g1215 ( 
.A1(n_1039),
.A2(n_1126),
.B1(n_1046),
.B2(n_1049),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_1141),
.A2(n_913),
.B(n_843),
.Y(n_1216)
);

CKINVDCx10_ASAP7_75t_R g1217 ( 
.A(n_1070),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1093),
.A2(n_876),
.B(n_971),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_1114),
.Y(n_1219)
);

INVx2_ASAP7_75t_SL g1220 ( 
.A(n_1128),
.Y(n_1220)
);

OAI21x1_ASAP7_75t_L g1221 ( 
.A1(n_1142),
.A2(n_843),
.B(n_846),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1033),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1178),
.A2(n_1159),
.B1(n_1149),
.B2(n_1164),
.Y(n_1223)
);

OA21x2_ASAP7_75t_L g1224 ( 
.A1(n_1077),
.A2(n_978),
.B(n_977),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_1114),
.Y(n_1225)
);

INVx6_ASAP7_75t_L g1226 ( 
.A(n_1181),
.Y(n_1226)
);

INVx2_ASAP7_75t_SL g1227 ( 
.A(n_1133),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_1142),
.A2(n_846),
.B(n_922),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1072),
.Y(n_1229)
);

NAND3xp33_ASAP7_75t_L g1230 ( 
.A(n_1081),
.B(n_870),
.C(n_911),
.Y(n_1230)
);

AO21x2_ASAP7_75t_L g1231 ( 
.A1(n_1144),
.A2(n_1117),
.B(n_1084),
.Y(n_1231)
);

HB1xp67_ASAP7_75t_L g1232 ( 
.A(n_1097),
.Y(n_1232)
);

AND2x2_ASAP7_75t_L g1233 ( 
.A(n_1118),
.B(n_969),
.Y(n_1233)
);

NOR2xp67_ASAP7_75t_L g1234 ( 
.A(n_1183),
.B(n_885),
.Y(n_1234)
);

OAI21xp5_ASAP7_75t_L g1235 ( 
.A1(n_1051),
.A2(n_969),
.B(n_912),
.Y(n_1235)
);

OAI21x1_ASAP7_75t_L g1236 ( 
.A1(n_1151),
.A2(n_892),
.B(n_939),
.Y(n_1236)
);

AND2x2_ASAP7_75t_L g1237 ( 
.A(n_1087),
.B(n_898),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1108),
.Y(n_1238)
);

NAND2x1p5_ASAP7_75t_L g1239 ( 
.A(n_1086),
.B(n_881),
.Y(n_1239)
);

OAI21xp5_ASAP7_75t_L g1240 ( 
.A1(n_1099),
.A2(n_1013),
.B(n_971),
.Y(n_1240)
);

AOI22xp33_ASAP7_75t_L g1241 ( 
.A1(n_1149),
.A2(n_965),
.B1(n_1012),
.B2(n_976),
.Y(n_1241)
);

INVx2_ASAP7_75t_L g1242 ( 
.A(n_1153),
.Y(n_1242)
);

NOR2xp67_ASAP7_75t_L g1243 ( 
.A(n_1184),
.B(n_939),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1151),
.A2(n_1157),
.B(n_1122),
.Y(n_1244)
);

AOI22xp33_ASAP7_75t_L g1245 ( 
.A1(n_1177),
.A2(n_1012),
.B1(n_976),
.B2(n_956),
.Y(n_1245)
);

AO21x1_ASAP7_75t_L g1246 ( 
.A1(n_1029),
.A2(n_950),
.B(n_931),
.Y(n_1246)
);

A2O1A1Ixp33_ASAP7_75t_L g1247 ( 
.A1(n_1179),
.A2(n_986),
.B(n_998),
.C(n_836),
.Y(n_1247)
);

NAND3x1_ASAP7_75t_L g1248 ( 
.A(n_1069),
.B(n_949),
.C(n_961),
.Y(n_1248)
);

O2A1O1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1096),
.A2(n_924),
.B(n_858),
.C(n_894),
.Y(n_1249)
);

OAI21x1_ASAP7_75t_L g1250 ( 
.A1(n_1157),
.A2(n_1122),
.B(n_1132),
.Y(n_1250)
);

OA21x2_ASAP7_75t_L g1251 ( 
.A1(n_1032),
.A2(n_950),
.B(n_985),
.Y(n_1251)
);

INVx2_ASAP7_75t_L g1252 ( 
.A(n_1174),
.Y(n_1252)
);

INVx1_ASAP7_75t_L g1253 ( 
.A(n_1037),
.Y(n_1253)
);

AO21x2_ASAP7_75t_L g1254 ( 
.A1(n_1099),
.A2(n_950),
.B(n_919),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1154),
.B(n_916),
.Y(n_1255)
);

OAI21x1_ASAP7_75t_L g1256 ( 
.A1(n_1132),
.A2(n_1011),
.B(n_973),
.Y(n_1256)
);

OA21x2_ASAP7_75t_L g1257 ( 
.A1(n_1032),
.A2(n_936),
.B(n_951),
.Y(n_1257)
);

INVx1_ASAP7_75t_SL g1258 ( 
.A(n_1067),
.Y(n_1258)
);

OAI22xp33_ASAP7_75t_L g1259 ( 
.A1(n_1167),
.A2(n_877),
.B1(n_845),
.B2(n_956),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1175),
.Y(n_1260)
);

NOR2x1_ASAP7_75t_SL g1261 ( 
.A(n_1140),
.B(n_863),
.Y(n_1261)
);

NAND2x1p5_ASAP7_75t_L g1262 ( 
.A(n_1181),
.B(n_863),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1054),
.Y(n_1263)
);

AOI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1120),
.A2(n_896),
.B1(n_931),
.B2(n_871),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1136),
.A2(n_1011),
.B(n_973),
.Y(n_1265)
);

OAI21x1_ASAP7_75t_L g1266 ( 
.A1(n_1136),
.A2(n_1011),
.B(n_973),
.Y(n_1266)
);

INVx3_ASAP7_75t_L g1267 ( 
.A(n_1026),
.Y(n_1267)
);

AND2x2_ASAP7_75t_L g1268 ( 
.A(n_1091),
.B(n_862),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_L g1269 ( 
.A1(n_1169),
.A2(n_877),
.B1(n_871),
.B2(n_945),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1059),
.Y(n_1270)
);

INVx5_ASAP7_75t_L g1271 ( 
.A(n_1140),
.Y(n_1271)
);

NAND2x1p5_ASAP7_75t_L g1272 ( 
.A(n_1171),
.B(n_863),
.Y(n_1272)
);

OA21x2_ASAP7_75t_L g1273 ( 
.A1(n_1041),
.A2(n_1011),
.B(n_1010),
.Y(n_1273)
);

OR2x2_ASAP7_75t_L g1274 ( 
.A(n_1091),
.B(n_871),
.Y(n_1274)
);

AOI21xp5_ASAP7_75t_SL g1275 ( 
.A1(n_1146),
.A2(n_844),
.B(n_847),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1061),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1062),
.Y(n_1277)
);

INVx2_ASAP7_75t_L g1278 ( 
.A(n_1073),
.Y(n_1278)
);

NOR2xp33_ASAP7_75t_L g1279 ( 
.A(n_1184),
.B(n_862),
.Y(n_1279)
);

NOR2xp33_ASAP7_75t_L g1280 ( 
.A(n_1047),
.B(n_968),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_1179),
.A2(n_945),
.B(n_1010),
.C(n_896),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1042),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1161),
.A2(n_973),
.B(n_847),
.Y(n_1283)
);

BUFx2_ASAP7_75t_L g1284 ( 
.A(n_1055),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1088),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1071),
.A2(n_847),
.B(n_863),
.Y(n_1286)
);

OAI22xp5_ASAP7_75t_L g1287 ( 
.A1(n_1026),
.A2(n_847),
.B1(n_928),
.B2(n_880),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1127),
.Y(n_1288)
);

OAI21x1_ASAP7_75t_SL g1289 ( 
.A1(n_1158),
.A2(n_883),
.B(n_880),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1131),
.Y(n_1290)
);

AO21x2_ASAP7_75t_L g1291 ( 
.A1(n_1053),
.A2(n_1057),
.B(n_1063),
.Y(n_1291)
);

AO32x2_ASAP7_75t_L g1292 ( 
.A1(n_1031),
.A2(n_961),
.A3(n_928),
.B1(n_880),
.B2(n_919),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1162),
.A2(n_877),
.B1(n_928),
.B2(n_880),
.Y(n_1293)
);

NAND2x1p5_ASAP7_75t_L g1294 ( 
.A(n_1171),
.B(n_928),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1185),
.Y(n_1295)
);

NOR2xp67_ASAP7_75t_L g1296 ( 
.A(n_1165),
.B(n_935),
.Y(n_1296)
);

AND2x2_ASAP7_75t_L g1297 ( 
.A(n_1096),
.B(n_1110),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1172),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1118),
.B(n_1056),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1161),
.A2(n_1066),
.B(n_1068),
.Y(n_1300)
);

INVx6_ASAP7_75t_L g1301 ( 
.A(n_1085),
.Y(n_1301)
);

OAI221xp5_ASAP7_75t_L g1302 ( 
.A1(n_1042),
.A2(n_935),
.B1(n_942),
.B2(n_883),
.C(n_44),
.Y(n_1302)
);

NAND2x1p5_ASAP7_75t_L g1303 ( 
.A(n_1171),
.B(n_37),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1127),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1041),
.A2(n_1180),
.B(n_1068),
.Y(n_1305)
);

OA21x2_ASAP7_75t_L g1306 ( 
.A1(n_1180),
.A2(n_1065),
.B(n_1168),
.Y(n_1306)
);

AND2x4_ASAP7_75t_L g1307 ( 
.A(n_1055),
.B(n_40),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1065),
.Y(n_1308)
);

AO21x2_ASAP7_75t_L g1309 ( 
.A1(n_1038),
.A2(n_41),
.B(n_48),
.Y(n_1309)
);

OAI21x1_ASAP7_75t_L g1310 ( 
.A1(n_1066),
.A2(n_48),
.B(n_49),
.Y(n_1310)
);

NAND2xp5_ASAP7_75t_L g1311 ( 
.A(n_1118),
.B(n_63),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1035),
.A2(n_1040),
.B1(n_1176),
.B2(n_1130),
.Y(n_1312)
);

NOR2x1_ASAP7_75t_R g1313 ( 
.A(n_1035),
.B(n_1040),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_1135),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1118),
.B(n_63),
.Y(n_1315)
);

OAI21x1_ASAP7_75t_L g1316 ( 
.A1(n_1090),
.A2(n_52),
.B(n_54),
.Y(n_1316)
);

OAI21xp5_ASAP7_75t_L g1317 ( 
.A1(n_1080),
.A2(n_56),
.B(n_57),
.Y(n_1317)
);

AOI22xp33_ASAP7_75t_L g1318 ( 
.A1(n_1035),
.A2(n_58),
.B1(n_62),
.B2(n_1040),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1043),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1112),
.B(n_1123),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_1085),
.Y(n_1321)
);

AOI22x1_ASAP7_75t_L g1322 ( 
.A1(n_1129),
.A2(n_1064),
.B1(n_1103),
.B2(n_1166),
.Y(n_1322)
);

OAI22xp5_ASAP7_75t_L g1323 ( 
.A1(n_1026),
.A2(n_1034),
.B1(n_1060),
.B2(n_1075),
.Y(n_1323)
);

INVx1_ASAP7_75t_L g1324 ( 
.A(n_1138),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1090),
.A2(n_1050),
.B(n_1043),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1176),
.A2(n_1170),
.B1(n_1075),
.B2(n_1060),
.Y(n_1326)
);

OAI21x1_ASAP7_75t_L g1327 ( 
.A1(n_1050),
.A2(n_1083),
.B(n_1168),
.Y(n_1327)
);

AO21x2_ASAP7_75t_L g1328 ( 
.A1(n_1163),
.A2(n_1082),
.B(n_1074),
.Y(n_1328)
);

OR2x6_ASAP7_75t_L g1329 ( 
.A(n_1034),
.B(n_1082),
.Y(n_1329)
);

AO31x2_ASAP7_75t_L g1330 ( 
.A1(n_1125),
.A2(n_1102),
.A3(n_1098),
.B(n_1105),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1147),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1034),
.A2(n_1143),
.B1(n_1127),
.B2(n_1113),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_1085),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1150),
.Y(n_1334)
);

INVx2_ASAP7_75t_L g1335 ( 
.A(n_1083),
.Y(n_1335)
);

INVx2_ASAP7_75t_SL g1336 ( 
.A(n_1106),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1155),
.Y(n_1337)
);

NOR2xp33_ASAP7_75t_L g1338 ( 
.A(n_1109),
.B(n_1139),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1052),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1155),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1155),
.Y(n_1341)
);

INVx1_ASAP7_75t_SL g1342 ( 
.A(n_1170),
.Y(n_1342)
);

O2A1O1Ixp5_ASAP7_75t_L g1343 ( 
.A1(n_1119),
.A2(n_1139),
.B(n_1160),
.C(n_1094),
.Y(n_1343)
);

OR2x2_ASAP7_75t_L g1344 ( 
.A(n_1052),
.B(n_1116),
.Y(n_1344)
);

AND2x4_ASAP7_75t_L g1345 ( 
.A(n_1119),
.B(n_1052),
.Y(n_1345)
);

OR2x2_ASAP7_75t_L g1346 ( 
.A(n_1052),
.B(n_1116),
.Y(n_1346)
);

AOI22xp5_ASAP7_75t_L g1347 ( 
.A1(n_1280),
.A2(n_1111),
.B1(n_1107),
.B2(n_1078),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1206),
.B(n_1101),
.Y(n_1348)
);

OR2x2_ASAP7_75t_L g1349 ( 
.A(n_1203),
.B(n_1116),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1213),
.A2(n_1078),
.B1(n_1074),
.B2(n_1111),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_SL g1351 ( 
.A1(n_1302),
.A2(n_1156),
.B1(n_1134),
.B2(n_1145),
.Y(n_1351)
);

BUFx2_ASAP7_75t_L g1352 ( 
.A(n_1255),
.Y(n_1352)
);

NOR2x1_ASAP7_75t_L g1353 ( 
.A(n_1196),
.B(n_1116),
.Y(n_1353)
);

INVx1_ASAP7_75t_L g1354 ( 
.A(n_1190),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1206),
.B(n_1100),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_L g1356 ( 
.A1(n_1213),
.A2(n_1100),
.B1(n_1297),
.B2(n_1223),
.Y(n_1356)
);

INVx2_ASAP7_75t_L g1357 ( 
.A(n_1238),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1214),
.B(n_1304),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1223),
.A2(n_1186),
.B1(n_1230),
.B2(n_1318),
.Y(n_1359)
);

AND2x6_ASAP7_75t_L g1360 ( 
.A(n_1345),
.B(n_1342),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_1242),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1318),
.A2(n_1241),
.B1(n_1210),
.B2(n_1317),
.Y(n_1362)
);

AOI22xp33_ASAP7_75t_L g1363 ( 
.A1(n_1241),
.A2(n_1188),
.B1(n_1298),
.B2(n_1245),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1215),
.B(n_1270),
.Y(n_1364)
);

INVx1_ASAP7_75t_L g1365 ( 
.A(n_1193),
.Y(n_1365)
);

NAND2xp5_ASAP7_75t_SL g1366 ( 
.A(n_1249),
.B(n_1259),
.Y(n_1366)
);

OAI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1208),
.A2(n_1264),
.B1(n_1295),
.B2(n_1280),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1214),
.B(n_1304),
.Y(n_1368)
);

AND2x2_ASAP7_75t_SL g1369 ( 
.A(n_1245),
.B(n_1293),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1198),
.Y(n_1370)
);

OAI22xp5_ASAP7_75t_L g1371 ( 
.A1(n_1275),
.A2(n_1247),
.B1(n_1207),
.B2(n_1281),
.Y(n_1371)
);

OAI22xp5_ASAP7_75t_L g1372 ( 
.A1(n_1247),
.A2(n_1281),
.B1(n_1293),
.B2(n_1333),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1252),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1253),
.Y(n_1374)
);

AOI22xp33_ASAP7_75t_L g1375 ( 
.A1(n_1191),
.A2(n_1237),
.B1(n_1269),
.B2(n_1309),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1252),
.Y(n_1376)
);

INVxp67_ASAP7_75t_SL g1377 ( 
.A(n_1232),
.Y(n_1377)
);

CKINVDCx5p33_ASAP7_75t_R g1378 ( 
.A(n_1217),
.Y(n_1378)
);

NAND2xp5_ASAP7_75t_L g1379 ( 
.A(n_1270),
.B(n_1278),
.Y(n_1379)
);

OAI22xp5_ASAP7_75t_L g1380 ( 
.A1(n_1333),
.A2(n_1271),
.B1(n_1211),
.B2(n_1263),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1276),
.B(n_1277),
.Y(n_1381)
);

AOI221xp5_ASAP7_75t_L g1382 ( 
.A1(n_1311),
.A2(n_1315),
.B1(n_1195),
.B2(n_1258),
.C(n_1220),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1307),
.B(n_1284),
.Y(n_1383)
);

BUFx3_ASAP7_75t_L g1384 ( 
.A(n_1282),
.Y(n_1384)
);

BUFx4f_ASAP7_75t_L g1385 ( 
.A(n_1194),
.Y(n_1385)
);

BUFx3_ASAP7_75t_L g1386 ( 
.A(n_1282),
.Y(n_1386)
);

OAI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1296),
.A2(n_1274),
.B1(n_1243),
.B2(n_1234),
.Y(n_1387)
);

NOR3xp33_ASAP7_75t_SL g1388 ( 
.A(n_1219),
.B(n_1225),
.C(n_1279),
.Y(n_1388)
);

BUFx6f_ASAP7_75t_L g1389 ( 
.A(n_1321),
.Y(n_1389)
);

INVx3_ASAP7_75t_L g1390 ( 
.A(n_1321),
.Y(n_1390)
);

OAI222xp33_ASAP7_75t_L g1391 ( 
.A1(n_1303),
.A2(n_1307),
.B1(n_1285),
.B2(n_1220),
.C1(n_1227),
.C2(n_1312),
.Y(n_1391)
);

INVx1_ASAP7_75t_L g1392 ( 
.A(n_1222),
.Y(n_1392)
);

OR2x6_ASAP7_75t_L g1393 ( 
.A(n_1289),
.B(n_1218),
.Y(n_1393)
);

INVx4_ASAP7_75t_L g1394 ( 
.A(n_1211),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1278),
.B(n_1227),
.Y(n_1395)
);

NAND2xp5_ASAP7_75t_L g1396 ( 
.A(n_1290),
.B(n_1336),
.Y(n_1396)
);

OAI22xp5_ASAP7_75t_L g1397 ( 
.A1(n_1211),
.A2(n_1271),
.B1(n_1307),
.B2(n_1299),
.Y(n_1397)
);

CKINVDCx5p33_ASAP7_75t_R g1398 ( 
.A(n_1200),
.Y(n_1398)
);

AND2x4_ASAP7_75t_L g1399 ( 
.A(n_1214),
.B(n_1268),
.Y(n_1399)
);

AOI22xp5_ASAP7_75t_L g1400 ( 
.A1(n_1248),
.A2(n_1312),
.B1(n_1279),
.B2(n_1254),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1229),
.Y(n_1401)
);

BUFx6f_ASAP7_75t_L g1402 ( 
.A(n_1321),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1321),
.Y(n_1403)
);

BUFx6f_ASAP7_75t_L g1404 ( 
.A(n_1301),
.Y(n_1404)
);

AND2x4_ASAP7_75t_L g1405 ( 
.A(n_1288),
.B(n_1211),
.Y(n_1405)
);

NAND3xp33_ASAP7_75t_L g1406 ( 
.A(n_1192),
.B(n_1240),
.C(n_1326),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1290),
.B(n_1336),
.Y(n_1407)
);

INVx4_ASAP7_75t_L g1408 ( 
.A(n_1271),
.Y(n_1408)
);

NOR2x1_ASAP7_75t_SL g1409 ( 
.A(n_1271),
.B(n_1329),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_1200),
.Y(n_1410)
);

CKINVDCx5p33_ASAP7_75t_R g1411 ( 
.A(n_1200),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1233),
.B(n_1301),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1286),
.A2(n_1320),
.B(n_1291),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1334),
.B(n_1314),
.Y(n_1414)
);

NOR3xp33_ASAP7_75t_SL g1415 ( 
.A(n_1219),
.B(n_1225),
.C(n_1338),
.Y(n_1415)
);

OAI22xp33_ASAP7_75t_L g1416 ( 
.A1(n_1303),
.A2(n_1194),
.B1(n_1235),
.B2(n_1288),
.Y(n_1416)
);

INVx1_ASAP7_75t_SL g1417 ( 
.A(n_1301),
.Y(n_1417)
);

INVx2_ASAP7_75t_SL g1418 ( 
.A(n_1226),
.Y(n_1418)
);

OAI22xp5_ASAP7_75t_L g1419 ( 
.A1(n_1326),
.A2(n_1248),
.B1(n_1331),
.B2(n_1324),
.Y(n_1419)
);

AOI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1309),
.A2(n_1233),
.B1(n_1254),
.B2(n_1246),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1339),
.A2(n_1340),
.B1(n_1337),
.B2(n_1341),
.Y(n_1421)
);

AOI22xp33_ASAP7_75t_SL g1422 ( 
.A1(n_1261),
.A2(n_1322),
.B1(n_1197),
.B2(n_1338),
.Y(n_1422)
);

CKINVDCx11_ASAP7_75t_R g1423 ( 
.A(n_1212),
.Y(n_1423)
);

AND2x4_ASAP7_75t_L g1424 ( 
.A(n_1212),
.B(n_1236),
.Y(n_1424)
);

INVxp33_ASAP7_75t_SL g1425 ( 
.A(n_1313),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1345),
.B(n_1226),
.Y(n_1426)
);

INVx2_ASAP7_75t_SL g1427 ( 
.A(n_1226),
.Y(n_1427)
);

BUFx6f_ASAP7_75t_L g1428 ( 
.A(n_1262),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1236),
.B(n_1292),
.Y(n_1429)
);

OAI21xp5_ASAP7_75t_L g1430 ( 
.A1(n_1343),
.A2(n_1323),
.B(n_1345),
.Y(n_1430)
);

OR2x2_ASAP7_75t_L g1431 ( 
.A(n_1272),
.B(n_1294),
.Y(n_1431)
);

AOI21xp5_ASAP7_75t_L g1432 ( 
.A1(n_1291),
.A2(n_1231),
.B(n_1266),
.Y(n_1432)
);

NAND3xp33_ASAP7_75t_SL g1433 ( 
.A(n_1239),
.B(n_1332),
.C(n_1262),
.Y(n_1433)
);

AND2x2_ASAP7_75t_L g1434 ( 
.A(n_1292),
.B(n_1339),
.Y(n_1434)
);

OR2x2_ASAP7_75t_L g1435 ( 
.A(n_1344),
.B(n_1346),
.Y(n_1435)
);

AOI21xp5_ASAP7_75t_L g1436 ( 
.A1(n_1231),
.A2(n_1265),
.B(n_1256),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1212),
.B(n_1267),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1199),
.Y(n_1438)
);

INVx4_ASAP7_75t_L g1439 ( 
.A(n_1267),
.Y(n_1439)
);

OR2x6_ASAP7_75t_L g1440 ( 
.A(n_1329),
.B(n_1239),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1199),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1187),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1310),
.Y(n_1443)
);

CKINVDCx16_ASAP7_75t_R g1444 ( 
.A(n_1329),
.Y(n_1444)
);

BUFx4f_ASAP7_75t_SL g1445 ( 
.A(n_1267),
.Y(n_1445)
);

AND2x2_ASAP7_75t_L g1446 ( 
.A(n_1292),
.B(n_1310),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1287),
.B(n_1330),
.Y(n_1447)
);

OR2x6_ASAP7_75t_L g1448 ( 
.A(n_1256),
.B(n_1265),
.Y(n_1448)
);

CKINVDCx8_ASAP7_75t_R g1449 ( 
.A(n_1273),
.Y(n_1449)
);

AND2x2_ASAP7_75t_L g1450 ( 
.A(n_1292),
.B(n_1316),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1273),
.Y(n_1451)
);

OAI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1308),
.A2(n_1273),
.B1(n_1319),
.B2(n_1335),
.Y(n_1452)
);

OAI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1308),
.A2(n_1319),
.B1(n_1257),
.B2(n_1224),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1283),
.A2(n_1327),
.B(n_1244),
.Y(n_1454)
);

AND2x4_ASAP7_75t_L g1455 ( 
.A(n_1266),
.B(n_1221),
.Y(n_1455)
);

OR2x2_ASAP7_75t_L g1456 ( 
.A(n_1330),
.B(n_1224),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1257),
.A2(n_1224),
.B1(n_1205),
.B2(n_1306),
.Y(n_1457)
);

INVx2_ASAP7_75t_L g1458 ( 
.A(n_1205),
.Y(n_1458)
);

AOI221xp5_ASAP7_75t_L g1459 ( 
.A1(n_1260),
.A2(n_1328),
.B1(n_1330),
.B2(n_1316),
.C(n_1205),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1251),
.A2(n_1257),
.B1(n_1306),
.B2(n_1305),
.Y(n_1460)
);

AND2x4_ASAP7_75t_L g1461 ( 
.A(n_1221),
.B(n_1228),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1251),
.A2(n_1306),
.B1(n_1305),
.B2(n_1330),
.Y(n_1462)
);

NOR2x1_ASAP7_75t_SL g1463 ( 
.A(n_1328),
.B(n_1228),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1209),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1283),
.A2(n_1327),
.B(n_1244),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1209),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1305),
.B(n_1251),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1189),
.Y(n_1468)
);

NAND2x1p5_ASAP7_75t_L g1469 ( 
.A(n_1216),
.B(n_1201),
.Y(n_1469)
);

NAND2xp5_ASAP7_75t_L g1470 ( 
.A(n_1201),
.B(n_1202),
.Y(n_1470)
);

OAI221xp5_ASAP7_75t_L g1471 ( 
.A1(n_1202),
.A2(n_1204),
.B1(n_1300),
.B2(n_1325),
.C(n_1216),
.Y(n_1471)
);

NAND2xp33_ASAP7_75t_L g1472 ( 
.A(n_1300),
.B(n_1204),
.Y(n_1472)
);

AOI22xp33_ASAP7_75t_SL g1473 ( 
.A1(n_1250),
.A2(n_675),
.B1(n_967),
.B2(n_674),
.Y(n_1473)
);

AOI222xp33_ASAP7_75t_L g1474 ( 
.A1(n_1250),
.A2(n_929),
.B1(n_675),
.B2(n_1182),
.C1(n_674),
.C2(n_997),
.Y(n_1474)
);

INVx2_ASAP7_75t_SL g1475 ( 
.A(n_1255),
.Y(n_1475)
);

INVx4_ASAP7_75t_L g1476 ( 
.A(n_1211),
.Y(n_1476)
);

BUFx2_ASAP7_75t_L g1477 ( 
.A(n_1255),
.Y(n_1477)
);

OAI21xp5_ASAP7_75t_L g1478 ( 
.A1(n_1317),
.A2(n_1028),
.B(n_675),
.Y(n_1478)
);

HB1xp67_ASAP7_75t_L g1479 ( 
.A(n_1232),
.Y(n_1479)
);

AND2x2_ASAP7_75t_L g1480 ( 
.A(n_1186),
.B(n_1206),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1186),
.B(n_1206),
.Y(n_1481)
);

AND2x4_ASAP7_75t_L g1482 ( 
.A(n_1214),
.B(n_1304),
.Y(n_1482)
);

INVx1_ASAP7_75t_L g1483 ( 
.A(n_1190),
.Y(n_1483)
);

OAI22xp5_ASAP7_75t_L g1484 ( 
.A1(n_1318),
.A2(n_675),
.B1(n_975),
.B2(n_1213),
.Y(n_1484)
);

AOI22xp33_ASAP7_75t_SL g1485 ( 
.A1(n_1302),
.A2(n_675),
.B1(n_967),
.B2(n_674),
.Y(n_1485)
);

AOI22xp5_ASAP7_75t_L g1486 ( 
.A1(n_1280),
.A2(n_675),
.B1(n_929),
.B2(n_674),
.Y(n_1486)
);

O2A1O1Ixp33_ASAP7_75t_L g1487 ( 
.A1(n_1249),
.A2(n_675),
.B(n_674),
.C(n_929),
.Y(n_1487)
);

BUFx6f_ASAP7_75t_L g1488 ( 
.A(n_1321),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1186),
.B(n_1206),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1190),
.Y(n_1490)
);

AOI22xp33_ASAP7_75t_SL g1491 ( 
.A1(n_1302),
.A2(n_675),
.B1(n_967),
.B2(n_674),
.Y(n_1491)
);

AOI221xp5_ASAP7_75t_L g1492 ( 
.A1(n_1484),
.A2(n_1487),
.B1(n_1478),
.B2(n_1362),
.C(n_1486),
.Y(n_1492)
);

OA21x2_ASAP7_75t_L g1493 ( 
.A1(n_1432),
.A2(n_1459),
.B(n_1413),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1354),
.Y(n_1494)
);

OAI211xp5_ASAP7_75t_SL g1495 ( 
.A1(n_1485),
.A2(n_1491),
.B(n_1474),
.C(n_1478),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1365),
.Y(n_1496)
);

BUFx6f_ASAP7_75t_L g1497 ( 
.A(n_1423),
.Y(n_1497)
);

AOI22xp33_ASAP7_75t_L g1498 ( 
.A1(n_1484),
.A2(n_1362),
.B1(n_1474),
.B2(n_1359),
.Y(n_1498)
);

OR2x6_ASAP7_75t_L g1499 ( 
.A(n_1440),
.B(n_1397),
.Y(n_1499)
);

AOI22xp33_ASAP7_75t_L g1500 ( 
.A1(n_1366),
.A2(n_1369),
.B1(n_1363),
.B2(n_1406),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1489),
.A2(n_1382),
.B1(n_1406),
.B2(n_1367),
.Y(n_1501)
);

AOI22xp5_ASAP7_75t_L g1502 ( 
.A1(n_1425),
.A2(n_1387),
.B1(n_1372),
.B2(n_1416),
.Y(n_1502)
);

OAI22xp33_ASAP7_75t_L g1503 ( 
.A1(n_1400),
.A2(n_1372),
.B1(n_1381),
.B2(n_1414),
.Y(n_1503)
);

AOI21xp33_ASAP7_75t_L g1504 ( 
.A1(n_1419),
.A2(n_1473),
.B(n_1375),
.Y(n_1504)
);

AOI221x1_ASAP7_75t_L g1505 ( 
.A1(n_1419),
.A2(n_1371),
.B1(n_1348),
.B2(n_1442),
.C(n_1397),
.Y(n_1505)
);

AOI22xp33_ASAP7_75t_L g1506 ( 
.A1(n_1356),
.A2(n_1477),
.B1(n_1352),
.B2(n_1371),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_SL g1507 ( 
.A1(n_1360),
.A2(n_1430),
.B1(n_1444),
.B2(n_1364),
.Y(n_1507)
);

AOI22xp33_ASAP7_75t_SL g1508 ( 
.A1(n_1360),
.A2(n_1430),
.B1(n_1364),
.B2(n_1380),
.Y(n_1508)
);

AOI21xp5_ASAP7_75t_L g1509 ( 
.A1(n_1436),
.A2(n_1472),
.B(n_1393),
.Y(n_1509)
);

A2O1A1Ixp33_ASAP7_75t_L g1510 ( 
.A1(n_1347),
.A2(n_1420),
.B(n_1415),
.C(n_1351),
.Y(n_1510)
);

INVx2_ASAP7_75t_SL g1511 ( 
.A(n_1384),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1383),
.B(n_1399),
.Y(n_1512)
);

INVxp67_ASAP7_75t_L g1513 ( 
.A(n_1377),
.Y(n_1513)
);

CKINVDCx6p67_ASAP7_75t_R g1514 ( 
.A(n_1386),
.Y(n_1514)
);

OAI211xp5_ASAP7_75t_L g1515 ( 
.A1(n_1479),
.A2(n_1348),
.B(n_1395),
.C(n_1422),
.Y(n_1515)
);

INVx1_ASAP7_75t_SL g1516 ( 
.A(n_1475),
.Y(n_1516)
);

OAI221xp5_ASAP7_75t_L g1517 ( 
.A1(n_1388),
.A2(n_1385),
.B1(n_1350),
.B2(n_1393),
.C(n_1417),
.Y(n_1517)
);

OAI22xp33_ASAP7_75t_L g1518 ( 
.A1(n_1374),
.A2(n_1379),
.B1(n_1483),
.B2(n_1490),
.Y(n_1518)
);

BUFx4f_ASAP7_75t_SL g1519 ( 
.A(n_1404),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1412),
.B(n_1358),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1370),
.Y(n_1521)
);

AND2x6_ASAP7_75t_SL g1522 ( 
.A(n_1398),
.B(n_1410),
.Y(n_1522)
);

NOR2xp33_ASAP7_75t_L g1523 ( 
.A(n_1368),
.B(n_1482),
.Y(n_1523)
);

OAI21xp5_ASAP7_75t_L g1524 ( 
.A1(n_1353),
.A2(n_1433),
.B(n_1349),
.Y(n_1524)
);

NAND3xp33_ASAP7_75t_L g1525 ( 
.A(n_1393),
.B(n_1355),
.C(n_1407),
.Y(n_1525)
);

AOI21xp33_ASAP7_75t_SL g1526 ( 
.A1(n_1378),
.A2(n_1411),
.B(n_1418),
.Y(n_1526)
);

OAI332xp33_ASAP7_75t_L g1527 ( 
.A1(n_1396),
.A2(n_1407),
.A3(n_1392),
.B1(n_1401),
.B2(n_1417),
.B3(n_1447),
.C1(n_1421),
.C2(n_1426),
.Y(n_1527)
);

CKINVDCx20_ASAP7_75t_R g1528 ( 
.A(n_1445),
.Y(n_1528)
);

AOI221xp5_ASAP7_75t_L g1529 ( 
.A1(n_1391),
.A2(n_1421),
.B1(n_1446),
.B2(n_1396),
.C(n_1450),
.Y(n_1529)
);

AOI221xp5_ASAP7_75t_L g1530 ( 
.A1(n_1462),
.A2(n_1453),
.B1(n_1452),
.B2(n_1443),
.C(n_1403),
.Y(n_1530)
);

AOI221xp5_ASAP7_75t_L g1531 ( 
.A1(n_1462),
.A2(n_1457),
.B1(n_1429),
.B2(n_1460),
.C(n_1451),
.Y(n_1531)
);

AND2x4_ASAP7_75t_L g1532 ( 
.A(n_1405),
.B(n_1440),
.Y(n_1532)
);

AOI222xp33_ASAP7_75t_L g1533 ( 
.A1(n_1434),
.A2(n_1409),
.B1(n_1361),
.B2(n_1373),
.C1(n_1376),
.C2(n_1357),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1404),
.A2(n_1427),
.B1(n_1390),
.B2(n_1437),
.Y(n_1534)
);

NOR3xp33_ASAP7_75t_L g1535 ( 
.A(n_1394),
.B(n_1476),
.C(n_1408),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1389),
.A2(n_1488),
.B1(n_1402),
.B2(n_1424),
.Y(n_1536)
);

OAI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1449),
.A2(n_1435),
.B1(n_1431),
.B2(n_1408),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1402),
.B(n_1488),
.Y(n_1538)
);

OAI22xp33_ASAP7_75t_L g1539 ( 
.A1(n_1394),
.A2(n_1476),
.B1(n_1428),
.B2(n_1439),
.Y(n_1539)
);

OAI221xp5_ASAP7_75t_L g1540 ( 
.A1(n_1471),
.A2(n_1456),
.B1(n_1469),
.B2(n_1470),
.C(n_1468),
.Y(n_1540)
);

OAI21x1_ASAP7_75t_L g1541 ( 
.A1(n_1454),
.A2(n_1465),
.B(n_1469),
.Y(n_1541)
);

AOI22xp33_ASAP7_75t_L g1542 ( 
.A1(n_1464),
.A2(n_1466),
.B1(n_1441),
.B2(n_1438),
.Y(n_1542)
);

OR2x2_ASAP7_75t_L g1543 ( 
.A(n_1467),
.B(n_1458),
.Y(n_1543)
);

OAI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1448),
.A2(n_1455),
.B1(n_1461),
.B2(n_1470),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1455),
.B(n_1461),
.Y(n_1545)
);

AND2x4_ASAP7_75t_L g1546 ( 
.A(n_1448),
.B(n_1463),
.Y(n_1546)
);

AOI21xp33_ASAP7_75t_L g1547 ( 
.A1(n_1460),
.A2(n_675),
.B(n_1487),
.Y(n_1547)
);

AOI221xp5_ASAP7_75t_L g1548 ( 
.A1(n_1448),
.A2(n_675),
.B1(n_674),
.B2(n_1484),
.C(n_1487),
.Y(n_1548)
);

AOI22xp33_ASAP7_75t_L g1549 ( 
.A1(n_1484),
.A2(n_929),
.B1(n_675),
.B2(n_1478),
.Y(n_1549)
);

AOI221xp5_ASAP7_75t_L g1550 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_674),
.B2(n_1487),
.C(n_1478),
.Y(n_1550)
);

NOR3xp33_ASAP7_75t_L g1551 ( 
.A(n_1487),
.B(n_675),
.C(n_929),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1485),
.A2(n_675),
.B1(n_1491),
.B2(n_1486),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1485),
.A2(n_675),
.B1(n_1491),
.B2(n_1486),
.Y(n_1553)
);

OR2x6_ASAP7_75t_L g1554 ( 
.A(n_1440),
.B(n_1397),
.Y(n_1554)
);

AOI22xp33_ASAP7_75t_L g1555 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_1362),
.B2(n_929),
.Y(n_1555)
);

NAND2xp5_ASAP7_75t_L g1556 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1354),
.Y(n_1557)
);

AND2x4_ASAP7_75t_L g1558 ( 
.A(n_1358),
.B(n_1368),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1478),
.A2(n_675),
.B(n_1218),
.Y(n_1559)
);

AOI22xp33_ASAP7_75t_SL g1560 ( 
.A1(n_1484),
.A2(n_1362),
.B1(n_675),
.B2(n_1369),
.Y(n_1560)
);

INVx4_ASAP7_75t_L g1561 ( 
.A(n_1423),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_SL g1562 ( 
.A1(n_1478),
.A2(n_675),
.B(n_1484),
.Y(n_1562)
);

OAI211xp5_ASAP7_75t_L g1563 ( 
.A1(n_1486),
.A2(n_675),
.B(n_674),
.C(n_1485),
.Y(n_1563)
);

AOI22xp5_ASAP7_75t_L g1564 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_929),
.B2(n_1486),
.Y(n_1564)
);

NAND2xp5_ASAP7_75t_L g1565 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1565)
);

AOI222xp33_ASAP7_75t_L g1566 ( 
.A1(n_1484),
.A2(n_929),
.B1(n_675),
.B2(n_1362),
.C1(n_1182),
.C2(n_456),
.Y(n_1566)
);

AOI222xp33_ASAP7_75t_L g1567 ( 
.A1(n_1484),
.A2(n_929),
.B1(n_675),
.B2(n_1362),
.C1(n_1182),
.C2(n_456),
.Y(n_1567)
);

BUFx12f_ASAP7_75t_L g1568 ( 
.A(n_1398),
.Y(n_1568)
);

OAI211xp5_ASAP7_75t_L g1569 ( 
.A1(n_1486),
.A2(n_675),
.B(n_674),
.C(n_1485),
.Y(n_1569)
);

AOI22xp33_ASAP7_75t_L g1570 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_1362),
.B2(n_929),
.Y(n_1570)
);

AOI222xp33_ASAP7_75t_L g1571 ( 
.A1(n_1484),
.A2(n_929),
.B1(n_675),
.B2(n_1362),
.C1(n_1182),
.C2(n_456),
.Y(n_1571)
);

OAI22xp5_ASAP7_75t_L g1572 ( 
.A1(n_1485),
.A2(n_675),
.B1(n_1491),
.B2(n_1486),
.Y(n_1572)
);

OAI211xp5_ASAP7_75t_L g1573 ( 
.A1(n_1486),
.A2(n_675),
.B(n_674),
.C(n_1485),
.Y(n_1573)
);

CKINVDCx5p33_ASAP7_75t_R g1574 ( 
.A(n_1378),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1575)
);

OAI221xp5_ASAP7_75t_L g1576 ( 
.A1(n_1486),
.A2(n_675),
.B1(n_1485),
.B2(n_1491),
.C(n_674),
.Y(n_1576)
);

AOI22xp33_ASAP7_75t_L g1577 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_1362),
.B2(n_929),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_674),
.B2(n_1487),
.C(n_1478),
.Y(n_1578)
);

O2A1O1Ixp33_ASAP7_75t_L g1579 ( 
.A1(n_1487),
.A2(n_675),
.B(n_1478),
.C(n_1484),
.Y(n_1579)
);

AOI22xp33_ASAP7_75t_L g1580 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_1362),
.B2(n_929),
.Y(n_1580)
);

OAI22xp5_ASAP7_75t_SL g1581 ( 
.A1(n_1485),
.A2(n_1491),
.B1(n_1302),
.B2(n_926),
.Y(n_1581)
);

OAI22xp5_ASAP7_75t_L g1582 ( 
.A1(n_1485),
.A2(n_675),
.B1(n_1491),
.B2(n_1486),
.Y(n_1582)
);

CKINVDCx5p33_ASAP7_75t_R g1583 ( 
.A(n_1378),
.Y(n_1583)
);

AOI33xp33_ASAP7_75t_L g1584 ( 
.A1(n_1485),
.A2(n_802),
.A3(n_513),
.B1(n_1110),
.B2(n_1491),
.B3(n_983),
.Y(n_1584)
);

OAI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1485),
.A2(n_675),
.B1(n_1491),
.B2(n_1486),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1485),
.A2(n_675),
.B1(n_1491),
.B2(n_1486),
.Y(n_1586)
);

AOI22xp33_ASAP7_75t_L g1587 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_1362),
.B2(n_929),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_SL g1588 ( 
.A1(n_1484),
.A2(n_1362),
.B1(n_675),
.B2(n_1369),
.Y(n_1588)
);

INVx4_ASAP7_75t_L g1589 ( 
.A(n_1423),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1590)
);

AOI22xp33_ASAP7_75t_L g1591 ( 
.A1(n_1484),
.A2(n_929),
.B1(n_675),
.B2(n_1478),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1480),
.B(n_1481),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_L g1593 ( 
.A1(n_1484),
.A2(n_675),
.B1(n_1362),
.B2(n_929),
.Y(n_1593)
);

AOI22xp33_ASAP7_75t_L g1594 ( 
.A1(n_1484),
.A2(n_929),
.B1(n_675),
.B2(n_1478),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1545),
.B(n_1543),
.Y(n_1595)
);

OR2x2_ASAP7_75t_L g1596 ( 
.A(n_1493),
.B(n_1544),
.Y(n_1596)
);

AND2x2_ASAP7_75t_L g1597 ( 
.A(n_1531),
.B(n_1493),
.Y(n_1597)
);

INVxp33_ASAP7_75t_L g1598 ( 
.A(n_1556),
.Y(n_1598)
);

AOI22xp33_ASAP7_75t_L g1599 ( 
.A1(n_1560),
.A2(n_1588),
.B1(n_1495),
.B2(n_1571),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1546),
.B(n_1542),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1541),
.Y(n_1601)
);

INVx3_ASAP7_75t_L g1602 ( 
.A(n_1546),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1494),
.Y(n_1603)
);

AND2x2_ASAP7_75t_L g1604 ( 
.A(n_1542),
.B(n_1499),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1496),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1559),
.B(n_1492),
.Y(n_1606)
);

AND2x4_ASAP7_75t_L g1607 ( 
.A(n_1554),
.B(n_1509),
.Y(n_1607)
);

AND2x2_ASAP7_75t_L g1608 ( 
.A(n_1554),
.B(n_1529),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1521),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1557),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1540),
.Y(n_1611)
);

OR2x2_ASAP7_75t_L g1612 ( 
.A(n_1524),
.B(n_1525),
.Y(n_1612)
);

INVx4_ASAP7_75t_L g1613 ( 
.A(n_1554),
.Y(n_1613)
);

BUFx2_ASAP7_75t_L g1614 ( 
.A(n_1530),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1518),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1505),
.B(n_1551),
.Y(n_1616)
);

OR2x2_ASAP7_75t_L g1617 ( 
.A(n_1537),
.B(n_1513),
.Y(n_1617)
);

NAND2xp5_ASAP7_75t_L g1618 ( 
.A(n_1551),
.B(n_1550),
.Y(n_1618)
);

AND2x2_ASAP7_75t_L g1619 ( 
.A(n_1508),
.B(n_1507),
.Y(n_1619)
);

INVxp33_ASAP7_75t_L g1620 ( 
.A(n_1565),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1578),
.B(n_1503),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1548),
.B(n_1579),
.Y(n_1622)
);

HB1xp67_ASAP7_75t_L g1623 ( 
.A(n_1532),
.Y(n_1623)
);

BUFx2_ASAP7_75t_L g1624 ( 
.A(n_1510),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1508),
.B(n_1507),
.Y(n_1625)
);

BUFx2_ASAP7_75t_L g1626 ( 
.A(n_1539),
.Y(n_1626)
);

INVx1_ASAP7_75t_L g1627 ( 
.A(n_1533),
.Y(n_1627)
);

HB1xp67_ASAP7_75t_L g1628 ( 
.A(n_1547),
.Y(n_1628)
);

BUFx12f_ASAP7_75t_L g1629 ( 
.A(n_1561),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1560),
.B(n_1588),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1538),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1515),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1564),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1498),
.B(n_1504),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1562),
.Y(n_1635)
);

AND2x2_ASAP7_75t_L g1636 ( 
.A(n_1500),
.B(n_1549),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1534),
.Y(n_1637)
);

AND2x2_ASAP7_75t_L g1638 ( 
.A(n_1549),
.B(n_1591),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1575),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1591),
.B(n_1594),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1629),
.Y(n_1641)
);

OAI22xp33_ASAP7_75t_L g1642 ( 
.A1(n_1624),
.A2(n_1576),
.B1(n_1552),
.B2(n_1586),
.Y(n_1642)
);

AND2x2_ASAP7_75t_L g1643 ( 
.A(n_1595),
.B(n_1592),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1605),
.Y(n_1644)
);

AOI221xp5_ASAP7_75t_L g1645 ( 
.A1(n_1624),
.A2(n_1581),
.B1(n_1572),
.B2(n_1553),
.C(n_1585),
.Y(n_1645)
);

INVx4_ASAP7_75t_R g1646 ( 
.A(n_1631),
.Y(n_1646)
);

OAI22xp5_ASAP7_75t_L g1647 ( 
.A1(n_1624),
.A2(n_1555),
.B1(n_1593),
.B2(n_1587),
.Y(n_1647)
);

AND2x2_ASAP7_75t_L g1648 ( 
.A(n_1595),
.B(n_1520),
.Y(n_1648)
);

OAI221xp5_ASAP7_75t_L g1649 ( 
.A1(n_1606),
.A2(n_1570),
.B1(n_1577),
.B2(n_1580),
.C(n_1567),
.Y(n_1649)
);

OAI211xp5_ASAP7_75t_L g1650 ( 
.A1(n_1599),
.A2(n_1566),
.B(n_1573),
.C(n_1569),
.Y(n_1650)
);

INVx2_ASAP7_75t_SL g1651 ( 
.A(n_1602),
.Y(n_1651)
);

AOI221xp5_ASAP7_75t_L g1652 ( 
.A1(n_1614),
.A2(n_1582),
.B1(n_1495),
.B2(n_1563),
.C(n_1594),
.Y(n_1652)
);

OAI211xp5_ASAP7_75t_L g1653 ( 
.A1(n_1599),
.A2(n_1501),
.B(n_1502),
.C(n_1506),
.Y(n_1653)
);

AOI22xp33_ASAP7_75t_L g1654 ( 
.A1(n_1634),
.A2(n_1501),
.B1(n_1506),
.B2(n_1584),
.Y(n_1654)
);

OR2x6_ASAP7_75t_L g1655 ( 
.A(n_1607),
.B(n_1497),
.Y(n_1655)
);

NAND3xp33_ASAP7_75t_L g1656 ( 
.A(n_1606),
.B(n_1517),
.C(n_1536),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1595),
.B(n_1590),
.Y(n_1657)
);

OAI22xp5_ASAP7_75t_L g1658 ( 
.A1(n_1621),
.A2(n_1589),
.B1(n_1561),
.B2(n_1497),
.Y(n_1658)
);

INVx4_ASAP7_75t_L g1659 ( 
.A(n_1629),
.Y(n_1659)
);

BUFx2_ASAP7_75t_L g1660 ( 
.A(n_1623),
.Y(n_1660)
);

NAND2xp5_ASAP7_75t_SL g1661 ( 
.A(n_1606),
.B(n_1535),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1639),
.B(n_1516),
.Y(n_1662)
);

NAND2xp5_ASAP7_75t_L g1663 ( 
.A(n_1639),
.B(n_1527),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1605),
.Y(n_1664)
);

AND2x2_ASAP7_75t_L g1665 ( 
.A(n_1595),
.B(n_1512),
.Y(n_1665)
);

AOI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1634),
.A2(n_1514),
.B1(n_1589),
.B2(n_1511),
.Y(n_1666)
);

NOR5xp2_ASAP7_75t_SL g1667 ( 
.A(n_1614),
.B(n_1522),
.C(n_1519),
.D(n_1497),
.E(n_1526),
.Y(n_1667)
);

OAI21x1_ASAP7_75t_L g1668 ( 
.A1(n_1601),
.A2(n_1535),
.B(n_1523),
.Y(n_1668)
);

INVxp67_ASAP7_75t_SL g1669 ( 
.A(n_1617),
.Y(n_1669)
);

NAND3xp33_ASAP7_75t_L g1670 ( 
.A(n_1618),
.B(n_1497),
.C(n_1558),
.Y(n_1670)
);

NAND2xp33_ASAP7_75t_R g1671 ( 
.A(n_1614),
.B(n_1626),
.Y(n_1671)
);

INVx1_ASAP7_75t_L g1672 ( 
.A(n_1605),
.Y(n_1672)
);

BUFx10_ASAP7_75t_L g1673 ( 
.A(n_1632),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1617),
.B(n_1574),
.Y(n_1674)
);

INVx1_ASAP7_75t_L g1675 ( 
.A(n_1609),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1603),
.Y(n_1676)
);

AND2x4_ASAP7_75t_L g1677 ( 
.A(n_1602),
.B(n_1528),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1609),
.Y(n_1678)
);

INVx1_ASAP7_75t_L g1679 ( 
.A(n_1609),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1610),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1623),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1618),
.B(n_1583),
.C(n_1519),
.Y(n_1682)
);

AND2x4_ASAP7_75t_L g1683 ( 
.A(n_1602),
.B(n_1568),
.Y(n_1683)
);

OAI22xp33_ASAP7_75t_L g1684 ( 
.A1(n_1621),
.A2(n_1622),
.B1(n_1630),
.B2(n_1618),
.Y(n_1684)
);

AO21x2_ASAP7_75t_L g1685 ( 
.A1(n_1616),
.A2(n_1622),
.B(n_1628),
.Y(n_1685)
);

NOR2xp67_ASAP7_75t_L g1686 ( 
.A(n_1651),
.B(n_1596),
.Y(n_1686)
);

AND2x2_ASAP7_75t_L g1687 ( 
.A(n_1651),
.B(n_1600),
.Y(n_1687)
);

BUFx3_ASAP7_75t_L g1688 ( 
.A(n_1641),
.Y(n_1688)
);

OR2x2_ASAP7_75t_L g1689 ( 
.A(n_1685),
.B(n_1596),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1669),
.B(n_1600),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1685),
.B(n_1596),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1676),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1644),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1664),
.Y(n_1694)
);

INVx1_ASAP7_75t_L g1695 ( 
.A(n_1672),
.Y(n_1695)
);

NOR2xp33_ASAP7_75t_R g1696 ( 
.A(n_1671),
.B(n_1629),
.Y(n_1696)
);

OR2x2_ASAP7_75t_L g1697 ( 
.A(n_1685),
.B(n_1596),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1675),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1597),
.Y(n_1699)
);

HB1xp67_ASAP7_75t_L g1700 ( 
.A(n_1678),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1679),
.B(n_1628),
.Y(n_1701)
);

NOR2xp67_ASAP7_75t_L g1702 ( 
.A(n_1670),
.B(n_1659),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1680),
.B(n_1615),
.Y(n_1703)
);

AND2x4_ASAP7_75t_SL g1704 ( 
.A(n_1673),
.B(n_1613),
.Y(n_1704)
);

INVx1_ASAP7_75t_L g1705 ( 
.A(n_1662),
.Y(n_1705)
);

INVx2_ASAP7_75t_SL g1706 ( 
.A(n_1646),
.Y(n_1706)
);

INVx2_ASAP7_75t_L g1707 ( 
.A(n_1668),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1660),
.Y(n_1708)
);

INVx2_ASAP7_75t_L g1709 ( 
.A(n_1668),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1681),
.Y(n_1710)
);

AND2x2_ASAP7_75t_L g1711 ( 
.A(n_1657),
.B(n_1597),
.Y(n_1711)
);

NAND2xp5_ASAP7_75t_L g1712 ( 
.A(n_1643),
.B(n_1615),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1655),
.B(n_1597),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1655),
.B(n_1597),
.Y(n_1714)
);

AND2x2_ASAP7_75t_L g1715 ( 
.A(n_1655),
.B(n_1604),
.Y(n_1715)
);

INVxp67_ASAP7_75t_L g1716 ( 
.A(n_1671),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1700),
.Y(n_1717)
);

AND2x2_ASAP7_75t_L g1718 ( 
.A(n_1699),
.B(n_1602),
.Y(n_1718)
);

OAI33xp33_ASAP7_75t_L g1719 ( 
.A1(n_1701),
.A2(n_1684),
.A3(n_1642),
.B1(n_1616),
.B2(n_1661),
.B3(n_1663),
.Y(n_1719)
);

INVx2_ASAP7_75t_L g1720 ( 
.A(n_1692),
.Y(n_1720)
);

AOI22xp33_ASAP7_75t_SL g1721 ( 
.A1(n_1696),
.A2(n_1650),
.B1(n_1619),
.B2(n_1625),
.Y(n_1721)
);

OR2x2_ASAP7_75t_L g1722 ( 
.A(n_1689),
.B(n_1612),
.Y(n_1722)
);

INVx1_ASAP7_75t_SL g1723 ( 
.A(n_1696),
.Y(n_1723)
);

OAI31xp33_ASAP7_75t_SL g1724 ( 
.A1(n_1715),
.A2(n_1645),
.A3(n_1653),
.B(n_1649),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1699),
.B(n_1711),
.Y(n_1725)
);

INVx1_ASAP7_75t_L g1726 ( 
.A(n_1700),
.Y(n_1726)
);

INVx1_ASAP7_75t_L g1727 ( 
.A(n_1693),
.Y(n_1727)
);

INVx2_ASAP7_75t_SL g1728 ( 
.A(n_1706),
.Y(n_1728)
);

INVx2_ASAP7_75t_SL g1729 ( 
.A(n_1706),
.Y(n_1729)
);

OR2x2_ASAP7_75t_L g1730 ( 
.A(n_1689),
.B(n_1612),
.Y(n_1730)
);

OAI21xp5_ASAP7_75t_L g1731 ( 
.A1(n_1716),
.A2(n_1622),
.B(n_1661),
.Y(n_1731)
);

OR2x2_ASAP7_75t_L g1732 ( 
.A(n_1689),
.B(n_1691),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1694),
.Y(n_1733)
);

INVxp67_ASAP7_75t_L g1734 ( 
.A(n_1712),
.Y(n_1734)
);

NOR2xp33_ASAP7_75t_L g1735 ( 
.A(n_1688),
.B(n_1629),
.Y(n_1735)
);

INVxp33_ASAP7_75t_L g1736 ( 
.A(n_1702),
.Y(n_1736)
);

OR2x2_ASAP7_75t_L g1737 ( 
.A(n_1691),
.B(n_1612),
.Y(n_1737)
);

INVx2_ASAP7_75t_SL g1738 ( 
.A(n_1706),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1711),
.B(n_1665),
.Y(n_1739)
);

AND2x4_ASAP7_75t_L g1740 ( 
.A(n_1686),
.B(n_1683),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1694),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1691),
.B(n_1612),
.Y(n_1742)
);

INVx1_ASAP7_75t_L g1743 ( 
.A(n_1693),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1711),
.B(n_1712),
.Y(n_1744)
);

OR2x2_ASAP7_75t_L g1745 ( 
.A(n_1697),
.B(n_1617),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1705),
.B(n_1611),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1694),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1716),
.B(n_1690),
.Y(n_1748)
);

INVxp67_ASAP7_75t_SL g1749 ( 
.A(n_1686),
.Y(n_1749)
);

INVx1_ASAP7_75t_L g1750 ( 
.A(n_1695),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1690),
.B(n_1648),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1690),
.B(n_1648),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1687),
.B(n_1607),
.Y(n_1753)
);

INVx1_ASAP7_75t_L g1754 ( 
.A(n_1698),
.Y(n_1754)
);

HB1xp67_ASAP7_75t_L g1755 ( 
.A(n_1748),
.Y(n_1755)
);

AND2x2_ASAP7_75t_L g1756 ( 
.A(n_1736),
.B(n_1713),
.Y(n_1756)
);

NAND3xp33_ASAP7_75t_L g1757 ( 
.A(n_1724),
.B(n_1652),
.C(n_1654),
.Y(n_1757)
);

INVxp67_ASAP7_75t_L g1758 ( 
.A(n_1731),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1734),
.B(n_1701),
.Y(n_1759)
);

INVx1_ASAP7_75t_L g1760 ( 
.A(n_1727),
.Y(n_1760)
);

INVxp67_ASAP7_75t_L g1761 ( 
.A(n_1746),
.Y(n_1761)
);

INVx2_ASAP7_75t_SL g1762 ( 
.A(n_1728),
.Y(n_1762)
);

NAND4xp25_ASAP7_75t_L g1763 ( 
.A(n_1721),
.B(n_1654),
.C(n_1621),
.D(n_1616),
.Y(n_1763)
);

INVx1_ASAP7_75t_L g1764 ( 
.A(n_1743),
.Y(n_1764)
);

INVxp67_ASAP7_75t_SL g1765 ( 
.A(n_1749),
.Y(n_1765)
);

INVx1_ASAP7_75t_L g1766 ( 
.A(n_1750),
.Y(n_1766)
);

OAI22xp5_ASAP7_75t_SL g1767 ( 
.A1(n_1723),
.A2(n_1682),
.B1(n_1658),
.B2(n_1666),
.Y(n_1767)
);

AND2x2_ASAP7_75t_L g1768 ( 
.A(n_1740),
.B(n_1713),
.Y(n_1768)
);

AND2x2_ASAP7_75t_SL g1769 ( 
.A(n_1740),
.B(n_1619),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1717),
.Y(n_1770)
);

AOI22x1_ASAP7_75t_L g1771 ( 
.A1(n_1719),
.A2(n_1641),
.B1(n_1632),
.B2(n_1659),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1722),
.B(n_1697),
.Y(n_1772)
);

NOR2xp33_ASAP7_75t_L g1773 ( 
.A(n_1735),
.B(n_1688),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1717),
.Y(n_1774)
);

INVxp67_ASAP7_75t_L g1775 ( 
.A(n_1748),
.Y(n_1775)
);

INVx2_ASAP7_75t_L g1776 ( 
.A(n_1720),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1720),
.Y(n_1777)
);

BUFx2_ASAP7_75t_L g1778 ( 
.A(n_1740),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1739),
.B(n_1753),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1733),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1726),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_SL g1782 ( 
.A(n_1728),
.B(n_1702),
.Y(n_1782)
);

AND2x2_ASAP7_75t_L g1783 ( 
.A(n_1739),
.B(n_1713),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1744),
.B(n_1722),
.Y(n_1784)
);

AO21x2_ASAP7_75t_L g1785 ( 
.A1(n_1732),
.A2(n_1697),
.B(n_1709),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1753),
.B(n_1714),
.Y(n_1786)
);

NAND2xp33_ASAP7_75t_R g1787 ( 
.A(n_1730),
.B(n_1667),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_SL g1788 ( 
.A(n_1729),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1733),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1729),
.Y(n_1790)
);

INVx1_ASAP7_75t_L g1791 ( 
.A(n_1741),
.Y(n_1791)
);

AND2x4_ASAP7_75t_SL g1792 ( 
.A(n_1738),
.B(n_1673),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1751),
.B(n_1714),
.Y(n_1793)
);

INVx3_ASAP7_75t_L g1794 ( 
.A(n_1718),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1730),
.B(n_1703),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1751),
.B(n_1714),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1752),
.B(n_1715),
.Y(n_1797)
);

AND2x2_ASAP7_75t_L g1798 ( 
.A(n_1769),
.B(n_1738),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1758),
.B(n_1771),
.Y(n_1799)
);

INVx2_ASAP7_75t_SL g1800 ( 
.A(n_1792),
.Y(n_1800)
);

INVx1_ASAP7_75t_L g1801 ( 
.A(n_1760),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1758),
.B(n_1752),
.Y(n_1802)
);

AOI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1757),
.A2(n_1647),
.B(n_1625),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1757),
.A2(n_1625),
.B(n_1619),
.Y(n_1804)
);

AOI222xp33_ASAP7_75t_L g1805 ( 
.A1(n_1767),
.A2(n_1634),
.B1(n_1619),
.B2(n_1625),
.C1(n_1636),
.C2(n_1632),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1760),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1764),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1764),
.Y(n_1808)
);

INVx1_ASAP7_75t_L g1809 ( 
.A(n_1766),
.Y(n_1809)
);

NOR3xp33_ASAP7_75t_SL g1810 ( 
.A(n_1787),
.B(n_1656),
.C(n_1667),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1766),
.Y(n_1811)
);

AND2x2_ASAP7_75t_L g1812 ( 
.A(n_1769),
.B(n_1778),
.Y(n_1812)
);

AOI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1763),
.A2(n_1634),
.B1(n_1630),
.B2(n_1636),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1771),
.B(n_1725),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1770),
.Y(n_1815)
);

INVxp67_ASAP7_75t_L g1816 ( 
.A(n_1765),
.Y(n_1816)
);

AOI322xp5_ASAP7_75t_L g1817 ( 
.A1(n_1769),
.A2(n_1636),
.A3(n_1630),
.B1(n_1638),
.B2(n_1608),
.C1(n_1640),
.C2(n_1633),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_SL g1818 ( 
.A1(n_1763),
.A2(n_1773),
.B(n_1775),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1770),
.Y(n_1819)
);

INVx1_ASAP7_75t_L g1820 ( 
.A(n_1774),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1767),
.B(n_1688),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1774),
.Y(n_1822)
);

INVx1_ASAP7_75t_L g1823 ( 
.A(n_1781),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1781),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1756),
.A2(n_1636),
.B1(n_1638),
.B2(n_1633),
.Y(n_1825)
);

AOI22xp33_ASAP7_75t_L g1826 ( 
.A1(n_1756),
.A2(n_1638),
.B1(n_1633),
.B2(n_1608),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1755),
.Y(n_1827)
);

INVx2_ASAP7_75t_L g1828 ( 
.A(n_1794),
.Y(n_1828)
);

AND2x2_ASAP7_75t_L g1829 ( 
.A(n_1778),
.B(n_1718),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1789),
.Y(n_1830)
);

AOI221xp5_ASAP7_75t_L g1831 ( 
.A1(n_1761),
.A2(n_1742),
.B1(n_1737),
.B2(n_1745),
.C(n_1732),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1789),
.Y(n_1832)
);

AOI22xp33_ASAP7_75t_L g1833 ( 
.A1(n_1782),
.A2(n_1638),
.B1(n_1608),
.B2(n_1635),
.Y(n_1833)
);

OR2x2_ASAP7_75t_L g1834 ( 
.A(n_1802),
.B(n_1759),
.Y(n_1834)
);

AOI31xp33_ASAP7_75t_L g1835 ( 
.A1(n_1821),
.A2(n_1790),
.A3(n_1762),
.B(n_1768),
.Y(n_1835)
);

CKINVDCx16_ASAP7_75t_R g1836 ( 
.A(n_1812),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1815),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1803),
.B(n_1797),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1818),
.B(n_1674),
.Y(n_1839)
);

OAI21xp33_ASAP7_75t_L g1840 ( 
.A1(n_1799),
.A2(n_1784),
.B(n_1759),
.Y(n_1840)
);

OR2x2_ASAP7_75t_L g1841 ( 
.A(n_1816),
.B(n_1784),
.Y(n_1841)
);

NAND4xp25_ASAP7_75t_L g1842 ( 
.A(n_1805),
.B(n_1790),
.C(n_1768),
.D(n_1742),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1804),
.B(n_1797),
.Y(n_1843)
);

OAI22xp5_ASAP7_75t_L g1844 ( 
.A1(n_1810),
.A2(n_1788),
.B1(n_1762),
.B2(n_1792),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1812),
.B(n_1798),
.Y(n_1845)
);

AOI32xp33_ASAP7_75t_L g1846 ( 
.A1(n_1821),
.A2(n_1813),
.A3(n_1814),
.B1(n_1798),
.B2(n_1833),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1817),
.B(n_1793),
.Y(n_1847)
);

AOI22xp33_ASAP7_75t_L g1848 ( 
.A1(n_1825),
.A2(n_1635),
.B1(n_1608),
.B2(n_1640),
.Y(n_1848)
);

OAI32xp33_ASAP7_75t_L g1849 ( 
.A1(n_1827),
.A2(n_1737),
.A3(n_1745),
.B1(n_1788),
.B2(n_1772),
.Y(n_1849)
);

A2O1A1Ixp33_ASAP7_75t_SL g1850 ( 
.A1(n_1827),
.A2(n_1777),
.B(n_1776),
.C(n_1780),
.Y(n_1850)
);

NAND2xp5_ASAP7_75t_L g1851 ( 
.A(n_1826),
.B(n_1793),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1815),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1820),
.Y(n_1853)
);

INVx1_ASAP7_75t_L g1854 ( 
.A(n_1820),
.Y(n_1854)
);

NOR3xp33_ASAP7_75t_L g1855 ( 
.A(n_1823),
.B(n_1659),
.C(n_1640),
.Y(n_1855)
);

AOI22xp33_ASAP7_75t_L g1856 ( 
.A1(n_1824),
.A2(n_1635),
.B1(n_1611),
.B2(n_1627),
.Y(n_1856)
);

INVx1_ASAP7_75t_SL g1857 ( 
.A(n_1800),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1806),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1800),
.B(n_1795),
.Y(n_1859)
);

INVx1_ASAP7_75t_L g1860 ( 
.A(n_1837),
.Y(n_1860)
);

O2A1O1Ixp33_ASAP7_75t_L g1861 ( 
.A1(n_1835),
.A2(n_1819),
.B(n_1822),
.C(n_1809),
.Y(n_1861)
);

O2A1O1Ixp33_ASAP7_75t_L g1862 ( 
.A1(n_1850),
.A2(n_1849),
.B(n_1839),
.C(n_1855),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1846),
.A2(n_1838),
.B(n_1840),
.C(n_1847),
.Y(n_1863)
);

XNOR2xp5_ASAP7_75t_L g1864 ( 
.A(n_1842),
.B(n_1677),
.Y(n_1864)
);

NAND2xp5_ASAP7_75t_SL g1865 ( 
.A(n_1836),
.B(n_1844),
.Y(n_1865)
);

NAND3xp33_ASAP7_75t_L g1866 ( 
.A(n_1855),
.B(n_1856),
.C(n_1841),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_R g1867 ( 
.A(n_1857),
.B(n_1801),
.Y(n_1867)
);

INVx1_ASAP7_75t_L g1868 ( 
.A(n_1852),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1845),
.B(n_1856),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1853),
.Y(n_1870)
);

INVx1_ASAP7_75t_L g1871 ( 
.A(n_1854),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1858),
.Y(n_1872)
);

INVx2_ASAP7_75t_L g1873 ( 
.A(n_1859),
.Y(n_1873)
);

NAND2x1_ASAP7_75t_L g1874 ( 
.A(n_1843),
.B(n_1829),
.Y(n_1874)
);

INVx1_ASAP7_75t_SL g1875 ( 
.A(n_1834),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1851),
.B(n_1829),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1848),
.B(n_1811),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1848),
.Y(n_1878)
);

XOR2x2_ASAP7_75t_L g1879 ( 
.A(n_1839),
.B(n_1677),
.Y(n_1879)
);

AOI221xp5_ASAP7_75t_SL g1880 ( 
.A1(n_1862),
.A2(n_1861),
.B1(n_1863),
.B2(n_1865),
.C(n_1878),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1873),
.Y(n_1881)
);

AO22x2_ASAP7_75t_L g1882 ( 
.A1(n_1865),
.A2(n_1807),
.B1(n_1806),
.B2(n_1808),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1873),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1860),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1876),
.B(n_1783),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1868),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1875),
.B(n_1828),
.Y(n_1887)
);

NOR2x1_ASAP7_75t_L g1888 ( 
.A(n_1866),
.B(n_1807),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1870),
.Y(n_1889)
);

AOI22xp5_ASAP7_75t_L g1890 ( 
.A1(n_1863),
.A2(n_1831),
.B1(n_1808),
.B2(n_1828),
.Y(n_1890)
);

INVx2_ASAP7_75t_SL g1891 ( 
.A(n_1867),
.Y(n_1891)
);

AOI211xp5_ASAP7_75t_L g1892 ( 
.A1(n_1880),
.A2(n_1867),
.B(n_1877),
.C(n_1869),
.Y(n_1892)
);

OAI211xp5_ASAP7_75t_L g1893 ( 
.A1(n_1888),
.A2(n_1874),
.B(n_1871),
.C(n_1872),
.Y(n_1893)
);

AOI22xp33_ASAP7_75t_SL g1894 ( 
.A1(n_1882),
.A2(n_1864),
.B1(n_1792),
.B2(n_1785),
.Y(n_1894)
);

NAND5xp2_ASAP7_75t_L g1895 ( 
.A(n_1890),
.B(n_1881),
.C(n_1887),
.D(n_1885),
.E(n_1886),
.Y(n_1895)
);

NAND3xp33_ASAP7_75t_L g1896 ( 
.A(n_1891),
.B(n_1832),
.C(n_1830),
.Y(n_1896)
);

AOI221xp5_ASAP7_75t_L g1897 ( 
.A1(n_1882),
.A2(n_1891),
.B1(n_1883),
.B2(n_1887),
.C(n_1884),
.Y(n_1897)
);

NOR3xp33_ASAP7_75t_L g1898 ( 
.A(n_1883),
.B(n_1879),
.C(n_1794),
.Y(n_1898)
);

NAND4xp25_ASAP7_75t_L g1899 ( 
.A(n_1889),
.B(n_1772),
.C(n_1677),
.D(n_1796),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1882),
.A2(n_1785),
.B1(n_1791),
.B2(n_1777),
.C(n_1776),
.Y(n_1900)
);

INVx1_ASAP7_75t_SL g1901 ( 
.A(n_1891),
.Y(n_1901)
);

AOI211xp5_ASAP7_75t_L g1902 ( 
.A1(n_1880),
.A2(n_1796),
.B(n_1783),
.C(n_1786),
.Y(n_1902)
);

NAND2xp5_ASAP7_75t_L g1903 ( 
.A(n_1901),
.B(n_1779),
.Y(n_1903)
);

AOI21xp5_ASAP7_75t_L g1904 ( 
.A1(n_1895),
.A2(n_1785),
.B(n_1776),
.Y(n_1904)
);

XNOR2xp5_ASAP7_75t_L g1905 ( 
.A(n_1892),
.B(n_1683),
.Y(n_1905)
);

INVx1_ASAP7_75t_SL g1906 ( 
.A(n_1894),
.Y(n_1906)
);

NOR3xp33_ASAP7_75t_L g1907 ( 
.A(n_1893),
.B(n_1794),
.C(n_1795),
.Y(n_1907)
);

NOR2xp67_ASAP7_75t_L g1908 ( 
.A(n_1896),
.B(n_1777),
.Y(n_1908)
);

NOR2xp33_ASAP7_75t_L g1909 ( 
.A(n_1903),
.B(n_1899),
.Y(n_1909)
);

INVx1_ASAP7_75t_L g1910 ( 
.A(n_1908),
.Y(n_1910)
);

NAND2xp5_ASAP7_75t_L g1911 ( 
.A(n_1906),
.B(n_1897),
.Y(n_1911)
);

AOI21xp5_ASAP7_75t_L g1912 ( 
.A1(n_1904),
.A2(n_1900),
.B(n_1898),
.Y(n_1912)
);

AND2x4_ASAP7_75t_L g1913 ( 
.A(n_1907),
.B(n_1786),
.Y(n_1913)
);

NAND4xp75_ASAP7_75t_L g1914 ( 
.A(n_1905),
.B(n_1902),
.C(n_1791),
.D(n_1780),
.Y(n_1914)
);

NOR2x1p5_ASAP7_75t_L g1915 ( 
.A(n_1914),
.B(n_1794),
.Y(n_1915)
);

NAND5xp2_ASAP7_75t_L g1916 ( 
.A(n_1909),
.B(n_1627),
.C(n_1715),
.D(n_1637),
.E(n_1779),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1910),
.Y(n_1917)
);

NOR2xp33_ASAP7_75t_SL g1918 ( 
.A(n_1913),
.B(n_1673),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1911),
.B(n_1780),
.Y(n_1919)
);

OR3x1_ASAP7_75t_L g1920 ( 
.A(n_1916),
.B(n_1912),
.C(n_1611),
.Y(n_1920)
);

NAND4xp75_ASAP7_75t_L g1921 ( 
.A(n_1917),
.B(n_1707),
.C(n_1709),
.D(n_1710),
.Y(n_1921)
);

NAND2xp5_ASAP7_75t_L g1922 ( 
.A(n_1915),
.B(n_1785),
.Y(n_1922)
);

OA21x2_ASAP7_75t_L g1923 ( 
.A1(n_1922),
.A2(n_1919),
.B(n_1918),
.Y(n_1923)
);

XOR2xp5_ASAP7_75t_L g1924 ( 
.A(n_1923),
.B(n_1920),
.Y(n_1924)
);

INVx1_ASAP7_75t_L g1925 ( 
.A(n_1924),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1924),
.Y(n_1926)
);

CKINVDCx20_ASAP7_75t_R g1927 ( 
.A(n_1925),
.Y(n_1927)
);

AOI211xp5_ASAP7_75t_L g1928 ( 
.A1(n_1926),
.A2(n_1923),
.B(n_1921),
.C(n_1709),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1927),
.A2(n_1754),
.B(n_1747),
.Y(n_1929)
);

HB1xp67_ASAP7_75t_L g1930 ( 
.A(n_1928),
.Y(n_1930)
);

AOI222xp33_ASAP7_75t_L g1931 ( 
.A1(n_1930),
.A2(n_1754),
.B1(n_1747),
.B2(n_1741),
.C1(n_1708),
.C2(n_1710),
.Y(n_1931)
);

OAI221xp5_ASAP7_75t_R g1932 ( 
.A1(n_1931),
.A2(n_1929),
.B1(n_1704),
.B2(n_1707),
.C(n_1708),
.Y(n_1932)
);

AOI211xp5_ASAP7_75t_L g1933 ( 
.A1(n_1932),
.A2(n_1707),
.B(n_1620),
.C(n_1598),
.Y(n_1933)
);


endmodule