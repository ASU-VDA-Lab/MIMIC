module fake_netlist_6_356_n_2623 (n_52, n_435, n_1, n_91, n_326, n_256, n_440, n_587, n_507, n_580, n_209, n_367, n_465, n_63, n_223, n_278, n_341, n_362, n_148, n_226, n_161, n_22, n_208, n_462, n_68, n_316, n_419, n_28, n_304, n_212, n_50, n_7, n_578, n_144, n_365, n_125, n_168, n_384, n_297, n_524, n_342, n_77, n_106, n_358, n_160, n_449, n_131, n_188, n_310, n_509, n_186, n_245, n_0, n_368, n_575, n_396, n_495, n_350, n_78, n_84, n_585, n_568, n_392, n_442, n_480, n_142, n_143, n_382, n_180, n_62, n_557, n_349, n_233, n_255, n_284, n_400, n_140, n_337, n_214, n_485, n_67, n_15, n_443, n_246, n_38, n_471, n_289, n_421, n_424, n_59, n_181, n_182, n_238, n_573, n_202, n_320, n_108, n_327, n_369, n_280, n_287, n_353, n_555, n_389, n_415, n_65, n_230, n_461, n_141, n_383, n_200, n_447, n_176, n_114, n_86, n_198, n_104, n_222, n_179, n_248, n_300, n_517, n_71, n_74, n_229, n_542, n_305, n_72, n_532, n_173, n_535, n_250, n_372, n_468, n_544, n_111, n_504, n_314, n_378, n_413, n_377, n_35, n_183, n_510, n_79, n_375, n_338, n_522, n_466, n_506, n_56, n_360, n_119, n_235, n_536, n_147, n_191, n_340, n_387, n_452, n_39, n_344, n_73, n_581, n_428, n_432, n_101, n_167, n_174, n_127, n_516, n_153, n_525, n_156, n_491, n_145, n_42, n_133, n_96, n_8, n_371, n_567, n_189, n_405, n_213, n_538, n_294, n_302, n_499, n_380, n_129, n_197, n_11, n_137, n_17, n_343, n_448, n_20, n_494, n_539, n_493, n_397, n_155, n_109, n_529, n_445, n_425, n_122, n_45, n_454, n_34, n_218, n_70, n_234, n_37, n_486, n_381, n_82, n_27, n_236, n_112, n_172, n_576, n_472, n_270, n_239, n_126, n_414, n_97, n_563, n_58, n_490, n_290, n_220, n_118, n_224, n_48, n_25, n_93, n_80, n_196, n_402, n_352, n_478, n_574, n_9, n_460, n_107, n_6, n_417, n_14, n_446, n_498, n_89, n_374, n_366, n_407, n_450, n_103, n_272, n_526, n_185, n_348, n_579, n_69, n_376, n_390, n_473, n_293, n_31, n_334, n_559, n_53, n_370, n_44, n_458, n_232, n_16, n_163, n_46, n_330, n_470, n_475, n_298, n_18, n_492, n_281, n_258, n_551, n_154, n_456, n_564, n_98, n_260, n_265, n_313, n_451, n_279, n_252, n_228, n_565, n_356, n_577, n_166, n_184, n_552, n_216, n_455, n_83, n_521, n_363, n_572, n_395, n_323, n_393, n_411, n_503, n_152, n_92, n_513, n_321, n_331, n_105, n_227, n_132, n_570, n_406, n_483, n_102, n_204, n_482, n_474, n_527, n_261, n_420, n_312, n_394, n_32, n_66, n_130, n_519, n_541, n_512, n_164, n_292, n_100, n_121, n_307, n_469, n_433, n_500, n_23, n_476, n_2, n_291, n_219, n_543, n_357, n_150, n_264, n_263, n_481, n_325, n_329, n_464, n_561, n_33, n_477, n_549, n_533, n_408, n_61, n_237, n_584, n_244, n_399, n_76, n_243, n_124, n_548, n_94, n_282, n_436, n_116, n_211, n_523, n_117, n_175, n_322, n_345, n_409, n_231, n_354, n_40, n_505, n_240, n_139, n_319, n_41, n_134, n_547, n_537, n_273, n_558, n_95, n_311, n_10, n_403, n_253, n_583, n_123, n_136, n_546, n_562, n_249, n_201, n_386, n_556, n_159, n_157, n_162, n_115, n_487, n_550, n_128, n_241, n_30, n_275, n_553, n_43, n_560, n_276, n_569, n_441, n_221, n_444, n_586, n_423, n_146, n_318, n_303, n_511, n_467, n_306, n_21, n_193, n_269, n_359, n_346, n_88, n_3, n_416, n_530, n_277, n_520, n_418, n_113, n_582, n_4, n_199, n_138, n_266, n_296, n_571, n_268, n_271, n_404, n_439, n_158, n_217, n_49, n_210, n_299, n_518, n_206, n_5, n_453, n_333, n_588, n_215, n_178, n_247, n_225, n_308, n_309, n_355, n_426, n_317, n_149, n_431, n_90, n_347, n_24, n_459, n_54, n_502, n_328, n_534, n_488, n_429, n_373, n_87, n_195, n_285, n_497, n_85, n_99, n_257, n_13, n_203, n_286, n_254, n_207, n_242, n_19, n_47, n_29, n_75, n_401, n_324, n_335, n_430, n_463, n_545, n_489, n_205, n_120, n_251, n_301, n_274, n_110, n_151, n_412, n_81, n_36, n_26, n_55, n_267, n_438, n_339, n_315, n_434, n_515, n_64, n_288, n_427, n_479, n_496, n_422, n_135, n_165, n_351, n_437, n_259, n_177, n_540, n_514, n_528, n_391, n_457, n_364, n_295, n_385, n_388, n_190, n_262, n_484, n_187, n_501, n_531, n_60, n_361, n_508, n_379, n_170, n_332, n_336, n_12, n_398, n_410, n_566, n_554, n_194, n_171, n_192, n_57, n_169, n_51, n_283, n_2623);

input n_52;
input n_435;
input n_1;
input n_91;
input n_326;
input n_256;
input n_440;
input n_587;
input n_507;
input n_580;
input n_209;
input n_367;
input n_465;
input n_63;
input n_223;
input n_278;
input n_341;
input n_362;
input n_148;
input n_226;
input n_161;
input n_22;
input n_208;
input n_462;
input n_68;
input n_316;
input n_419;
input n_28;
input n_304;
input n_212;
input n_50;
input n_7;
input n_578;
input n_144;
input n_365;
input n_125;
input n_168;
input n_384;
input n_297;
input n_524;
input n_342;
input n_77;
input n_106;
input n_358;
input n_160;
input n_449;
input n_131;
input n_188;
input n_310;
input n_509;
input n_186;
input n_245;
input n_0;
input n_368;
input n_575;
input n_396;
input n_495;
input n_350;
input n_78;
input n_84;
input n_585;
input n_568;
input n_392;
input n_442;
input n_480;
input n_142;
input n_143;
input n_382;
input n_180;
input n_62;
input n_557;
input n_349;
input n_233;
input n_255;
input n_284;
input n_400;
input n_140;
input n_337;
input n_214;
input n_485;
input n_67;
input n_15;
input n_443;
input n_246;
input n_38;
input n_471;
input n_289;
input n_421;
input n_424;
input n_59;
input n_181;
input n_182;
input n_238;
input n_573;
input n_202;
input n_320;
input n_108;
input n_327;
input n_369;
input n_280;
input n_287;
input n_353;
input n_555;
input n_389;
input n_415;
input n_65;
input n_230;
input n_461;
input n_141;
input n_383;
input n_200;
input n_447;
input n_176;
input n_114;
input n_86;
input n_198;
input n_104;
input n_222;
input n_179;
input n_248;
input n_300;
input n_517;
input n_71;
input n_74;
input n_229;
input n_542;
input n_305;
input n_72;
input n_532;
input n_173;
input n_535;
input n_250;
input n_372;
input n_468;
input n_544;
input n_111;
input n_504;
input n_314;
input n_378;
input n_413;
input n_377;
input n_35;
input n_183;
input n_510;
input n_79;
input n_375;
input n_338;
input n_522;
input n_466;
input n_506;
input n_56;
input n_360;
input n_119;
input n_235;
input n_536;
input n_147;
input n_191;
input n_340;
input n_387;
input n_452;
input n_39;
input n_344;
input n_73;
input n_581;
input n_428;
input n_432;
input n_101;
input n_167;
input n_174;
input n_127;
input n_516;
input n_153;
input n_525;
input n_156;
input n_491;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_371;
input n_567;
input n_189;
input n_405;
input n_213;
input n_538;
input n_294;
input n_302;
input n_499;
input n_380;
input n_129;
input n_197;
input n_11;
input n_137;
input n_17;
input n_343;
input n_448;
input n_20;
input n_494;
input n_539;
input n_493;
input n_397;
input n_155;
input n_109;
input n_529;
input n_445;
input n_425;
input n_122;
input n_45;
input n_454;
input n_34;
input n_218;
input n_70;
input n_234;
input n_37;
input n_486;
input n_381;
input n_82;
input n_27;
input n_236;
input n_112;
input n_172;
input n_576;
input n_472;
input n_270;
input n_239;
input n_126;
input n_414;
input n_97;
input n_563;
input n_58;
input n_490;
input n_290;
input n_220;
input n_118;
input n_224;
input n_48;
input n_25;
input n_93;
input n_80;
input n_196;
input n_402;
input n_352;
input n_478;
input n_574;
input n_9;
input n_460;
input n_107;
input n_6;
input n_417;
input n_14;
input n_446;
input n_498;
input n_89;
input n_374;
input n_366;
input n_407;
input n_450;
input n_103;
input n_272;
input n_526;
input n_185;
input n_348;
input n_579;
input n_69;
input n_376;
input n_390;
input n_473;
input n_293;
input n_31;
input n_334;
input n_559;
input n_53;
input n_370;
input n_44;
input n_458;
input n_232;
input n_16;
input n_163;
input n_46;
input n_330;
input n_470;
input n_475;
input n_298;
input n_18;
input n_492;
input n_281;
input n_258;
input n_551;
input n_154;
input n_456;
input n_564;
input n_98;
input n_260;
input n_265;
input n_313;
input n_451;
input n_279;
input n_252;
input n_228;
input n_565;
input n_356;
input n_577;
input n_166;
input n_184;
input n_552;
input n_216;
input n_455;
input n_83;
input n_521;
input n_363;
input n_572;
input n_395;
input n_323;
input n_393;
input n_411;
input n_503;
input n_152;
input n_92;
input n_513;
input n_321;
input n_331;
input n_105;
input n_227;
input n_132;
input n_570;
input n_406;
input n_483;
input n_102;
input n_204;
input n_482;
input n_474;
input n_527;
input n_261;
input n_420;
input n_312;
input n_394;
input n_32;
input n_66;
input n_130;
input n_519;
input n_541;
input n_512;
input n_164;
input n_292;
input n_100;
input n_121;
input n_307;
input n_469;
input n_433;
input n_500;
input n_23;
input n_476;
input n_2;
input n_291;
input n_219;
input n_543;
input n_357;
input n_150;
input n_264;
input n_263;
input n_481;
input n_325;
input n_329;
input n_464;
input n_561;
input n_33;
input n_477;
input n_549;
input n_533;
input n_408;
input n_61;
input n_237;
input n_584;
input n_244;
input n_399;
input n_76;
input n_243;
input n_124;
input n_548;
input n_94;
input n_282;
input n_436;
input n_116;
input n_211;
input n_523;
input n_117;
input n_175;
input n_322;
input n_345;
input n_409;
input n_231;
input n_354;
input n_40;
input n_505;
input n_240;
input n_139;
input n_319;
input n_41;
input n_134;
input n_547;
input n_537;
input n_273;
input n_558;
input n_95;
input n_311;
input n_10;
input n_403;
input n_253;
input n_583;
input n_123;
input n_136;
input n_546;
input n_562;
input n_249;
input n_201;
input n_386;
input n_556;
input n_159;
input n_157;
input n_162;
input n_115;
input n_487;
input n_550;
input n_128;
input n_241;
input n_30;
input n_275;
input n_553;
input n_43;
input n_560;
input n_276;
input n_569;
input n_441;
input n_221;
input n_444;
input n_586;
input n_423;
input n_146;
input n_318;
input n_303;
input n_511;
input n_467;
input n_306;
input n_21;
input n_193;
input n_269;
input n_359;
input n_346;
input n_88;
input n_3;
input n_416;
input n_530;
input n_277;
input n_520;
input n_418;
input n_113;
input n_582;
input n_4;
input n_199;
input n_138;
input n_266;
input n_296;
input n_571;
input n_268;
input n_271;
input n_404;
input n_439;
input n_158;
input n_217;
input n_49;
input n_210;
input n_299;
input n_518;
input n_206;
input n_5;
input n_453;
input n_333;
input n_588;
input n_215;
input n_178;
input n_247;
input n_225;
input n_308;
input n_309;
input n_355;
input n_426;
input n_317;
input n_149;
input n_431;
input n_90;
input n_347;
input n_24;
input n_459;
input n_54;
input n_502;
input n_328;
input n_534;
input n_488;
input n_429;
input n_373;
input n_87;
input n_195;
input n_285;
input n_497;
input n_85;
input n_99;
input n_257;
input n_13;
input n_203;
input n_286;
input n_254;
input n_207;
input n_242;
input n_19;
input n_47;
input n_29;
input n_75;
input n_401;
input n_324;
input n_335;
input n_430;
input n_463;
input n_545;
input n_489;
input n_205;
input n_120;
input n_251;
input n_301;
input n_274;
input n_110;
input n_151;
input n_412;
input n_81;
input n_36;
input n_26;
input n_55;
input n_267;
input n_438;
input n_339;
input n_315;
input n_434;
input n_515;
input n_64;
input n_288;
input n_427;
input n_479;
input n_496;
input n_422;
input n_135;
input n_165;
input n_351;
input n_437;
input n_259;
input n_177;
input n_540;
input n_514;
input n_528;
input n_391;
input n_457;
input n_364;
input n_295;
input n_385;
input n_388;
input n_190;
input n_262;
input n_484;
input n_187;
input n_501;
input n_531;
input n_60;
input n_361;
input n_508;
input n_379;
input n_170;
input n_332;
input n_336;
input n_12;
input n_398;
input n_410;
input n_566;
input n_554;
input n_194;
input n_171;
input n_192;
input n_57;
input n_169;
input n_51;
input n_283;

output n_2623;

wire n_992;
wire n_2542;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_2576;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_1212;
wire n_726;
wire n_2157;
wire n_2332;
wire n_700;
wire n_1307;
wire n_2003;
wire n_1038;
wire n_1581;
wire n_1003;
wire n_1237;
wire n_1061;
wire n_2353;
wire n_2534;
wire n_1357;
wire n_1853;
wire n_783;
wire n_2451;
wire n_1738;
wire n_2243;
wire n_798;
wire n_1575;
wire n_1854;
wire n_2324;
wire n_1923;
wire n_1342;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_2260;
wire n_1708;
wire n_677;
wire n_805;
wire n_1151;
wire n_1739;
wire n_2051;
wire n_2317;
wire n_1380;
wire n_2359;
wire n_1402;
wire n_2557;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_2405;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1991;
wire n_2570;
wire n_2179;
wire n_2386;
wire n_1724;
wire n_1032;
wire n_2336;
wire n_1247;
wire n_1547;
wire n_2521;
wire n_1553;
wire n_893;
wire n_1099;
wire n_2491;
wire n_1264;
wire n_1192;
wire n_1844;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_2211;
wire n_1370;
wire n_1786;
wire n_2382;
wire n_2291;
wire n_830;
wire n_2299;
wire n_873;
wire n_1371;
wire n_1285;
wire n_1985;
wire n_2184;
wire n_1803;
wire n_1172;
wire n_852;
wire n_2509;
wire n_2513;
wire n_1590;
wire n_1532;
wire n_2313;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_1711;
wire n_2247;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_2344;
wire n_1579;
wire n_2365;
wire n_2470;
wire n_2321;
wire n_1263;
wire n_2019;
wire n_836;
wire n_2074;
wire n_2447;
wire n_2129;
wire n_2340;
wire n_1261;
wire n_945;
wire n_2286;
wire n_1649;
wire n_2094;
wire n_2018;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_2356;
wire n_2399;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_2013;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_2044;
wire n_1954;
wire n_1735;
wire n_2510;
wire n_1541;
wire n_1300;
wire n_641;
wire n_2480;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_2212;
wire n_758;
wire n_1455;
wire n_2418;
wire n_1163;
wire n_1180;
wire n_2256;
wire n_2582;
wire n_943;
wire n_1798;
wire n_1550;
wire n_1591;
wire n_772;
wire n_1344;
wire n_2495;
wire n_666;
wire n_940;
wire n_770;
wire n_1781;
wire n_1971;
wire n_2090;
wire n_2058;
wire n_2603;
wire n_2173;
wire n_2004;
wire n_1106;
wire n_886;
wire n_1471;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_2394;
wire n_2108;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_2124;
wire n_2378;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_2155;
wire n_1445;
wire n_2364;
wire n_2551;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_1231;
wire n_2599;
wire n_1978;
wire n_2085;
wire n_917;
wire n_2370;
wire n_2612;
wire n_907;
wire n_1446;
wire n_2591;
wire n_659;
wire n_1815;
wire n_2214;
wire n_913;
wire n_1658;
wire n_2593;
wire n_808;
wire n_867;
wire n_1230;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_2613;
wire n_1333;
wire n_2496;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_2011;
wire n_2277;
wire n_1558;
wire n_1732;
wire n_2300;
wire n_699;
wire n_1986;
wire n_2397;
wire n_824;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_2113;
wire n_1918;
wire n_2190;
wire n_1843;
wire n_619;
wire n_2268;
wire n_1367;
wire n_1336;
wire n_813;
wire n_1909;
wire n_2080;
wire n_1481;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_2104;
wire n_645;
wire n_1381;
wire n_1699;
wire n_916;
wire n_2093;
wire n_2207;
wire n_1970;
wire n_608;
wire n_2101;
wire n_630;
wire n_2059;
wire n_2198;
wire n_2073;
wire n_2273;
wire n_2546;
wire n_792;
wire n_2522;
wire n_1328;
wire n_1957;
wire n_2616;
wire n_1907;
wire n_2529;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_982;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_932;
wire n_1876;
wire n_1895;
wire n_2123;
wire n_1697;
wire n_2143;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_993;
wire n_689;
wire n_2031;
wire n_2130;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_2228;
wire n_1988;
wire n_1278;
wire n_2455;
wire n_2469;
wire n_1064;
wire n_1396;
wire n_634;
wire n_2355;
wire n_966;
wire n_764;
wire n_1663;
wire n_2009;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_2245;
wire n_2068;
wire n_1107;
wire n_2457;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_2580;
wire n_882;
wire n_2176;
wire n_2072;
wire n_1354;
wire n_1875;
wire n_1865;
wire n_2459;
wire n_1701;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_1563;
wire n_1912;
wire n_2434;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_1167;
wire n_1359;
wire n_2428;
wire n_674;
wire n_871;
wire n_922;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_2028;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_1165;
wire n_702;
wire n_2008;
wire n_2192;
wire n_2254;
wire n_2345;
wire n_1926;
wire n_1175;
wire n_1386;
wire n_2311;
wire n_1896;
wire n_1747;
wire n_1012;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_2350;
wire n_2453;
wire n_2193;
wire n_1655;
wire n_835;
wire n_928;
wire n_1214;
wire n_1801;
wire n_690;
wire n_850;
wire n_1886;
wire n_2092;
wire n_2347;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_2514;
wire n_2206;
wire n_604;
wire n_2319;
wire n_2519;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_2467;
wire n_2602;
wire n_2468;
wire n_1124;
wire n_1624;
wire n_2096;
wire n_1965;
wire n_2476;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_1082;
wire n_1317;
wire n_593;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_2377;
wire n_701;
wire n_2178;
wire n_950;
wire n_2036;
wire n_2152;
wire n_1709;
wire n_2411;
wire n_2525;
wire n_1825;
wire n_2393;
wire n_1757;
wire n_1796;
wire n_1792;
wire n_891;
wire n_2067;
wire n_2136;
wire n_2409;
wire n_2082;
wire n_2252;
wire n_1412;
wire n_2497;
wire n_949;
wire n_1630;
wire n_678;
wire n_2075;
wire n_2194;
wire n_2619;
wire n_1987;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_2271;
wire n_1008;
wire n_760;
wire n_1546;
wire n_2583;
wire n_590;
wire n_2606;
wire n_2279;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_1990;
wire n_2391;
wire n_2431;
wire n_694;
wire n_2150;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_2078;
wire n_595;
wire n_627;
wire n_1767;
wire n_1779;
wire n_1465;
wire n_2622;
wire n_1858;
wire n_1044;
wire n_2165;
wire n_2133;
wire n_1712;
wire n_1391;
wire n_1523;
wire n_2558;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_2349;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_815;
wire n_1100;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_2493;
wire n_673;
wire n_2230;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_2145;
wire n_1968;
wire n_898;
wire n_1952;
wire n_865;
wire n_2573;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_2535;
wire n_1364;
wire n_2436;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_2151;
wire n_1451;
wire n_963;
wire n_639;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_2341;
wire n_685;
wire n_1765;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_2537;
wire n_2554;
wire n_996;
wire n_1308;
wire n_2089;
wire n_1376;
wire n_1513;
wire n_791;
wire n_1913;
wire n_837;
wire n_2097;
wire n_2170;
wire n_1488;
wire n_1808;
wire n_948;
wire n_2517;
wire n_704;
wire n_2148;
wire n_977;
wire n_2339;
wire n_1005;
wire n_1947;
wire n_1788;
wire n_1999;
wire n_622;
wire n_2590;
wire n_1469;
wire n_2060;
wire n_2608;
wire n_1838;
wire n_1835;
wire n_1766;
wire n_1776;
wire n_1959;
wire n_2002;
wire n_2138;
wire n_765;
wire n_987;
wire n_1492;
wire n_2414;
wire n_1340;
wire n_1771;
wire n_2316;
wire n_631;
wire n_720;
wire n_842;
wire n_2262;
wire n_1707;
wire n_2239;
wire n_1432;
wire n_2208;
wire n_843;
wire n_656;
wire n_989;
wire n_2604;
wire n_2407;
wire n_1277;
wire n_797;
wire n_1473;
wire n_2191;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_2574;
wire n_899;
wire n_738;
wire n_2012;
wire n_1304;
wire n_1035;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_2134;
wire n_1529;
wire n_2335;
wire n_2473;
wire n_1022;
wire n_614;
wire n_2069;
wire n_2307;
wire n_2362;
wire n_684;
wire n_2539;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_2297;
wire n_1181;
wire n_2119;
wire n_1822;
wire n_947;
wire n_1117;
wire n_2489;
wire n_1087;
wire n_1448;
wire n_1992;
wire n_648;
wire n_657;
wire n_1049;
wire n_2445;
wire n_2057;
wire n_2103;
wire n_2605;
wire n_1666;
wire n_1505;
wire n_803;
wire n_1717;
wire n_926;
wire n_1817;
wire n_2449;
wire n_927;
wire n_2610;
wire n_1849;
wire n_919;
wire n_1698;
wire n_2231;
wire n_929;
wire n_2520;
wire n_1228;
wire n_1568;
wire n_1490;
wire n_2372;
wire n_777;
wire n_1299;
wire n_1183;
wire n_1436;
wire n_2251;
wire n_1384;
wire n_2494;
wire n_2501;
wire n_2238;
wire n_2368;
wire n_1070;
wire n_2403;
wire n_998;
wire n_717;
wire n_1665;
wire n_2524;
wire n_1383;
wire n_2460;
wire n_1178;
wire n_2127;
wire n_1424;
wire n_2338;
wire n_1073;
wire n_1000;
wire n_796;
wire n_1195;
wire n_2137;
wire n_1626;
wire n_1507;
wire n_2482;
wire n_2532;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_2481;
wire n_912;
wire n_1857;
wire n_1519;
wire n_2144;
wire n_745;
wire n_1284;
wire n_1604;
wire n_2296;
wire n_2424;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_2354;
wire n_2589;
wire n_1395;
wire n_2110;
wire n_2199;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_931;
wire n_1021;
wire n_683;
wire n_1207;
wire n_811;
wire n_2442;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_2064;
wire n_880;
wire n_2053;
wire n_2259;
wire n_2121;
wire n_2545;
wire n_889;
wire n_2432;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_2294;
wire n_1363;
wire n_2581;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_2218;
wire n_2435;
wire n_954;
wire n_864;
wire n_2504;
wire n_1110;
wire n_2213;
wire n_1410;
wire n_2389;
wire n_1440;
wire n_2132;
wire n_2063;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_1483;
wire n_1834;
wire n_2331;
wire n_1372;
wire n_2292;
wire n_2330;
wire n_1457;
wire n_1719;
wire n_1339;
wire n_1787;
wire n_2475;
wire n_2511;
wire n_1993;
wire n_2281;
wire n_1427;
wire n_2416;
wire n_2617;
wire n_1466;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_1141;
wire n_1268;
wire n_1939;
wire n_2030;
wire n_1769;
wire n_1220;
wire n_2323;
wire n_1893;
wire n_2209;
wire n_2301;
wire n_2387;
wire n_1755;
wire n_1602;
wire n_2421;
wire n_1136;
wire n_2618;
wire n_2025;
wire n_2357;
wire n_2464;
wire n_1125;
wire n_970;
wire n_2488;
wire n_2224;
wire n_1980;
wire n_1159;
wire n_995;
wire n_642;
wire n_2329;
wire n_1092;
wire n_2237;
wire n_1060;
wire n_1951;
wire n_2250;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_2115;
wire n_2410;
wire n_2552;
wire n_1053;
wire n_2374;
wire n_1681;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_2596;
wire n_2274;
wire n_775;
wire n_651;
wire n_1153;
wire n_1618;
wire n_1531;
wire n_1185;
wire n_2384;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_2585;
wire n_2621;
wire n_1653;
wire n_2352;
wire n_1679;
wire n_1625;
wire n_2601;
wire n_2160;
wire n_1453;
wire n_2146;
wire n_2226;
wire n_2131;
wire n_2502;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_2556;
wire n_1315;
wire n_1647;
wire n_2575;
wire n_1224;
wire n_2306;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_2462;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_1617;
wire n_1470;
wire n_2550;
wire n_1243;
wire n_848;
wire n_1096;
wire n_2249;
wire n_1091;
wire n_1917;
wire n_2000;
wire n_1580;
wire n_2227;
wire n_2270;
wire n_1425;
wire n_1881;
wire n_1267;
wire n_1281;
wire n_1806;
wire n_983;
wire n_2023;
wire n_2572;
wire n_2204;
wire n_1520;
wire n_2159;
wire n_906;
wire n_1390;
wire n_688;
wire n_2289;
wire n_1077;
wire n_1733;
wire n_2315;
wire n_1419;
wire n_1731;
wire n_2158;
wire n_2087;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_2135;
wire n_1645;
wire n_1832;
wire n_1687;
wire n_1439;
wire n_2328;
wire n_1323;
wire n_2202;
wire n_858;
wire n_2049;
wire n_1331;
wire n_613;
wire n_736;
wire n_956;
wire n_960;
wire n_2276;
wire n_663;
wire n_856;
wire n_2100;
wire n_778;
wire n_1668;
wire n_1134;
wire n_1129;
wire n_602;
wire n_1696;
wire n_1995;
wire n_1594;
wire n_2181;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_2379;
wire n_1905;
wire n_2016;
wire n_2343;
wire n_793;
wire n_1593;
wire n_762;
wire n_1202;
wire n_1030;
wire n_1937;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_2515;
wire n_1744;
wire n_828;
wire n_2139;
wire n_2142;
wire n_607;
wire n_1551;
wire n_2448;
wire n_1103;
wire n_2555;
wire n_2219;
wire n_1203;
wire n_820;
wire n_2327;
wire n_951;
wire n_2201;
wire n_952;
wire n_725;
wire n_999;
wire n_1254;
wire n_2420;
wire n_994;
wire n_2263;
wire n_2304;
wire n_1508;
wire n_2487;
wire n_732;
wire n_974;
wire n_2240;
wire n_2278;
wire n_2538;
wire n_724;
wire n_2597;
wire n_2375;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_1871;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_1549;
wire n_1510;
wire n_892;
wire n_768;
wire n_1468;
wire n_1859;
wire n_2102;
wire n_2563;
wire n_1095;
wire n_2024;
wire n_1595;
wire n_2156;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_2598;
wire n_597;
wire n_1270;
wire n_2549;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_2153;
wire n_2544;
wire n_2381;
wire n_1847;
wire n_2052;
wire n_2302;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_923;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_2526;
wire n_2423;
wire n_1057;
wire n_2548;
wire n_603;
wire n_991;
wire n_1657;
wire n_1126;
wire n_2412;
wire n_1997;
wire n_710;
wire n_1108;
wire n_1818;
wire n_2439;
wire n_2404;
wire n_1182;
wire n_1298;
wire n_2559;
wire n_2177;
wire n_2595;
wire n_2088;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_2061;
wire n_1686;
wire n_2337;
wire n_2401;
wire n_1356;
wire n_1589;
wire n_2309;
wire n_2607;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_2452;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_2499;
wire n_1622;
wire n_1586;
wire n_2543;
wire n_2264;
wire n_1694;
wire n_1535;
wire n_2486;
wire n_2571;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_1983;
wire n_1938;
wire n_2498;
wire n_2220;
wire n_2577;
wire n_1262;
wire n_2472;
wire n_1891;
wire n_2171;
wire n_1213;
wire n_2235;
wire n_1350;
wire n_1673;
wire n_2232;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_2392;
wire n_2037;
wire n_2298;
wire n_782;
wire n_2326;
wire n_1539;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_2305;
wire n_2120;
wire n_1472;
wire n_2050;
wire n_2373;
wire n_2164;
wire n_2402;
wire n_2225;
wire n_1081;
wire n_1870;
wire n_1692;
wire n_1084;
wire n_800;
wire n_1171;
wire n_2169;
wire n_2371;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_2006;
wire n_1491;
wire n_2187;
wire n_662;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_2244;
wire n_2586;
wire n_1684;
wire n_921;
wire n_2446;
wire n_1346;
wire n_711;
wire n_1642;
wire n_1352;
wire n_937;
wire n_2257;
wire n_1682;
wire n_2017;
wire n_1695;
wire n_1828;
wire n_2046;
wire n_2272;
wire n_2200;
wire n_650;
wire n_1046;
wire n_2560;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_2376;
wire n_1406;
wire n_1332;
wire n_624;
wire n_962;
wire n_1041;
wire n_2346;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_2342;
wire n_2167;
wire n_2084;
wire n_2541;
wire n_654;
wire n_2518;
wire n_2458;
wire n_1222;
wire n_599;
wire n_776;
wire n_1823;
wire n_2479;
wire n_1974;
wire n_2456;
wire n_1720;
wire n_2527;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_1341;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_2314;
wire n_942;
wire n_1524;
wire n_2229;
wire n_1964;
wire n_2288;
wire n_1920;
wire n_2099;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_2007;
wire n_2039;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_2258;
wire n_1640;
wire n_804;
wire n_1846;
wire n_2406;
wire n_2390;
wire n_806;
wire n_959;
wire n_879;
wire n_2310;
wire n_2506;
wire n_2141;
wire n_2562;
wire n_1343;
wire n_1522;
wire n_1782;
wire n_2383;
wire n_1676;
wire n_833;
wire n_1830;
wire n_2351;
wire n_1567;
wire n_1319;
wire n_707;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_2536;
wire n_2196;
wire n_1633;
wire n_2195;
wire n_787;
wire n_2172;
wire n_1416;
wire n_1528;
wire n_2293;
wire n_1146;
wire n_2021;
wire n_2454;
wire n_2114;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_2125;
wire n_2026;
wire n_1282;
wire n_2561;
wire n_2567;
wire n_2322;
wire n_652;
wire n_2154;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_2533;
wire n_1758;
wire n_2283;
wire n_2422;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_2361;
wire n_1373;
wire n_1292;
wire n_2266;
wire n_2427;
wire n_1029;
wire n_1447;
wire n_2388;
wire n_2056;
wire n_790;
wire n_2611;
wire n_1706;
wire n_1498;
wire n_2417;
wire n_1210;
wire n_1248;
wire n_1556;
wire n_902;
wire n_2189;
wire n_2246;
wire n_1047;
wire n_1984;
wire n_2236;
wire n_1385;
wire n_1269;
wire n_1931;
wire n_2083;
wire n_672;
wire n_2441;
wire n_1257;
wire n_1751;
wire n_1375;
wire n_1941;
wire n_2128;
wire n_655;
wire n_1045;
wire n_706;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_2398;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_1804;
wire n_1727;
wire n_2508;
wire n_1019;
wire n_636;
wire n_2054;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_2062;
wire n_2041;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_2070;
wire n_2588;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_2484;
wire n_2348;
wire n_2614;
wire n_2126;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_2253;
wire n_2366;
wire n_646;
wire n_1098;
wire n_1329;
wire n_2045;
wire n_817;
wire n_2261;
wire n_2216;
wire n_2210;
wire n_897;
wire n_846;
wire n_2066;
wire n_841;
wire n_1476;
wire n_2516;
wire n_1001;
wire n_1800;
wire n_2241;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_1191;
wire n_1826;
wire n_1023;
wire n_1882;
wire n_1118;
wire n_1076;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_2369;
wire n_1592;
wire n_855;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_853;
wire n_695;
wire n_1542;
wire n_2587;
wire n_875;
wire n_680;
wire n_1678;
wire n_2569;
wire n_661;
wire n_2400;
wire n_1716;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_2122;
wire n_2109;
wire n_1435;
wire n_969;
wire n_988;
wire n_2140;
wire n_1065;
wire n_2507;
wire n_1401;
wire n_2358;
wire n_1255;
wire n_1516;
wire n_1536;
wire n_2163;
wire n_2186;
wire n_2029;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_1074;
wire n_698;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_955;
wire n_739;
wire n_1379;
wire n_2528;
wire n_1338;
wire n_1097;
wire n_2395;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_769;
wire n_2380;
wire n_676;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_2295;
wire n_814;
wire n_1643;
wire n_2020;
wire n_2500;
wire n_2269;
wire n_1729;
wire n_669;
wire n_2290;
wire n_2048;
wire n_2005;
wire n_747;
wire n_2565;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_691;
wire n_2076;
wire n_1408;
wire n_1196;
wire n_1598;
wire n_863;
wire n_2175;
wire n_601;
wire n_2182;
wire n_1283;
wire n_2385;
wire n_918;
wire n_748;
wire n_1114;
wire n_1848;
wire n_1147;
wire n_763;
wire n_1785;
wire n_1754;
wire n_2149;
wire n_2396;
wire n_1506;
wire n_2584;
wire n_1652;
wire n_1812;
wire n_957;
wire n_1994;
wire n_895;
wire n_866;
wire n_1227;
wire n_2450;
wire n_2485;
wire n_2284;
wire n_2566;
wire n_2287;
wire n_744;
wire n_971;
wire n_946;
wire n_1303;
wire n_761;
wire n_1205;
wire n_2492;
wire n_1258;
wire n_2438;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_2463;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_2180;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_844;
wire n_1017;
wire n_2117;
wire n_2234;
wire n_1083;
wire n_1561;
wire n_930;
wire n_888;
wire n_2275;
wire n_1112;
wire n_2465;
wire n_2620;
wire n_2081;
wire n_2168;
wire n_2568;
wire n_2022;
wire n_1945;
wire n_2203;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_2112;
wire n_2255;
wire n_1464;
wire n_653;
wire n_1737;
wire n_2430;
wire n_1414;
wire n_908;
wire n_752;
wire n_944;
wire n_2034;
wire n_1028;
wire n_2106;
wire n_2265;
wire n_2615;
wire n_1922;
wire n_2032;
wire n_1011;
wire n_2474;
wire n_1566;
wire n_1215;
wire n_2444;
wire n_839;
wire n_2437;
wire n_708;
wire n_1973;
wire n_2267;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_2205;
wire n_1104;
wire n_1058;
wire n_854;
wire n_2312;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_2242;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_2222;
wire n_712;
wire n_1276;
wire n_2015;
wire n_2118;
wire n_2111;
wire n_2466;
wire n_2530;
wire n_1148;
wire n_2188;
wire n_2505;
wire n_1989;
wire n_1161;
wire n_2609;
wire n_1085;
wire n_2014;
wire n_2042;
wire n_1239;
wire n_771;
wire n_1584;
wire n_2425;
wire n_924;
wire n_1582;
wire n_2318;
wire n_2408;
wire n_1149;
wire n_1184;
wire n_2483;
wire n_719;
wire n_1972;
wire n_2592;
wire n_1525;
wire n_2594;
wire n_1585;
wire n_1851;
wire n_1799;
wire n_1090;
wire n_2147;
wire n_2564;
wire n_592;
wire n_1816;
wire n_2503;
wire n_2433;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_984;
wire n_2600;
wire n_1829;
wire n_2035;
wire n_1450;
wire n_1638;
wire n_868;
wire n_859;
wire n_2033;
wire n_735;
wire n_1789;
wire n_2531;
wire n_1770;
wire n_878;
wire n_620;
wire n_2523;
wire n_1218;
wire n_2413;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_1144;
wire n_2071;
wire n_2429;
wire n_985;
wire n_2233;
wire n_2440;
wire n_997;
wire n_1710;
wire n_2161;
wire n_1301;
wire n_802;
wire n_980;
wire n_1306;
wire n_2010;
wire n_2282;
wire n_1651;
wire n_1198;
wire n_2360;
wire n_2047;
wire n_2095;
wire n_1609;
wire n_2174;
wire n_2334;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1998;
wire n_1574;
wire n_2426;
wire n_2490;
wire n_756;
wire n_2303;
wire n_1619;
wire n_2478;
wire n_1981;
wire n_2285;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_1552;
wire n_1996;
wire n_2367;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_2043;
wire n_1480;
wire n_1158;
wire n_2248;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_2363;
wire n_2578;
wire n_849;
wire n_753;
wire n_1753;
wire n_2471;
wire n_2540;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_2197;
wire n_2217;
wire n_2065;
wire n_861;
wire n_857;
wire n_967;
wire n_2215;
wire n_2461;
wire n_2001;
wire n_2107;
wire n_1884;
wire n_2040;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_2221;
wire n_1260;
wire n_1819;
wire n_2055;
wire n_1010;
wire n_2553;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_2038;
wire n_812;
wire n_1131;
wire n_1761;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_2477;
wire n_1557;
wire n_1888;
wire n_2280;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_2325;
wire n_670;
wire n_1850;
wire n_1898;
wire n_2443;
wire n_2308;
wire n_2162;
wire n_1868;
wire n_2333;
wire n_2079;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_2512;
wire n_1365;
wire n_1417;
wire n_1242;
wire n_2185;
wire n_2086;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_2166;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_2077;
wire n_784;
wire n_1059;
wire n_1197;
wire n_2579;
wire n_722;
wire n_862;
wire n_2105;
wire n_2098;
wire n_1423;
wire n_1935;
wire n_2027;
wire n_2223;
wire n_2091;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_2547;
wire n_2415;
wire n_900;
wire n_1449;
wire n_827;
wire n_1025;
wire n_2419;
wire n_2116;
wire n_2320;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_2183;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

CKINVDCx5p33_ASAP7_75t_R g589 ( 
.A(n_453),
.Y(n_589)
);

CKINVDCx5p33_ASAP7_75t_R g590 ( 
.A(n_583),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_140),
.Y(n_591)
);

CKINVDCx5p33_ASAP7_75t_R g592 ( 
.A(n_472),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_31),
.Y(n_593)
);

CKINVDCx5p33_ASAP7_75t_R g594 ( 
.A(n_326),
.Y(n_594)
);

CKINVDCx5p33_ASAP7_75t_R g595 ( 
.A(n_223),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_70),
.Y(n_596)
);

CKINVDCx5p33_ASAP7_75t_R g597 ( 
.A(n_493),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_54),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_559),
.Y(n_599)
);

CKINVDCx14_ASAP7_75t_R g600 ( 
.A(n_83),
.Y(n_600)
);

CKINVDCx20_ASAP7_75t_R g601 ( 
.A(n_522),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_206),
.Y(n_602)
);

BUFx2_ASAP7_75t_L g603 ( 
.A(n_263),
.Y(n_603)
);

CKINVDCx5p33_ASAP7_75t_R g604 ( 
.A(n_564),
.Y(n_604)
);

CKINVDCx5p33_ASAP7_75t_R g605 ( 
.A(n_6),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_474),
.Y(n_606)
);

INVx2_ASAP7_75t_SL g607 ( 
.A(n_357),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_127),
.Y(n_608)
);

INVx2_ASAP7_75t_SL g609 ( 
.A(n_113),
.Y(n_609)
);

BUFx5_ASAP7_75t_L g610 ( 
.A(n_366),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_217),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_301),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_469),
.Y(n_613)
);

BUFx10_ASAP7_75t_L g614 ( 
.A(n_262),
.Y(n_614)
);

BUFx6f_ASAP7_75t_L g615 ( 
.A(n_314),
.Y(n_615)
);

CKINVDCx5p33_ASAP7_75t_R g616 ( 
.A(n_452),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_510),
.Y(n_617)
);

CKINVDCx5p33_ASAP7_75t_R g618 ( 
.A(n_247),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_91),
.Y(n_619)
);

CKINVDCx20_ASAP7_75t_R g620 ( 
.A(n_87),
.Y(n_620)
);

CKINVDCx20_ASAP7_75t_R g621 ( 
.A(n_198),
.Y(n_621)
);

CKINVDCx14_ASAP7_75t_R g622 ( 
.A(n_254),
.Y(n_622)
);

BUFx2_ASAP7_75t_L g623 ( 
.A(n_459),
.Y(n_623)
);

CKINVDCx5p33_ASAP7_75t_R g624 ( 
.A(n_446),
.Y(n_624)
);

INVx1_ASAP7_75t_SL g625 ( 
.A(n_34),
.Y(n_625)
);

BUFx2_ASAP7_75t_L g626 ( 
.A(n_498),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_154),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_376),
.Y(n_628)
);

CKINVDCx5p33_ASAP7_75t_R g629 ( 
.A(n_388),
.Y(n_629)
);

CKINVDCx5p33_ASAP7_75t_R g630 ( 
.A(n_7),
.Y(n_630)
);

CKINVDCx5p33_ASAP7_75t_R g631 ( 
.A(n_9),
.Y(n_631)
);

CKINVDCx5p33_ASAP7_75t_R g632 ( 
.A(n_439),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_273),
.Y(n_633)
);

INVxp67_ASAP7_75t_L g634 ( 
.A(n_192),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_14),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_430),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_514),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_263),
.Y(n_638)
);

BUFx5_ASAP7_75t_L g639 ( 
.A(n_267),
.Y(n_639)
);

CKINVDCx20_ASAP7_75t_R g640 ( 
.A(n_404),
.Y(n_640)
);

INVx1_ASAP7_75t_L g641 ( 
.A(n_22),
.Y(n_641)
);

CKINVDCx5p33_ASAP7_75t_R g642 ( 
.A(n_310),
.Y(n_642)
);

BUFx10_ASAP7_75t_L g643 ( 
.A(n_417),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_282),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_228),
.Y(n_645)
);

CKINVDCx5p33_ASAP7_75t_R g646 ( 
.A(n_548),
.Y(n_646)
);

CKINVDCx5p33_ASAP7_75t_R g647 ( 
.A(n_396),
.Y(n_647)
);

INVx2_ASAP7_75t_L g648 ( 
.A(n_232),
.Y(n_648)
);

CKINVDCx5p33_ASAP7_75t_R g649 ( 
.A(n_27),
.Y(n_649)
);

CKINVDCx5p33_ASAP7_75t_R g650 ( 
.A(n_495),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_200),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_355),
.Y(n_652)
);

CKINVDCx5p33_ASAP7_75t_R g653 ( 
.A(n_95),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_328),
.Y(n_654)
);

CKINVDCx5p33_ASAP7_75t_R g655 ( 
.A(n_454),
.Y(n_655)
);

CKINVDCx5p33_ASAP7_75t_R g656 ( 
.A(n_35),
.Y(n_656)
);

CKINVDCx5p33_ASAP7_75t_R g657 ( 
.A(n_107),
.Y(n_657)
);

CKINVDCx5p33_ASAP7_75t_R g658 ( 
.A(n_303),
.Y(n_658)
);

CKINVDCx20_ASAP7_75t_R g659 ( 
.A(n_254),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_456),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_48),
.Y(n_661)
);

CKINVDCx5p33_ASAP7_75t_R g662 ( 
.A(n_323),
.Y(n_662)
);

CKINVDCx5p33_ASAP7_75t_R g663 ( 
.A(n_257),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_188),
.Y(n_664)
);

CKINVDCx5p33_ASAP7_75t_R g665 ( 
.A(n_495),
.Y(n_665)
);

INVx2_ASAP7_75t_L g666 ( 
.A(n_516),
.Y(n_666)
);

INVx1_ASAP7_75t_SL g667 ( 
.A(n_135),
.Y(n_667)
);

CKINVDCx5p33_ASAP7_75t_R g668 ( 
.A(n_380),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_563),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_253),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_441),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_170),
.Y(n_672)
);

CKINVDCx5p33_ASAP7_75t_R g673 ( 
.A(n_503),
.Y(n_673)
);

CKINVDCx5p33_ASAP7_75t_R g674 ( 
.A(n_446),
.Y(n_674)
);

CKINVDCx5p33_ASAP7_75t_R g675 ( 
.A(n_24),
.Y(n_675)
);

CKINVDCx5p33_ASAP7_75t_R g676 ( 
.A(n_437),
.Y(n_676)
);

BUFx3_ASAP7_75t_L g677 ( 
.A(n_524),
.Y(n_677)
);

INVx1_ASAP7_75t_SL g678 ( 
.A(n_251),
.Y(n_678)
);

CKINVDCx5p33_ASAP7_75t_R g679 ( 
.A(n_463),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_182),
.Y(n_680)
);

CKINVDCx5p33_ASAP7_75t_R g681 ( 
.A(n_570),
.Y(n_681)
);

CKINVDCx5p33_ASAP7_75t_R g682 ( 
.A(n_214),
.Y(n_682)
);

INVx1_ASAP7_75t_L g683 ( 
.A(n_407),
.Y(n_683)
);

CKINVDCx5p33_ASAP7_75t_R g684 ( 
.A(n_402),
.Y(n_684)
);

CKINVDCx5p33_ASAP7_75t_R g685 ( 
.A(n_508),
.Y(n_685)
);

CKINVDCx5p33_ASAP7_75t_R g686 ( 
.A(n_315),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_63),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_34),
.Y(n_688)
);

CKINVDCx5p33_ASAP7_75t_R g689 ( 
.A(n_519),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_496),
.Y(n_690)
);

INVx1_ASAP7_75t_SL g691 ( 
.A(n_507),
.Y(n_691)
);

CKINVDCx20_ASAP7_75t_R g692 ( 
.A(n_575),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_216),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_285),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_338),
.Y(n_695)
);

CKINVDCx5p33_ASAP7_75t_R g696 ( 
.A(n_578),
.Y(n_696)
);

CKINVDCx16_ASAP7_75t_R g697 ( 
.A(n_463),
.Y(n_697)
);

CKINVDCx5p33_ASAP7_75t_R g698 ( 
.A(n_297),
.Y(n_698)
);

CKINVDCx5p33_ASAP7_75t_R g699 ( 
.A(n_58),
.Y(n_699)
);

INVx1_ASAP7_75t_L g700 ( 
.A(n_452),
.Y(n_700)
);

INVx1_ASAP7_75t_SL g701 ( 
.A(n_467),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_586),
.Y(n_702)
);

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_498),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_474),
.Y(n_704)
);

CKINVDCx5p33_ASAP7_75t_R g705 ( 
.A(n_356),
.Y(n_705)
);

CKINVDCx5p33_ASAP7_75t_R g706 ( 
.A(n_353),
.Y(n_706)
);

CKINVDCx5p33_ASAP7_75t_R g707 ( 
.A(n_291),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_577),
.Y(n_708)
);

CKINVDCx14_ASAP7_75t_R g709 ( 
.A(n_103),
.Y(n_709)
);

CKINVDCx5p33_ASAP7_75t_R g710 ( 
.A(n_381),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_126),
.Y(n_711)
);

INVx2_ASAP7_75t_L g712 ( 
.A(n_386),
.Y(n_712)
);

CKINVDCx20_ASAP7_75t_R g713 ( 
.A(n_366),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_380),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_9),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_456),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_269),
.Y(n_717)
);

CKINVDCx5p33_ASAP7_75t_R g718 ( 
.A(n_282),
.Y(n_718)
);

CKINVDCx16_ASAP7_75t_R g719 ( 
.A(n_481),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_119),
.Y(n_720)
);

INVx1_ASAP7_75t_SL g721 ( 
.A(n_445),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_287),
.Y(n_722)
);

INVx1_ASAP7_75t_L g723 ( 
.A(n_432),
.Y(n_723)
);

CKINVDCx5p33_ASAP7_75t_R g724 ( 
.A(n_417),
.Y(n_724)
);

CKINVDCx5p33_ASAP7_75t_R g725 ( 
.A(n_402),
.Y(n_725)
);

INVx2_ASAP7_75t_L g726 ( 
.A(n_243),
.Y(n_726)
);

CKINVDCx5p33_ASAP7_75t_R g727 ( 
.A(n_333),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_258),
.Y(n_728)
);

INVx2_ASAP7_75t_SL g729 ( 
.A(n_587),
.Y(n_729)
);

INVx2_ASAP7_75t_SL g730 ( 
.A(n_87),
.Y(n_730)
);

CKINVDCx20_ASAP7_75t_R g731 ( 
.A(n_433),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_180),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_473),
.Y(n_733)
);

CKINVDCx5p33_ASAP7_75t_R g734 ( 
.A(n_323),
.Y(n_734)
);

CKINVDCx20_ASAP7_75t_R g735 ( 
.A(n_262),
.Y(n_735)
);

CKINVDCx5p33_ASAP7_75t_R g736 ( 
.A(n_491),
.Y(n_736)
);

CKINVDCx5p33_ASAP7_75t_R g737 ( 
.A(n_545),
.Y(n_737)
);

CKINVDCx16_ASAP7_75t_R g738 ( 
.A(n_45),
.Y(n_738)
);

INVx2_ASAP7_75t_SL g739 ( 
.A(n_235),
.Y(n_739)
);

INVx3_ASAP7_75t_L g740 ( 
.A(n_135),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_264),
.Y(n_741)
);

INVx2_ASAP7_75t_SL g742 ( 
.A(n_115),
.Y(n_742)
);

CKINVDCx5p33_ASAP7_75t_R g743 ( 
.A(n_472),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_151),
.Y(n_744)
);

INVx1_ASAP7_75t_L g745 ( 
.A(n_574),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_424),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_20),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_434),
.Y(n_748)
);

CKINVDCx5p33_ASAP7_75t_R g749 ( 
.A(n_45),
.Y(n_749)
);

BUFx6f_ASAP7_75t_L g750 ( 
.A(n_175),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_62),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_40),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_462),
.Y(n_753)
);

CKINVDCx20_ASAP7_75t_R g754 ( 
.A(n_492),
.Y(n_754)
);

CKINVDCx5p33_ASAP7_75t_R g755 ( 
.A(n_156),
.Y(n_755)
);

CKINVDCx5p33_ASAP7_75t_R g756 ( 
.A(n_203),
.Y(n_756)
);

INVx1_ASAP7_75t_L g757 ( 
.A(n_334),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_409),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_221),
.Y(n_759)
);

INVx1_ASAP7_75t_L g760 ( 
.A(n_485),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_3),
.Y(n_761)
);

BUFx6f_ASAP7_75t_L g762 ( 
.A(n_408),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_66),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_2),
.Y(n_764)
);

CKINVDCx5p33_ASAP7_75t_R g765 ( 
.A(n_211),
.Y(n_765)
);

CKINVDCx5p33_ASAP7_75t_R g766 ( 
.A(n_147),
.Y(n_766)
);

CKINVDCx5p33_ASAP7_75t_R g767 ( 
.A(n_156),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_107),
.Y(n_768)
);

INVx1_ASAP7_75t_L g769 ( 
.A(n_239),
.Y(n_769)
);

CKINVDCx5p33_ASAP7_75t_R g770 ( 
.A(n_555),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_579),
.Y(n_771)
);

BUFx2_ASAP7_75t_L g772 ( 
.A(n_252),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_59),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_357),
.Y(n_774)
);

CKINVDCx16_ASAP7_75t_R g775 ( 
.A(n_486),
.Y(n_775)
);

CKINVDCx5p33_ASAP7_75t_R g776 ( 
.A(n_354),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_378),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_118),
.Y(n_778)
);

CKINVDCx16_ASAP7_75t_R g779 ( 
.A(n_65),
.Y(n_779)
);

INVx1_ASAP7_75t_L g780 ( 
.A(n_435),
.Y(n_780)
);

CKINVDCx14_ASAP7_75t_R g781 ( 
.A(n_73),
.Y(n_781)
);

CKINVDCx5p33_ASAP7_75t_R g782 ( 
.A(n_521),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_192),
.Y(n_783)
);

CKINVDCx20_ASAP7_75t_R g784 ( 
.A(n_269),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_405),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_272),
.Y(n_786)
);

CKINVDCx16_ASAP7_75t_R g787 ( 
.A(n_77),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_208),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_557),
.Y(n_789)
);

CKINVDCx20_ASAP7_75t_R g790 ( 
.A(n_488),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_335),
.Y(n_791)
);

CKINVDCx5p33_ASAP7_75t_R g792 ( 
.A(n_313),
.Y(n_792)
);

BUFx5_ASAP7_75t_L g793 ( 
.A(n_41),
.Y(n_793)
);

CKINVDCx5p33_ASAP7_75t_R g794 ( 
.A(n_529),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_410),
.Y(n_795)
);

BUFx5_ASAP7_75t_L g796 ( 
.A(n_356),
.Y(n_796)
);

CKINVDCx20_ASAP7_75t_R g797 ( 
.A(n_326),
.Y(n_797)
);

INVx2_ASAP7_75t_L g798 ( 
.A(n_487),
.Y(n_798)
);

INVx1_ASAP7_75t_L g799 ( 
.A(n_484),
.Y(n_799)
);

CKINVDCx5p33_ASAP7_75t_R g800 ( 
.A(n_333),
.Y(n_800)
);

CKINVDCx5p33_ASAP7_75t_R g801 ( 
.A(n_389),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_363),
.Y(n_802)
);

CKINVDCx5p33_ASAP7_75t_R g803 ( 
.A(n_331),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_470),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_230),
.Y(n_805)
);

INVx1_ASAP7_75t_SL g806 ( 
.A(n_136),
.Y(n_806)
);

BUFx10_ASAP7_75t_L g807 ( 
.A(n_489),
.Y(n_807)
);

CKINVDCx20_ASAP7_75t_R g808 ( 
.A(n_65),
.Y(n_808)
);

CKINVDCx5p33_ASAP7_75t_R g809 ( 
.A(n_55),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_412),
.Y(n_810)
);

CKINVDCx5p33_ASAP7_75t_R g811 ( 
.A(n_292),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_539),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_271),
.Y(n_813)
);

INVx2_ASAP7_75t_L g814 ( 
.A(n_359),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_260),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_350),
.Y(n_816)
);

BUFx5_ASAP7_75t_L g817 ( 
.A(n_295),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_490),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_83),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_230),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_89),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_404),
.Y(n_822)
);

BUFx3_ASAP7_75t_L g823 ( 
.A(n_414),
.Y(n_823)
);

CKINVDCx5p33_ASAP7_75t_R g824 ( 
.A(n_600),
.Y(n_824)
);

INVx2_ASAP7_75t_L g825 ( 
.A(n_610),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_610),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_610),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_610),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_610),
.Y(n_829)
);

BUFx3_ASAP7_75t_L g830 ( 
.A(n_677),
.Y(n_830)
);

INVx4_ASAP7_75t_R g831 ( 
.A(n_677),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_610),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_610),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_639),
.Y(n_834)
);

BUFx3_ASAP7_75t_L g835 ( 
.A(n_708),
.Y(n_835)
);

CKINVDCx16_ASAP7_75t_R g836 ( 
.A(n_697),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_639),
.Y(n_837)
);

INVxp33_ASAP7_75t_L g838 ( 
.A(n_603),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_639),
.Y(n_839)
);

INVx2_ASAP7_75t_L g840 ( 
.A(n_639),
.Y(n_840)
);

CKINVDCx5p33_ASAP7_75t_R g841 ( 
.A(n_622),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_709),
.Y(n_842)
);

CKINVDCx20_ASAP7_75t_R g843 ( 
.A(n_620),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_639),
.Y(n_844)
);

INVx2_ASAP7_75t_L g845 ( 
.A(n_639),
.Y(n_845)
);

BUFx6f_ASAP7_75t_L g846 ( 
.A(n_708),
.Y(n_846)
);

INVx1_ASAP7_75t_L g847 ( 
.A(n_639),
.Y(n_847)
);

BUFx5_ASAP7_75t_L g848 ( 
.A(n_599),
.Y(n_848)
);

BUFx2_ASAP7_75t_L g849 ( 
.A(n_623),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_793),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_793),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_793),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_793),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_793),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_793),
.Y(n_855)
);

INVx1_ASAP7_75t_SL g856 ( 
.A(n_626),
.Y(n_856)
);

HB1xp67_ASAP7_75t_L g857 ( 
.A(n_719),
.Y(n_857)
);

INVx1_ASAP7_75t_L g858 ( 
.A(n_793),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_796),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_781),
.Y(n_860)
);

INVx2_ASAP7_75t_SL g861 ( 
.A(n_661),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_796),
.Y(n_862)
);

INVxp67_ASAP7_75t_SL g863 ( 
.A(n_740),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_796),
.Y(n_864)
);

HB1xp67_ASAP7_75t_L g865 ( 
.A(n_738),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_796),
.Y(n_866)
);

INVx1_ASAP7_75t_L g867 ( 
.A(n_796),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_796),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_796),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_817),
.Y(n_870)
);

INVxp33_ASAP7_75t_L g871 ( 
.A(n_772),
.Y(n_871)
);

CKINVDCx20_ASAP7_75t_R g872 ( 
.A(n_620),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_817),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_817),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_817),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_817),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_817),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_621),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_817),
.Y(n_879)
);

CKINVDCx16_ASAP7_75t_R g880 ( 
.A(n_775),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_740),
.Y(n_881)
);

CKINVDCx16_ASAP7_75t_R g882 ( 
.A(n_779),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_615),
.Y(n_883)
);

CKINVDCx16_ASAP7_75t_R g884 ( 
.A(n_787),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_740),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_615),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_823),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_823),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_661),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_615),
.Y(n_890)
);

HB1xp67_ASAP7_75t_L g891 ( 
.A(n_608),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_615),
.Y(n_892)
);

INVx1_ASAP7_75t_L g893 ( 
.A(n_750),
.Y(n_893)
);

INVxp67_ASAP7_75t_SL g894 ( 
.A(n_750),
.Y(n_894)
);

CKINVDCx16_ASAP7_75t_R g895 ( 
.A(n_601),
.Y(n_895)
);

INVxp67_ASAP7_75t_SL g896 ( 
.A(n_750),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_750),
.Y(n_897)
);

INVx2_ASAP7_75t_L g898 ( 
.A(n_762),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_762),
.Y(n_899)
);

INVx1_ASAP7_75t_L g900 ( 
.A(n_762),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_762),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_591),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_598),
.Y(n_903)
);

CKINVDCx16_ASAP7_75t_R g904 ( 
.A(n_692),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_606),
.Y(n_905)
);

INVxp33_ASAP7_75t_L g906 ( 
.A(n_619),
.Y(n_906)
);

CKINVDCx14_ASAP7_75t_R g907 ( 
.A(n_614),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_633),
.Y(n_908)
);

CKINVDCx5p33_ASAP7_75t_R g909 ( 
.A(n_589),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_611),
.Y(n_910)
);

INVxp67_ASAP7_75t_L g911 ( 
.A(n_614),
.Y(n_911)
);

CKINVDCx5p33_ASAP7_75t_R g912 ( 
.A(n_592),
.Y(n_912)
);

INVxp33_ASAP7_75t_L g913 ( 
.A(n_636),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_638),
.Y(n_914)
);

INVx1_ASAP7_75t_L g915 ( 
.A(n_641),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_644),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_611),
.Y(n_917)
);

INVx1_ASAP7_75t_L g918 ( 
.A(n_648),
.Y(n_918)
);

BUFx6f_ASAP7_75t_L g919 ( 
.A(n_666),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_621),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_648),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_660),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_660),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_651),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_919),
.Y(n_925)
);

AND2x2_ASAP7_75t_L g926 ( 
.A(n_863),
.B(n_607),
.Y(n_926)
);

INVx3_ASAP7_75t_L g927 ( 
.A(n_919),
.Y(n_927)
);

INVx3_ASAP7_75t_L g928 ( 
.A(n_919),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_895),
.Y(n_929)
);

NOR2xp33_ASAP7_75t_SL g930 ( 
.A(n_856),
.B(n_692),
.Y(n_930)
);

NOR2xp67_ASAP7_75t_L g931 ( 
.A(n_826),
.B(n_729),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_886),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_919),
.Y(n_933)
);

NOR2x1_ASAP7_75t_L g934 ( 
.A(n_883),
.B(n_666),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_919),
.Y(n_935)
);

AND2x2_ASAP7_75t_L g936 ( 
.A(n_830),
.B(n_607),
.Y(n_936)
);

AND2x4_ASAP7_75t_L g937 ( 
.A(n_894),
.B(n_729),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_886),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_896),
.B(n_669),
.Y(n_939)
);

INVx4_ASAP7_75t_L g940 ( 
.A(n_846),
.Y(n_940)
);

INVx3_ASAP7_75t_L g941 ( 
.A(n_825),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_899),
.B(n_669),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_830),
.B(n_637),
.Y(n_943)
);

AND2x4_ASAP7_75t_L g944 ( 
.A(n_846),
.B(n_745),
.Y(n_944)
);

BUFx6f_ASAP7_75t_L g945 ( 
.A(n_892),
.Y(n_945)
);

BUFx6f_ASAP7_75t_L g946 ( 
.A(n_892),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_835),
.B(n_771),
.Y(n_947)
);

NOR2xp33_ASAP7_75t_L g948 ( 
.A(n_824),
.B(n_691),
.Y(n_948)
);

AND2x4_ASAP7_75t_L g949 ( 
.A(n_846),
.B(n_789),
.Y(n_949)
);

INVx5_ASAP7_75t_L g950 ( 
.A(n_846),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_835),
.B(n_609),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_883),
.Y(n_952)
);

AND2x4_ASAP7_75t_L g953 ( 
.A(n_846),
.B(n_693),
.Y(n_953)
);

BUFx3_ASAP7_75t_L g954 ( 
.A(n_887),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_861),
.B(n_590),
.Y(n_955)
);

INVx5_ASAP7_75t_L g956 ( 
.A(n_825),
.Y(n_956)
);

CKINVDCx5p33_ASAP7_75t_R g957 ( 
.A(n_824),
.Y(n_957)
);

INVx1_ASAP7_75t_L g958 ( 
.A(n_898),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_861),
.B(n_604),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_841),
.B(n_614),
.Y(n_960)
);

AND2x4_ASAP7_75t_L g961 ( 
.A(n_881),
.B(n_693),
.Y(n_961)
);

BUFx6f_ASAP7_75t_L g962 ( 
.A(n_898),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_840),
.Y(n_963)
);

NOR2xp33_ASAP7_75t_SL g964 ( 
.A(n_836),
.B(n_640),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_890),
.Y(n_965)
);

AND2x6_ASAP7_75t_L g966 ( 
.A(n_840),
.B(n_712),
.Y(n_966)
);

BUFx6f_ASAP7_75t_L g967 ( 
.A(n_845),
.Y(n_967)
);

NOR2xp33_ASAP7_75t_L g968 ( 
.A(n_841),
.B(n_617),
.Y(n_968)
);

CKINVDCx6p67_ASAP7_75t_R g969 ( 
.A(n_880),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_845),
.Y(n_970)
);

INVx1_ASAP7_75t_L g971 ( 
.A(n_893),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_862),
.Y(n_972)
);

AND2x4_ASAP7_75t_L g973 ( 
.A(n_885),
.B(n_712),
.Y(n_973)
);

NOR2xp33_ASAP7_75t_SL g974 ( 
.A(n_882),
.B(n_640),
.Y(n_974)
);

AND2x4_ASAP7_75t_L g975 ( 
.A(n_897),
.B(n_900),
.Y(n_975)
);

BUFx6f_ASAP7_75t_L g976 ( 
.A(n_862),
.Y(n_976)
);

AND2x4_ASAP7_75t_L g977 ( 
.A(n_901),
.B(n_726),
.Y(n_977)
);

BUFx6f_ASAP7_75t_L g978 ( 
.A(n_869),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_SL g979 ( 
.A(n_842),
.B(n_643),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_910),
.Y(n_980)
);

NOR2x1_ASAP7_75t_L g981 ( 
.A(n_826),
.B(n_652),
.Y(n_981)
);

BUFx12f_ASAP7_75t_L g982 ( 
.A(n_842),
.Y(n_982)
);

NOR2xp33_ASAP7_75t_L g983 ( 
.A(n_860),
.B(n_646),
.Y(n_983)
);

BUFx6f_ASAP7_75t_L g984 ( 
.A(n_869),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_910),
.Y(n_985)
);

NOR2xp33_ASAP7_75t_L g986 ( 
.A(n_860),
.B(n_673),
.Y(n_986)
);

INVx5_ASAP7_75t_L g987 ( 
.A(n_848),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_888),
.B(n_609),
.Y(n_988)
);

BUFx12f_ASAP7_75t_L g989 ( 
.A(n_909),
.Y(n_989)
);

INVx1_ASAP7_75t_L g990 ( 
.A(n_833),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_953),
.Y(n_991)
);

BUFx6f_ASAP7_75t_L g992 ( 
.A(n_933),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_953),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_933),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_937),
.B(n_848),
.Y(n_995)
);

HB1xp67_ASAP7_75t_L g996 ( 
.A(n_936),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_932),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_937),
.B(n_848),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_953),
.Y(n_999)
);

INVxp67_ASAP7_75t_L g1000 ( 
.A(n_930),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_933),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_932),
.Y(n_1002)
);

HB1xp67_ASAP7_75t_L g1003 ( 
.A(n_936),
.Y(n_1003)
);

AND2x2_ASAP7_75t_L g1004 ( 
.A(n_926),
.B(n_951),
.Y(n_1004)
);

BUFx6f_ASAP7_75t_L g1005 ( 
.A(n_933),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_981),
.B(n_902),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_990),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_954),
.Y(n_1008)
);

AND2x2_ASAP7_75t_L g1009 ( 
.A(n_926),
.B(n_889),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_938),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_948),
.B(n_909),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_954),
.Y(n_1012)
);

NOR2xp33_ASAP7_75t_L g1013 ( 
.A(n_968),
.B(n_912),
.Y(n_1013)
);

BUFx6f_ASAP7_75t_L g1014 ( 
.A(n_933),
.Y(n_1014)
);

AOI22xp5_ASAP7_75t_L g1015 ( 
.A1(n_983),
.A2(n_912),
.B1(n_884),
.B2(n_907),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_937),
.B(n_944),
.Y(n_1016)
);

AND2x2_ASAP7_75t_L g1017 ( 
.A(n_951),
.B(n_917),
.Y(n_1017)
);

AND2x6_ASAP7_75t_L g1018 ( 
.A(n_981),
.B(n_944),
.Y(n_1018)
);

INVx2_ASAP7_75t_L g1019 ( 
.A(n_938),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_963),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_986),
.B(n_838),
.Y(n_1021)
);

HB1xp67_ASAP7_75t_L g1022 ( 
.A(n_955),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_975),
.Y(n_1023)
);

NAND2xp5_ASAP7_75t_L g1024 ( 
.A(n_944),
.B(n_848),
.Y(n_1024)
);

INVxp67_ASAP7_75t_L g1025 ( 
.A(n_964),
.Y(n_1025)
);

BUFx6f_ASAP7_75t_L g1026 ( 
.A(n_935),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_949),
.Y(n_1027)
);

BUFx6f_ASAP7_75t_L g1028 ( 
.A(n_935),
.Y(n_1028)
);

BUFx2_ASAP7_75t_L g1029 ( 
.A(n_959),
.Y(n_1029)
);

BUFx6f_ASAP7_75t_L g1030 ( 
.A(n_935),
.Y(n_1030)
);

INVx2_ASAP7_75t_L g1031 ( 
.A(n_963),
.Y(n_1031)
);

XOR2xp5_ASAP7_75t_L g1032 ( 
.A(n_929),
.B(n_843),
.Y(n_1032)
);

CKINVDCx8_ASAP7_75t_R g1033 ( 
.A(n_957),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_952),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_965),
.Y(n_1035)
);

INVx2_ASAP7_75t_L g1036 ( 
.A(n_970),
.Y(n_1036)
);

NOR2xp33_ASAP7_75t_L g1037 ( 
.A(n_960),
.B(n_871),
.Y(n_1037)
);

INVx3_ASAP7_75t_L g1038 ( 
.A(n_935),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_971),
.Y(n_1039)
);

INVx3_ASAP7_75t_L g1040 ( 
.A(n_935),
.Y(n_1040)
);

XNOR2xp5_ASAP7_75t_L g1041 ( 
.A(n_979),
.B(n_843),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_971),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_970),
.Y(n_1043)
);

AND2x4_ASAP7_75t_L g1044 ( 
.A(n_977),
.B(n_903),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_940),
.B(n_848),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_941),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_941),
.Y(n_1047)
);

INVx3_ASAP7_75t_L g1048 ( 
.A(n_967),
.Y(n_1048)
);

BUFx6f_ASAP7_75t_L g1049 ( 
.A(n_967),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_941),
.Y(n_1050)
);

OAI21x1_ASAP7_75t_L g1051 ( 
.A1(n_934),
.A2(n_828),
.B(n_827),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_967),
.Y(n_1052)
);

INVx3_ASAP7_75t_L g1053 ( 
.A(n_967),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_940),
.B(n_925),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_925),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_967),
.Y(n_1056)
);

BUFx6f_ASAP7_75t_L g1057 ( 
.A(n_972),
.Y(n_1057)
);

BUFx6f_ASAP7_75t_L g1058 ( 
.A(n_972),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_925),
.Y(n_1059)
);

NOR2xp33_ASAP7_75t_L g1060 ( 
.A(n_943),
.B(n_857),
.Y(n_1060)
);

AND2x4_ASAP7_75t_L g1061 ( 
.A(n_977),
.B(n_905),
.Y(n_1061)
);

AND2x2_ASAP7_75t_L g1062 ( 
.A(n_988),
.B(n_917),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_977),
.B(n_908),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_972),
.Y(n_1064)
);

AND2x4_ASAP7_75t_L g1065 ( 
.A(n_961),
.B(n_914),
.Y(n_1065)
);

NAND2x1_ASAP7_75t_L g1066 ( 
.A(n_966),
.B(n_831),
.Y(n_1066)
);

BUFx6f_ASAP7_75t_L g1067 ( 
.A(n_972),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_982),
.Y(n_1068)
);

INVx2_ASAP7_75t_L g1069 ( 
.A(n_972),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_988),
.B(n_918),
.Y(n_1070)
);

AOI22xp5_ASAP7_75t_L g1071 ( 
.A1(n_974),
.A2(n_865),
.B1(n_989),
.B2(n_849),
.Y(n_1071)
);

INVx2_ASAP7_75t_L g1072 ( 
.A(n_1031),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_991),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_993),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1011),
.B(n_904),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_SL g1076 ( 
.A(n_995),
.B(n_931),
.Y(n_1076)
);

INVx2_ASAP7_75t_L g1077 ( 
.A(n_1031),
.Y(n_1077)
);

NOR3xp33_ASAP7_75t_L g1078 ( 
.A(n_1037),
.B(n_911),
.C(n_891),
.Y(n_1078)
);

INVx2_ASAP7_75t_L g1079 ( 
.A(n_1036),
.Y(n_1079)
);

NAND2xp5_ASAP7_75t_SL g1080 ( 
.A(n_998),
.B(n_931),
.Y(n_1080)
);

INVx4_ASAP7_75t_L g1081 ( 
.A(n_1049),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_1036),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_993),
.Y(n_1083)
);

NAND2xp33_ASAP7_75t_L g1084 ( 
.A(n_1018),
.B(n_966),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_999),
.Y(n_1085)
);

INVx1_ASAP7_75t_L g1086 ( 
.A(n_999),
.Y(n_1086)
);

AOI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_1004),
.A2(n_942),
.B1(n_939),
.B2(n_989),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_1033),
.Y(n_1088)
);

NOR2xp33_ASAP7_75t_L g1089 ( 
.A(n_1013),
.B(n_982),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_1033),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1016),
.B(n_928),
.Y(n_1091)
);

OAI22xp33_ASAP7_75t_L g1092 ( 
.A1(n_1029),
.A2(n_947),
.B1(n_969),
.B2(n_849),
.Y(n_1092)
);

NOR2xp33_ASAP7_75t_L g1093 ( 
.A(n_1021),
.B(n_969),
.Y(n_1093)
);

INVxp67_ASAP7_75t_SL g1094 ( 
.A(n_1049),
.Y(n_1094)
);

OR2x2_ASAP7_75t_L g1095 ( 
.A(n_1000),
.B(n_625),
.Y(n_1095)
);

NAND3xp33_ASAP7_75t_L g1096 ( 
.A(n_1060),
.B(n_594),
.C(n_593),
.Y(n_1096)
);

NAND2xp5_ASAP7_75t_SL g1097 ( 
.A(n_1004),
.B(n_976),
.Y(n_1097)
);

CKINVDCx6p67_ASAP7_75t_R g1098 ( 
.A(n_1068),
.Y(n_1098)
);

BUFx2_ASAP7_75t_L g1099 ( 
.A(n_1025),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_1023),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_1017),
.B(n_961),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_1029),
.B(n_976),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_1043),
.Y(n_1103)
);

INVx1_ASAP7_75t_SL g1104 ( 
.A(n_1032),
.Y(n_1104)
);

INVx3_ASAP7_75t_L g1105 ( 
.A(n_1043),
.Y(n_1105)
);

AOI22xp33_ASAP7_75t_L g1106 ( 
.A1(n_1018),
.A2(n_966),
.B1(n_848),
.B2(n_832),
.Y(n_1106)
);

INVx2_ASAP7_75t_L g1107 ( 
.A(n_997),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_SL g1108 ( 
.A(n_1006),
.B(n_976),
.Y(n_1108)
);

INVx2_ASAP7_75t_L g1109 ( 
.A(n_997),
.Y(n_1109)
);

XNOR2xp5_ASAP7_75t_L g1110 ( 
.A(n_1032),
.B(n_872),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_1027),
.Y(n_1111)
);

INVx2_ASAP7_75t_L g1112 ( 
.A(n_1002),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_SL g1113 ( 
.A(n_1006),
.B(n_976),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_1002),
.Y(n_1114)
);

INVx2_ASAP7_75t_SL g1115 ( 
.A(n_1017),
.Y(n_1115)
);

INVxp33_ASAP7_75t_L g1116 ( 
.A(n_1009),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_SL g1117 ( 
.A(n_1006),
.B(n_976),
.Y(n_1117)
);

INVx2_ASAP7_75t_L g1118 ( 
.A(n_1010),
.Y(n_1118)
);

INVxp67_ASAP7_75t_SL g1119 ( 
.A(n_1049),
.Y(n_1119)
);

BUFx6f_ASAP7_75t_L g1120 ( 
.A(n_1066),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_1035),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1010),
.Y(n_1122)
);

INVx2_ASAP7_75t_L g1123 ( 
.A(n_1019),
.Y(n_1123)
);

INVxp67_ASAP7_75t_SL g1124 ( 
.A(n_1049),
.Y(n_1124)
);

AOI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1022),
.A2(n_966),
.B1(n_685),
.B2(n_689),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_1039),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_996),
.B(n_872),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_1042),
.Y(n_1128)
);

INVx2_ASAP7_75t_SL g1129 ( 
.A(n_1003),
.Y(n_1129)
);

BUFx10_ASAP7_75t_L g1130 ( 
.A(n_1065),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_1020),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_1034),
.Y(n_1132)
);

NOR2xp33_ASAP7_75t_L g1133 ( 
.A(n_1008),
.B(n_878),
.Y(n_1133)
);

INVx2_ASAP7_75t_L g1134 ( 
.A(n_1020),
.Y(n_1134)
);

NAND2xp33_ASAP7_75t_SL g1135 ( 
.A(n_1009),
.B(n_659),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_SL g1136 ( 
.A(n_1024),
.B(n_1007),
.Y(n_1136)
);

INVxp33_ASAP7_75t_L g1137 ( 
.A(n_1062),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_1012),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1018),
.B(n_928),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_1065),
.Y(n_1140)
);

INVx1_ASAP7_75t_L g1141 ( 
.A(n_1065),
.Y(n_1141)
);

INVx5_ASAP7_75t_L g1142 ( 
.A(n_1018),
.Y(n_1142)
);

NAND2xp5_ASAP7_75t_SL g1143 ( 
.A(n_1064),
.B(n_978),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1044),
.Y(n_1144)
);

INVx3_ASAP7_75t_L g1145 ( 
.A(n_1064),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_1015),
.B(n_878),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1044),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1018),
.B(n_927),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_1046),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_1046),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_1044),
.Y(n_1151)
);

NAND2xp5_ASAP7_75t_L g1152 ( 
.A(n_1052),
.B(n_927),
.Y(n_1152)
);

INVx2_ASAP7_75t_L g1153 ( 
.A(n_1047),
.Y(n_1153)
);

AOI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1062),
.A2(n_966),
.B1(n_696),
.B2(n_702),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_1061),
.Y(n_1155)
);

NAND2xp5_ASAP7_75t_SL g1156 ( 
.A(n_1069),
.B(n_1055),
.Y(n_1156)
);

INVx4_ASAP7_75t_L g1157 ( 
.A(n_1049),
.Y(n_1157)
);

NAND2xp5_ASAP7_75t_L g1158 ( 
.A(n_1069),
.B(n_928),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1070),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_L g1160 ( 
.A1(n_1070),
.A2(n_966),
.B1(n_737),
.B2(n_770),
.Y(n_1160)
);

INVx2_ASAP7_75t_L g1161 ( 
.A(n_1047),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1048),
.B(n_1053),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_1050),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_1061),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_1050),
.Y(n_1165)
);

INVx2_ASAP7_75t_L g1166 ( 
.A(n_1059),
.Y(n_1166)
);

INVx2_ASAP7_75t_SL g1167 ( 
.A(n_1061),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_SL g1168 ( 
.A(n_1054),
.B(n_978),
.Y(n_1168)
);

NOR2xp33_ASAP7_75t_L g1169 ( 
.A(n_1071),
.B(n_920),
.Y(n_1169)
);

NAND2xp5_ASAP7_75t_SL g1170 ( 
.A(n_1063),
.B(n_978),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_1051),
.Y(n_1171)
);

INVx3_ASAP7_75t_L g1172 ( 
.A(n_1048),
.Y(n_1172)
);

NAND2xp5_ASAP7_75t_L g1173 ( 
.A(n_1048),
.B(n_978),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_1051),
.Y(n_1174)
);

NOR2xp33_ASAP7_75t_SL g1175 ( 
.A(n_1068),
.B(n_659),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1038),
.Y(n_1176)
);

INVx2_ASAP7_75t_L g1177 ( 
.A(n_1038),
.Y(n_1177)
);

NAND2xp5_ASAP7_75t_L g1178 ( 
.A(n_1053),
.B(n_978),
.Y(n_1178)
);

NAND2xp5_ASAP7_75t_L g1179 ( 
.A(n_1053),
.B(n_984),
.Y(n_1179)
);

INVx2_ASAP7_75t_L g1180 ( 
.A(n_1040),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_1040),
.Y(n_1181)
);

INVx2_ASAP7_75t_L g1182 ( 
.A(n_1040),
.Y(n_1182)
);

NAND3xp33_ASAP7_75t_L g1183 ( 
.A(n_1041),
.B(n_596),
.C(n_595),
.Y(n_1183)
);

INVx2_ASAP7_75t_L g1184 ( 
.A(n_1056),
.Y(n_1184)
);

INVx2_ASAP7_75t_SL g1185 ( 
.A(n_1056),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_992),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1057),
.Y(n_1187)
);

INVx2_ASAP7_75t_L g1188 ( 
.A(n_1057),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_992),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_992),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_1057),
.B(n_984),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_L g1192 ( 
.A(n_1067),
.B(n_984),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_992),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_1066),
.B(n_961),
.Y(n_1194)
);

NOR2xp33_ASAP7_75t_L g1195 ( 
.A(n_1041),
.B(n_906),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_1088),
.Y(n_1196)
);

INVx1_ASAP7_75t_L g1197 ( 
.A(n_1073),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1074),
.Y(n_1198)
);

AND2x2_ASAP7_75t_L g1199 ( 
.A(n_1137),
.B(n_913),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1083),
.Y(n_1200)
);

INVx1_ASAP7_75t_L g1201 ( 
.A(n_1085),
.Y(n_1201)
);

AND2x2_ASAP7_75t_L g1202 ( 
.A(n_1116),
.B(n_973),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_SL g1203 ( 
.A(n_1142),
.B(n_713),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_1086),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_1163),
.Y(n_1205)
);

INVx2_ASAP7_75t_SL g1206 ( 
.A(n_1095),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_1163),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1165),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1165),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_1088),
.Y(n_1210)
);

CKINVDCx20_ASAP7_75t_R g1211 ( 
.A(n_1090),
.Y(n_1211)
);

NOR2xp33_ASAP7_75t_L g1212 ( 
.A(n_1075),
.B(n_713),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1116),
.B(n_973),
.Y(n_1213)
);

AND2x2_ASAP7_75t_SL g1214 ( 
.A(n_1146),
.B(n_726),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_1072),
.Y(n_1215)
);

INVxp67_ASAP7_75t_L g1216 ( 
.A(n_1101),
.Y(n_1216)
);

AND2x2_ASAP7_75t_L g1217 ( 
.A(n_1159),
.B(n_643),
.Y(n_1217)
);

XNOR2x2_ASAP7_75t_L g1218 ( 
.A(n_1110),
.B(n_667),
.Y(n_1218)
);

XOR2xp5_ASAP7_75t_L g1219 ( 
.A(n_1090),
.B(n_1087),
.Y(n_1219)
);

AND2x2_ASAP7_75t_L g1220 ( 
.A(n_1159),
.B(n_1115),
.Y(n_1220)
);

NOR2xp33_ASAP7_75t_L g1221 ( 
.A(n_1129),
.B(n_731),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1129),
.B(n_731),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1111),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_1131),
.Y(n_1224)
);

AND2x6_ASAP7_75t_L g1225 ( 
.A(n_1171),
.B(n_1045),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1131),
.Y(n_1226)
);

NOR2xp33_ASAP7_75t_L g1227 ( 
.A(n_1099),
.B(n_735),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1134),
.Y(n_1228)
);

INVx1_ASAP7_75t_L g1229 ( 
.A(n_1134),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_1098),
.Y(n_1230)
);

INVx1_ASAP7_75t_L g1231 ( 
.A(n_1100),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_1072),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1132),
.Y(n_1233)
);

INVxp33_ASAP7_75t_L g1234 ( 
.A(n_1195),
.Y(n_1234)
);

XOR2xp5_ASAP7_75t_L g1235 ( 
.A(n_1183),
.B(n_735),
.Y(n_1235)
);

INVx1_ASAP7_75t_L g1236 ( 
.A(n_1121),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_1130),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1167),
.B(n_915),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1126),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1128),
.Y(n_1240)
);

INVx1_ASAP7_75t_L g1241 ( 
.A(n_1149),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1149),
.Y(n_1242)
);

NOR2xp33_ASAP7_75t_L g1243 ( 
.A(n_1115),
.B(n_1089),
.Y(n_1243)
);

AND2x2_ASAP7_75t_L g1244 ( 
.A(n_1101),
.B(n_643),
.Y(n_1244)
);

NOR2xp33_ASAP7_75t_L g1245 ( 
.A(n_1135),
.B(n_754),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1150),
.Y(n_1246)
);

BUFx6f_ASAP7_75t_L g1247 ( 
.A(n_1130),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1150),
.Y(n_1248)
);

AND2x2_ASAP7_75t_L g1249 ( 
.A(n_1078),
.B(n_807),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1153),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1104),
.B(n_678),
.Y(n_1251)
);

INVx2_ASAP7_75t_SL g1252 ( 
.A(n_1138),
.Y(n_1252)
);

XOR2xp5_ASAP7_75t_L g1253 ( 
.A(n_1096),
.B(n_754),
.Y(n_1253)
);

AND2x2_ASAP7_75t_L g1254 ( 
.A(n_1127),
.B(n_807),
.Y(n_1254)
);

INVx1_ASAP7_75t_L g1255 ( 
.A(n_1153),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1161),
.Y(n_1256)
);

AND2x4_ASAP7_75t_L g1257 ( 
.A(n_1167),
.B(n_916),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1135),
.B(n_784),
.Y(n_1258)
);

NOR2xp67_ASAP7_75t_L g1259 ( 
.A(n_1093),
.B(n_924),
.Y(n_1259)
);

CKINVDCx20_ASAP7_75t_R g1260 ( 
.A(n_1098),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1161),
.Y(n_1261)
);

AND2x2_ASAP7_75t_L g1262 ( 
.A(n_1133),
.B(n_807),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1166),
.Y(n_1263)
);

INVx2_ASAP7_75t_L g1264 ( 
.A(n_1077),
.Y(n_1264)
);

INVx1_ASAP7_75t_L g1265 ( 
.A(n_1166),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1077),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1079),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1079),
.Y(n_1268)
);

BUFx5_ASAP7_75t_L g1269 ( 
.A(n_1174),
.Y(n_1269)
);

INVx1_ASAP7_75t_L g1270 ( 
.A(n_1082),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1082),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1136),
.B(n_1097),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1103),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1103),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1107),
.Y(n_1275)
);

AND2x4_ASAP7_75t_L g1276 ( 
.A(n_1140),
.B(n_918),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1107),
.Y(n_1277)
);

XOR2xp5_ASAP7_75t_L g1278 ( 
.A(n_1125),
.B(n_784),
.Y(n_1278)
);

INVx2_ASAP7_75t_L g1279 ( 
.A(n_1109),
.Y(n_1279)
);

NAND2xp33_ASAP7_75t_SL g1280 ( 
.A(n_1141),
.B(n_790),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_L g1281 ( 
.A(n_1136),
.B(n_1057),
.Y(n_1281)
);

NOR2xp33_ASAP7_75t_SL g1282 ( 
.A(n_1142),
.B(n_790),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1109),
.Y(n_1283)
);

NOR2xp33_ASAP7_75t_L g1284 ( 
.A(n_1102),
.B(n_797),
.Y(n_1284)
);

NOR2xp67_ASAP7_75t_L g1285 ( 
.A(n_1144),
.B(n_681),
.Y(n_1285)
);

XOR2x2_ASAP7_75t_L g1286 ( 
.A(n_1169),
.B(n_701),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_1112),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1112),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1114),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1114),
.Y(n_1290)
);

NAND2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1142),
.B(n_1057),
.Y(n_1291)
);

NOR2xp33_ASAP7_75t_L g1292 ( 
.A(n_1102),
.B(n_797),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1118),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1118),
.Y(n_1294)
);

XNOR2xp5_ASAP7_75t_L g1295 ( 
.A(n_1092),
.B(n_808),
.Y(n_1295)
);

NAND2x1p5_ASAP7_75t_L g1296 ( 
.A(n_1142),
.B(n_1058),
.Y(n_1296)
);

INVx1_ASAP7_75t_L g1297 ( 
.A(n_1122),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1122),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1123),
.Y(n_1299)
);

AND2x2_ASAP7_75t_L g1300 ( 
.A(n_1147),
.B(n_721),
.Y(n_1300)
);

NOR2xp67_ASAP7_75t_L g1301 ( 
.A(n_1151),
.B(n_782),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1155),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1164),
.B(n_808),
.Y(n_1303)
);

INVx1_ASAP7_75t_L g1304 ( 
.A(n_1105),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1175),
.B(n_1058),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1105),
.Y(n_1306)
);

NOR2xp33_ASAP7_75t_L g1307 ( 
.A(n_1108),
.B(n_806),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1184),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1184),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_1145),
.Y(n_1310)
);

INVxp67_ASAP7_75t_SL g1311 ( 
.A(n_1094),
.Y(n_1311)
);

NAND2x1p5_ASAP7_75t_L g1312 ( 
.A(n_1194),
.B(n_1058),
.Y(n_1312)
);

XNOR2xp5_ASAP7_75t_L g1313 ( 
.A(n_1154),
.B(n_794),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1108),
.B(n_634),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1113),
.B(n_1058),
.Y(n_1315)
);

NOR2xp33_ASAP7_75t_L g1316 ( 
.A(n_1113),
.B(n_1067),
.Y(n_1316)
);

INVx2_ASAP7_75t_L g1317 ( 
.A(n_1145),
.Y(n_1317)
);

NOR2xp33_ASAP7_75t_L g1318 ( 
.A(n_1117),
.B(n_1067),
.Y(n_1318)
);

NAND2xp33_ASAP7_75t_R g1319 ( 
.A(n_1139),
.B(n_812),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1177),
.Y(n_1320)
);

CKINVDCx20_ASAP7_75t_R g1321 ( 
.A(n_1117),
.Y(n_1321)
);

CKINVDCx20_ASAP7_75t_R g1322 ( 
.A(n_1170),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1177),
.Y(n_1323)
);

INVx2_ASAP7_75t_SL g1324 ( 
.A(n_1194),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_L g1325 ( 
.A(n_1091),
.B(n_1067),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_1180),
.Y(n_1326)
);

XOR2xp5_ASAP7_75t_L g1327 ( 
.A(n_1160),
.B(n_502),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1170),
.B(n_1067),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1180),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1182),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1182),
.Y(n_1331)
);

INVx1_ASAP7_75t_L g1332 ( 
.A(n_1176),
.Y(n_1332)
);

NAND2xp33_ASAP7_75t_SL g1333 ( 
.A(n_1120),
.B(n_730),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_1181),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1172),
.Y(n_1335)
);

XNOR2xp5_ASAP7_75t_L g1336 ( 
.A(n_1076),
.B(n_608),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1172),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1148),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1172),
.Y(n_1339)
);

XNOR2xp5_ASAP7_75t_L g1340 ( 
.A(n_1080),
.B(n_612),
.Y(n_1340)
);

CKINVDCx5p33_ASAP7_75t_R g1341 ( 
.A(n_1120),
.Y(n_1341)
);

XOR2x2_ASAP7_75t_L g1342 ( 
.A(n_1080),
.B(n_1),
.Y(n_1342)
);

INVx2_ASAP7_75t_L g1343 ( 
.A(n_1185),
.Y(n_1343)
);

AND2x4_ASAP7_75t_L g1344 ( 
.A(n_1120),
.B(n_921),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1185),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1106),
.B(n_922),
.Y(n_1346)
);

AND2x2_ASAP7_75t_SL g1347 ( 
.A(n_1084),
.B(n_791),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1152),
.Y(n_1348)
);

CKINVDCx20_ASAP7_75t_R g1349 ( 
.A(n_1156),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1156),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_1120),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1187),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1187),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1158),
.Y(n_1354)
);

NAND2xp5_ASAP7_75t_L g1355 ( 
.A(n_1188),
.B(n_1119),
.Y(n_1355)
);

INVx3_ASAP7_75t_L g1356 ( 
.A(n_1188),
.Y(n_1356)
);

INVx2_ASAP7_75t_SL g1357 ( 
.A(n_1162),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_1186),
.Y(n_1358)
);

NAND2xp5_ASAP7_75t_L g1359 ( 
.A(n_1124),
.B(n_848),
.Y(n_1359)
);

INVx4_ASAP7_75t_L g1360 ( 
.A(n_1081),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1189),
.Y(n_1361)
);

NOR2xp33_ASAP7_75t_L g1362 ( 
.A(n_1190),
.B(n_597),
.Y(n_1362)
);

XNOR2xp5_ASAP7_75t_L g1363 ( 
.A(n_1168),
.B(n_612),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1193),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1084),
.B(n_922),
.Y(n_1365)
);

INVx3_ASAP7_75t_R g1366 ( 
.A(n_1143),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1173),
.Y(n_1367)
);

AND2x2_ASAP7_75t_L g1368 ( 
.A(n_1168),
.B(n_923),
.Y(n_1368)
);

CKINVDCx20_ASAP7_75t_R g1369 ( 
.A(n_1178),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1179),
.Y(n_1370)
);

NAND2xp5_ASAP7_75t_L g1371 ( 
.A(n_1081),
.B(n_984),
.Y(n_1371)
);

XNOR2x2_ASAP7_75t_L g1372 ( 
.A(n_1191),
.B(n_670),
.Y(n_1372)
);

AND2x2_ASAP7_75t_L g1373 ( 
.A(n_1199),
.B(n_923),
.Y(n_1373)
);

NAND2xp5_ASAP7_75t_SL g1374 ( 
.A(n_1214),
.B(n_1081),
.Y(n_1374)
);

INVx2_ASAP7_75t_L g1375 ( 
.A(n_1215),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1232),
.Y(n_1376)
);

NOR3xp33_ASAP7_75t_L g1377 ( 
.A(n_1212),
.B(n_739),
.C(n_730),
.Y(n_1377)
);

NOR2xp33_ASAP7_75t_L g1378 ( 
.A(n_1212),
.B(n_1157),
.Y(n_1378)
);

OAI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1203),
.A2(n_739),
.B1(n_742),
.B2(n_675),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1234),
.B(n_1243),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1205),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1216),
.B(n_1192),
.Y(n_1382)
);

NOR2xp67_ASAP7_75t_L g1383 ( 
.A(n_1206),
.B(n_504),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1264),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1272),
.B(n_1338),
.Y(n_1385)
);

INVx2_ASAP7_75t_L g1386 ( 
.A(n_1277),
.Y(n_1386)
);

NAND2xp5_ASAP7_75t_SL g1387 ( 
.A(n_1203),
.B(n_1001),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1272),
.B(n_829),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_SL g1389 ( 
.A(n_1282),
.B(n_994),
.Y(n_1389)
);

INVx2_ASAP7_75t_SL g1390 ( 
.A(n_1251),
.Y(n_1390)
);

INVx2_ASAP7_75t_SL g1391 ( 
.A(n_1369),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1360),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1207),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1208),
.Y(n_1394)
);

NAND2xp5_ASAP7_75t_L g1395 ( 
.A(n_1220),
.B(n_980),
.Y(n_1395)
);

NOR2xp33_ASAP7_75t_L g1396 ( 
.A(n_1227),
.B(n_602),
.Y(n_1396)
);

NAND3xp33_ASAP7_75t_L g1397 ( 
.A(n_1295),
.B(n_613),
.C(n_605),
.Y(n_1397)
);

OAI22xp5_ASAP7_75t_L g1398 ( 
.A1(n_1341),
.A2(n_742),
.B1(n_798),
.B2(n_791),
.Y(n_1398)
);

NOR2xp33_ASAP7_75t_L g1399 ( 
.A(n_1227),
.B(n_616),
.Y(n_1399)
);

INVxp67_ASAP7_75t_SL g1400 ( 
.A(n_1311),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1307),
.B(n_980),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1351),
.A2(n_804),
.B1(n_813),
.B2(n_798),
.Y(n_1402)
);

INVxp67_ASAP7_75t_L g1403 ( 
.A(n_1221),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1279),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1284),
.A2(n_866),
.B1(n_867),
.B2(n_864),
.Y(n_1405)
);

NOR2xp67_ASAP7_75t_L g1406 ( 
.A(n_1259),
.B(n_1252),
.Y(n_1406)
);

NAND2xp5_ASAP7_75t_L g1407 ( 
.A(n_1307),
.B(n_985),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1314),
.B(n_1202),
.Y(n_1408)
);

INVx1_ASAP7_75t_L g1409 ( 
.A(n_1209),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1213),
.B(n_958),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1311),
.B(n_958),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1224),
.Y(n_1412)
);

INVxp67_ASAP7_75t_L g1413 ( 
.A(n_1221),
.Y(n_1413)
);

NAND2xp5_ASAP7_75t_L g1414 ( 
.A(n_1354),
.B(n_994),
.Y(n_1414)
);

INVx2_ASAP7_75t_SL g1415 ( 
.A(n_1217),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1300),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1226),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1228),
.Y(n_1418)
);

AND2x4_ASAP7_75t_L g1419 ( 
.A(n_1237),
.B(n_671),
.Y(n_1419)
);

INVx2_ASAP7_75t_SL g1420 ( 
.A(n_1244),
.Y(n_1420)
);

NAND2xp33_ASAP7_75t_SL g1421 ( 
.A(n_1322),
.B(n_675),
.Y(n_1421)
);

INVx2_ASAP7_75t_L g1422 ( 
.A(n_1289),
.Y(n_1422)
);

INVxp67_ASAP7_75t_L g1423 ( 
.A(n_1222),
.Y(n_1423)
);

NAND2xp5_ASAP7_75t_L g1424 ( 
.A(n_1197),
.B(n_1001),
.Y(n_1424)
);

NAND2xp5_ASAP7_75t_L g1425 ( 
.A(n_1198),
.B(n_1001),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1290),
.Y(n_1426)
);

AND2x2_ASAP7_75t_L g1427 ( 
.A(n_1284),
.B(n_618),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1229),
.Y(n_1428)
);

AOI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1292),
.A2(n_870),
.B1(n_873),
.B2(n_868),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1241),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1200),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1242),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1338),
.B(n_875),
.Y(n_1433)
);

AND2x4_ASAP7_75t_L g1434 ( 
.A(n_1237),
.B(n_672),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1292),
.B(n_624),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1222),
.B(n_1245),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1201),
.B(n_1005),
.Y(n_1437)
);

BUFx4f_ASAP7_75t_L g1438 ( 
.A(n_1247),
.Y(n_1438)
);

NOR2xp33_ASAP7_75t_L g1439 ( 
.A(n_1245),
.B(n_627),
.Y(n_1439)
);

BUFx8_ASAP7_75t_L g1440 ( 
.A(n_1249),
.Y(n_1440)
);

INVx1_ASAP7_75t_L g1441 ( 
.A(n_1204),
.Y(n_1441)
);

BUFx6f_ASAP7_75t_L g1442 ( 
.A(n_1247),
.Y(n_1442)
);

NOR2xp33_ASAP7_75t_L g1443 ( 
.A(n_1258),
.B(n_628),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1246),
.Y(n_1444)
);

BUFx3_ASAP7_75t_L g1445 ( 
.A(n_1196),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1258),
.B(n_821),
.Y(n_1446)
);

AO221x1_ASAP7_75t_L g1447 ( 
.A1(n_1247),
.A2(n_687),
.B1(n_688),
.B2(n_683),
.C(n_680),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1248),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1262),
.B(n_629),
.Y(n_1449)
);

NAND2xp5_ASAP7_75t_SL g1450 ( 
.A(n_1324),
.B(n_1014),
.Y(n_1450)
);

NAND2xp5_ASAP7_75t_SL g1451 ( 
.A(n_1238),
.B(n_1257),
.Y(n_1451)
);

AND2x4_ASAP7_75t_L g1452 ( 
.A(n_1238),
.B(n_690),
.Y(n_1452)
);

AOI22xp5_ASAP7_75t_L g1453 ( 
.A1(n_1321),
.A2(n_1026),
.B1(n_1028),
.B2(n_1014),
.Y(n_1453)
);

INVx2_ASAP7_75t_SL g1454 ( 
.A(n_1210),
.Y(n_1454)
);

NOR2xp33_ASAP7_75t_L g1455 ( 
.A(n_1278),
.B(n_630),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1223),
.B(n_1026),
.Y(n_1456)
);

INVx3_ASAP7_75t_L g1457 ( 
.A(n_1312),
.Y(n_1457)
);

OAI22xp5_ASAP7_75t_L g1458 ( 
.A1(n_1347),
.A2(n_813),
.B1(n_814),
.B2(n_804),
.Y(n_1458)
);

AOI22xp5_ASAP7_75t_L g1459 ( 
.A1(n_1349),
.A2(n_1028),
.B1(n_1030),
.B2(n_1026),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1250),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1348),
.B(n_1350),
.Y(n_1461)
);

NOR2xp33_ASAP7_75t_L g1462 ( 
.A(n_1303),
.B(n_631),
.Y(n_1462)
);

O2A1O1Ixp5_ASAP7_75t_L g1463 ( 
.A1(n_1333),
.A2(n_814),
.B(n_876),
.C(n_874),
.Y(n_1463)
);

INVx3_ASAP7_75t_L g1464 ( 
.A(n_1312),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1303),
.B(n_1254),
.Y(n_1465)
);

AOI22xp5_ASAP7_75t_L g1466 ( 
.A1(n_1280),
.A2(n_1319),
.B1(n_1285),
.B2(n_1301),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1231),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1255),
.Y(n_1468)
);

INVx3_ASAP7_75t_L g1469 ( 
.A(n_1344),
.Y(n_1469)
);

NOR2xp33_ASAP7_75t_SL g1470 ( 
.A(n_1230),
.B(n_821),
.Y(n_1470)
);

A2O1A1Ixp33_ASAP7_75t_L g1471 ( 
.A1(n_1302),
.A2(n_695),
.B(n_700),
.C(n_694),
.Y(n_1471)
);

NOR2xp67_ASAP7_75t_L g1472 ( 
.A(n_1233),
.B(n_505),
.Y(n_1472)
);

NAND2xp5_ASAP7_75t_L g1473 ( 
.A(n_1236),
.B(n_1028),
.Y(n_1473)
);

AND2x2_ASAP7_75t_L g1474 ( 
.A(n_1336),
.B(n_632),
.Y(n_1474)
);

NAND2xp5_ASAP7_75t_L g1475 ( 
.A(n_1239),
.B(n_1240),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1340),
.B(n_635),
.Y(n_1476)
);

AOI22xp5_ASAP7_75t_L g1477 ( 
.A1(n_1305),
.A2(n_1030),
.B1(n_879),
.B2(n_877),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_SL g1478 ( 
.A(n_1363),
.B(n_950),
.Y(n_1478)
);

NAND2xp5_ASAP7_75t_SL g1479 ( 
.A(n_1313),
.B(n_950),
.Y(n_1479)
);

NAND2xp5_ASAP7_75t_L g1480 ( 
.A(n_1357),
.B(n_642),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1256),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_SL g1482 ( 
.A(n_1362),
.B(n_1276),
.Y(n_1482)
);

NAND2xp5_ASAP7_75t_L g1483 ( 
.A(n_1367),
.B(n_645),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1276),
.Y(n_1484)
);

INVx1_ASAP7_75t_SL g1485 ( 
.A(n_1211),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1218),
.Y(n_1486)
);

NAND2xp5_ASAP7_75t_L g1487 ( 
.A(n_1370),
.B(n_833),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1253),
.B(n_647),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1286),
.B(n_649),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1266),
.Y(n_1490)
);

BUFx6f_ASAP7_75t_SL g1491 ( 
.A(n_1344),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_SL g1492 ( 
.A(n_1263),
.B(n_1265),
.Y(n_1492)
);

INVx2_ASAP7_75t_L g1493 ( 
.A(n_1261),
.Y(n_1493)
);

OAI22xp5_ASAP7_75t_L g1494 ( 
.A1(n_1327),
.A2(n_720),
.B1(n_723),
.B2(n_717),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1365),
.B(n_834),
.Y(n_1495)
);

INVx2_ASAP7_75t_SL g1496 ( 
.A(n_1342),
.Y(n_1496)
);

NAND2x1p5_ASAP7_75t_L g1497 ( 
.A(n_1356),
.B(n_1335),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1267),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1368),
.B(n_834),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1268),
.Y(n_1500)
);

AOI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1219),
.A2(n_1346),
.B1(n_1235),
.B2(n_1345),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1270),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1343),
.B(n_837),
.Y(n_1503)
);

BUFx8_ASAP7_75t_L g1504 ( 
.A(n_1332),
.Y(n_1504)
);

NAND2xp33_ASAP7_75t_L g1505 ( 
.A(n_1269),
.B(n_650),
.Y(n_1505)
);

NAND2xp5_ASAP7_75t_SL g1506 ( 
.A(n_1269),
.B(n_1334),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1271),
.B(n_837),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1273),
.B(n_839),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1274),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1275),
.Y(n_1510)
);

AND2x6_ASAP7_75t_L g1511 ( 
.A(n_1315),
.B(n_732),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1283),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1287),
.Y(n_1513)
);

INVx2_ASAP7_75t_SL g1514 ( 
.A(n_1260),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1328),
.A2(n_1316),
.B1(n_1318),
.B2(n_1315),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1288),
.Y(n_1516)
);

INVx3_ASAP7_75t_L g1517 ( 
.A(n_1291),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1293),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1294),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1297),
.B(n_653),
.Y(n_1520)
);

NAND2xp5_ASAP7_75t_L g1521 ( 
.A(n_1298),
.B(n_654),
.Y(n_1521)
);

INVx2_ASAP7_75t_L g1522 ( 
.A(n_1299),
.Y(n_1522)
);

NAND2xp33_ASAP7_75t_L g1523 ( 
.A(n_1358),
.B(n_655),
.Y(n_1523)
);

INVx2_ASAP7_75t_SL g1524 ( 
.A(n_1372),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1325),
.B(n_656),
.Y(n_1525)
);

NOR2xp33_ASAP7_75t_L g1526 ( 
.A(n_1361),
.B(n_657),
.Y(n_1526)
);

NAND2xp5_ASAP7_75t_L g1527 ( 
.A(n_1355),
.B(n_658),
.Y(n_1527)
);

BUFx5_ASAP7_75t_L g1528 ( 
.A(n_1225),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_L g1529 ( 
.A(n_1364),
.B(n_662),
.Y(n_1529)
);

NAND2xp33_ASAP7_75t_L g1530 ( 
.A(n_1291),
.B(n_1296),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1308),
.Y(n_1531)
);

NAND2xp5_ASAP7_75t_L g1532 ( 
.A(n_1355),
.B(n_663),
.Y(n_1532)
);

NAND2xp5_ASAP7_75t_L g1533 ( 
.A(n_1316),
.B(n_664),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1318),
.B(n_665),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_L g1535 ( 
.A(n_1366),
.B(n_668),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_1309),
.Y(n_1536)
);

INVx8_ASAP7_75t_L g1537 ( 
.A(n_1225),
.Y(n_1537)
);

NOR2xp33_ASAP7_75t_L g1538 ( 
.A(n_1337),
.B(n_674),
.Y(n_1538)
);

NOR2xp33_ASAP7_75t_L g1539 ( 
.A(n_1339),
.B(n_676),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1320),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1323),
.A2(n_844),
.B1(n_847),
.B2(n_839),
.Y(n_1541)
);

CKINVDCx20_ASAP7_75t_R g1542 ( 
.A(n_1352),
.Y(n_1542)
);

NOR2xp33_ASAP7_75t_L g1543 ( 
.A(n_1353),
.B(n_679),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1326),
.A2(n_847),
.B1(n_850),
.B2(n_844),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_SL g1545 ( 
.A(n_1310),
.B(n_682),
.Y(n_1545)
);

NOR2xp33_ASAP7_75t_L g1546 ( 
.A(n_1356),
.B(n_684),
.Y(n_1546)
);

BUFx2_ASAP7_75t_L g1547 ( 
.A(n_1329),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_SL g1548 ( 
.A(n_1317),
.B(n_686),
.Y(n_1548)
);

INVx2_ASAP7_75t_L g1549 ( 
.A(n_1330),
.Y(n_1549)
);

NAND2xp5_ASAP7_75t_L g1550 ( 
.A(n_1281),
.B(n_850),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1281),
.B(n_851),
.Y(n_1551)
);

NAND2xp5_ASAP7_75t_SL g1552 ( 
.A(n_1380),
.B(n_1304),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1436),
.B(n_1359),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1408),
.B(n_1331),
.Y(n_1554)
);

OAI22xp5_ASAP7_75t_L g1555 ( 
.A1(n_1400),
.A2(n_1296),
.B1(n_1371),
.B2(n_1306),
.Y(n_1555)
);

AND2x2_ASAP7_75t_L g1556 ( 
.A(n_1427),
.B(n_698),
.Y(n_1556)
);

INVx2_ASAP7_75t_SL g1557 ( 
.A(n_1438),
.Y(n_1557)
);

NAND2xp5_ASAP7_75t_L g1558 ( 
.A(n_1465),
.B(n_1225),
.Y(n_1558)
);

AOI21xp5_ASAP7_75t_L g1559 ( 
.A1(n_1495),
.A2(n_987),
.B(n_984),
.Y(n_1559)
);

AOI21xp5_ASAP7_75t_L g1560 ( 
.A1(n_1482),
.A2(n_987),
.B(n_956),
.Y(n_1560)
);

INVx2_ASAP7_75t_L g1561 ( 
.A(n_1430),
.Y(n_1561)
);

AOI21xp5_ASAP7_75t_L g1562 ( 
.A1(n_1505),
.A2(n_987),
.B(n_956),
.Y(n_1562)
);

AO21x1_ASAP7_75t_L g1563 ( 
.A1(n_1378),
.A2(n_741),
.B(n_733),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1530),
.A2(n_987),
.B(n_956),
.Y(n_1564)
);

INVx1_ASAP7_75t_SL g1565 ( 
.A(n_1390),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1515),
.A2(n_703),
.B1(n_704),
.B2(n_699),
.Y(n_1566)
);

INVx8_ASAP7_75t_L g1567 ( 
.A(n_1491),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_SL g1568 ( 
.A(n_1501),
.B(n_705),
.Y(n_1568)
);

AO21x1_ASAP7_75t_L g1569 ( 
.A1(n_1435),
.A2(n_748),
.B(n_746),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1467),
.Y(n_1570)
);

OAI21xp33_ASAP7_75t_L g1571 ( 
.A1(n_1439),
.A2(n_1443),
.B(n_1462),
.Y(n_1571)
);

BUFx2_ASAP7_75t_L g1572 ( 
.A(n_1542),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1385),
.B(n_1225),
.Y(n_1573)
);

AOI21xp5_ASAP7_75t_L g1574 ( 
.A1(n_1388),
.A2(n_956),
.B(n_852),
.Y(n_1574)
);

BUFx2_ASAP7_75t_L g1575 ( 
.A(n_1391),
.Y(n_1575)
);

O2A1O1Ixp33_ASAP7_75t_L g1576 ( 
.A1(n_1396),
.A2(n_753),
.B(n_757),
.C(n_751),
.Y(n_1576)
);

O2A1O1Ixp33_ASAP7_75t_L g1577 ( 
.A1(n_1399),
.A2(n_760),
.B(n_764),
.C(n_759),
.Y(n_1577)
);

AOI21xp5_ASAP7_75t_L g1578 ( 
.A1(n_1499),
.A2(n_956),
.B(n_852),
.Y(n_1578)
);

INVx3_ASAP7_75t_L g1579 ( 
.A(n_1392),
.Y(n_1579)
);

A2O1A1Ixp33_ASAP7_75t_L g1580 ( 
.A1(n_1449),
.A2(n_1377),
.B(n_1413),
.C(n_1403),
.Y(n_1580)
);

AOI21xp5_ASAP7_75t_L g1581 ( 
.A1(n_1374),
.A2(n_853),
.B(n_851),
.Y(n_1581)
);

AOI22xp33_ASAP7_75t_L g1582 ( 
.A1(n_1397),
.A2(n_818),
.B1(n_822),
.B2(n_816),
.Y(n_1582)
);

AOI22xp33_ASAP7_75t_L g1583 ( 
.A1(n_1486),
.A2(n_1474),
.B1(n_1476),
.B2(n_1524),
.Y(n_1583)
);

O2A1O1Ixp33_ASAP7_75t_L g1584 ( 
.A1(n_1423),
.A2(n_773),
.B(n_774),
.C(n_769),
.Y(n_1584)
);

BUFx4f_ASAP7_75t_L g1585 ( 
.A(n_1442),
.Y(n_1585)
);

NAND2xp5_ASAP7_75t_L g1586 ( 
.A(n_1385),
.B(n_780),
.Y(n_1586)
);

OAI21xp5_ASAP7_75t_L g1587 ( 
.A1(n_1533),
.A2(n_854),
.B(n_853),
.Y(n_1587)
);

INVxp67_ASAP7_75t_L g1588 ( 
.A(n_1416),
.Y(n_1588)
);

OAI21xp5_ASAP7_75t_L g1589 ( 
.A1(n_1534),
.A2(n_858),
.B(n_855),
.Y(n_1589)
);

INVx2_ASAP7_75t_L g1590 ( 
.A(n_1432),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1461),
.A2(n_859),
.B(n_858),
.Y(n_1591)
);

NOR2xp33_ASAP7_75t_L g1592 ( 
.A(n_1488),
.B(n_706),
.Y(n_1592)
);

AO21x2_ASAP7_75t_L g1593 ( 
.A1(n_1506),
.A2(n_859),
.B(n_799),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1373),
.B(n_786),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1527),
.B(n_810),
.Y(n_1595)
);

OAI321xp33_ASAP7_75t_L g1596 ( 
.A1(n_1379),
.A2(n_714),
.A3(n_710),
.B1(n_715),
.B2(n_711),
.C(n_707),
.Y(n_1596)
);

INVx2_ASAP7_75t_L g1597 ( 
.A(n_1444),
.Y(n_1597)
);

INVx1_ASAP7_75t_L g1598 ( 
.A(n_1431),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1532),
.B(n_716),
.Y(n_1599)
);

NAND2xp33_ASAP7_75t_L g1600 ( 
.A(n_1442),
.B(n_718),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1448),
.Y(n_1601)
);

AOI21xp5_ASAP7_75t_L g1602 ( 
.A1(n_1550),
.A2(n_946),
.B(n_945),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1451),
.B(n_722),
.Y(n_1603)
);

INVx3_ASAP7_75t_L g1604 ( 
.A(n_1392),
.Y(n_1604)
);

AOI21xp5_ASAP7_75t_L g1605 ( 
.A1(n_1551),
.A2(n_946),
.B(n_945),
.Y(n_1605)
);

NAND2xp33_ASAP7_75t_L g1606 ( 
.A(n_1511),
.B(n_724),
.Y(n_1606)
);

AND2x2_ASAP7_75t_L g1607 ( 
.A(n_1446),
.B(n_725),
.Y(n_1607)
);

OR2x2_ASAP7_75t_SL g1608 ( 
.A(n_1483),
.B(n_1484),
.Y(n_1608)
);

AOI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1415),
.A2(n_728),
.B1(n_734),
.B2(n_727),
.Y(n_1609)
);

AOI21xp5_ASAP7_75t_L g1610 ( 
.A1(n_1551),
.A2(n_962),
.B(n_946),
.Y(n_1610)
);

AO21x1_ASAP7_75t_L g1611 ( 
.A1(n_1387),
.A2(n_4),
.B(n_2),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1475),
.B(n_736),
.Y(n_1612)
);

NOR2xp33_ASAP7_75t_L g1613 ( 
.A(n_1455),
.B(n_743),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1441),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_L g1615 ( 
.A(n_1525),
.B(n_744),
.Y(n_1615)
);

NOR2xp67_ASAP7_75t_L g1616 ( 
.A(n_1420),
.B(n_506),
.Y(n_1616)
);

NOR3xp33_ASAP7_75t_L g1617 ( 
.A(n_1489),
.B(n_749),
.C(n_747),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1460),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_L g1619 ( 
.A(n_1395),
.B(n_752),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_L g1620 ( 
.A1(n_1389),
.A2(n_962),
.B(n_511),
.Y(n_1620)
);

NOR2xp33_ASAP7_75t_L g1621 ( 
.A(n_1496),
.B(n_755),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1490),
.Y(n_1622)
);

AOI21xp5_ASAP7_75t_L g1623 ( 
.A1(n_1487),
.A2(n_512),
.B(n_509),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1401),
.B(n_756),
.Y(n_1624)
);

OAI22xp5_ASAP7_75t_L g1625 ( 
.A1(n_1469),
.A2(n_761),
.B1(n_763),
.B2(n_758),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1407),
.A2(n_515),
.B(n_513),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1411),
.A2(n_518),
.B(n_517),
.Y(n_1627)
);

INVx2_ASAP7_75t_SL g1628 ( 
.A(n_1445),
.Y(n_1628)
);

NOR2xp33_ASAP7_75t_R g1629 ( 
.A(n_1454),
.B(n_520),
.Y(n_1629)
);

INVx3_ASAP7_75t_SL g1630 ( 
.A(n_1485),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1466),
.A2(n_766),
.B(n_767),
.C(n_765),
.Y(n_1631)
);

BUFx6f_ASAP7_75t_L g1632 ( 
.A(n_1419),
.Y(n_1632)
);

NAND2x1p5_ASAP7_75t_L g1633 ( 
.A(n_1469),
.B(n_527),
.Y(n_1633)
);

NAND2xp5_ASAP7_75t_SL g1634 ( 
.A(n_1406),
.B(n_768),
.Y(n_1634)
);

INVx3_ASAP7_75t_L g1635 ( 
.A(n_1517),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_SL g1636 ( 
.A(n_1470),
.B(n_776),
.Y(n_1636)
);

AO21x1_ASAP7_75t_L g1637 ( 
.A1(n_1458),
.A2(n_5),
.B(n_4),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_SL g1638 ( 
.A(n_1470),
.B(n_777),
.Y(n_1638)
);

AND2x2_ASAP7_75t_L g1639 ( 
.A(n_1452),
.B(n_778),
.Y(n_1639)
);

INVx1_ASAP7_75t_SL g1640 ( 
.A(n_1485),
.Y(n_1640)
);

A2O1A1Ixp33_ASAP7_75t_L g1641 ( 
.A1(n_1535),
.A2(n_1529),
.B(n_1526),
.C(n_1543),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1468),
.Y(n_1642)
);

INVx2_ASAP7_75t_L g1643 ( 
.A(n_1481),
.Y(n_1643)
);

INVx8_ASAP7_75t_L g1644 ( 
.A(n_1491),
.Y(n_1644)
);

INVx2_ASAP7_75t_L g1645 ( 
.A(n_1493),
.Y(n_1645)
);

AOI21xp5_ASAP7_75t_L g1646 ( 
.A1(n_1410),
.A2(n_525),
.B(n_523),
.Y(n_1646)
);

AOI21xp5_ASAP7_75t_L g1647 ( 
.A1(n_1433),
.A2(n_528),
.B(n_526),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1433),
.B(n_783),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1498),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1419),
.Y(n_1650)
);

AND2x4_ASAP7_75t_L g1651 ( 
.A(n_1547),
.B(n_530),
.Y(n_1651)
);

CKINVDCx10_ASAP7_75t_R g1652 ( 
.A(n_1440),
.Y(n_1652)
);

NAND3xp33_ASAP7_75t_L g1653 ( 
.A(n_1494),
.B(n_788),
.C(n_785),
.Y(n_1653)
);

CKINVDCx5p33_ASAP7_75t_R g1654 ( 
.A(n_1440),
.Y(n_1654)
);

INVx2_ASAP7_75t_L g1655 ( 
.A(n_1509),
.Y(n_1655)
);

AOI21xp5_ASAP7_75t_L g1656 ( 
.A1(n_1414),
.A2(n_532),
.B(n_531),
.Y(n_1656)
);

BUFx2_ASAP7_75t_L g1657 ( 
.A(n_1434),
.Y(n_1657)
);

OAI21xp5_ASAP7_75t_L g1658 ( 
.A1(n_1382),
.A2(n_795),
.B(n_792),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1452),
.B(n_800),
.Y(n_1659)
);

BUFx6f_ASAP7_75t_L g1660 ( 
.A(n_1434),
.Y(n_1660)
);

OAI21xp5_ASAP7_75t_L g1661 ( 
.A1(n_1492),
.A2(n_802),
.B(n_801),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1546),
.B(n_803),
.Y(n_1662)
);

NOR2xp33_ASAP7_75t_R g1663 ( 
.A(n_1421),
.B(n_1514),
.Y(n_1663)
);

NAND2xp5_ASAP7_75t_L g1664 ( 
.A(n_1538),
.B(n_805),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_L g1665 ( 
.A(n_1539),
.B(n_809),
.Y(n_1665)
);

OR2x6_ASAP7_75t_L g1666 ( 
.A(n_1537),
.B(n_533),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1507),
.A2(n_535),
.B(n_534),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1500),
.Y(n_1668)
);

CKINVDCx20_ASAP7_75t_R g1669 ( 
.A(n_1479),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1520),
.B(n_811),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1521),
.B(n_815),
.Y(n_1671)
);

AOI21xp5_ASAP7_75t_L g1672 ( 
.A1(n_1507),
.A2(n_537),
.B(n_536),
.Y(n_1672)
);

OAI21xp5_ASAP7_75t_L g1673 ( 
.A1(n_1503),
.A2(n_820),
.B(n_819),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1502),
.Y(n_1674)
);

AOI21xp5_ASAP7_75t_L g1675 ( 
.A1(n_1508),
.A2(n_540),
.B(n_538),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1480),
.B(n_0),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1478),
.B(n_0),
.Y(n_1677)
);

AOI21xp5_ASAP7_75t_L g1678 ( 
.A1(n_1508),
.A2(n_542),
.B(n_541),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1523),
.A2(n_544),
.B(n_543),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1517),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_SL g1681 ( 
.A(n_1472),
.B(n_1383),
.Y(n_1681)
);

NAND3xp33_ASAP7_75t_L g1682 ( 
.A(n_1494),
.B(n_5),
.C(n_6),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1522),
.Y(n_1683)
);

OAI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1503),
.A2(n_547),
.B(n_546),
.Y(n_1684)
);

OAI22xp5_ASAP7_75t_L g1685 ( 
.A1(n_1459),
.A2(n_10),
.B1(n_7),
.B2(n_8),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1545),
.B(n_8),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_SL g1687 ( 
.A(n_1428),
.B(n_10),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1510),
.Y(n_1688)
);

AOI21xp33_ASAP7_75t_L g1689 ( 
.A1(n_1548),
.A2(n_11),
.B(n_12),
.Y(n_1689)
);

OAI22xp5_ASAP7_75t_L g1690 ( 
.A1(n_1453),
.A2(n_13),
.B1(n_11),
.B2(n_12),
.Y(n_1690)
);

NOR2x1_ASAP7_75t_L g1691 ( 
.A(n_1457),
.B(n_549),
.Y(n_1691)
);

AOI22xp5_ASAP7_75t_L g1692 ( 
.A1(n_1447),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_SL g1693 ( 
.A(n_1504),
.B(n_15),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1471),
.B(n_16),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1531),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1381),
.B(n_17),
.Y(n_1696)
);

INVx2_ASAP7_75t_SL g1697 ( 
.A(n_1504),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1512),
.Y(n_1698)
);

A2O1A1Ixp33_ASAP7_75t_L g1699 ( 
.A1(n_1463),
.A2(n_19),
.B(n_17),
.C(n_18),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1513),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1398),
.B(n_18),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1424),
.A2(n_1437),
.B(n_1425),
.Y(n_1702)
);

INVx3_ASAP7_75t_L g1703 ( 
.A(n_1464),
.Y(n_1703)
);

NOR2xp33_ASAP7_75t_L g1704 ( 
.A(n_1398),
.B(n_19),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1393),
.B(n_21),
.Y(n_1705)
);

NAND2xp5_ASAP7_75t_L g1706 ( 
.A(n_1394),
.B(n_21),
.Y(n_1706)
);

OAI21xp5_ASAP7_75t_L g1707 ( 
.A1(n_1541),
.A2(n_551),
.B(n_550),
.Y(n_1707)
);

BUFx6f_ASAP7_75t_L g1708 ( 
.A(n_1537),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1409),
.B(n_22),
.Y(n_1709)
);

AOI21xp5_ASAP7_75t_L g1710 ( 
.A1(n_1456),
.A2(n_553),
.B(n_552),
.Y(n_1710)
);

OR2x6_ASAP7_75t_L g1711 ( 
.A(n_1537),
.B(n_554),
.Y(n_1711)
);

BUFx12f_ASAP7_75t_L g1712 ( 
.A(n_1511),
.Y(n_1712)
);

INVx3_ASAP7_75t_L g1713 ( 
.A(n_1464),
.Y(n_1713)
);

AOI21xp5_ASAP7_75t_L g1714 ( 
.A1(n_1473),
.A2(n_558),
.B(n_556),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1516),
.Y(n_1715)
);

OAI21xp33_ASAP7_75t_L g1716 ( 
.A1(n_1402),
.A2(n_23),
.B(n_24),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1518),
.Y(n_1717)
);

AOI21xp5_ASAP7_75t_L g1718 ( 
.A1(n_1450),
.A2(n_561),
.B(n_560),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1412),
.B(n_23),
.Y(n_1719)
);

NOR2xp33_ASAP7_75t_L g1720 ( 
.A(n_1571),
.B(n_1375),
.Y(n_1720)
);

OAI21xp5_ASAP7_75t_L g1721 ( 
.A1(n_1571),
.A2(n_1477),
.B(n_1429),
.Y(n_1721)
);

O2A1O1Ixp33_ASAP7_75t_L g1722 ( 
.A1(n_1641),
.A2(n_1580),
.B(n_1592),
.C(n_1613),
.Y(n_1722)
);

NOR2xp33_ASAP7_75t_L g1723 ( 
.A(n_1640),
.B(n_1376),
.Y(n_1723)
);

BUFx3_ASAP7_75t_L g1724 ( 
.A(n_1567),
.Y(n_1724)
);

INVx3_ASAP7_75t_L g1725 ( 
.A(n_1708),
.Y(n_1725)
);

NOR3xp33_ASAP7_75t_L g1726 ( 
.A(n_1664),
.B(n_1458),
.C(n_1418),
.Y(n_1726)
);

NAND2xp5_ASAP7_75t_L g1727 ( 
.A(n_1553),
.B(n_1417),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_SL g1728 ( 
.A(n_1583),
.B(n_1549),
.Y(n_1728)
);

NOR2xp33_ASAP7_75t_L g1729 ( 
.A(n_1630),
.B(n_1384),
.Y(n_1729)
);

OAI22xp5_ASAP7_75t_L g1730 ( 
.A1(n_1608),
.A2(n_1519),
.B1(n_1540),
.B2(n_1536),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1554),
.B(n_1386),
.Y(n_1731)
);

O2A1O1Ixp33_ASAP7_75t_SL g1732 ( 
.A1(n_1681),
.A2(n_1422),
.B(n_1426),
.C(n_1404),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1556),
.B(n_1405),
.Y(n_1733)
);

INVx1_ASAP7_75t_SL g1734 ( 
.A(n_1565),
.Y(n_1734)
);

AO21x1_ASAP7_75t_L g1735 ( 
.A1(n_1685),
.A2(n_1497),
.B(n_1544),
.Y(n_1735)
);

NAND2xp5_ASAP7_75t_SL g1736 ( 
.A(n_1632),
.B(n_1497),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1570),
.Y(n_1737)
);

INVx1_ASAP7_75t_SL g1738 ( 
.A(n_1572),
.Y(n_1738)
);

A2O1A1Ixp33_ASAP7_75t_L g1739 ( 
.A1(n_1707),
.A2(n_1528),
.B(n_26),
.C(n_25),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1662),
.B(n_562),
.Y(n_1740)
);

INVx1_ASAP7_75t_L g1741 ( 
.A(n_1598),
.Y(n_1741)
);

INVx1_ASAP7_75t_SL g1742 ( 
.A(n_1575),
.Y(n_1742)
);

INVx2_ASAP7_75t_L g1743 ( 
.A(n_1561),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_SL g1744 ( 
.A(n_1632),
.B(n_28),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1648),
.B(n_29),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1624),
.B(n_1586),
.Y(n_1746)
);

CKINVDCx6p67_ASAP7_75t_R g1747 ( 
.A(n_1652),
.Y(n_1747)
);

AND2x6_ASAP7_75t_L g1748 ( 
.A(n_1691),
.B(n_565),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1590),
.Y(n_1749)
);

AOI22xp5_ASAP7_75t_L g1750 ( 
.A1(n_1617),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_1750)
);

CKINVDCx10_ASAP7_75t_R g1751 ( 
.A(n_1652),
.Y(n_1751)
);

O2A1O1Ixp33_ASAP7_75t_L g1752 ( 
.A1(n_1576),
.A2(n_33),
.B(n_30),
.C(n_32),
.Y(n_1752)
);

INVxp67_ASAP7_75t_L g1753 ( 
.A(n_1639),
.Y(n_1753)
);

BUFx6f_ASAP7_75t_L g1754 ( 
.A(n_1585),
.Y(n_1754)
);

NOR3xp33_ASAP7_75t_L g1755 ( 
.A(n_1665),
.B(n_32),
.C(n_33),
.Y(n_1755)
);

INVx2_ASAP7_75t_L g1756 ( 
.A(n_1597),
.Y(n_1756)
);

AOI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1587),
.A2(n_588),
.B(n_567),
.Y(n_1757)
);

NAND2xp5_ASAP7_75t_SL g1758 ( 
.A(n_1632),
.B(n_1650),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1601),
.Y(n_1759)
);

O2A1O1Ixp33_ASAP7_75t_L g1760 ( 
.A1(n_1577),
.A2(n_37),
.B(n_35),
.C(n_36),
.Y(n_1760)
);

O2A1O1Ixp33_ASAP7_75t_SL g1761 ( 
.A1(n_1699),
.A2(n_38),
.B(n_36),
.C(n_37),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_L g1762 ( 
.A(n_1588),
.B(n_566),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1614),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1595),
.B(n_38),
.Y(n_1764)
);

AOI21xp5_ASAP7_75t_L g1765 ( 
.A1(n_1589),
.A2(n_569),
.B(n_568),
.Y(n_1765)
);

AND2x4_ASAP7_75t_SL g1766 ( 
.A(n_1651),
.B(n_571),
.Y(n_1766)
);

NOR2xp33_ASAP7_75t_SL g1767 ( 
.A(n_1654),
.B(n_572),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_SL g1768 ( 
.A(n_1650),
.B(n_39),
.Y(n_1768)
);

NAND2xp5_ASAP7_75t_L g1769 ( 
.A(n_1619),
.B(n_39),
.Y(n_1769)
);

HB1xp67_ASAP7_75t_L g1770 ( 
.A(n_1657),
.Y(n_1770)
);

A2O1A1Ixp33_ASAP7_75t_L g1771 ( 
.A1(n_1686),
.A2(n_42),
.B(n_40),
.C(n_41),
.Y(n_1771)
);

A2O1A1Ixp33_ASAP7_75t_SL g1772 ( 
.A1(n_1701),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_1772)
);

AOI21xp5_ASAP7_75t_L g1773 ( 
.A1(n_1564),
.A2(n_1702),
.B(n_1562),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1599),
.B(n_573),
.Y(n_1774)
);

O2A1O1Ixp33_ASAP7_75t_L g1775 ( 
.A1(n_1704),
.A2(n_46),
.B(n_43),
.C(n_44),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_SL g1776 ( 
.A(n_1650),
.B(n_46),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1569),
.A2(n_49),
.B1(n_47),
.B2(n_48),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_L g1778 ( 
.A(n_1621),
.B(n_576),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_L g1779 ( 
.A(n_1594),
.B(n_47),
.Y(n_1779)
);

A2O1A1Ixp33_ASAP7_75t_L g1780 ( 
.A1(n_1676),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_1780)
);

NAND2xp5_ASAP7_75t_L g1781 ( 
.A(n_1607),
.B(n_50),
.Y(n_1781)
);

BUFx6f_ASAP7_75t_L g1782 ( 
.A(n_1585),
.Y(n_1782)
);

INVx2_ASAP7_75t_L g1783 ( 
.A(n_1618),
.Y(n_1783)
);

NOR2xp33_ASAP7_75t_L g1784 ( 
.A(n_1628),
.B(n_580),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1622),
.Y(n_1785)
);

NAND3xp33_ASAP7_75t_L g1786 ( 
.A(n_1682),
.B(n_52),
.C(n_53),
.Y(n_1786)
);

AOI21xp5_ASAP7_75t_L g1787 ( 
.A1(n_1684),
.A2(n_585),
.B(n_582),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1649),
.Y(n_1788)
);

INVx2_ASAP7_75t_L g1789 ( 
.A(n_1642),
.Y(n_1789)
);

AND2x2_ASAP7_75t_L g1790 ( 
.A(n_1659),
.B(n_54),
.Y(n_1790)
);

INVx2_ASAP7_75t_L g1791 ( 
.A(n_1643),
.Y(n_1791)
);

NOR2xp33_ASAP7_75t_L g1792 ( 
.A(n_1615),
.B(n_581),
.Y(n_1792)
);

NOR2xp33_ASAP7_75t_L g1793 ( 
.A(n_1568),
.B(n_584),
.Y(n_1793)
);

A2O1A1Ixp33_ASAP7_75t_L g1794 ( 
.A1(n_1596),
.A2(n_1716),
.B(n_1631),
.C(n_1658),
.Y(n_1794)
);

AND2x2_ASAP7_75t_L g1795 ( 
.A(n_1694),
.B(n_55),
.Y(n_1795)
);

CKINVDCx5p33_ASAP7_75t_R g1796 ( 
.A(n_1663),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1612),
.B(n_56),
.Y(n_1797)
);

O2A1O1Ixp33_ASAP7_75t_SL g1798 ( 
.A1(n_1558),
.A2(n_58),
.B(n_56),
.C(n_57),
.Y(n_1798)
);

AOI22xp5_ASAP7_75t_L g1799 ( 
.A1(n_1716),
.A2(n_60),
.B1(n_57),
.B2(n_59),
.Y(n_1799)
);

INVx4_ASAP7_75t_L g1800 ( 
.A(n_1567),
.Y(n_1800)
);

A2O1A1Ixp33_ASAP7_75t_L g1801 ( 
.A1(n_1679),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1801)
);

AOI21xp5_ASAP7_75t_L g1802 ( 
.A1(n_1573),
.A2(n_501),
.B(n_61),
.Y(n_1802)
);

NAND2xp5_ASAP7_75t_L g1803 ( 
.A(n_1670),
.B(n_1671),
.Y(n_1803)
);

AOI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1555),
.A2(n_63),
.B(n_64),
.Y(n_1804)
);

OA22x2_ASAP7_75t_L g1805 ( 
.A1(n_1692),
.A2(n_67),
.B1(n_64),
.B2(n_66),
.Y(n_1805)
);

AOI21xp5_ASAP7_75t_L g1806 ( 
.A1(n_1559),
.A2(n_501),
.B(n_67),
.Y(n_1806)
);

AOI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1669),
.A2(n_70),
.B1(n_68),
.B2(n_69),
.Y(n_1807)
);

INVx1_ASAP7_75t_L g1808 ( 
.A(n_1668),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1660),
.A2(n_73),
.B1(n_71),
.B2(n_72),
.Y(n_1809)
);

AOI21xp5_ASAP7_75t_L g1810 ( 
.A1(n_1602),
.A2(n_500),
.B(n_74),
.Y(n_1810)
);

NOR2xp33_ASAP7_75t_L g1811 ( 
.A(n_1636),
.B(n_75),
.Y(n_1811)
);

BUFx6f_ASAP7_75t_L g1812 ( 
.A(n_1567),
.Y(n_1812)
);

AOI21xp5_ASAP7_75t_L g1813 ( 
.A1(n_1605),
.A2(n_500),
.B(n_76),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1674),
.Y(n_1814)
);

NOR2xp33_ASAP7_75t_L g1815 ( 
.A(n_1638),
.B(n_77),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_SL g1816 ( 
.A(n_1660),
.B(n_78),
.Y(n_1816)
);

CKINVDCx5p33_ASAP7_75t_R g1817 ( 
.A(n_1644),
.Y(n_1817)
);

NAND2xp5_ASAP7_75t_L g1818 ( 
.A(n_1660),
.B(n_78),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1610),
.A2(n_499),
.B(n_79),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1645),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1677),
.A2(n_1690),
.B1(n_1606),
.B2(n_1712),
.Y(n_1821)
);

NAND3xp33_ASAP7_75t_L g1822 ( 
.A(n_1653),
.B(n_79),
.C(n_80),
.Y(n_1822)
);

BUFx12f_ASAP7_75t_L g1823 ( 
.A(n_1697),
.Y(n_1823)
);

NOR2xp33_ASAP7_75t_L g1824 ( 
.A(n_1651),
.B(n_80),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1609),
.B(n_81),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1688),
.Y(n_1826)
);

O2A1O1Ixp33_ASAP7_75t_L g1827 ( 
.A1(n_1566),
.A2(n_1689),
.B(n_1687),
.C(n_1584),
.Y(n_1827)
);

CKINVDCx16_ASAP7_75t_R g1828 ( 
.A(n_1629),
.Y(n_1828)
);

AOI22xp5_ASAP7_75t_L g1829 ( 
.A1(n_1634),
.A2(n_84),
.B1(n_81),
.B2(n_82),
.Y(n_1829)
);

INVx1_ASAP7_75t_L g1830 ( 
.A(n_1698),
.Y(n_1830)
);

OAI22x1_ASAP7_75t_L g1831 ( 
.A1(n_1693),
.A2(n_88),
.B1(n_85),
.B2(n_86),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1673),
.B(n_85),
.Y(n_1832)
);

INVx1_ASAP7_75t_L g1833 ( 
.A(n_1700),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1655),
.Y(n_1834)
);

AND2x6_ASAP7_75t_L g1835 ( 
.A(n_1708),
.B(n_86),
.Y(n_1835)
);

NAND2xp5_ASAP7_75t_L g1836 ( 
.A(n_1552),
.B(n_88),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1683),
.B(n_89),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1695),
.B(n_90),
.Y(n_1838)
);

NOR2xp33_ASAP7_75t_L g1839 ( 
.A(n_1603),
.B(n_90),
.Y(n_1839)
);

OR2x6_ASAP7_75t_SL g1840 ( 
.A(n_1696),
.B(n_499),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1715),
.B(n_1717),
.Y(n_1841)
);

AOI21xp5_ASAP7_75t_L g1842 ( 
.A1(n_1574),
.A2(n_91),
.B(n_92),
.Y(n_1842)
);

OAI22xp5_ASAP7_75t_L g1843 ( 
.A1(n_1609),
.A2(n_94),
.B1(n_92),
.B2(n_93),
.Y(n_1843)
);

INVx3_ASAP7_75t_SL g1844 ( 
.A(n_1644),
.Y(n_1844)
);

OAI22x1_ASAP7_75t_L g1845 ( 
.A1(n_1557),
.A2(n_95),
.B1(n_93),
.B2(n_94),
.Y(n_1845)
);

NAND2xp33_ASAP7_75t_L g1846 ( 
.A(n_1708),
.B(n_96),
.Y(n_1846)
);

OR2x6_ASAP7_75t_SL g1847 ( 
.A(n_1705),
.B(n_497),
.Y(n_1847)
);

INVx5_ASAP7_75t_L g1848 ( 
.A(n_1644),
.Y(n_1848)
);

AOI22xp5_ASAP7_75t_L g1849 ( 
.A1(n_1600),
.A2(n_98),
.B1(n_96),
.B2(n_97),
.Y(n_1849)
);

AOI22xp5_ASAP7_75t_L g1850 ( 
.A1(n_1616),
.A2(n_99),
.B1(n_97),
.B2(n_98),
.Y(n_1850)
);

AO21x1_ASAP7_75t_L g1851 ( 
.A1(n_1626),
.A2(n_99),
.B(n_100),
.Y(n_1851)
);

NOR2xp33_ASAP7_75t_L g1852 ( 
.A(n_1706),
.B(n_100),
.Y(n_1852)
);

NAND2xp33_ASAP7_75t_SL g1853 ( 
.A(n_1709),
.B(n_101),
.Y(n_1853)
);

INVx3_ASAP7_75t_L g1854 ( 
.A(n_1703),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1719),
.B(n_102),
.Y(n_1855)
);

AOI21xp5_ASAP7_75t_L g1856 ( 
.A1(n_1578),
.A2(n_104),
.B(n_105),
.Y(n_1856)
);

AOI22xp33_ASAP7_75t_L g1857 ( 
.A1(n_1563),
.A2(n_106),
.B1(n_104),
.B2(n_105),
.Y(n_1857)
);

AO21x1_ASAP7_75t_L g1858 ( 
.A1(n_1647),
.A2(n_106),
.B(n_108),
.Y(n_1858)
);

OAI21xp33_ASAP7_75t_L g1859 ( 
.A1(n_1582),
.A2(n_1661),
.B(n_1625),
.Y(n_1859)
);

NAND2xp5_ASAP7_75t_L g1860 ( 
.A(n_1591),
.B(n_108),
.Y(n_1860)
);

AOI21xp5_ASAP7_75t_L g1861 ( 
.A1(n_1646),
.A2(n_109),
.B(n_110),
.Y(n_1861)
);

CKINVDCx11_ASAP7_75t_R g1862 ( 
.A(n_1666),
.Y(n_1862)
);

O2A1O1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1637),
.A2(n_111),
.B(n_109),
.C(n_110),
.Y(n_1863)
);

INVx3_ASAP7_75t_L g1864 ( 
.A(n_1703),
.Y(n_1864)
);

O2A1O1Ixp33_ASAP7_75t_L g1865 ( 
.A1(n_1611),
.A2(n_1623),
.B(n_1627),
.C(n_1667),
.Y(n_1865)
);

AOI21xp5_ASAP7_75t_L g1866 ( 
.A1(n_1620),
.A2(n_111),
.B(n_112),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1713),
.B(n_112),
.Y(n_1867)
);

AO21x1_ASAP7_75t_L g1868 ( 
.A1(n_1672),
.A2(n_114),
.B(n_116),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1579),
.B(n_116),
.Y(n_1869)
);

AOI22xp33_ASAP7_75t_SL g1870 ( 
.A1(n_1666),
.A2(n_119),
.B1(n_117),
.B2(n_118),
.Y(n_1870)
);

AOI21xp5_ASAP7_75t_L g1871 ( 
.A1(n_1675),
.A2(n_117),
.B(n_120),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1579),
.B(n_120),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1722),
.A2(n_1678),
.B(n_1656),
.Y(n_1873)
);

AOI21xp5_ASAP7_75t_L g1874 ( 
.A1(n_1773),
.A2(n_1714),
.B(n_1710),
.Y(n_1874)
);

OAI21xp5_ASAP7_75t_L g1875 ( 
.A1(n_1794),
.A2(n_1581),
.B(n_1718),
.Y(n_1875)
);

OAI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1821),
.A2(n_1666),
.B1(n_1711),
.B2(n_1604),
.Y(n_1876)
);

AOI21xp5_ASAP7_75t_L g1877 ( 
.A1(n_1865),
.A2(n_1787),
.B(n_1765),
.Y(n_1877)
);

BUFx6f_ASAP7_75t_L g1878 ( 
.A(n_1754),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1743),
.Y(n_1879)
);

NOR2xp33_ASAP7_75t_L g1880 ( 
.A(n_1803),
.B(n_1635),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1795),
.B(n_1711),
.Y(n_1881)
);

BUFx2_ASAP7_75t_L g1882 ( 
.A(n_1770),
.Y(n_1882)
);

AOI21xp5_ASAP7_75t_L g1883 ( 
.A1(n_1757),
.A2(n_1711),
.B(n_1604),
.Y(n_1883)
);

NAND3x1_ASAP7_75t_L g1884 ( 
.A(n_1755),
.B(n_1680),
.C(n_1635),
.Y(n_1884)
);

BUFx3_ASAP7_75t_L g1885 ( 
.A(n_1812),
.Y(n_1885)
);

AOI21xp5_ASAP7_75t_L g1886 ( 
.A1(n_1721),
.A2(n_1593),
.B(n_1560),
.Y(n_1886)
);

OAI21xp5_ASAP7_75t_SL g1887 ( 
.A1(n_1750),
.A2(n_1633),
.B(n_1680),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1737),
.Y(n_1888)
);

AND2x4_ASAP7_75t_L g1889 ( 
.A(n_1848),
.B(n_1593),
.Y(n_1889)
);

NOR2xp33_ASAP7_75t_L g1890 ( 
.A(n_1738),
.B(n_121),
.Y(n_1890)
);

NAND3x1_ASAP7_75t_L g1891 ( 
.A(n_1807),
.B(n_121),
.C(n_122),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1746),
.B(n_497),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1749),
.Y(n_1893)
);

OR2x2_ASAP7_75t_L g1894 ( 
.A(n_1841),
.B(n_123),
.Y(n_1894)
);

CKINVDCx5p33_ASAP7_75t_R g1895 ( 
.A(n_1751),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1727),
.B(n_124),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1741),
.B(n_125),
.Y(n_1897)
);

NAND2x1p5_ASAP7_75t_L g1898 ( 
.A(n_1848),
.B(n_126),
.Y(n_1898)
);

AO31x2_ASAP7_75t_L g1899 ( 
.A1(n_1739),
.A2(n_129),
.A3(n_127),
.B(n_128),
.Y(n_1899)
);

NOR2x1_ASAP7_75t_R g1900 ( 
.A(n_1862),
.B(n_128),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1720),
.B(n_130),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1731),
.B(n_1832),
.Y(n_1902)
);

AND2x4_ASAP7_75t_L g1903 ( 
.A(n_1848),
.B(n_1800),
.Y(n_1903)
);

OAI22xp5_ASAP7_75t_L g1904 ( 
.A1(n_1799),
.A2(n_133),
.B1(n_131),
.B2(n_132),
.Y(n_1904)
);

AO21x1_ASAP7_75t_L g1905 ( 
.A1(n_1863),
.A2(n_134),
.B(n_137),
.Y(n_1905)
);

AO31x2_ASAP7_75t_L g1906 ( 
.A1(n_1868),
.A2(n_140),
.A3(n_138),
.B(n_139),
.Y(n_1906)
);

OAI21x1_ASAP7_75t_L g1907 ( 
.A1(n_1806),
.A2(n_139),
.B(n_141),
.Y(n_1907)
);

BUFx2_ASAP7_75t_L g1908 ( 
.A(n_1742),
.Y(n_1908)
);

AOI21xp5_ASAP7_75t_L g1909 ( 
.A1(n_1859),
.A2(n_141),
.B(n_142),
.Y(n_1909)
);

OAI21xp5_ASAP7_75t_L g1910 ( 
.A1(n_1827),
.A2(n_142),
.B(n_143),
.Y(n_1910)
);

AOI21xp5_ASAP7_75t_L g1911 ( 
.A1(n_1861),
.A2(n_143),
.B(n_144),
.Y(n_1911)
);

NAND3xp33_ASAP7_75t_L g1912 ( 
.A(n_1811),
.B(n_144),
.C(n_145),
.Y(n_1912)
);

O2A1O1Ixp5_ASAP7_75t_L g1913 ( 
.A1(n_1851),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1913)
);

NAND2xp5_ASAP7_75t_L g1914 ( 
.A(n_1852),
.B(n_146),
.Y(n_1914)
);

AO31x2_ASAP7_75t_L g1915 ( 
.A1(n_1858),
.A2(n_150),
.A3(n_148),
.B(n_149),
.Y(n_1915)
);

INVx1_ASAP7_75t_L g1916 ( 
.A(n_1763),
.Y(n_1916)
);

BUFx8_ASAP7_75t_L g1917 ( 
.A(n_1823),
.Y(n_1917)
);

OAI21xp5_ASAP7_75t_L g1918 ( 
.A1(n_1871),
.A2(n_152),
.B(n_153),
.Y(n_1918)
);

NAND3x1_ASAP7_75t_L g1919 ( 
.A(n_1815),
.B(n_153),
.C(n_154),
.Y(n_1919)
);

OAI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1801),
.A2(n_155),
.B(n_157),
.Y(n_1920)
);

AOI21xp5_ASAP7_75t_L g1921 ( 
.A1(n_1740),
.A2(n_155),
.B(n_157),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1800),
.B(n_158),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1730),
.B(n_158),
.Y(n_1923)
);

OAI21x1_ASAP7_75t_L g1924 ( 
.A1(n_1866),
.A2(n_159),
.B(n_160),
.Y(n_1924)
);

NAND4xp25_ASAP7_75t_L g1925 ( 
.A(n_1839),
.B(n_161),
.C(n_159),
.D(n_160),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_L g1926 ( 
.A(n_1756),
.B(n_496),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1732),
.A2(n_161),
.B(n_162),
.Y(n_1927)
);

OAI21x1_ASAP7_75t_L g1928 ( 
.A1(n_1810),
.A2(n_162),
.B(n_163),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1785),
.Y(n_1929)
);

OAI21x1_ASAP7_75t_L g1930 ( 
.A1(n_1813),
.A2(n_164),
.B(n_165),
.Y(n_1930)
);

OAI21xp33_ASAP7_75t_L g1931 ( 
.A1(n_1771),
.A2(n_164),
.B(n_165),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1726),
.A2(n_166),
.B(n_167),
.Y(n_1932)
);

INVx2_ASAP7_75t_SL g1933 ( 
.A(n_1812),
.Y(n_1933)
);

NOR2x1_ASAP7_75t_L g1934 ( 
.A(n_1822),
.B(n_166),
.Y(n_1934)
);

CKINVDCx5p33_ASAP7_75t_R g1935 ( 
.A(n_1751),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1774),
.B(n_167),
.Y(n_1936)
);

CKINVDCx11_ASAP7_75t_R g1937 ( 
.A(n_1747),
.Y(n_1937)
);

BUFx6f_ASAP7_75t_L g1938 ( 
.A(n_1754),
.Y(n_1938)
);

AOI21x1_ASAP7_75t_L g1939 ( 
.A1(n_1804),
.A2(n_168),
.B(n_169),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1788),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1736),
.A2(n_168),
.B(n_169),
.Y(n_1941)
);

INVx1_ASAP7_75t_L g1942 ( 
.A(n_1808),
.Y(n_1942)
);

AOI21xp5_ASAP7_75t_SL g1943 ( 
.A1(n_1778),
.A2(n_170),
.B(n_171),
.Y(n_1943)
);

OAI21x1_ASAP7_75t_L g1944 ( 
.A1(n_1819),
.A2(n_171),
.B(n_172),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1792),
.B(n_172),
.Y(n_1945)
);

AO31x2_ASAP7_75t_L g1946 ( 
.A1(n_1735),
.A2(n_1856),
.A3(n_1814),
.B(n_1830),
.Y(n_1946)
);

INVx5_ASAP7_75t_L g1947 ( 
.A(n_1748),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1828),
.A2(n_175),
.B1(n_173),
.B2(n_174),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_SL g1949 ( 
.A1(n_1775),
.A2(n_173),
.B(n_174),
.Y(n_1949)
);

OAI21x1_ASAP7_75t_L g1950 ( 
.A1(n_1842),
.A2(n_176),
.B(n_177),
.Y(n_1950)
);

OAI21xp5_ASAP7_75t_L g1951 ( 
.A1(n_1786),
.A2(n_176),
.B(n_177),
.Y(n_1951)
);

OAI21x1_ASAP7_75t_L g1952 ( 
.A1(n_1802),
.A2(n_178),
.B(n_179),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_L g1953 ( 
.A(n_1759),
.B(n_494),
.Y(n_1953)
);

INVxp67_ASAP7_75t_SL g1954 ( 
.A(n_1723),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1753),
.A2(n_180),
.B1(n_178),
.B2(n_179),
.Y(n_1955)
);

OAI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1825),
.A2(n_183),
.B1(n_181),
.B2(n_182),
.Y(n_1956)
);

OAI21xp5_ASAP7_75t_L g1957 ( 
.A1(n_1752),
.A2(n_181),
.B(n_183),
.Y(n_1957)
);

NAND2xp5_ASAP7_75t_SL g1958 ( 
.A(n_1733),
.B(n_184),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1783),
.B(n_494),
.Y(n_1959)
);

OAI21x1_ASAP7_75t_L g1960 ( 
.A1(n_1854),
.A2(n_184),
.B(n_185),
.Y(n_1960)
);

A2O1A1Ixp33_ASAP7_75t_L g1961 ( 
.A1(n_1760),
.A2(n_187),
.B(n_185),
.C(n_186),
.Y(n_1961)
);

NAND3x1_ASAP7_75t_L g1962 ( 
.A(n_1849),
.B(n_186),
.C(n_187),
.Y(n_1962)
);

O2A1O1Ixp33_ASAP7_75t_SL g1963 ( 
.A1(n_1772),
.A2(n_190),
.B(n_188),
.C(n_189),
.Y(n_1963)
);

INVx2_ASAP7_75t_SL g1964 ( 
.A(n_1812),
.Y(n_1964)
);

NOR2xp33_ASAP7_75t_L g1965 ( 
.A(n_1734),
.B(n_189),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1789),
.B(n_190),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1791),
.B(n_1820),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1834),
.B(n_493),
.Y(n_1968)
);

OAI21xp5_ASAP7_75t_L g1969 ( 
.A1(n_1860),
.A2(n_191),
.B(n_193),
.Y(n_1969)
);

INVx1_ASAP7_75t_L g1970 ( 
.A(n_1826),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_L g1971 ( 
.A(n_1728),
.B(n_191),
.Y(n_1971)
);

AOI21xp5_ASAP7_75t_L g1972 ( 
.A1(n_1761),
.A2(n_193),
.B(n_194),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_L g1973 ( 
.A(n_1836),
.B(n_1855),
.Y(n_1973)
);

OAI21xp33_ASAP7_75t_L g1974 ( 
.A1(n_1829),
.A2(n_1780),
.B(n_1777),
.Y(n_1974)
);

OAI21x1_ASAP7_75t_L g1975 ( 
.A1(n_1854),
.A2(n_194),
.B(n_195),
.Y(n_1975)
);

NOR2x1_ASAP7_75t_L g1976 ( 
.A(n_1864),
.B(n_195),
.Y(n_1976)
);

OAI22xp5_ASAP7_75t_L g1977 ( 
.A1(n_1870),
.A2(n_198),
.B1(n_196),
.B2(n_197),
.Y(n_1977)
);

INVx5_ASAP7_75t_L g1978 ( 
.A(n_1947),
.Y(n_1978)
);

BUFx2_ASAP7_75t_L g1979 ( 
.A(n_1882),
.Y(n_1979)
);

AOI21xp5_ASAP7_75t_SL g1980 ( 
.A1(n_1910),
.A2(n_1805),
.B(n_1793),
.Y(n_1980)
);

INVx3_ASAP7_75t_SL g1981 ( 
.A(n_1895),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1888),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1954),
.B(n_1729),
.Y(n_1983)
);

NOR2xp33_ASAP7_75t_L g1984 ( 
.A(n_1902),
.B(n_1797),
.Y(n_1984)
);

HB1xp67_ASAP7_75t_L g1985 ( 
.A(n_1946),
.Y(n_1985)
);

INVx5_ASAP7_75t_L g1986 ( 
.A(n_1947),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_L g1987 ( 
.A(n_1888),
.B(n_1833),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1916),
.Y(n_1988)
);

INVx3_ASAP7_75t_L g1989 ( 
.A(n_1903),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1916),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1881),
.B(n_1790),
.Y(n_1991)
);

INVx3_ASAP7_75t_SL g1992 ( 
.A(n_1935),
.Y(n_1992)
);

INVx4_ASAP7_75t_L g1993 ( 
.A(n_1903),
.Y(n_1993)
);

AND2x4_ASAP7_75t_L g1994 ( 
.A(n_1929),
.B(n_1940),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1929),
.B(n_1745),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1940),
.B(n_1764),
.Y(n_1996)
);

CKINVDCx16_ASAP7_75t_R g1997 ( 
.A(n_1885),
.Y(n_1997)
);

AOI22xp5_ASAP7_75t_L g1998 ( 
.A1(n_1974),
.A2(n_1853),
.B1(n_1846),
.B2(n_1843),
.Y(n_1998)
);

BUFx8_ASAP7_75t_L g1999 ( 
.A(n_1878),
.Y(n_1999)
);

INVx1_ASAP7_75t_SL g2000 ( 
.A(n_1908),
.Y(n_2000)
);

HB1xp67_ASAP7_75t_L g2001 ( 
.A(n_1946),
.Y(n_2001)
);

INVx2_ASAP7_75t_L g2002 ( 
.A(n_1942),
.Y(n_2002)
);

INVx2_ASAP7_75t_SL g2003 ( 
.A(n_1878),
.Y(n_2003)
);

BUFx3_ASAP7_75t_L g2004 ( 
.A(n_1917),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1880),
.B(n_1824),
.Y(n_2005)
);

BUFx3_ASAP7_75t_L g2006 ( 
.A(n_1917),
.Y(n_2006)
);

AOI21xp5_ASAP7_75t_L g2007 ( 
.A1(n_1877),
.A2(n_1798),
.B(n_1766),
.Y(n_2007)
);

OR2x2_ASAP7_75t_L g2008 ( 
.A(n_1942),
.B(n_1818),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1970),
.B(n_1769),
.Y(n_2009)
);

INVx1_ASAP7_75t_L g2010 ( 
.A(n_1970),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_L g2011 ( 
.A(n_1973),
.B(n_1779),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1946),
.Y(n_2012)
);

INVx2_ASAP7_75t_L g2013 ( 
.A(n_1879),
.Y(n_2013)
);

INVx2_ASAP7_75t_L g2014 ( 
.A(n_1893),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1967),
.Y(n_2015)
);

AND2x2_ASAP7_75t_L g2016 ( 
.A(n_1894),
.B(n_1867),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1901),
.B(n_1758),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1926),
.Y(n_2018)
);

OR2x6_ASAP7_75t_L g2019 ( 
.A(n_1883),
.B(n_1724),
.Y(n_2019)
);

BUFx3_ASAP7_75t_L g2020 ( 
.A(n_1878),
.Y(n_2020)
);

BUFx2_ASAP7_75t_L g2021 ( 
.A(n_1933),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1947),
.B(n_1889),
.Y(n_2022)
);

CKINVDCx5p33_ASAP7_75t_R g2023 ( 
.A(n_1937),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1953),
.Y(n_2024)
);

BUFx6f_ASAP7_75t_L g2025 ( 
.A(n_1938),
.Y(n_2025)
);

INVx3_ASAP7_75t_L g2026 ( 
.A(n_1938),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1906),
.Y(n_2027)
);

BUFx6f_ASAP7_75t_L g2028 ( 
.A(n_1938),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_SL g2029 ( 
.A(n_1900),
.B(n_1796),
.Y(n_2029)
);

BUFx6f_ASAP7_75t_L g2030 ( 
.A(n_1964),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_L g2031 ( 
.A(n_1915),
.B(n_1837),
.Y(n_2031)
);

AOI21xp5_ASAP7_75t_L g2032 ( 
.A1(n_1874),
.A2(n_1857),
.B(n_1768),
.Y(n_2032)
);

AND2x2_ASAP7_75t_L g2033 ( 
.A(n_1897),
.B(n_1781),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1922),
.Y(n_2034)
);

OAI22xp5_ASAP7_75t_L g2035 ( 
.A1(n_1919),
.A2(n_1840),
.B1(n_1847),
.B2(n_1809),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1896),
.B(n_1838),
.Y(n_2036)
);

INVx3_ASAP7_75t_L g2037 ( 
.A(n_1922),
.Y(n_2037)
);

AOI22xp33_ASAP7_75t_L g2038 ( 
.A1(n_1931),
.A2(n_1831),
.B1(n_1845),
.B2(n_1850),
.Y(n_2038)
);

OAI21xp5_ASAP7_75t_L g2039 ( 
.A1(n_1873),
.A2(n_1776),
.B(n_1744),
.Y(n_2039)
);

AND2x4_ASAP7_75t_L g2040 ( 
.A(n_1976),
.B(n_1725),
.Y(n_2040)
);

INVx4_ASAP7_75t_L g2041 ( 
.A(n_1898),
.Y(n_2041)
);

AOI21xp5_ASAP7_75t_L g2042 ( 
.A1(n_1886),
.A2(n_1816),
.B(n_1767),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1891),
.A2(n_1912),
.B1(n_1962),
.B2(n_1904),
.Y(n_2043)
);

NOR2xp33_ASAP7_75t_L g2044 ( 
.A(n_1892),
.B(n_1762),
.Y(n_2044)
);

AOI21xp5_ASAP7_75t_L g2045 ( 
.A1(n_1875),
.A2(n_1872),
.B(n_1869),
.Y(n_2045)
);

INVx6_ASAP7_75t_L g2046 ( 
.A(n_1999),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_L g2047 ( 
.A(n_1994),
.B(n_1899),
.Y(n_2047)
);

AOI22xp5_ASAP7_75t_L g2048 ( 
.A1(n_2043),
.A2(n_1957),
.B1(n_1876),
.B2(n_1905),
.Y(n_2048)
);

BUFx4f_ASAP7_75t_SL g2049 ( 
.A(n_1981),
.Y(n_2049)
);

AOI22xp33_ASAP7_75t_L g2050 ( 
.A1(n_2043),
.A2(n_1920),
.B1(n_1918),
.B2(n_1925),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_SL g2051 ( 
.A1(n_2035),
.A2(n_1969),
.B1(n_1951),
.B2(n_1977),
.Y(n_2051)
);

OAI22xp33_ASAP7_75t_L g2052 ( 
.A1(n_1998),
.A2(n_1972),
.B1(n_1909),
.B2(n_1923),
.Y(n_2052)
);

BUFx2_ASAP7_75t_SL g2053 ( 
.A(n_2004),
.Y(n_2053)
);

INVx1_ASAP7_75t_L g2054 ( 
.A(n_1994),
.Y(n_2054)
);

OAI22xp5_ASAP7_75t_L g2055 ( 
.A1(n_2038),
.A2(n_2035),
.B1(n_1980),
.B2(n_1961),
.Y(n_2055)
);

AO22x1_ASAP7_75t_L g2056 ( 
.A1(n_1978),
.A2(n_1934),
.B1(n_1835),
.B2(n_1844),
.Y(n_2056)
);

INVx6_ASAP7_75t_SL g2057 ( 
.A(n_2019),
.Y(n_2057)
);

BUFx6f_ASAP7_75t_L g2058 ( 
.A(n_2025),
.Y(n_2058)
);

OAI22xp5_ASAP7_75t_L g2059 ( 
.A1(n_2038),
.A2(n_1943),
.B1(n_1914),
.B2(n_1936),
.Y(n_2059)
);

AOI22xp33_ASAP7_75t_SL g2060 ( 
.A1(n_2039),
.A2(n_2044),
.B1(n_2007),
.B2(n_1949),
.Y(n_2060)
);

OAI22xp5_ASAP7_75t_L g2061 ( 
.A1(n_1984),
.A2(n_1945),
.B1(n_1884),
.B2(n_1958),
.Y(n_2061)
);

OAI22xp5_ASAP7_75t_L g2062 ( 
.A1(n_1984),
.A2(n_1956),
.B1(n_1921),
.B2(n_1932),
.Y(n_2062)
);

OAI22xp33_ASAP7_75t_L g2063 ( 
.A1(n_2007),
.A2(n_1971),
.B1(n_1948),
.B2(n_1927),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_2002),
.Y(n_2064)
);

INVx6_ASAP7_75t_L g2065 ( 
.A(n_1999),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_2025),
.Y(n_2066)
);

INVx1_ASAP7_75t_SL g2067 ( 
.A(n_2000),
.Y(n_2067)
);

INVx4_ASAP7_75t_L g2068 ( 
.A(n_2025),
.Y(n_2068)
);

INVx2_ASAP7_75t_L g2069 ( 
.A(n_1982),
.Y(n_2069)
);

INVx2_ASAP7_75t_L g2070 ( 
.A(n_1988),
.Y(n_2070)
);

INVx2_ASAP7_75t_L g2071 ( 
.A(n_1990),
.Y(n_2071)
);

INVx3_ASAP7_75t_L g2072 ( 
.A(n_1993),
.Y(n_2072)
);

INVx2_ASAP7_75t_L g2073 ( 
.A(n_2010),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_2023),
.Y(n_2074)
);

INVx6_ASAP7_75t_L g2075 ( 
.A(n_1978),
.Y(n_2075)
);

INVx4_ASAP7_75t_L g2076 ( 
.A(n_2028),
.Y(n_2076)
);

CKINVDCx5p33_ASAP7_75t_R g2077 ( 
.A(n_1981),
.Y(n_2077)
);

INVx3_ASAP7_75t_L g2078 ( 
.A(n_1993),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1987),
.Y(n_2079)
);

INVx2_ASAP7_75t_L g2080 ( 
.A(n_1987),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_2013),
.Y(n_2081)
);

AOI22xp33_ASAP7_75t_L g2082 ( 
.A1(n_2042),
.A2(n_1911),
.B1(n_1835),
.B2(n_1748),
.Y(n_2082)
);

CKINVDCx11_ASAP7_75t_R g2083 ( 
.A(n_1992),
.Y(n_2083)
);

BUFx2_ASAP7_75t_L g2084 ( 
.A(n_1989),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2014),
.Y(n_2085)
);

INVx6_ASAP7_75t_L g2086 ( 
.A(n_1978),
.Y(n_2086)
);

CKINVDCx6p67_ASAP7_75t_R g2087 ( 
.A(n_1992),
.Y(n_2087)
);

INVx6_ASAP7_75t_L g2088 ( 
.A(n_1978),
.Y(n_2088)
);

OR2x2_ASAP7_75t_L g2089 ( 
.A(n_1979),
.B(n_1899),
.Y(n_2089)
);

BUFx12f_ASAP7_75t_L g2090 ( 
.A(n_2006),
.Y(n_2090)
);

BUFx8_ASAP7_75t_L g2091 ( 
.A(n_2028),
.Y(n_2091)
);

INVx2_ASAP7_75t_L g2092 ( 
.A(n_2015),
.Y(n_2092)
);

AOI22xp33_ASAP7_75t_SL g2093 ( 
.A1(n_2039),
.A2(n_1835),
.B1(n_1890),
.B2(n_1952),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2047),
.B(n_2027),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_2069),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_L g2096 ( 
.A(n_2079),
.B(n_2080),
.Y(n_2096)
);

INVxp67_ASAP7_75t_L g2097 ( 
.A(n_2054),
.Y(n_2097)
);

INVx2_ASAP7_75t_L g2098 ( 
.A(n_2070),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2047),
.B(n_1985),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_SL g2100 ( 
.A1(n_2055),
.A2(n_1784),
.B(n_1965),
.C(n_2045),
.Y(n_2100)
);

INVx3_ASAP7_75t_L g2101 ( 
.A(n_2075),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_2084),
.B(n_2001),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_2081),
.B(n_2045),
.Y(n_2103)
);

O2A1O1Ixp33_ASAP7_75t_L g2104 ( 
.A1(n_2055),
.A2(n_1963),
.B(n_1955),
.C(n_2042),
.Y(n_2104)
);

AND2x4_ASAP7_75t_SL g2105 ( 
.A(n_2087),
.B(n_2019),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_2085),
.B(n_1995),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2071),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_2073),
.Y(n_2108)
);

OR2x2_ASAP7_75t_L g2109 ( 
.A(n_2089),
.B(n_2001),
.Y(n_2109)
);

OR2x6_ASAP7_75t_L g2110 ( 
.A(n_2075),
.B(n_2019),
.Y(n_2110)
);

AND2x2_ASAP7_75t_L g2111 ( 
.A(n_2092),
.B(n_2064),
.Y(n_2111)
);

HB1xp67_ASAP7_75t_L g2112 ( 
.A(n_2067),
.Y(n_2112)
);

O2A1O1Ixp33_ASAP7_75t_L g2113 ( 
.A1(n_2059),
.A2(n_1913),
.B(n_2036),
.C(n_2031),
.Y(n_2113)
);

CKINVDCx5p33_ASAP7_75t_R g2114 ( 
.A(n_2083),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_2072),
.B(n_2012),
.Y(n_2115)
);

OAI22xp5_ASAP7_75t_L g2116 ( 
.A1(n_2050),
.A2(n_1983),
.B1(n_2032),
.B2(n_2036),
.Y(n_2116)
);

AOI22xp33_ASAP7_75t_L g2117 ( 
.A1(n_2116),
.A2(n_2051),
.B1(n_2048),
.B2(n_2059),
.Y(n_2117)
);

INVx2_ASAP7_75t_L g2118 ( 
.A(n_2095),
.Y(n_2118)
);

AOI22xp33_ASAP7_75t_SL g2119 ( 
.A1(n_2116),
.A2(n_2061),
.B1(n_2062),
.B2(n_2041),
.Y(n_2119)
);

NOR2x1_ASAP7_75t_SL g2120 ( 
.A(n_2110),
.B(n_1986),
.Y(n_2120)
);

AND2x2_ASAP7_75t_L g2121 ( 
.A(n_2101),
.B(n_2072),
.Y(n_2121)
);

AND2x4_ASAP7_75t_L g2122 ( 
.A(n_2110),
.B(n_2078),
.Y(n_2122)
);

INVx1_ASAP7_75t_SL g2123 ( 
.A(n_2114),
.Y(n_2123)
);

AOI22xp33_ASAP7_75t_L g2124 ( 
.A1(n_2103),
.A2(n_2051),
.B1(n_2062),
.B2(n_2052),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2095),
.Y(n_2125)
);

NOR3xp33_ASAP7_75t_SL g2126 ( 
.A(n_2113),
.B(n_2077),
.C(n_2074),
.Y(n_2126)
);

BUFx2_ASAP7_75t_L g2127 ( 
.A(n_2110),
.Y(n_2127)
);

INVx2_ASAP7_75t_L g2128 ( 
.A(n_2095),
.Y(n_2128)
);

INVx3_ASAP7_75t_L g2129 ( 
.A(n_2122),
.Y(n_2129)
);

OA21x2_ASAP7_75t_L g2130 ( 
.A1(n_2127),
.A2(n_2099),
.B(n_2094),
.Y(n_2130)
);

AO21x2_ASAP7_75t_L g2131 ( 
.A1(n_2120),
.A2(n_2100),
.B(n_2063),
.Y(n_2131)
);

BUFx6f_ASAP7_75t_L g2132 ( 
.A(n_2127),
.Y(n_2132)
);

AO21x2_ASAP7_75t_L g2133 ( 
.A1(n_2120),
.A2(n_2063),
.B(n_2012),
.Y(n_2133)
);

INVx2_ASAP7_75t_L g2134 ( 
.A(n_2118),
.Y(n_2134)
);

AO21x2_ASAP7_75t_L g2135 ( 
.A1(n_2118),
.A2(n_2052),
.B(n_2115),
.Y(n_2135)
);

INVx2_ASAP7_75t_L g2136 ( 
.A(n_2125),
.Y(n_2136)
);

INVx2_ASAP7_75t_L g2137 ( 
.A(n_2132),
.Y(n_2137)
);

INVxp33_ASAP7_75t_L g2138 ( 
.A(n_2132),
.Y(n_2138)
);

INVx2_ASAP7_75t_L g2139 ( 
.A(n_2132),
.Y(n_2139)
);

AOI22xp33_ASAP7_75t_L g2140 ( 
.A1(n_2131),
.A2(n_2117),
.B1(n_2119),
.B2(n_2124),
.Y(n_2140)
);

AOI21x1_ASAP7_75t_L g2141 ( 
.A1(n_2134),
.A2(n_2121),
.B(n_2125),
.Y(n_2141)
);

OR2x2_ASAP7_75t_L g2142 ( 
.A(n_2132),
.B(n_2094),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2129),
.B(n_2121),
.Y(n_2143)
);

INVx1_ASAP7_75t_L g2144 ( 
.A(n_2134),
.Y(n_2144)
);

INVx1_ASAP7_75t_L g2145 ( 
.A(n_2134),
.Y(n_2145)
);

AND2x2_ASAP7_75t_L g2146 ( 
.A(n_2129),
.B(n_2132),
.Y(n_2146)
);

OAI22xp5_ASAP7_75t_L g2147 ( 
.A1(n_2140),
.A2(n_2126),
.B1(n_2060),
.B2(n_2093),
.Y(n_2147)
);

INVx4_ASAP7_75t_L g2148 ( 
.A(n_2137),
.Y(n_2148)
);

AND2x2_ASAP7_75t_L g2149 ( 
.A(n_2146),
.B(n_2143),
.Y(n_2149)
);

INVx2_ASAP7_75t_L g2150 ( 
.A(n_2146),
.Y(n_2150)
);

AOI221xp5_ASAP7_75t_L g2151 ( 
.A1(n_2138),
.A2(n_2132),
.B1(n_2131),
.B2(n_2135),
.C(n_2104),
.Y(n_2151)
);

INVx1_ASAP7_75t_L g2152 ( 
.A(n_2145),
.Y(n_2152)
);

BUFx3_ASAP7_75t_L g2153 ( 
.A(n_2137),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2141),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2144),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_2139),
.B(n_2129),
.Y(n_2156)
);

AOI22xp33_ASAP7_75t_L g2157 ( 
.A1(n_2139),
.A2(n_2131),
.B1(n_2132),
.B2(n_2133),
.Y(n_2157)
);

AND2x4_ASAP7_75t_L g2158 ( 
.A(n_2143),
.B(n_2129),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2158),
.Y(n_2159)
);

AND2x2_ASAP7_75t_L g2160 ( 
.A(n_2149),
.B(n_2132),
.Y(n_2160)
);

INVx1_ASAP7_75t_L g2161 ( 
.A(n_2152),
.Y(n_2161)
);

INVx1_ASAP7_75t_L g2162 ( 
.A(n_2152),
.Y(n_2162)
);

AND2x2_ASAP7_75t_L g2163 ( 
.A(n_2149),
.B(n_2129),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2158),
.B(n_2150),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2158),
.B(n_2142),
.Y(n_2165)
);

INVx2_ASAP7_75t_L g2166 ( 
.A(n_2158),
.Y(n_2166)
);

INVx3_ASAP7_75t_L g2167 ( 
.A(n_2156),
.Y(n_2167)
);

AND2x2_ASAP7_75t_L g2168 ( 
.A(n_2160),
.B(n_2150),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_2160),
.B(n_2153),
.Y(n_2169)
);

NOR2xp33_ASAP7_75t_SL g2170 ( 
.A(n_2164),
.B(n_2159),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_2167),
.Y(n_2171)
);

OR2x2_ASAP7_75t_L g2172 ( 
.A(n_2171),
.B(n_2168),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_L g2173 ( 
.A(n_2169),
.B(n_2170),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_2170),
.Y(n_2174)
);

INVxp67_ASAP7_75t_L g2175 ( 
.A(n_2170),
.Y(n_2175)
);

OAI32xp33_ASAP7_75t_L g2176 ( 
.A1(n_2175),
.A2(n_2157),
.A3(n_2154),
.B1(n_2166),
.B2(n_2159),
.Y(n_2176)
);

INVx1_ASAP7_75t_L g2177 ( 
.A(n_2172),
.Y(n_2177)
);

AOI211xp5_ASAP7_75t_L g2178 ( 
.A1(n_2174),
.A2(n_2151),
.B(n_2147),
.C(n_2164),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_2173),
.B(n_2166),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_L g2180 ( 
.A(n_2175),
.B(n_2165),
.Y(n_2180)
);

NAND2xp5_ASAP7_75t_L g2181 ( 
.A(n_2175),
.B(n_2165),
.Y(n_2181)
);

NOR2xp33_ASAP7_75t_L g2182 ( 
.A(n_2180),
.B(n_2123),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_2177),
.B(n_2167),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_2181),
.B(n_2167),
.Y(n_2184)
);

NOR2xp33_ASAP7_75t_L g2185 ( 
.A(n_2179),
.B(n_2090),
.Y(n_2185)
);

INVx1_ASAP7_75t_SL g2186 ( 
.A(n_2176),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_2178),
.A2(n_2163),
.B1(n_2131),
.B2(n_2154),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_2180),
.B(n_2049),
.Y(n_2188)
);

INVx2_ASAP7_75t_L g2189 ( 
.A(n_2180),
.Y(n_2189)
);

INVx3_ASAP7_75t_L g2190 ( 
.A(n_2177),
.Y(n_2190)
);

AND2x2_ASAP7_75t_L g2191 ( 
.A(n_2177),
.B(n_2163),
.Y(n_2191)
);

INVx1_ASAP7_75t_SL g2192 ( 
.A(n_2191),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2184),
.Y(n_2193)
);

OAI322xp33_ASAP7_75t_L g2194 ( 
.A1(n_2186),
.A2(n_2161),
.A3(n_2162),
.B1(n_2148),
.B2(n_2154),
.C1(n_2155),
.C2(n_2142),
.Y(n_2194)
);

OAI21xp5_ASAP7_75t_SL g2195 ( 
.A1(n_2187),
.A2(n_2156),
.B(n_2155),
.Y(n_2195)
);

OAI22xp5_ASAP7_75t_L g2196 ( 
.A1(n_2189),
.A2(n_2153),
.B1(n_2148),
.B2(n_2156),
.Y(n_2196)
);

NOR2xp33_ASAP7_75t_L g2197 ( 
.A(n_2190),
.B(n_2148),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2183),
.Y(n_2198)
);

NOR2xp33_ASAP7_75t_L g2199 ( 
.A(n_2190),
.B(n_2053),
.Y(n_2199)
);

OAI321xp33_ASAP7_75t_L g2200 ( 
.A1(n_2182),
.A2(n_2145),
.A3(n_2144),
.B1(n_2141),
.B2(n_2061),
.C(n_2110),
.Y(n_2200)
);

NOR2xp33_ASAP7_75t_L g2201 ( 
.A(n_2188),
.B(n_2029),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2185),
.Y(n_2202)
);

OAI22xp5_ASAP7_75t_L g2203 ( 
.A1(n_2186),
.A2(n_2112),
.B1(n_2130),
.B2(n_2046),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_2191),
.Y(n_2204)
);

AOI22xp5_ASAP7_75t_L g2205 ( 
.A1(n_2199),
.A2(n_2131),
.B1(n_2046),
.B2(n_2065),
.Y(n_2205)
);

OAI22xp33_ASAP7_75t_L g2206 ( 
.A1(n_2192),
.A2(n_2130),
.B1(n_2046),
.B2(n_2065),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_2204),
.B(n_2130),
.Y(n_2207)
);

NOR2xp33_ASAP7_75t_SL g2208 ( 
.A(n_2194),
.B(n_1817),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_2193),
.A2(n_2133),
.B1(n_2135),
.B2(n_2065),
.Y(n_2209)
);

OR2x2_ASAP7_75t_L g2210 ( 
.A(n_2203),
.B(n_2130),
.Y(n_2210)
);

INVx1_ASAP7_75t_L g2211 ( 
.A(n_2197),
.Y(n_2211)
);

AOI221xp5_ASAP7_75t_SL g2212 ( 
.A1(n_2196),
.A2(n_2136),
.B1(n_2134),
.B2(n_1941),
.C(n_2011),
.Y(n_2212)
);

AND2x2_ASAP7_75t_L g2213 ( 
.A(n_2198),
.B(n_2201),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2195),
.Y(n_2214)
);

NOR2x1_ASAP7_75t_R g2215 ( 
.A(n_2202),
.B(n_2041),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_2200),
.Y(n_2216)
);

AOI221xp5_ASAP7_75t_L g2217 ( 
.A1(n_2194),
.A2(n_2135),
.B1(n_2133),
.B2(n_2136),
.C(n_2056),
.Y(n_2217)
);

A2O1A1Ixp33_ASAP7_75t_L g2218 ( 
.A1(n_2197),
.A2(n_2136),
.B(n_2105),
.C(n_2011),
.Y(n_2218)
);

INVx1_ASAP7_75t_L g2219 ( 
.A(n_2204),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2219),
.Y(n_2220)
);

INVx2_ASAP7_75t_SL g2221 ( 
.A(n_2207),
.Y(n_2221)
);

INVx2_ASAP7_75t_L g2222 ( 
.A(n_2210),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2214),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2208),
.B(n_2135),
.Y(n_2224)
);

NOR2x1_ASAP7_75t_L g2225 ( 
.A(n_2211),
.B(n_2133),
.Y(n_2225)
);

INVx1_ASAP7_75t_L g2226 ( 
.A(n_2213),
.Y(n_2226)
);

NOR2xp33_ASAP7_75t_L g2227 ( 
.A(n_2215),
.B(n_2130),
.Y(n_2227)
);

AND2x2_ASAP7_75t_L g2228 ( 
.A(n_2216),
.B(n_2130),
.Y(n_2228)
);

NAND2xp5_ASAP7_75t_L g2229 ( 
.A(n_2212),
.B(n_2135),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2206),
.B(n_2218),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_2217),
.B(n_2136),
.Y(n_2231)
);

INVx1_ASAP7_75t_L g2232 ( 
.A(n_2205),
.Y(n_2232)
);

AOI22xp33_ASAP7_75t_L g2233 ( 
.A1(n_2209),
.A2(n_2133),
.B1(n_2101),
.B2(n_2105),
.Y(n_2233)
);

AOI21xp33_ASAP7_75t_L g2234 ( 
.A1(n_2223),
.A2(n_1966),
.B(n_1959),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_2222),
.Y(n_2235)
);

INVx2_ASAP7_75t_SL g2236 ( 
.A(n_2220),
.Y(n_2236)
);

AOI22xp5_ASAP7_75t_L g2237 ( 
.A1(n_2228),
.A2(n_2122),
.B1(n_1835),
.B2(n_2101),
.Y(n_2237)
);

NOR3x1_ASAP7_75t_L g2238 ( 
.A(n_2230),
.B(n_1968),
.C(n_1960),
.Y(n_2238)
);

NAND2xp5_ASAP7_75t_L g2239 ( 
.A(n_2226),
.B(n_2033),
.Y(n_2239)
);

NOR2xp33_ASAP7_75t_SL g2240 ( 
.A(n_2221),
.B(n_1754),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_2231),
.Y(n_2241)
);

NAND2xp5_ASAP7_75t_L g2242 ( 
.A(n_2232),
.B(n_2128),
.Y(n_2242)
);

INVx1_ASAP7_75t_L g2243 ( 
.A(n_2231),
.Y(n_2243)
);

NAND3xp33_ASAP7_75t_L g2244 ( 
.A(n_2227),
.B(n_1782),
.C(n_2091),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2229),
.Y(n_2245)
);

NAND3xp33_ASAP7_75t_SL g2246 ( 
.A(n_2224),
.B(n_2060),
.C(n_2093),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_L g2247 ( 
.A(n_2233),
.B(n_1782),
.C(n_2091),
.Y(n_2247)
);

NAND2xp5_ASAP7_75t_L g2248 ( 
.A(n_2225),
.B(n_2128),
.Y(n_2248)
);

NAND2xp5_ASAP7_75t_L g2249 ( 
.A(n_2228),
.B(n_2016),
.Y(n_2249)
);

OR2x2_ASAP7_75t_L g2250 ( 
.A(n_2223),
.B(n_2101),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2221),
.Y(n_2251)
);

AOI21xp5_ASAP7_75t_L g2252 ( 
.A1(n_2221),
.A2(n_2009),
.B(n_1995),
.Y(n_2252)
);

OAI211xp5_ASAP7_75t_L g2253 ( 
.A1(n_2223),
.A2(n_1782),
.B(n_2082),
.C(n_199),
.Y(n_2253)
);

NOR3xp33_ASAP7_75t_L g2254 ( 
.A(n_2226),
.B(n_1997),
.C(n_1991),
.Y(n_2254)
);

NOR2xp33_ASAP7_75t_L g2255 ( 
.A(n_2223),
.B(n_196),
.Y(n_2255)
);

AOI211x1_ASAP7_75t_L g2256 ( 
.A1(n_2247),
.A2(n_1939),
.B(n_2005),
.C(n_1996),
.Y(n_2256)
);

NAND3x1_ASAP7_75t_L g2257 ( 
.A(n_2255),
.B(n_2235),
.C(n_2241),
.Y(n_2257)
);

NAND2xp5_ASAP7_75t_L g2258 ( 
.A(n_2251),
.B(n_2018),
.Y(n_2258)
);

NAND4xp25_ASAP7_75t_L g2259 ( 
.A(n_2244),
.B(n_2122),
.C(n_2017),
.D(n_1725),
.Y(n_2259)
);

NOR3xp33_ASAP7_75t_L g2260 ( 
.A(n_2236),
.B(n_2243),
.C(n_2245),
.Y(n_2260)
);

OAI22xp5_ASAP7_75t_L g2261 ( 
.A1(n_2237),
.A2(n_2122),
.B1(n_2105),
.B2(n_2097),
.Y(n_2261)
);

NAND3xp33_ASAP7_75t_L g2262 ( 
.A(n_2240),
.B(n_197),
.C(n_199),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2254),
.B(n_2024),
.Y(n_2263)
);

NAND4xp25_ASAP7_75t_L g2264 ( 
.A(n_2250),
.B(n_202),
.C(n_200),
.D(n_201),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2249),
.B(n_201),
.Y(n_2265)
);

NAND2xp5_ASAP7_75t_L g2266 ( 
.A(n_2239),
.B(n_202),
.Y(n_2266)
);

NOR2xp33_ASAP7_75t_L g2267 ( 
.A(n_2253),
.B(n_203),
.Y(n_2267)
);

AOI211xp5_ASAP7_75t_L g2268 ( 
.A1(n_2242),
.A2(n_2246),
.B(n_2234),
.C(n_2248),
.Y(n_2268)
);

NAND2xp33_ASAP7_75t_SL g2269 ( 
.A(n_2238),
.B(n_2028),
.Y(n_2269)
);

INVxp67_ASAP7_75t_L g2270 ( 
.A(n_2252),
.Y(n_2270)
);

AOI21xp5_ASAP7_75t_L g2271 ( 
.A1(n_2251),
.A2(n_1996),
.B(n_2032),
.Y(n_2271)
);

INVx1_ASAP7_75t_SL g2272 ( 
.A(n_2250),
.Y(n_2272)
);

NAND4xp25_ASAP7_75t_L g2273 ( 
.A(n_2244),
.B(n_206),
.C(n_204),
.D(n_205),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2251),
.Y(n_2274)
);

AOI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2251),
.A2(n_1950),
.B(n_1907),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2247),
.A2(n_2099),
.B1(n_2109),
.B2(n_2110),
.Y(n_2276)
);

OAI321xp33_ASAP7_75t_L g2277 ( 
.A1(n_2244),
.A2(n_2109),
.A3(n_2003),
.B1(n_2021),
.B2(n_2115),
.C(n_2030),
.Y(n_2277)
);

INVx1_ASAP7_75t_L g2278 ( 
.A(n_2251),
.Y(n_2278)
);

NAND2xp5_ASAP7_75t_L g2279 ( 
.A(n_2255),
.B(n_204),
.Y(n_2279)
);

INVx1_ASAP7_75t_L g2280 ( 
.A(n_2251),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2251),
.Y(n_2281)
);

NOR2xp33_ASAP7_75t_SL g2282 ( 
.A(n_2251),
.B(n_2068),
.Y(n_2282)
);

AOI22xp33_ASAP7_75t_L g2283 ( 
.A1(n_2251),
.A2(n_2076),
.B1(n_2068),
.B2(n_2057),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2255),
.B(n_205),
.Y(n_2284)
);

NOR3xp33_ASAP7_75t_L g2285 ( 
.A(n_2251),
.B(n_1975),
.C(n_207),
.Y(n_2285)
);

NOR3xp33_ASAP7_75t_L g2286 ( 
.A(n_2251),
.B(n_207),
.C(n_208),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2251),
.Y(n_2287)
);

INVx1_ASAP7_75t_L g2288 ( 
.A(n_2251),
.Y(n_2288)
);

NAND3xp33_ASAP7_75t_L g2289 ( 
.A(n_2251),
.B(n_209),
.C(n_210),
.Y(n_2289)
);

INVx1_ASAP7_75t_L g2290 ( 
.A(n_2251),
.Y(n_2290)
);

NAND5xp2_ASAP7_75t_L g2291 ( 
.A(n_2235),
.B(n_1887),
.C(n_211),
.D(n_209),
.E(n_210),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2251),
.Y(n_2292)
);

O2A1O1Ixp33_ASAP7_75t_L g2293 ( 
.A1(n_2274),
.A2(n_2278),
.B(n_2281),
.C(n_2280),
.Y(n_2293)
);

NOR2x1_ASAP7_75t_L g2294 ( 
.A(n_2289),
.B(n_2264),
.Y(n_2294)
);

AOI211xp5_ASAP7_75t_L g2295 ( 
.A1(n_2273),
.A2(n_214),
.B(n_212),
.C(n_213),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_2282),
.B(n_212),
.Y(n_2296)
);

NAND4xp25_ASAP7_75t_L g2297 ( 
.A(n_2287),
.B(n_216),
.C(n_213),
.D(n_215),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2288),
.B(n_215),
.Y(n_2298)
);

NAND4xp25_ASAP7_75t_L g2299 ( 
.A(n_2290),
.B(n_219),
.C(n_217),
.D(n_218),
.Y(n_2299)
);

NOR2xp33_ASAP7_75t_L g2300 ( 
.A(n_2292),
.B(n_218),
.Y(n_2300)
);

AND4x1_ASAP7_75t_L g2301 ( 
.A(n_2286),
.B(n_221),
.C(n_219),
.D(n_220),
.Y(n_2301)
);

OAI22xp33_ASAP7_75t_L g2302 ( 
.A1(n_2272),
.A2(n_2075),
.B1(n_2088),
.B2(n_2086),
.Y(n_2302)
);

NOR2xp33_ASAP7_75t_L g2303 ( 
.A(n_2279),
.B(n_220),
.Y(n_2303)
);

NOR2xp33_ASAP7_75t_L g2304 ( 
.A(n_2284),
.B(n_222),
.Y(n_2304)
);

NOR2xp33_ASAP7_75t_L g2305 ( 
.A(n_2265),
.B(n_222),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_SL g2306 ( 
.A(n_2262),
.B(n_2076),
.Y(n_2306)
);

NOR3xp33_ASAP7_75t_L g2307 ( 
.A(n_2266),
.B(n_223),
.C(n_224),
.Y(n_2307)
);

NOR3xp33_ASAP7_75t_L g2308 ( 
.A(n_2267),
.B(n_224),
.C(n_225),
.Y(n_2308)
);

OAI21xp33_ASAP7_75t_L g2309 ( 
.A1(n_2259),
.A2(n_2102),
.B(n_2020),
.Y(n_2309)
);

NOR2xp67_ASAP7_75t_L g2310 ( 
.A(n_2270),
.B(n_225),
.Y(n_2310)
);

NOR3xp33_ASAP7_75t_L g2311 ( 
.A(n_2260),
.B(n_226),
.C(n_227),
.Y(n_2311)
);

NOR2x1_ASAP7_75t_L g2312 ( 
.A(n_2291),
.B(n_226),
.Y(n_2312)
);

NAND2xp5_ASAP7_75t_SL g2313 ( 
.A(n_2283),
.B(n_2040),
.Y(n_2313)
);

NAND4xp25_ASAP7_75t_SL g2314 ( 
.A(n_2268),
.B(n_2106),
.C(n_2102),
.D(n_2096),
.Y(n_2314)
);

NAND2xp5_ASAP7_75t_L g2315 ( 
.A(n_2257),
.B(n_227),
.Y(n_2315)
);

AOI21xp5_ASAP7_75t_L g2316 ( 
.A1(n_2258),
.A2(n_228),
.B(n_229),
.Y(n_2316)
);

O2A1O1Ixp33_ASAP7_75t_L g2317 ( 
.A1(n_2263),
.A2(n_232),
.B(n_229),
.C(n_231),
.Y(n_2317)
);

AOI21xp5_ASAP7_75t_L g2318 ( 
.A1(n_2269),
.A2(n_2271),
.B(n_2261),
.Y(n_2318)
);

NOR4xp25_ASAP7_75t_L g2319 ( 
.A(n_2277),
.B(n_234),
.C(n_231),
.D(n_233),
.Y(n_2319)
);

INVxp67_ASAP7_75t_SL g2320 ( 
.A(n_2285),
.Y(n_2320)
);

NOR3xp33_ASAP7_75t_L g2321 ( 
.A(n_2275),
.B(n_233),
.C(n_234),
.Y(n_2321)
);

NAND4xp25_ASAP7_75t_L g2322 ( 
.A(n_2256),
.B(n_237),
.C(n_235),
.D(n_236),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2276),
.B(n_236),
.Y(n_2323)
);

NAND4xp25_ASAP7_75t_L g2324 ( 
.A(n_2282),
.B(n_239),
.C(n_237),
.D(n_238),
.Y(n_2324)
);

OAI21xp5_ASAP7_75t_SL g2325 ( 
.A1(n_2292),
.A2(n_2040),
.B(n_238),
.Y(n_2325)
);

NAND4xp25_ASAP7_75t_L g2326 ( 
.A(n_2282),
.B(n_242),
.C(n_240),
.D(n_241),
.Y(n_2326)
);

NAND4xp75_ASAP7_75t_L g2327 ( 
.A(n_2274),
.B(n_242),
.C(n_240),
.D(n_241),
.Y(n_2327)
);

NAND2xp5_ASAP7_75t_L g2328 ( 
.A(n_2274),
.B(n_243),
.Y(n_2328)
);

NOR3xp33_ASAP7_75t_L g2329 ( 
.A(n_2292),
.B(n_244),
.C(n_245),
.Y(n_2329)
);

AOI22xp5_ASAP7_75t_L g2330 ( 
.A1(n_2306),
.A2(n_1748),
.B1(n_2088),
.B2(n_2086),
.Y(n_2330)
);

OAI21xp33_ASAP7_75t_L g2331 ( 
.A1(n_2312),
.A2(n_2078),
.B(n_2037),
.Y(n_2331)
);

NAND4xp25_ASAP7_75t_L g2332 ( 
.A(n_2293),
.B(n_246),
.C(n_244),
.D(n_245),
.Y(n_2332)
);

NOR2xp67_ASAP7_75t_L g2333 ( 
.A(n_2324),
.B(n_246),
.Y(n_2333)
);

NAND2xp5_ASAP7_75t_SL g2334 ( 
.A(n_2319),
.B(n_2030),
.Y(n_2334)
);

AND3x2_ASAP7_75t_L g2335 ( 
.A(n_2329),
.B(n_247),
.C(n_248),
.Y(n_2335)
);

NOR2xp33_ASAP7_75t_L g2336 ( 
.A(n_2301),
.B(n_248),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_SL g2337 ( 
.A(n_2310),
.B(n_2030),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2300),
.B(n_249),
.Y(n_2338)
);

NOR2x1_ASAP7_75t_L g2339 ( 
.A(n_2327),
.B(n_249),
.Y(n_2339)
);

NAND3xp33_ASAP7_75t_SL g2340 ( 
.A(n_2311),
.B(n_2315),
.C(n_2295),
.Y(n_2340)
);

NAND4xp25_ASAP7_75t_L g2341 ( 
.A(n_2294),
.B(n_252),
.C(n_250),
.D(n_251),
.Y(n_2341)
);

AND2x2_ASAP7_75t_L g2342 ( 
.A(n_2308),
.B(n_2111),
.Y(n_2342)
);

NOR3xp33_ASAP7_75t_L g2343 ( 
.A(n_2303),
.B(n_2304),
.C(n_2305),
.Y(n_2343)
);

AOI22xp5_ASAP7_75t_L g2344 ( 
.A1(n_2307),
.A2(n_1748),
.B1(n_2088),
.B2(n_2086),
.Y(n_2344)
);

NAND2xp5_ASAP7_75t_L g2345 ( 
.A(n_2296),
.B(n_250),
.Y(n_2345)
);

NOR2xp33_ASAP7_75t_L g2346 ( 
.A(n_2297),
.B(n_253),
.Y(n_2346)
);

OAI21xp33_ASAP7_75t_L g2347 ( 
.A1(n_2309),
.A2(n_2037),
.B(n_2034),
.Y(n_2347)
);

AOI22xp5_ASAP7_75t_L g2348 ( 
.A1(n_2313),
.A2(n_2066),
.B1(n_2058),
.B2(n_2026),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2298),
.Y(n_2349)
);

OAI211xp5_ASAP7_75t_L g2350 ( 
.A1(n_2325),
.A2(n_257),
.B(n_255),
.C(n_256),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2328),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2323),
.Y(n_2352)
);

NAND3xp33_ASAP7_75t_L g2353 ( 
.A(n_2317),
.B(n_2316),
.C(n_2326),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2299),
.Y(n_2354)
);

NOR3xp33_ASAP7_75t_L g2355 ( 
.A(n_2320),
.B(n_255),
.C(n_256),
.Y(n_2355)
);

NOR4xp25_ASAP7_75t_L g2356 ( 
.A(n_2322),
.B(n_260),
.C(n_258),
.D(n_259),
.Y(n_2356)
);

NAND5xp2_ASAP7_75t_L g2357 ( 
.A(n_2318),
.B(n_264),
.C(n_259),
.D(n_261),
.E(n_265),
.Y(n_2357)
);

NOR2xp33_ASAP7_75t_L g2358 ( 
.A(n_2302),
.B(n_261),
.Y(n_2358)
);

O2A1O1Ixp5_ASAP7_75t_L g2359 ( 
.A1(n_2321),
.A2(n_267),
.B(n_265),
.C(n_266),
.Y(n_2359)
);

HB1xp67_ASAP7_75t_L g2360 ( 
.A(n_2314),
.Y(n_2360)
);

NAND3xp33_ASAP7_75t_L g2361 ( 
.A(n_2311),
.B(n_266),
.C(n_268),
.Y(n_2361)
);

NOR3xp33_ASAP7_75t_SL g2362 ( 
.A(n_2315),
.B(n_268),
.C(n_270),
.Y(n_2362)
);

AOI21xp5_ASAP7_75t_L g2363 ( 
.A1(n_2293),
.A2(n_270),
.B(n_271),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2315),
.Y(n_2364)
);

NAND3xp33_ASAP7_75t_SL g2365 ( 
.A(n_2293),
.B(n_272),
.C(n_273),
.Y(n_2365)
);

A2O1A1Ixp33_ASAP7_75t_L g2366 ( 
.A1(n_2293),
.A2(n_276),
.B(n_274),
.C(n_275),
.Y(n_2366)
);

NAND3xp33_ASAP7_75t_L g2367 ( 
.A(n_2311),
.B(n_274),
.C(n_275),
.Y(n_2367)
);

AOI211xp5_ASAP7_75t_L g2368 ( 
.A1(n_2293),
.A2(n_278),
.B(n_276),
.C(n_277),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_2301),
.B(n_277),
.Y(n_2369)
);

NAND4xp25_ASAP7_75t_SL g2370 ( 
.A(n_2293),
.B(n_280),
.C(n_278),
.D(n_279),
.Y(n_2370)
);

NAND3xp33_ASAP7_75t_SL g2371 ( 
.A(n_2293),
.B(n_279),
.C(n_280),
.Y(n_2371)
);

NAND3xp33_ASAP7_75t_L g2372 ( 
.A(n_2311),
.B(n_281),
.C(n_283),
.Y(n_2372)
);

NAND5xp2_ASAP7_75t_L g2373 ( 
.A(n_2293),
.B(n_281),
.C(n_283),
.D(n_284),
.E(n_285),
.Y(n_2373)
);

NAND2xp5_ASAP7_75t_SL g2374 ( 
.A(n_2319),
.B(n_2058),
.Y(n_2374)
);

O2A1O1Ixp33_ASAP7_75t_L g2375 ( 
.A1(n_2315),
.A2(n_287),
.B(n_284),
.C(n_286),
.Y(n_2375)
);

NAND2xp5_ASAP7_75t_L g2376 ( 
.A(n_2310),
.B(n_286),
.Y(n_2376)
);

NAND2xp5_ASAP7_75t_L g2377 ( 
.A(n_2310),
.B(n_288),
.Y(n_2377)
);

NOR4xp25_ASAP7_75t_L g2378 ( 
.A(n_2293),
.B(n_290),
.C(n_288),
.D(n_289),
.Y(n_2378)
);

NOR3x1_ASAP7_75t_L g2379 ( 
.A(n_2325),
.B(n_289),
.C(n_290),
.Y(n_2379)
);

AOI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2293),
.A2(n_291),
.B(n_292),
.Y(n_2380)
);

NAND3x1_ASAP7_75t_L g2381 ( 
.A(n_2315),
.B(n_293),
.C(n_294),
.Y(n_2381)
);

NOR3xp33_ASAP7_75t_L g2382 ( 
.A(n_2293),
.B(n_293),
.C(n_294),
.Y(n_2382)
);

NAND5xp2_ASAP7_75t_L g2383 ( 
.A(n_2293),
.B(n_295),
.C(n_296),
.D(n_297),
.E(n_298),
.Y(n_2383)
);

NOR2xp33_ASAP7_75t_L g2384 ( 
.A(n_2301),
.B(n_296),
.Y(n_2384)
);

NAND2xp5_ASAP7_75t_L g2385 ( 
.A(n_2310),
.B(n_298),
.Y(n_2385)
);

NOR2x1_ASAP7_75t_L g2386 ( 
.A(n_2327),
.B(n_299),
.Y(n_2386)
);

NAND3xp33_ASAP7_75t_L g2387 ( 
.A(n_2311),
.B(n_299),
.C(n_300),
.Y(n_2387)
);

HB1xp67_ASAP7_75t_L g2388 ( 
.A(n_2370),
.Y(n_2388)
);

OAI211xp5_ASAP7_75t_L g2389 ( 
.A1(n_2378),
.A2(n_302),
.B(n_300),
.C(n_301),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2335),
.B(n_302),
.Y(n_2390)
);

AOI211xp5_ASAP7_75t_L g2391 ( 
.A1(n_2350),
.A2(n_305),
.B(n_303),
.C(n_304),
.Y(n_2391)
);

HB1xp67_ASAP7_75t_L g2392 ( 
.A(n_2339),
.Y(n_2392)
);

AOI22xp5_ASAP7_75t_SL g2393 ( 
.A1(n_2383),
.A2(n_2026),
.B1(n_2066),
.B2(n_2058),
.Y(n_2393)
);

OR2x2_ASAP7_75t_L g2394 ( 
.A(n_2357),
.B(n_304),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_R g2395 ( 
.A(n_2365),
.B(n_305),
.Y(n_2395)
);

NAND2xp5_ASAP7_75t_L g2396 ( 
.A(n_2356),
.B(n_306),
.Y(n_2396)
);

NAND2xp33_ASAP7_75t_L g2397 ( 
.A(n_2381),
.B(n_2066),
.Y(n_2397)
);

CKINVDCx16_ASAP7_75t_R g2398 ( 
.A(n_2371),
.Y(n_2398)
);

XNOR2xp5_ASAP7_75t_L g2399 ( 
.A(n_2332),
.B(n_306),
.Y(n_2399)
);

OAI221xp5_ASAP7_75t_L g2400 ( 
.A1(n_2382),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.C(n_310),
.Y(n_2400)
);

INVx1_ASAP7_75t_L g2401 ( 
.A(n_2376),
.Y(n_2401)
);

OAI221xp5_ASAP7_75t_L g2402 ( 
.A1(n_2368),
.A2(n_307),
.B1(n_308),
.B2(n_309),
.C(n_311),
.Y(n_2402)
);

A2O1A1Ixp33_ASAP7_75t_L g2403 ( 
.A1(n_2375),
.A2(n_313),
.B(n_311),
.C(n_312),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2362),
.B(n_2111),
.Y(n_2404)
);

HB1xp67_ASAP7_75t_L g2405 ( 
.A(n_2386),
.Y(n_2405)
);

BUFx6f_ASAP7_75t_L g2406 ( 
.A(n_2364),
.Y(n_2406)
);

AOI21xp5_ASAP7_75t_L g2407 ( 
.A1(n_2377),
.A2(n_312),
.B(n_314),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_2385),
.Y(n_2408)
);

NOR2xp33_ASAP7_75t_R g2409 ( 
.A(n_2340),
.B(n_315),
.Y(n_2409)
);

O2A1O1Ixp33_ASAP7_75t_L g2410 ( 
.A1(n_2366),
.A2(n_318),
.B(n_316),
.C(n_317),
.Y(n_2410)
);

INVx1_ASAP7_75t_SL g2411 ( 
.A(n_2338),
.Y(n_2411)
);

INVx2_ASAP7_75t_L g2412 ( 
.A(n_2379),
.Y(n_2412)
);

AND2x4_ASAP7_75t_L g2413 ( 
.A(n_2337),
.B(n_316),
.Y(n_2413)
);

AOI22xp5_ASAP7_75t_L g2414 ( 
.A1(n_2333),
.A2(n_2034),
.B1(n_2108),
.B2(n_2107),
.Y(n_2414)
);

NAND2x1_ASAP7_75t_L g2415 ( 
.A(n_2336),
.B(n_317),
.Y(n_2415)
);

AOI22xp5_ASAP7_75t_L g2416 ( 
.A1(n_2346),
.A2(n_2108),
.B1(n_2107),
.B2(n_2098),
.Y(n_2416)
);

HB1xp67_ASAP7_75t_L g2417 ( 
.A(n_2369),
.Y(n_2417)
);

INVx1_ASAP7_75t_L g2418 ( 
.A(n_2384),
.Y(n_2418)
);

NOR2x1_ASAP7_75t_L g2419 ( 
.A(n_2383),
.B(n_318),
.Y(n_2419)
);

INVx2_ASAP7_75t_L g2420 ( 
.A(n_2359),
.Y(n_2420)
);

A2O1A1Ixp33_ASAP7_75t_L g2421 ( 
.A1(n_2363),
.A2(n_321),
.B(n_319),
.C(n_320),
.Y(n_2421)
);

AOI22xp5_ASAP7_75t_L g2422 ( 
.A1(n_2374),
.A2(n_2098),
.B1(n_1986),
.B2(n_1928),
.Y(n_2422)
);

NOR2xp33_ASAP7_75t_R g2423 ( 
.A(n_2354),
.B(n_319),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2373),
.B(n_320),
.Y(n_2424)
);

XOR2xp5_ASAP7_75t_L g2425 ( 
.A(n_2341),
.B(n_321),
.Y(n_2425)
);

NAND3xp33_ASAP7_75t_L g2426 ( 
.A(n_2380),
.B(n_322),
.C(n_324),
.Y(n_2426)
);

NAND2xp5_ASAP7_75t_L g2427 ( 
.A(n_2355),
.B(n_322),
.Y(n_2427)
);

OAI21xp5_ASAP7_75t_L g2428 ( 
.A1(n_2387),
.A2(n_1944),
.B(n_1930),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2342),
.B(n_2098),
.Y(n_2429)
);

O2A1O1Ixp33_ASAP7_75t_L g2430 ( 
.A1(n_2360),
.A2(n_327),
.B(n_324),
.C(n_325),
.Y(n_2430)
);

AOI221xp5_ASAP7_75t_L g2431 ( 
.A1(n_2358),
.A2(n_2334),
.B1(n_2367),
.B2(n_2361),
.C(n_2372),
.Y(n_2431)
);

OR2x2_ASAP7_75t_L g2432 ( 
.A(n_2345),
.B(n_325),
.Y(n_2432)
);

AOI21xp5_ASAP7_75t_L g2433 ( 
.A1(n_2353),
.A2(n_2351),
.B(n_2349),
.Y(n_2433)
);

OAI21xp33_ASAP7_75t_L g2434 ( 
.A1(n_2331),
.A2(n_2008),
.B(n_1924),
.Y(n_2434)
);

NAND4xp75_ASAP7_75t_L g2435 ( 
.A(n_2352),
.B(n_329),
.C(n_327),
.D(n_328),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_R g2436 ( 
.A(n_2343),
.B(n_329),
.Y(n_2436)
);

INVx1_ASAP7_75t_L g2437 ( 
.A(n_2344),
.Y(n_2437)
);

INVx1_ASAP7_75t_L g2438 ( 
.A(n_2348),
.Y(n_2438)
);

INVx1_ASAP7_75t_L g2439 ( 
.A(n_2347),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2330),
.B(n_330),
.Y(n_2440)
);

NOR2xp33_ASAP7_75t_R g2441 ( 
.A(n_2365),
.B(n_330),
.Y(n_2441)
);

OAI322xp33_ASAP7_75t_L g2442 ( 
.A1(n_2374),
.A2(n_331),
.A3(n_332),
.B1(n_334),
.B2(n_335),
.C1(n_336),
.C2(n_337),
.Y(n_2442)
);

INVx1_ASAP7_75t_SL g2443 ( 
.A(n_2335),
.Y(n_2443)
);

NOR2x1_ASAP7_75t_L g2444 ( 
.A(n_2383),
.B(n_332),
.Y(n_2444)
);

NOR2x1p5_ASAP7_75t_L g2445 ( 
.A(n_2415),
.B(n_336),
.Y(n_2445)
);

NOR3xp33_ASAP7_75t_SL g2446 ( 
.A(n_2398),
.B(n_337),
.C(n_338),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_SL g2447 ( 
.A(n_2419),
.B(n_339),
.Y(n_2447)
);

OR2x2_ASAP7_75t_L g2448 ( 
.A(n_2394),
.B(n_339),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2444),
.Y(n_2449)
);

NAND4xp75_ASAP7_75t_L g2450 ( 
.A(n_2433),
.B(n_340),
.C(n_341),
.D(n_342),
.Y(n_2450)
);

INVx1_ASAP7_75t_L g2451 ( 
.A(n_2390),
.Y(n_2451)
);

INVx1_ASAP7_75t_L g2452 ( 
.A(n_2396),
.Y(n_2452)
);

INVx3_ASAP7_75t_L g2453 ( 
.A(n_2413),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2393),
.B(n_1989),
.Y(n_2454)
);

INVx1_ASAP7_75t_SL g2455 ( 
.A(n_2423),
.Y(n_2455)
);

NAND4xp75_ASAP7_75t_L g2456 ( 
.A(n_2407),
.B(n_340),
.C(n_341),
.D(n_342),
.Y(n_2456)
);

INVx1_ASAP7_75t_L g2457 ( 
.A(n_2399),
.Y(n_2457)
);

NAND4xp75_ASAP7_75t_L g2458 ( 
.A(n_2427),
.B(n_343),
.C(n_344),
.D(n_345),
.Y(n_2458)
);

NAND4xp75_ASAP7_75t_L g2459 ( 
.A(n_2418),
.B(n_343),
.C(n_344),
.D(n_345),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2435),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_2443),
.B(n_346),
.Y(n_2461)
);

OR2x2_ASAP7_75t_L g2462 ( 
.A(n_2426),
.B(n_346),
.Y(n_2462)
);

INVx1_ASAP7_75t_L g2463 ( 
.A(n_2425),
.Y(n_2463)
);

OAI211xp5_ASAP7_75t_SL g2464 ( 
.A1(n_2431),
.A2(n_347),
.B(n_348),
.C(n_349),
.Y(n_2464)
);

AND2x4_ASAP7_75t_L g2465 ( 
.A(n_2413),
.B(n_347),
.Y(n_2465)
);

INVx2_ASAP7_75t_SL g2466 ( 
.A(n_2432),
.Y(n_2466)
);

NOR3xp33_ASAP7_75t_L g2467 ( 
.A(n_2412),
.B(n_348),
.C(n_349),
.Y(n_2467)
);

AND2x4_ASAP7_75t_L g2468 ( 
.A(n_2404),
.B(n_350),
.Y(n_2468)
);

NAND4xp75_ASAP7_75t_L g2469 ( 
.A(n_2438),
.B(n_351),
.C(n_352),
.D(n_353),
.Y(n_2469)
);

INVxp67_ASAP7_75t_L g2470 ( 
.A(n_2424),
.Y(n_2470)
);

NOR2xp67_ASAP7_75t_L g2471 ( 
.A(n_2389),
.B(n_351),
.Y(n_2471)
);

NAND4xp75_ASAP7_75t_L g2472 ( 
.A(n_2401),
.B(n_352),
.C(n_354),
.D(n_355),
.Y(n_2472)
);

NOR2x1_ASAP7_75t_SL g2473 ( 
.A(n_2420),
.B(n_1986),
.Y(n_2473)
);

XNOR2xp5_ASAP7_75t_L g2474 ( 
.A(n_2391),
.B(n_358),
.Y(n_2474)
);

NAND4xp75_ASAP7_75t_L g2475 ( 
.A(n_2408),
.B(n_2437),
.C(n_2440),
.D(n_2439),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2406),
.Y(n_2476)
);

XNOR2xp5_ASAP7_75t_L g2477 ( 
.A(n_2388),
.B(n_358),
.Y(n_2477)
);

AND2x4_ASAP7_75t_L g2478 ( 
.A(n_2392),
.B(n_359),
.Y(n_2478)
);

INVx1_ASAP7_75t_L g2479 ( 
.A(n_2397),
.Y(n_2479)
);

XNOR2xp5_ASAP7_75t_L g2480 ( 
.A(n_2417),
.B(n_360),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_2405),
.Y(n_2481)
);

NOR2x1_ASAP7_75t_L g2482 ( 
.A(n_2442),
.B(n_360),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2430),
.Y(n_2483)
);

NOR2x1p5_ASAP7_75t_L g2484 ( 
.A(n_2406),
.B(n_361),
.Y(n_2484)
);

HB1xp67_ASAP7_75t_L g2485 ( 
.A(n_2436),
.Y(n_2485)
);

INVx1_ASAP7_75t_L g2486 ( 
.A(n_2410),
.Y(n_2486)
);

NOR2xp33_ASAP7_75t_L g2487 ( 
.A(n_2402),
.B(n_361),
.Y(n_2487)
);

INVx1_ASAP7_75t_L g2488 ( 
.A(n_2403),
.Y(n_2488)
);

INVx1_ASAP7_75t_L g2489 ( 
.A(n_2421),
.Y(n_2489)
);

INVx1_ASAP7_75t_L g2490 ( 
.A(n_2406),
.Y(n_2490)
);

NAND4xp75_ASAP7_75t_L g2491 ( 
.A(n_2409),
.B(n_362),
.C(n_363),
.D(n_364),
.Y(n_2491)
);

NAND4xp75_ASAP7_75t_L g2492 ( 
.A(n_2429),
.B(n_362),
.C(n_364),
.D(n_365),
.Y(n_2492)
);

NAND4xp25_ASAP7_75t_L g2493 ( 
.A(n_2461),
.B(n_2471),
.C(n_2487),
.D(n_2448),
.Y(n_2493)
);

NOR2x1_ASAP7_75t_L g2494 ( 
.A(n_2484),
.B(n_2450),
.Y(n_2494)
);

AOI211xp5_ASAP7_75t_L g2495 ( 
.A1(n_2464),
.A2(n_2400),
.B(n_2395),
.C(n_2441),
.Y(n_2495)
);

NAND3xp33_ASAP7_75t_SL g2496 ( 
.A(n_2490),
.B(n_2411),
.C(n_2414),
.Y(n_2496)
);

NAND3xp33_ASAP7_75t_L g2497 ( 
.A(n_2446),
.B(n_2416),
.C(n_2434),
.Y(n_2497)
);

NOR2x1_ASAP7_75t_L g2498 ( 
.A(n_2469),
.B(n_2428),
.Y(n_2498)
);

INVx1_ASAP7_75t_SL g2499 ( 
.A(n_2465),
.Y(n_2499)
);

AOI211xp5_ASAP7_75t_L g2500 ( 
.A1(n_2447),
.A2(n_2422),
.B(n_367),
.C(n_368),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2477),
.Y(n_2501)
);

OAI211xp5_ASAP7_75t_SL g2502 ( 
.A1(n_2481),
.A2(n_365),
.B(n_367),
.C(n_368),
.Y(n_2502)
);

NOR3xp33_ASAP7_75t_SL g2503 ( 
.A(n_2475),
.B(n_369),
.C(n_370),
.Y(n_2503)
);

NOR3xp33_ASAP7_75t_SL g2504 ( 
.A(n_2449),
.B(n_2479),
.C(n_2483),
.Y(n_2504)
);

NOR2x1p5_ASAP7_75t_L g2505 ( 
.A(n_2491),
.B(n_369),
.Y(n_2505)
);

NOR5xp2_ASAP7_75t_L g2506 ( 
.A(n_2485),
.B(n_370),
.C(n_371),
.D(n_372),
.E(n_373),
.Y(n_2506)
);

NAND3xp33_ASAP7_75t_SL g2507 ( 
.A(n_2476),
.B(n_371),
.C(n_372),
.Y(n_2507)
);

XNOR2xp5_ASAP7_75t_L g2508 ( 
.A(n_2474),
.B(n_373),
.Y(n_2508)
);

AND3x1_ASAP7_75t_L g2509 ( 
.A(n_2453),
.B(n_374),
.C(n_375),
.Y(n_2509)
);

NOR2x1_ASAP7_75t_L g2510 ( 
.A(n_2445),
.B(n_374),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_L g2511 ( 
.A(n_2465),
.B(n_376),
.Y(n_2511)
);

INVxp67_ASAP7_75t_L g2512 ( 
.A(n_2458),
.Y(n_2512)
);

NAND4xp25_ASAP7_75t_L g2513 ( 
.A(n_2482),
.B(n_377),
.C(n_378),
.D(n_379),
.Y(n_2513)
);

NAND2xp5_ASAP7_75t_L g2514 ( 
.A(n_2467),
.B(n_2468),
.Y(n_2514)
);

NOR3xp33_ASAP7_75t_L g2515 ( 
.A(n_2470),
.B(n_377),
.C(n_379),
.Y(n_2515)
);

NAND3xp33_ASAP7_75t_SL g2516 ( 
.A(n_2455),
.B(n_381),
.C(n_382),
.Y(n_2516)
);

NOR3xp33_ASAP7_75t_L g2517 ( 
.A(n_2451),
.B(n_382),
.C(n_383),
.Y(n_2517)
);

NOR3xp33_ASAP7_75t_L g2518 ( 
.A(n_2488),
.B(n_383),
.C(n_384),
.Y(n_2518)
);

AO22x2_ASAP7_75t_L g2519 ( 
.A1(n_2456),
.A2(n_384),
.B1(n_385),
.B2(n_386),
.Y(n_2519)
);

NOR3xp33_ASAP7_75t_L g2520 ( 
.A(n_2452),
.B(n_385),
.C(n_387),
.Y(n_2520)
);

INVx1_ASAP7_75t_L g2521 ( 
.A(n_2480),
.Y(n_2521)
);

INVx1_ASAP7_75t_L g2522 ( 
.A(n_2473),
.Y(n_2522)
);

INVx5_ASAP7_75t_L g2523 ( 
.A(n_2466),
.Y(n_2523)
);

NOR3xp33_ASAP7_75t_SL g2524 ( 
.A(n_2486),
.B(n_387),
.C(n_388),
.Y(n_2524)
);

NOR3xp33_ASAP7_75t_L g2525 ( 
.A(n_2457),
.B(n_389),
.C(n_390),
.Y(n_2525)
);

NAND4xp25_ASAP7_75t_L g2526 ( 
.A(n_2460),
.B(n_2463),
.C(n_2468),
.D(n_2462),
.Y(n_2526)
);

NOR4xp75_ASAP7_75t_L g2527 ( 
.A(n_2492),
.B(n_390),
.C(n_391),
.D(n_392),
.Y(n_2527)
);

NAND5xp2_ASAP7_75t_L g2528 ( 
.A(n_2489),
.B(n_391),
.C(n_392),
.D(n_393),
.E(n_394),
.Y(n_2528)
);

NOR5xp2_ASAP7_75t_L g2529 ( 
.A(n_2472),
.B(n_393),
.C(n_394),
.D(n_395),
.E(n_396),
.Y(n_2529)
);

NAND5xp2_ASAP7_75t_L g2530 ( 
.A(n_2454),
.B(n_395),
.C(n_397),
.D(n_398),
.E(n_399),
.Y(n_2530)
);

INVxp67_ASAP7_75t_L g2531 ( 
.A(n_2459),
.Y(n_2531)
);

BUFx2_ASAP7_75t_L g2532 ( 
.A(n_2509),
.Y(n_2532)
);

INVx1_ASAP7_75t_SL g2533 ( 
.A(n_2511),
.Y(n_2533)
);

BUFx2_ASAP7_75t_L g2534 ( 
.A(n_2519),
.Y(n_2534)
);

INVx2_ASAP7_75t_L g2535 ( 
.A(n_2505),
.Y(n_2535)
);

NAND4xp25_ASAP7_75t_L g2536 ( 
.A(n_2513),
.B(n_2494),
.C(n_2526),
.D(n_2495),
.Y(n_2536)
);

CKINVDCx5p33_ASAP7_75t_R g2537 ( 
.A(n_2504),
.Y(n_2537)
);

OR2x2_ASAP7_75t_L g2538 ( 
.A(n_2530),
.B(n_2478),
.Y(n_2538)
);

BUFx2_ASAP7_75t_L g2539 ( 
.A(n_2510),
.Y(n_2539)
);

BUFx2_ASAP7_75t_L g2540 ( 
.A(n_2503),
.Y(n_2540)
);

CKINVDCx20_ASAP7_75t_R g2541 ( 
.A(n_2508),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2527),
.Y(n_2542)
);

NOR2xp67_ASAP7_75t_L g2543 ( 
.A(n_2528),
.B(n_2478),
.Y(n_2543)
);

CKINVDCx5p33_ASAP7_75t_R g2544 ( 
.A(n_2499),
.Y(n_2544)
);

CKINVDCx5p33_ASAP7_75t_R g2545 ( 
.A(n_2523),
.Y(n_2545)
);

CKINVDCx5p33_ASAP7_75t_R g2546 ( 
.A(n_2523),
.Y(n_2546)
);

CKINVDCx5p33_ASAP7_75t_R g2547 ( 
.A(n_2501),
.Y(n_2547)
);

INVx1_ASAP7_75t_L g2548 ( 
.A(n_2524),
.Y(n_2548)
);

INVx1_ASAP7_75t_L g2549 ( 
.A(n_2507),
.Y(n_2549)
);

OAI221xp5_ASAP7_75t_L g2550 ( 
.A1(n_2531),
.A2(n_397),
.B1(n_398),
.B2(n_399),
.C(n_400),
.Y(n_2550)
);

XNOR2x1_ASAP7_75t_L g2551 ( 
.A(n_2521),
.B(n_400),
.Y(n_2551)
);

CKINVDCx5p33_ASAP7_75t_R g2552 ( 
.A(n_2512),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2516),
.Y(n_2553)
);

BUFx2_ASAP7_75t_L g2554 ( 
.A(n_2522),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2498),
.B(n_2022),
.Y(n_2555)
);

NAND2x1_ASAP7_75t_L g2556 ( 
.A(n_2529),
.B(n_401),
.Y(n_2556)
);

OAI322xp33_ASAP7_75t_L g2557 ( 
.A1(n_2556),
.A2(n_2514),
.A3(n_2497),
.B1(n_2500),
.B2(n_2496),
.C1(n_2493),
.C2(n_2506),
.Y(n_2557)
);

OAI322xp33_ASAP7_75t_L g2558 ( 
.A1(n_2538),
.A2(n_2502),
.A3(n_2525),
.B1(n_2518),
.B2(n_2520),
.C1(n_2517),
.C2(n_2515),
.Y(n_2558)
);

AOI322xp5_ASAP7_75t_L g2559 ( 
.A1(n_2555),
.A2(n_401),
.A3(n_403),
.B1(n_405),
.B2(n_406),
.C1(n_407),
.C2(n_408),
.Y(n_2559)
);

AOI32xp33_ASAP7_75t_L g2560 ( 
.A1(n_2554),
.A2(n_403),
.A3(n_406),
.B1(n_409),
.B2(n_410),
.Y(n_2560)
);

AOI32xp33_ASAP7_75t_L g2561 ( 
.A1(n_2542),
.A2(n_411),
.A3(n_412),
.B1(n_413),
.B2(n_415),
.Y(n_2561)
);

AOI322xp5_ASAP7_75t_L g2562 ( 
.A1(n_2553),
.A2(n_411),
.A3(n_413),
.B1(n_415),
.B2(n_416),
.C1(n_418),
.C2(n_419),
.Y(n_2562)
);

INVxp67_ASAP7_75t_L g2563 ( 
.A(n_2551),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2545),
.Y(n_2564)
);

OAI221xp5_ASAP7_75t_L g2565 ( 
.A1(n_2546),
.A2(n_416),
.B1(n_418),
.B2(n_419),
.C(n_420),
.Y(n_2565)
);

AOI221xp5_ASAP7_75t_L g2566 ( 
.A1(n_2537),
.A2(n_420),
.B1(n_421),
.B2(n_422),
.C(n_423),
.Y(n_2566)
);

NOR2x1p5_ASAP7_75t_L g2567 ( 
.A(n_2548),
.B(n_421),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2534),
.Y(n_2568)
);

OAI322xp33_ASAP7_75t_SL g2569 ( 
.A1(n_2544),
.A2(n_422),
.A3(n_423),
.B1(n_424),
.B2(n_425),
.C1(n_426),
.C2(n_427),
.Y(n_2569)
);

AOI221xp5_ASAP7_75t_SL g2570 ( 
.A1(n_2536),
.A2(n_425),
.B1(n_426),
.B2(n_427),
.C(n_428),
.Y(n_2570)
);

AOI211x1_ASAP7_75t_L g2571 ( 
.A1(n_2536),
.A2(n_428),
.B(n_429),
.C(n_430),
.Y(n_2571)
);

INVx1_ASAP7_75t_SL g2572 ( 
.A(n_2532),
.Y(n_2572)
);

INVx1_ASAP7_75t_SL g2573 ( 
.A(n_2539),
.Y(n_2573)
);

OAI211xp5_ASAP7_75t_SL g2574 ( 
.A1(n_2549),
.A2(n_2533),
.B(n_2535),
.C(n_2552),
.Y(n_2574)
);

AOI322xp5_ASAP7_75t_L g2575 ( 
.A1(n_2540),
.A2(n_429),
.A3(n_431),
.B1(n_432),
.B2(n_433),
.C1(n_434),
.C2(n_435),
.Y(n_2575)
);

AOI221xp5_ASAP7_75t_L g2576 ( 
.A1(n_2547),
.A2(n_431),
.B1(n_436),
.B2(n_437),
.C(n_438),
.Y(n_2576)
);

OAI22xp5_ASAP7_75t_L g2577 ( 
.A1(n_2568),
.A2(n_2543),
.B1(n_2541),
.B2(n_2550),
.Y(n_2577)
);

OAI22x1_ASAP7_75t_L g2578 ( 
.A1(n_2567),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_2578)
);

NOR4xp25_ASAP7_75t_L g2579 ( 
.A(n_2557),
.B(n_440),
.C(n_441),
.D(n_442),
.Y(n_2579)
);

AOI31xp33_ASAP7_75t_L g2580 ( 
.A1(n_2572),
.A2(n_2573),
.A3(n_2563),
.B(n_2564),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2571),
.Y(n_2581)
);

AO22x2_ASAP7_75t_L g2582 ( 
.A1(n_2570),
.A2(n_440),
.B1(n_442),
.B2(n_443),
.Y(n_2582)
);

INVx2_ASAP7_75t_L g2583 ( 
.A(n_2565),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2558),
.Y(n_2584)
);

BUFx2_ASAP7_75t_L g2585 ( 
.A(n_2566),
.Y(n_2585)
);

INVx1_ASAP7_75t_L g2586 ( 
.A(n_2574),
.Y(n_2586)
);

AND4x2_ASAP7_75t_L g2587 ( 
.A(n_2576),
.B(n_443),
.C(n_444),
.D(n_445),
.Y(n_2587)
);

AO22x2_ASAP7_75t_L g2588 ( 
.A1(n_2560),
.A2(n_444),
.B1(n_447),
.B2(n_448),
.Y(n_2588)
);

XNOR2x1_ASAP7_75t_SL g2589 ( 
.A(n_2582),
.B(n_2569),
.Y(n_2589)
);

NAND5xp2_ASAP7_75t_L g2590 ( 
.A(n_2586),
.B(n_2561),
.C(n_2559),
.D(n_2562),
.E(n_2575),
.Y(n_2590)
);

XOR2xp5_ASAP7_75t_L g2591 ( 
.A(n_2577),
.B(n_447),
.Y(n_2591)
);

NOR2xp33_ASAP7_75t_L g2592 ( 
.A(n_2581),
.B(n_448),
.Y(n_2592)
);

OAI221xp5_ASAP7_75t_L g2593 ( 
.A1(n_2579),
.A2(n_449),
.B1(n_450),
.B2(n_451),
.C(n_453),
.Y(n_2593)
);

XNOR2xp5_ASAP7_75t_L g2594 ( 
.A(n_2584),
.B(n_449),
.Y(n_2594)
);

NAND2xp5_ASAP7_75t_L g2595 ( 
.A(n_2588),
.B(n_450),
.Y(n_2595)
);

INVx1_ASAP7_75t_L g2596 ( 
.A(n_2594),
.Y(n_2596)
);

OAI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2591),
.A2(n_2580),
.B1(n_2583),
.B2(n_2585),
.Y(n_2597)
);

OAI22x1_ASAP7_75t_L g2598 ( 
.A1(n_2592),
.A2(n_2595),
.B1(n_2589),
.B2(n_2590),
.Y(n_2598)
);

O2A1O1Ixp33_ASAP7_75t_SL g2599 ( 
.A1(n_2593),
.A2(n_2587),
.B(n_2578),
.C(n_455),
.Y(n_2599)
);

INVx2_ASAP7_75t_L g2600 ( 
.A(n_2594),
.Y(n_2600)
);

AND2x4_ASAP7_75t_L g2601 ( 
.A(n_2592),
.B(n_451),
.Y(n_2601)
);

OAI22xp5_ASAP7_75t_L g2602 ( 
.A1(n_2596),
.A2(n_454),
.B1(n_455),
.B2(n_457),
.Y(n_2602)
);

BUFx2_ASAP7_75t_L g2603 ( 
.A(n_2601),
.Y(n_2603)
);

AO22x1_ASAP7_75t_L g2604 ( 
.A1(n_2600),
.A2(n_457),
.B1(n_458),
.B2(n_459),
.Y(n_2604)
);

INVx1_ASAP7_75t_L g2605 ( 
.A(n_2599),
.Y(n_2605)
);

OAI22xp5_ASAP7_75t_SL g2606 ( 
.A1(n_2605),
.A2(n_2598),
.B1(n_2597),
.B2(n_461),
.Y(n_2606)
);

OAI22xp5_ASAP7_75t_SL g2607 ( 
.A1(n_2603),
.A2(n_458),
.B1(n_460),
.B2(n_461),
.Y(n_2607)
);

AOI22xp5_ASAP7_75t_L g2608 ( 
.A1(n_2602),
.A2(n_460),
.B1(n_462),
.B2(n_464),
.Y(n_2608)
);

INVx2_ASAP7_75t_L g2609 ( 
.A(n_2604),
.Y(n_2609)
);

OAI21x1_ASAP7_75t_SL g2610 ( 
.A1(n_2605),
.A2(n_464),
.B(n_465),
.Y(n_2610)
);

AOI21xp5_ASAP7_75t_L g2611 ( 
.A1(n_2606),
.A2(n_465),
.B(n_466),
.Y(n_2611)
);

NOR2xp67_ASAP7_75t_L g2612 ( 
.A(n_2609),
.B(n_466),
.Y(n_2612)
);

OAI22x1_ASAP7_75t_L g2613 ( 
.A1(n_2608),
.A2(n_467),
.B1(n_468),
.B2(n_469),
.Y(n_2613)
);

AOI22xp5_ASAP7_75t_L g2614 ( 
.A1(n_2607),
.A2(n_468),
.B1(n_470),
.B2(n_471),
.Y(n_2614)
);

OAI22xp5_ASAP7_75t_L g2615 ( 
.A1(n_2614),
.A2(n_2610),
.B1(n_473),
.B2(n_475),
.Y(n_2615)
);

AOI22xp5_ASAP7_75t_L g2616 ( 
.A1(n_2613),
.A2(n_471),
.B1(n_475),
.B2(n_476),
.Y(n_2616)
);

OAI22xp5_ASAP7_75t_L g2617 ( 
.A1(n_2611),
.A2(n_476),
.B1(n_477),
.B2(n_478),
.Y(n_2617)
);

NAND2xp5_ASAP7_75t_SL g2618 ( 
.A(n_2616),
.B(n_2612),
.Y(n_2618)
);

OA21x2_ASAP7_75t_L g2619 ( 
.A1(n_2617),
.A2(n_477),
.B(n_478),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2618),
.Y(n_2620)
);

AOI221xp5_ASAP7_75t_L g2621 ( 
.A1(n_2620),
.A2(n_2615),
.B1(n_2619),
.B2(n_482),
.C(n_483),
.Y(n_2621)
);

AOI21xp5_ASAP7_75t_L g2622 ( 
.A1(n_2621),
.A2(n_479),
.B(n_480),
.Y(n_2622)
);

AOI211xp5_ASAP7_75t_L g2623 ( 
.A1(n_2622),
.A2(n_479),
.B(n_480),
.C(n_482),
.Y(n_2623)
);


endmodule