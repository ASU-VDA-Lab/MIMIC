module fake_netlist_6_3706_n_1781 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1781);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1781;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_1738;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1009;
wire n_1743;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1704;
wire n_1078;
wire n_250;
wire n_544;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1697;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_210;
wire n_1069;
wire n_1664;
wire n_1722;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_1214;
wire n_928;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_1709;
wire n_1757;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1033;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_627;
wire n_297;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_1766;
wire n_1776;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_927;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_527;
wire n_474;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1769;
wire n_1220;
wire n_556;
wire n_162;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1267;
wire n_1281;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_171;
wire n_1764;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_1768;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_750;
wire n_1115;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1373;
wire n_1292;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_1725;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_545;
wire n_489;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_22),
.Y(n_155)
);

CKINVDCx5p33_ASAP7_75t_R g156 ( 
.A(n_38),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_3),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_138),
.Y(n_158)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_53),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_115),
.Y(n_160)
);

BUFx3_ASAP7_75t_L g161 ( 
.A(n_21),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_134),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_103),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_0),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_130),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_42),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_111),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_14),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_74),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_71),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_87),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_67),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_28),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_136),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_13),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_76),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_121),
.Y(n_178)
);

CKINVDCx5p33_ASAP7_75t_R g179 ( 
.A(n_9),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_122),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_52),
.Y(n_181)
);

INVx3_ASAP7_75t_L g182 ( 
.A(n_83),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_63),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_70),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_91),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx3_ASAP7_75t_L g187 ( 
.A(n_106),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_59),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g189 ( 
.A(n_34),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_82),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_96),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_0),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_52),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_23),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_109),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_2),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_101),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_100),
.Y(n_199)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_47),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_29),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_80),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_99),
.Y(n_203)
);

BUFx10_ASAP7_75t_L g204 ( 
.A(n_108),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_26),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_104),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_4),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_3),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_154),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_128),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_9),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_65),
.Y(n_212)
);

BUFx3_ASAP7_75t_L g213 ( 
.A(n_90),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_43),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_141),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_22),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_28),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_88),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_7),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_94),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_23),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_86),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g223 ( 
.A(n_7),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_143),
.Y(n_224)
);

BUFx5_ASAP7_75t_L g225 ( 
.A(n_133),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_75),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_129),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_93),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_69),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_151),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_142),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_27),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_20),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_42),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_18),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_81),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_84),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_14),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_57),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_32),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_19),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_18),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_89),
.Y(n_243)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_30),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_124),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_73),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_98),
.Y(n_247)
);

BUFx8_ASAP7_75t_SL g248 ( 
.A(n_92),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_112),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_16),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_120),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_58),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_113),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_119),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_146),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_62),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_72),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_5),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_144),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_132),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_10),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_54),
.Y(n_263)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_135),
.Y(n_264)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_77),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_153),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_60),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_39),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_50),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g270 ( 
.A(n_39),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_79),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_102),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_148),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_20),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_40),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_149),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_12),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_48),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_66),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_41),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_15),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_5),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_13),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g284 ( 
.A(n_78),
.Y(n_284)
);

INVx2_ASAP7_75t_SL g285 ( 
.A(n_51),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_34),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_32),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_36),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_140),
.Y(n_289)
);

BUFx10_ASAP7_75t_L g290 ( 
.A(n_21),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_27),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g292 ( 
.A(n_36),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_43),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_26),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_116),
.Y(n_295)
);

CKINVDCx5p33_ASAP7_75t_R g296 ( 
.A(n_16),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_55),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_110),
.Y(n_298)
);

BUFx10_ASAP7_75t_L g299 ( 
.A(n_38),
.Y(n_299)
);

BUFx3_ASAP7_75t_L g300 ( 
.A(n_123),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_147),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_30),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_127),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_49),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_118),
.Y(n_305)
);

INVx2_ASAP7_75t_SL g306 ( 
.A(n_50),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_56),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_248),
.Y(n_308)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_182),
.B(n_1),
.Y(n_309)
);

HB1xp67_ASAP7_75t_L g310 ( 
.A(n_189),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g311 ( 
.A(n_159),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_175),
.Y(n_312)
);

INVxp67_ASAP7_75t_SL g313 ( 
.A(n_187),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_182),
.B(n_1),
.Y(n_314)
);

INVx2_ASAP7_75t_L g315 ( 
.A(n_223),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_223),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_177),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_223),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_223),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g320 ( 
.A(n_287),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_223),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_178),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_180),
.Y(n_323)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_183),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_186),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_223),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_223),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_223),
.B(n_2),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_209),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_188),
.Y(n_331)
);

INVxp67_ASAP7_75t_SL g332 ( 
.A(n_187),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_198),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_195),
.Y(n_334)
);

NOR2xp67_ASAP7_75t_L g335 ( 
.A(n_182),
.B(n_6),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_199),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_228),
.Y(n_337)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_264),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_255),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_195),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_195),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_212),
.B(n_6),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_195),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_195),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_258),
.Y(n_345)
);

INVxp67_ASAP7_75t_SL g346 ( 
.A(n_213),
.Y(n_346)
);

XOR2x2_ASAP7_75t_L g347 ( 
.A(n_285),
.B(n_8),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_263),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_221),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_161),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_161),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_212),
.B(n_8),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_202),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_265),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_221),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_221),
.Y(n_356)
);

CKINVDCx20_ASAP7_75t_R g357 ( 
.A(n_267),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_221),
.Y(n_358)
);

INVxp67_ASAP7_75t_L g359 ( 
.A(n_290),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_221),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_247),
.B(n_10),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_206),
.Y(n_362)
);

NAND2xp33_ASAP7_75t_R g363 ( 
.A(n_158),
.B(n_11),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_244),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_244),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_244),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_244),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_215),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_218),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_244),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_276),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_270),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_270),
.Y(n_373)
);

INVxp67_ASAP7_75t_SL g374 ( 
.A(n_213),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_270),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_220),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_270),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_270),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_193),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_224),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_193),
.Y(n_381)
);

BUFx2_ASAP7_75t_L g382 ( 
.A(n_157),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_157),
.Y(n_383)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_315),
.Y(n_384)
);

BUFx6f_ASAP7_75t_L g385 ( 
.A(n_315),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_316),
.Y(n_386)
);

NOR2xp33_ASAP7_75t_L g387 ( 
.A(n_314),
.B(n_160),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_316),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_318),
.Y(n_389)
);

INVx3_ASAP7_75t_L g390 ( 
.A(n_318),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_334),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_334),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_340),
.Y(n_394)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_309),
.B(n_285),
.Y(n_395)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_319),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_313),
.B(n_300),
.Y(n_397)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_332),
.B(n_300),
.Y(n_398)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_321),
.Y(n_399)
);

INVxp33_ASAP7_75t_SL g400 ( 
.A(n_312),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_382),
.Y(n_401)
);

NOR2xp33_ASAP7_75t_SL g402 ( 
.A(n_335),
.B(n_306),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_346),
.B(n_247),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_321),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_340),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_341),
.Y(n_406)
);

INVx3_ASAP7_75t_L g407 ( 
.A(n_327),
.Y(n_407)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_327),
.Y(n_408)
);

AND2x4_ASAP7_75t_L g409 ( 
.A(n_341),
.B(n_303),
.Y(n_409)
);

INVx2_ASAP7_75t_L g410 ( 
.A(n_328),
.Y(n_410)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_328),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_343),
.Y(n_412)
);

INVx2_ASAP7_75t_L g413 ( 
.A(n_343),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_374),
.B(n_303),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_344),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_344),
.Y(n_416)
);

BUFx6f_ASAP7_75t_L g417 ( 
.A(n_349),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_349),
.Y(n_418)
);

AND2x2_ASAP7_75t_L g419 ( 
.A(n_350),
.B(n_163),
.Y(n_419)
);

AND2x2_ASAP7_75t_SL g420 ( 
.A(n_329),
.B(n_271),
.Y(n_420)
);

BUFx6f_ASAP7_75t_L g421 ( 
.A(n_355),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_355),
.B(n_165),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_356),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_356),
.Y(n_424)
);

INVx2_ASAP7_75t_L g425 ( 
.A(n_358),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g427 ( 
.A1(n_347),
.A2(n_240),
.B1(n_294),
.B2(n_211),
.Y(n_427)
);

INVx2_ASAP7_75t_L g428 ( 
.A(n_360),
.Y(n_428)
);

INVx2_ASAP7_75t_L g429 ( 
.A(n_360),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_364),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_365),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_365),
.B(n_366),
.Y(n_433)
);

INVx3_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_367),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_367),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_370),
.Y(n_437)
);

BUFx6f_ASAP7_75t_L g438 ( 
.A(n_370),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_351),
.B(n_167),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_372),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g441 ( 
.A(n_372),
.B(n_171),
.Y(n_441)
);

CKINVDCx5p33_ASAP7_75t_R g442 ( 
.A(n_380),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_373),
.Y(n_443)
);

BUFx6f_ASAP7_75t_L g444 ( 
.A(n_373),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_375),
.Y(n_445)
);

BUFx2_ASAP7_75t_L g446 ( 
.A(n_359),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_375),
.B(n_184),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_377),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_377),
.Y(n_449)
);

HB1xp67_ASAP7_75t_L g450 ( 
.A(n_382),
.Y(n_450)
);

AND2x2_ASAP7_75t_L g451 ( 
.A(n_378),
.B(n_185),
.Y(n_451)
);

INVx2_ASAP7_75t_L g452 ( 
.A(n_378),
.Y(n_452)
);

INVx1_ASAP7_75t_SL g453 ( 
.A(n_446),
.Y(n_453)
);

BUFx3_ASAP7_75t_L g454 ( 
.A(n_451),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_390),
.Y(n_455)
);

NAND2xp33_ASAP7_75t_R g456 ( 
.A(n_446),
.B(n_383),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_384),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

INVx2_ASAP7_75t_SL g459 ( 
.A(n_397),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_SL g460 ( 
.A(n_387),
.B(n_338),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_384),
.Y(n_461)
);

AND3x2_ASAP7_75t_L g462 ( 
.A(n_395),
.B(n_352),
.C(n_342),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_387),
.B(n_317),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_390),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_450),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_400),
.B(n_322),
.Y(n_466)
);

NAND2x1p5_ASAP7_75t_L g467 ( 
.A(n_420),
.B(n_190),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_400),
.B(n_325),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

BUFx3_ASAP7_75t_L g470 ( 
.A(n_451),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_390),
.Y(n_471)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_384),
.Y(n_472)
);

INVxp33_ASAP7_75t_L g473 ( 
.A(n_450),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_390),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_384),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_384),
.Y(n_476)
);

INVx2_ASAP7_75t_L g477 ( 
.A(n_388),
.Y(n_477)
);

INVx1_ASAP7_75t_SL g478 ( 
.A(n_442),
.Y(n_478)
);

INVxp33_ASAP7_75t_L g479 ( 
.A(n_446),
.Y(n_479)
);

INVx1_ASAP7_75t_SL g480 ( 
.A(n_442),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_407),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_403),
.B(n_331),
.Y(n_482)
);

INVx2_ASAP7_75t_SL g483 ( 
.A(n_397),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_395),
.B(n_333),
.Y(n_484)
);

BUFx3_ASAP7_75t_L g485 ( 
.A(n_451),
.Y(n_485)
);

OAI21xp33_ASAP7_75t_SL g486 ( 
.A1(n_420),
.A2(n_361),
.B(n_306),
.Y(n_486)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_401),
.A2(n_347),
.B1(n_363),
.B2(n_166),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_403),
.B(n_336),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_403),
.B(n_353),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_388),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_403),
.B(n_362),
.Y(n_491)
);

AO22x2_ASAP7_75t_L g492 ( 
.A1(n_401),
.A2(n_235),
.B1(n_302),
.B2(n_208),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_395),
.B(n_368),
.Y(n_493)
);

INVx1_ASAP7_75t_SL g494 ( 
.A(n_397),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_407),
.Y(n_495)
);

AND2x2_ASAP7_75t_L g496 ( 
.A(n_414),
.B(n_381),
.Y(n_496)
);

INVx1_ASAP7_75t_SL g497 ( 
.A(n_397),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_414),
.B(n_369),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_L g499 ( 
.A(n_414),
.B(n_376),
.Y(n_499)
);

INVx3_ASAP7_75t_L g500 ( 
.A(n_385),
.Y(n_500)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_398),
.Y(n_501)
);

NAND2xp33_ASAP7_75t_L g502 ( 
.A(n_414),
.B(n_271),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_407),
.Y(n_503)
);

INVx2_ASAP7_75t_SL g504 ( 
.A(n_398),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_402),
.B(n_308),
.Y(n_505)
);

INVx3_ASAP7_75t_L g506 ( 
.A(n_385),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_402),
.B(n_204),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_402),
.A2(n_166),
.B1(n_168),
.B2(n_164),
.Y(n_508)
);

INVx2_ASAP7_75t_L g509 ( 
.A(n_388),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_398),
.B(n_204),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_407),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_388),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_398),
.B(n_420),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_407),
.Y(n_514)
);

BUFx6f_ASAP7_75t_L g515 ( 
.A(n_385),
.Y(n_515)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_419),
.B(n_310),
.Y(n_516)
);

AND2x2_ASAP7_75t_L g517 ( 
.A(n_419),
.B(n_379),
.Y(n_517)
);

OAI22xp33_ASAP7_75t_L g518 ( 
.A1(n_427),
.A2(n_194),
.B1(n_269),
.B2(n_268),
.Y(n_518)
);

INVx2_ASAP7_75t_L g519 ( 
.A(n_388),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_407),
.Y(n_520)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_389),
.Y(n_521)
);

INVx2_ASAP7_75t_L g522 ( 
.A(n_389),
.Y(n_522)
);

INVx2_ASAP7_75t_L g523 ( 
.A(n_389),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_389),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_389),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_393),
.Y(n_526)
);

AND2x6_ASAP7_75t_L g527 ( 
.A(n_451),
.B(n_271),
.Y(n_527)
);

INVx4_ASAP7_75t_L g528 ( 
.A(n_385),
.Y(n_528)
);

INVx2_ASAP7_75t_SL g529 ( 
.A(n_419),
.Y(n_529)
);

INVx4_ASAP7_75t_L g530 ( 
.A(n_385),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_393),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g532 ( 
.A(n_419),
.B(n_320),
.Y(n_532)
);

BUFx6f_ASAP7_75t_L g533 ( 
.A(n_385),
.Y(n_533)
);

INVx1_ASAP7_75t_SL g534 ( 
.A(n_439),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_393),
.Y(n_535)
);

AND2x2_ASAP7_75t_L g536 ( 
.A(n_439),
.B(n_379),
.Y(n_536)
);

BUFx4f_ASAP7_75t_L g537 ( 
.A(n_420),
.Y(n_537)
);

BUFx3_ASAP7_75t_L g538 ( 
.A(n_439),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_420),
.B(n_245),
.Y(n_539)
);

INVx2_ASAP7_75t_SL g540 ( 
.A(n_439),
.Y(n_540)
);

OR2x2_ASAP7_75t_L g541 ( 
.A(n_422),
.B(n_324),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_385),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_393),
.B(n_396),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_393),
.Y(n_544)
);

OAI22xp33_ASAP7_75t_L g545 ( 
.A1(n_427),
.A2(n_181),
.B1(n_197),
.B2(n_201),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_396),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_396),
.Y(n_547)
);

INVx2_ASAP7_75t_L g548 ( 
.A(n_396),
.Y(n_548)
);

AND3x1_ASAP7_75t_L g549 ( 
.A(n_427),
.B(n_235),
.C(n_208),
.Y(n_549)
);

CKINVDCx5p33_ASAP7_75t_R g550 ( 
.A(n_409),
.Y(n_550)
);

INVx2_ASAP7_75t_L g551 ( 
.A(n_396),
.Y(n_551)
);

INVx1_ASAP7_75t_SL g552 ( 
.A(n_422),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_399),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_399),
.Y(n_554)
);

BUFx6f_ASAP7_75t_L g555 ( 
.A(n_385),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_399),
.B(n_284),
.Y(n_556)
);

INVx2_ASAP7_75t_L g557 ( 
.A(n_399),
.Y(n_557)
);

INVx3_ASAP7_75t_L g558 ( 
.A(n_385),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_399),
.Y(n_559)
);

AND2x6_ASAP7_75t_L g560 ( 
.A(n_408),
.B(n_271),
.Y(n_560)
);

NAND2xp33_ASAP7_75t_SL g561 ( 
.A(n_422),
.B(n_164),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_408),
.B(n_410),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_385),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_408),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_408),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_408),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_410),
.Y(n_567)
);

INVx1_ASAP7_75t_SL g568 ( 
.A(n_441),
.Y(n_568)
);

AND3x1_ASAP7_75t_L g569 ( 
.A(n_441),
.B(n_302),
.C(n_176),
.Y(n_569)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_410),
.B(n_226),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_410),
.Y(n_571)
);

BUFx6f_ASAP7_75t_L g572 ( 
.A(n_404),
.Y(n_572)
);

AND2x2_ASAP7_75t_L g573 ( 
.A(n_409),
.B(n_381),
.Y(n_573)
);

AO22x2_ASAP7_75t_L g574 ( 
.A1(n_409),
.A2(n_234),
.B1(n_275),
.B2(n_262),
.Y(n_574)
);

INVx5_ASAP7_75t_L g575 ( 
.A(n_404),
.Y(n_575)
);

INVx2_ASAP7_75t_L g576 ( 
.A(n_410),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_411),
.B(n_229),
.Y(n_577)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_411),
.B(n_230),
.Y(n_578)
);

INVx2_ASAP7_75t_L g579 ( 
.A(n_411),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_411),
.B(n_231),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_411),
.B(n_239),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_409),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_391),
.B(n_392),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_391),
.B(n_243),
.Y(n_584)
);

NOR3xp33_ASAP7_75t_SL g585 ( 
.A(n_441),
.B(n_173),
.C(n_168),
.Y(n_585)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_424),
.Y(n_586)
);

XNOR2xp5_ASAP7_75t_L g587 ( 
.A(n_409),
.B(n_311),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_424),
.Y(n_588)
);

BUFx3_ASAP7_75t_L g589 ( 
.A(n_409),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_391),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_424),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_392),
.Y(n_592)
);

INVx4_ASAP7_75t_SL g593 ( 
.A(n_404),
.Y(n_593)
);

AND2x4_ASAP7_75t_L g594 ( 
.A(n_409),
.B(n_191),
.Y(n_594)
);

INVx2_ASAP7_75t_L g595 ( 
.A(n_424),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_425),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_447),
.B(n_371),
.Y(n_597)
);

INVx3_ASAP7_75t_L g598 ( 
.A(n_404),
.Y(n_598)
);

AND3x2_ASAP7_75t_L g599 ( 
.A(n_447),
.B(n_200),
.C(n_242),
.Y(n_599)
);

NOR3xp33_ASAP7_75t_L g600 ( 
.A(n_447),
.B(n_256),
.C(n_155),
.Y(n_600)
);

NOR2x1p5_ASAP7_75t_L g601 ( 
.A(n_433),
.B(n_173),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_552),
.B(n_404),
.Y(n_602)
);

AOI22xp33_ASAP7_75t_L g603 ( 
.A1(n_513),
.A2(n_192),
.B1(n_196),
.B2(n_203),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_552),
.B(n_404),
.Y(n_604)
);

A2O1A1Ixp33_ASAP7_75t_L g605 ( 
.A1(n_486),
.A2(n_304),
.B(n_259),
.C(n_216),
.Y(n_605)
);

INVxp67_ASAP7_75t_L g606 ( 
.A(n_456),
.Y(n_606)
);

AND2x2_ASAP7_75t_L g607 ( 
.A(n_497),
.B(n_323),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_568),
.B(n_404),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_590),
.Y(n_609)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_463),
.B(n_326),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_573),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_459),
.B(n_404),
.Y(n_612)
);

OR2x2_ASAP7_75t_L g613 ( 
.A(n_453),
.B(n_465),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_537),
.B(n_404),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_590),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_573),
.Y(n_616)
);

BUFx6f_ASAP7_75t_L g617 ( 
.A(n_589),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_L g618 ( 
.A(n_459),
.B(n_404),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_454),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_483),
.B(n_386),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_454),
.Y(n_621)
);

NAND2xp5_ASAP7_75t_SL g622 ( 
.A(n_537),
.B(n_271),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_483),
.B(n_386),
.Y(n_623)
);

NAND2xp5_ASAP7_75t_L g624 ( 
.A(n_501),
.B(n_386),
.Y(n_624)
);

NAND3xp33_ASAP7_75t_L g625 ( 
.A(n_516),
.B(n_179),
.C(n_156),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_501),
.B(n_386),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_497),
.B(n_330),
.Y(n_627)
);

CKINVDCx5p33_ASAP7_75t_R g628 ( 
.A(n_478),
.Y(n_628)
);

AOI22xp5_ASAP7_75t_L g629 ( 
.A1(n_494),
.A2(n_348),
.B1(n_354),
.B2(n_357),
.Y(n_629)
);

NOR2xp33_ASAP7_75t_L g630 ( 
.A(n_597),
.B(n_482),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_504),
.B(n_386),
.Y(n_631)
);

CKINVDCx11_ASAP7_75t_R g632 ( 
.A(n_480),
.Y(n_632)
);

OA21x2_ASAP7_75t_L g633 ( 
.A1(n_543),
.A2(n_394),
.B(n_392),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_592),
.Y(n_634)
);

INVx8_ASAP7_75t_L g635 ( 
.A(n_550),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_470),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_504),
.B(n_386),
.Y(n_637)
);

AND2x2_ASAP7_75t_L g638 ( 
.A(n_534),
.B(n_337),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_539),
.B(n_386),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_L g640 ( 
.A(n_529),
.B(n_386),
.Y(n_640)
);

OAI22xp5_ASAP7_75t_L g641 ( 
.A1(n_537),
.A2(n_345),
.B1(n_339),
.B2(n_227),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_470),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_SL g643 ( 
.A(n_486),
.B(n_272),
.Y(n_643)
);

NOR2xp33_ASAP7_75t_L g644 ( 
.A(n_488),
.B(n_489),
.Y(n_644)
);

INVxp67_ASAP7_75t_SL g645 ( 
.A(n_485),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_529),
.B(n_386),
.Y(n_646)
);

INVx8_ASAP7_75t_L g647 ( 
.A(n_550),
.Y(n_647)
);

NOR2xp33_ASAP7_75t_L g648 ( 
.A(n_491),
.B(n_158),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_592),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_485),
.Y(n_650)
);

INVx4_ASAP7_75t_L g651 ( 
.A(n_515),
.Y(n_651)
);

CKINVDCx5p33_ASAP7_75t_R g652 ( 
.A(n_505),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_589),
.Y(n_653)
);

NAND2xp5_ASAP7_75t_L g654 ( 
.A(n_540),
.B(n_386),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_540),
.B(n_467),
.Y(n_655)
);

NOR3xp33_ASAP7_75t_L g656 ( 
.A(n_460),
.B(n_278),
.C(n_250),
.Y(n_656)
);

NAND2xp33_ASAP7_75t_L g657 ( 
.A(n_467),
.B(n_225),
.Y(n_657)
);

AOI22xp33_ASAP7_75t_L g658 ( 
.A1(n_467),
.A2(n_298),
.B1(n_307),
.B2(n_210),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_586),
.Y(n_659)
);

INVxp33_ASAP7_75t_L g660 ( 
.A(n_532),
.Y(n_660)
);

NAND2xp5_ASAP7_75t_SL g661 ( 
.A(n_582),
.B(n_272),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_SL g662 ( 
.A(n_582),
.B(n_272),
.Y(n_662)
);

NAND2xp5_ASAP7_75t_L g663 ( 
.A(n_498),
.B(n_386),
.Y(n_663)
);

O2A1O1Ixp5_ASAP7_75t_L g664 ( 
.A1(n_570),
.A2(n_394),
.B(n_449),
.C(n_412),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_SL g665 ( 
.A(n_538),
.B(n_272),
.Y(n_665)
);

OAI21xp5_ASAP7_75t_L g666 ( 
.A1(n_563),
.A2(n_433),
.B(n_434),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_538),
.B(n_272),
.Y(n_667)
);

NOR2xp67_ASAP7_75t_L g668 ( 
.A(n_541),
.B(n_433),
.Y(n_668)
);

NAND2xp5_ASAP7_75t_L g669 ( 
.A(n_499),
.B(n_394),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_SL g670 ( 
.A(n_455),
.B(n_225),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_SL g671 ( 
.A(n_455),
.B(n_458),
.Y(n_671)
);

HB1xp67_ASAP7_75t_L g672 ( 
.A(n_465),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_458),
.B(n_225),
.Y(n_673)
);

NOR2xp67_ASAP7_75t_L g674 ( 
.A(n_541),
.B(n_246),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_517),
.Y(n_675)
);

O2A1O1Ixp33_ASAP7_75t_L g676 ( 
.A1(n_502),
.A2(n_415),
.B(n_449),
.C(n_412),
.Y(n_676)
);

AOI22xp33_ASAP7_75t_L g677 ( 
.A1(n_594),
.A2(n_295),
.B1(n_237),
.B2(n_222),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_517),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_572),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_496),
.B(n_405),
.Y(n_680)
);

NAND2xp33_ASAP7_75t_L g681 ( 
.A(n_527),
.B(n_225),
.Y(n_681)
);

OR2x2_ASAP7_75t_L g682 ( 
.A(n_453),
.B(n_238),
.Y(n_682)
);

O2A1O1Ixp5_ASAP7_75t_L g683 ( 
.A1(n_577),
.A2(n_580),
.B(n_581),
.C(n_578),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_464),
.B(n_225),
.Y(n_684)
);

INVx2_ASAP7_75t_L g685 ( 
.A(n_586),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_536),
.Y(n_686)
);

AND2x6_ASAP7_75t_L g687 ( 
.A(n_464),
.B(n_236),
.Y(n_687)
);

NAND2xp5_ASAP7_75t_SL g688 ( 
.A(n_469),
.B(n_471),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_588),
.Y(n_689)
);

NOR2xp67_ASAP7_75t_L g690 ( 
.A(n_466),
.B(n_468),
.Y(n_690)
);

INVx1_ASAP7_75t_L g691 ( 
.A(n_536),
.Y(n_691)
);

INVx2_ASAP7_75t_L g692 ( 
.A(n_588),
.Y(n_692)
);

NOR2xp67_ASAP7_75t_L g693 ( 
.A(n_587),
.B(n_249),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_496),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_462),
.B(n_469),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_471),
.B(n_405),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_474),
.Y(n_697)
);

OAI22xp33_ASAP7_75t_L g698 ( 
.A1(n_479),
.A2(n_291),
.B1(n_293),
.B2(n_238),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_591),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_L g700 ( 
.A(n_473),
.B(n_162),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_474),
.B(n_405),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_481),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_591),
.Y(n_703)
);

BUFx2_ASAP7_75t_L g704 ( 
.A(n_587),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_481),
.B(n_406),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_595),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_SL g707 ( 
.A(n_495),
.B(n_225),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_495),
.B(n_406),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_L g709 ( 
.A(n_503),
.B(n_406),
.Y(n_709)
);

AND2x2_ASAP7_75t_L g710 ( 
.A(n_487),
.B(n_290),
.Y(n_710)
);

INVx2_ASAP7_75t_SL g711 ( 
.A(n_601),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_503),
.B(n_412),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_511),
.B(n_415),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_595),
.Y(n_714)
);

AND2x2_ASAP7_75t_SL g715 ( 
.A(n_549),
.B(n_415),
.Y(n_715)
);

INVx1_ASAP7_75t_L g716 ( 
.A(n_511),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_596),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_596),
.Y(n_718)
);

INVx1_ASAP7_75t_L g719 ( 
.A(n_514),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_514),
.B(n_430),
.Y(n_720)
);

INVx2_ASAP7_75t_L g721 ( 
.A(n_477),
.Y(n_721)
);

INVx1_ASAP7_75t_L g722 ( 
.A(n_520),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_SL g723 ( 
.A(n_520),
.B(n_225),
.Y(n_723)
);

INVx1_ASAP7_75t_L g724 ( 
.A(n_583),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_601),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_594),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_484),
.B(n_493),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_SL g728 ( 
.A(n_594),
.B(n_225),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_556),
.B(n_430),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_SL g730 ( 
.A(n_594),
.B(n_251),
.Y(n_730)
);

NAND2xp5_ASAP7_75t_L g731 ( 
.A(n_584),
.B(n_430),
.Y(n_731)
);

INVx3_ASAP7_75t_L g732 ( 
.A(n_515),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_487),
.B(n_290),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_477),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_502),
.B(n_432),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_521),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_598),
.B(n_432),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_521),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_598),
.B(n_432),
.Y(n_739)
);

INVx8_ASAP7_75t_L g740 ( 
.A(n_527),
.Y(n_740)
);

INVx2_ASAP7_75t_L g741 ( 
.A(n_490),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_510),
.B(n_507),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_490),
.Y(n_743)
);

AOI22xp5_ASAP7_75t_L g744 ( 
.A1(n_561),
.A2(n_266),
.B1(n_252),
.B2(n_253),
.Y(n_744)
);

OAI22xp5_ASAP7_75t_L g745 ( 
.A1(n_508),
.A2(n_170),
.B1(n_169),
.B2(n_162),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_598),
.B(n_437),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_509),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_525),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_500),
.B(n_506),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_515),
.B(n_254),
.Y(n_750)
);

BUFx3_ASAP7_75t_L g751 ( 
.A(n_515),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_509),
.Y(n_752)
);

BUFx3_ASAP7_75t_L g753 ( 
.A(n_515),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_533),
.B(n_555),
.Y(n_754)
);

NAND3xp33_ASAP7_75t_L g755 ( 
.A(n_508),
.B(n_232),
.C(n_205),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_L g756 ( 
.A(n_527),
.B(n_169),
.Y(n_756)
);

OAI22xp33_ASAP7_75t_L g757 ( 
.A1(n_518),
.A2(n_545),
.B1(n_291),
.B2(n_296),
.Y(n_757)
);

NAND2xp5_ASAP7_75t_L g758 ( 
.A(n_500),
.B(n_437),
.Y(n_758)
);

NOR2xp33_ASAP7_75t_L g759 ( 
.A(n_599),
.B(n_170),
.Y(n_759)
);

BUFx6f_ASAP7_75t_L g760 ( 
.A(n_572),
.Y(n_760)
);

NOR2xp33_ASAP7_75t_L g761 ( 
.A(n_528),
.B(n_172),
.Y(n_761)
);

INVx2_ASAP7_75t_SL g762 ( 
.A(n_492),
.Y(n_762)
);

A2O1A1Ixp33_ASAP7_75t_L g763 ( 
.A1(n_600),
.A2(n_293),
.B(n_296),
.C(n_283),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_492),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_SL g765 ( 
.A(n_533),
.B(n_257),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_500),
.B(n_506),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_506),
.B(n_437),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_525),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_542),
.B(n_440),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_512),
.Y(n_770)
);

AOI22xp5_ASAP7_75t_L g771 ( 
.A1(n_574),
.A2(n_279),
.B1(n_260),
.B2(n_261),
.Y(n_771)
);

BUFx2_ASAP7_75t_R g772 ( 
.A(n_549),
.Y(n_772)
);

HB1xp67_ASAP7_75t_L g773 ( 
.A(n_492),
.Y(n_773)
);

OR2x2_ASAP7_75t_L g774 ( 
.A(n_512),
.B(n_207),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_651),
.A2(n_528),
.B(n_530),
.Y(n_775)
);

NOR2xp33_ASAP7_75t_L g776 ( 
.A(n_660),
.B(n_528),
.Y(n_776)
);

INVx4_ASAP7_75t_L g777 ( 
.A(n_617),
.Y(n_777)
);

OAI21xp5_ASAP7_75t_L g778 ( 
.A1(n_605),
.A2(n_562),
.B(n_531),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_630),
.B(n_585),
.Y(n_779)
);

OAI21xp5_ASAP7_75t_L g780 ( 
.A1(n_605),
.A2(n_531),
.B(n_535),
.Y(n_780)
);

OAI21xp5_ASAP7_75t_L g781 ( 
.A1(n_643),
.A2(n_553),
.B(n_535),
.Y(n_781)
);

AOI21xp5_ASAP7_75t_L g782 ( 
.A1(n_651),
.A2(n_530),
.B(n_533),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_SL g783 ( 
.A(n_644),
.B(n_569),
.Y(n_783)
);

OAI321xp33_ASAP7_75t_L g784 ( 
.A1(n_757),
.A2(n_492),
.A3(n_569),
.B1(n_449),
.B2(n_440),
.C(n_443),
.Y(n_784)
);

AOI21xp5_ASAP7_75t_L g785 ( 
.A1(n_651),
.A2(n_530),
.B(n_533),
.Y(n_785)
);

AOI21xp33_ASAP7_75t_L g786 ( 
.A1(n_660),
.A2(n_574),
.B(n_559),
.Y(n_786)
);

OAI21xp33_ASAP7_75t_L g787 ( 
.A1(n_700),
.A2(n_288),
.B(n_286),
.Y(n_787)
);

AOI21x1_ASAP7_75t_L g788 ( 
.A1(n_614),
.A2(n_553),
.B(n_559),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_609),
.Y(n_789)
);

AOI21xp5_ASAP7_75t_L g790 ( 
.A1(n_614),
.A2(n_533),
.B(n_555),
.Y(n_790)
);

NOR2xp33_ASAP7_75t_L g791 ( 
.A(n_652),
.B(n_606),
.Y(n_791)
);

AND2x4_ASAP7_75t_L g792 ( 
.A(n_675),
.B(n_678),
.Y(n_792)
);

AO21x1_ASAP7_75t_L g793 ( 
.A1(n_622),
.A2(n_567),
.B(n_571),
.Y(n_793)
);

OAI21xp5_ASAP7_75t_L g794 ( 
.A1(n_643),
.A2(n_564),
.B(n_567),
.Y(n_794)
);

AOI21xp5_ASAP7_75t_L g795 ( 
.A1(n_657),
.A2(n_555),
.B(n_542),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_724),
.B(n_564),
.Y(n_796)
);

AOI22xp5_ASAP7_75t_L g797 ( 
.A1(n_727),
.A2(n_742),
.B1(n_695),
.B2(n_645),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_668),
.B(n_542),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_669),
.B(n_558),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_657),
.A2(n_555),
.B(n_558),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_SL g801 ( 
.A(n_617),
.B(n_172),
.Y(n_801)
);

AOI21xp5_ASAP7_75t_L g802 ( 
.A1(n_655),
.A2(n_555),
.B(n_558),
.Y(n_802)
);

INVx3_ASAP7_75t_L g803 ( 
.A(n_617),
.Y(n_803)
);

AND2x4_ASAP7_75t_SL g804 ( 
.A(n_672),
.B(n_204),
.Y(n_804)
);

OAI21xp5_ASAP7_75t_L g805 ( 
.A1(n_683),
.A2(n_571),
.B(n_579),
.Y(n_805)
);

AOI21xp5_ASAP7_75t_L g806 ( 
.A1(n_655),
.A2(n_572),
.B(n_575),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_617),
.Y(n_807)
);

OAI21x1_ASAP7_75t_L g808 ( 
.A1(n_749),
.A2(n_524),
.B(n_579),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_613),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_608),
.B(n_519),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_615),
.Y(n_811)
);

O2A1O1Ixp33_ASAP7_75t_L g812 ( 
.A1(n_773),
.A2(n_526),
.B(n_576),
.C(n_519),
.Y(n_812)
);

BUFx6f_ASAP7_75t_L g813 ( 
.A(n_679),
.Y(n_813)
);

AOI21xp5_ASAP7_75t_L g814 ( 
.A1(n_663),
.A2(n_572),
.B(n_575),
.Y(n_814)
);

AOI21x1_ASAP7_75t_L g815 ( 
.A1(n_754),
.A2(n_524),
.B(n_576),
.Y(n_815)
);

INVxp67_ASAP7_75t_L g816 ( 
.A(n_682),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_634),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_610),
.B(n_174),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_607),
.B(n_574),
.Y(n_819)
);

AOI21xp5_ASAP7_75t_L g820 ( 
.A1(n_602),
.A2(n_572),
.B(n_575),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_627),
.B(n_574),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_634),
.Y(n_822)
);

NOR2xp33_ASAP7_75t_SL g823 ( 
.A(n_628),
.B(n_174),
.Y(n_823)
);

NOR2xp33_ASAP7_75t_L g824 ( 
.A(n_638),
.B(n_297),
.Y(n_824)
);

AND2x2_ASAP7_75t_L g825 ( 
.A(n_694),
.B(n_299),
.Y(n_825)
);

AND2x4_ASAP7_75t_L g826 ( 
.A(n_686),
.B(n_593),
.Y(n_826)
);

OAI321xp33_ASAP7_75t_L g827 ( 
.A1(n_763),
.A2(n_443),
.A3(n_440),
.B1(n_299),
.B2(n_425),
.C(n_426),
.Y(n_827)
);

BUFx2_ASAP7_75t_L g828 ( 
.A(n_629),
.Y(n_828)
);

AOI22xp5_ASAP7_75t_L g829 ( 
.A1(n_611),
.A2(n_527),
.B1(n_289),
.B2(n_273),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_762),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_604),
.B(n_522),
.Y(n_831)
);

INVx1_ASAP7_75t_L g832 ( 
.A(n_649),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_639),
.A2(n_575),
.B(n_522),
.Y(n_833)
);

AOI21xp5_ASAP7_75t_L g834 ( 
.A1(n_754),
.A2(n_575),
.B(n_548),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_648),
.B(n_523),
.Y(n_835)
);

AND2x2_ASAP7_75t_L g836 ( 
.A(n_674),
.B(n_299),
.Y(n_836)
);

AOI21xp5_ASAP7_75t_L g837 ( 
.A1(n_751),
.A2(n_575),
.B(n_548),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_649),
.Y(n_838)
);

AND2x4_ASAP7_75t_L g839 ( 
.A(n_691),
.B(n_593),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_751),
.A2(n_547),
.B(n_566),
.Y(n_840)
);

OAI321xp33_ASAP7_75t_L g841 ( 
.A1(n_763),
.A2(n_443),
.A3(n_426),
.B1(n_428),
.B2(n_425),
.C(n_452),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_SL g842 ( 
.A(n_690),
.B(n_297),
.Y(n_842)
);

OAI22xp5_ASAP7_75t_L g843 ( 
.A1(n_764),
.A2(n_277),
.B1(n_281),
.B2(n_280),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_753),
.A2(n_547),
.B(n_566),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_753),
.A2(n_546),
.B(n_565),
.Y(n_845)
);

INVx1_ASAP7_75t_L g846 ( 
.A(n_697),
.Y(n_846)
);

HB1xp67_ASAP7_75t_L g847 ( 
.A(n_725),
.Y(n_847)
);

AND2x4_ASAP7_75t_L g848 ( 
.A(n_619),
.B(n_593),
.Y(n_848)
);

OAI21xp5_ASAP7_75t_L g849 ( 
.A1(n_664),
.A2(n_546),
.B(n_565),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_621),
.B(n_523),
.Y(n_850)
);

INVx3_ASAP7_75t_L g851 ( 
.A(n_653),
.Y(n_851)
);

AND2x4_ASAP7_75t_L g852 ( 
.A(n_636),
.B(n_642),
.Y(n_852)
);

OAI21xp5_ASAP7_75t_L g853 ( 
.A1(n_622),
.A2(n_544),
.B(n_526),
.Y(n_853)
);

AND2x2_ASAP7_75t_L g854 ( 
.A(n_710),
.B(n_214),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_SL g855 ( 
.A(n_650),
.B(n_301),
.Y(n_855)
);

BUFx6f_ASAP7_75t_L g856 ( 
.A(n_679),
.Y(n_856)
);

AOI21xp5_ASAP7_75t_L g857 ( 
.A1(n_612),
.A2(n_551),
.B(n_544),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_618),
.A2(n_551),
.B(n_554),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_620),
.A2(n_557),
.B(n_554),
.Y(n_859)
);

BUFx3_ASAP7_75t_L g860 ( 
.A(n_632),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_623),
.A2(n_557),
.B(n_461),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_733),
.B(n_217),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_616),
.A2(n_527),
.B1(n_301),
.B2(n_305),
.Y(n_863)
);

BUFx3_ASAP7_75t_L g864 ( 
.A(n_632),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_641),
.B(n_305),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_731),
.B(n_457),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_624),
.A2(n_457),
.B(n_461),
.Y(n_867)
);

NOR2xp33_ASAP7_75t_L g868 ( 
.A(n_625),
.B(n_219),
.Y(n_868)
);

BUFx2_ASAP7_75t_L g869 ( 
.A(n_704),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_680),
.B(n_472),
.Y(n_870)
);

AOI21xp5_ASAP7_75t_L g871 ( 
.A1(n_626),
.A2(n_472),
.B(n_475),
.Y(n_871)
);

O2A1O1Ixp5_ASAP7_75t_L g872 ( 
.A1(n_665),
.A2(n_476),
.B(n_475),
.C(n_434),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_711),
.B(n_233),
.Y(n_873)
);

NOR2xp33_ASAP7_75t_L g874 ( 
.A(n_745),
.B(n_241),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_702),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_653),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_631),
.A2(n_476),
.B(n_413),
.Y(n_877)
);

AND2x2_ASAP7_75t_L g878 ( 
.A(n_693),
.B(n_282),
.Y(n_878)
);

NOR2xp33_ASAP7_75t_L g879 ( 
.A(n_715),
.B(n_274),
.Y(n_879)
);

OAI22xp5_ASAP7_75t_L g880 ( 
.A1(n_603),
.A2(n_434),
.B1(n_418),
.B2(n_448),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_SL g881 ( 
.A(n_715),
.B(n_593),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_729),
.B(n_527),
.Y(n_882)
);

AOI21xp5_ASAP7_75t_L g883 ( 
.A1(n_637),
.A2(n_431),
.B(n_416),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_761),
.B(n_716),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_698),
.B(n_11),
.Y(n_885)
);

AND2x2_ASAP7_75t_L g886 ( 
.A(n_759),
.B(n_656),
.Y(n_886)
);

NOR2xp67_ASAP7_75t_L g887 ( 
.A(n_755),
.B(n_117),
.Y(n_887)
);

O2A1O1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_665),
.A2(n_434),
.B(n_452),
.C(n_428),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_771),
.B(n_744),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_766),
.A2(n_431),
.B(n_416),
.Y(n_890)
);

BUFx2_ASAP7_75t_L g891 ( 
.A(n_774),
.Y(n_891)
);

INVx4_ASAP7_75t_L g892 ( 
.A(n_635),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_640),
.A2(n_431),
.B(n_416),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_635),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_719),
.Y(n_895)
);

BUFx6f_ASAP7_75t_L g896 ( 
.A(n_679),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_635),
.B(n_417),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_722),
.B(n_658),
.Y(n_898)
);

NOR3xp33_ASAP7_75t_L g899 ( 
.A(n_730),
.B(n_434),
.C(n_452),
.Y(n_899)
);

A2O1A1Ixp33_ASAP7_75t_L g900 ( 
.A1(n_726),
.A2(n_434),
.B(n_448),
.C(n_418),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_646),
.A2(n_429),
.B(n_416),
.Y(n_901)
);

A2O1A1Ixp33_ASAP7_75t_L g902 ( 
.A1(n_654),
.A2(n_429),
.B(n_418),
.C(n_435),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_736),
.B(n_527),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_635),
.B(n_417),
.Y(n_904)
);

INVx2_ASAP7_75t_L g905 ( 
.A(n_659),
.Y(n_905)
);

AND2x2_ASAP7_75t_L g906 ( 
.A(n_772),
.B(n_425),
.Y(n_906)
);

BUFx6f_ASAP7_75t_L g907 ( 
.A(n_679),
.Y(n_907)
);

AOI21xp5_ASAP7_75t_L g908 ( 
.A1(n_666),
.A2(n_429),
.B(n_416),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_760),
.A2(n_431),
.B(n_418),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_647),
.Y(n_910)
);

OAI22xp5_ASAP7_75t_L g911 ( 
.A1(n_677),
.A2(n_431),
.B1(n_413),
.B2(n_418),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_738),
.B(n_426),
.Y(n_912)
);

OAI21xp5_ASAP7_75t_L g913 ( 
.A1(n_671),
.A2(n_688),
.B(n_705),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_748),
.B(n_426),
.Y(n_914)
);

AOI33xp33_ASAP7_75t_L g915 ( 
.A1(n_768),
.A2(n_452),
.A3(n_428),
.B1(n_429),
.B2(n_435),
.B3(n_413),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_L g916 ( 
.A(n_667),
.B(n_428),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_659),
.Y(n_917)
);

AOI21xp33_ASAP7_75t_L g918 ( 
.A1(n_667),
.A2(n_413),
.B(n_429),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_685),
.Y(n_919)
);

AOI22xp5_ASAP7_75t_L g920 ( 
.A1(n_647),
.A2(n_560),
.B1(n_448),
.B2(n_445),
.Y(n_920)
);

AOI21xp5_ASAP7_75t_L g921 ( 
.A1(n_760),
.A2(n_436),
.B(n_448),
.Y(n_921)
);

OAI21xp5_ASAP7_75t_L g922 ( 
.A1(n_671),
.A2(n_560),
.B(n_448),
.Y(n_922)
);

INVx3_ASAP7_75t_L g923 ( 
.A(n_732),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_688),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_760),
.A2(n_435),
.B(n_445),
.Y(n_925)
);

BUFx2_ASAP7_75t_L g926 ( 
.A(n_647),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_L g927 ( 
.A(n_685),
.B(n_435),
.Y(n_927)
);

AOI21xp5_ASAP7_75t_L g928 ( 
.A1(n_760),
.A2(n_435),
.B(n_445),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_689),
.B(n_436),
.Y(n_929)
);

AOI21xp5_ASAP7_75t_L g930 ( 
.A1(n_750),
.A2(n_436),
.B(n_445),
.Y(n_930)
);

INVx2_ASAP7_75t_L g931 ( 
.A(n_689),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_692),
.B(n_436),
.Y(n_932)
);

AOI21xp5_ASAP7_75t_L g933 ( 
.A1(n_750),
.A2(n_436),
.B(n_445),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_692),
.B(n_413),
.Y(n_934)
);

INVx2_ASAP7_75t_L g935 ( 
.A(n_699),
.Y(n_935)
);

AOI21xp5_ASAP7_75t_L g936 ( 
.A1(n_765),
.A2(n_444),
.B(n_438),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_765),
.A2(n_444),
.B(n_438),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_699),
.B(n_444),
.Y(n_938)
);

BUFx5_ASAP7_75t_L g939 ( 
.A(n_687),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_703),
.Y(n_940)
);

O2A1O1Ixp33_ASAP7_75t_L g941 ( 
.A1(n_670),
.A2(n_12),
.B(n_15),
.C(n_17),
.Y(n_941)
);

A2O1A1Ixp33_ASAP7_75t_L g942 ( 
.A1(n_730),
.A2(n_417),
.B(n_421),
.C(n_423),
.Y(n_942)
);

NAND2x1p5_ASAP7_75t_L g943 ( 
.A(n_732),
.B(n_417),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_647),
.B(n_732),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_670),
.A2(n_723),
.B(n_673),
.C(n_684),
.Y(n_945)
);

OAI21xp5_ASAP7_75t_L g946 ( 
.A1(n_696),
.A2(n_560),
.B(n_444),
.Y(n_946)
);

OAI21xp5_ASAP7_75t_L g947 ( 
.A1(n_701),
.A2(n_560),
.B(n_444),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_758),
.A2(n_444),
.B(n_438),
.Y(n_948)
);

OR2x6_ASAP7_75t_L g949 ( 
.A(n_740),
.B(n_417),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_703),
.B(n_444),
.Y(n_950)
);

BUFx2_ASAP7_75t_L g951 ( 
.A(n_687),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_706),
.B(n_444),
.Y(n_952)
);

NAND2x1_ASAP7_75t_L g953 ( 
.A(n_721),
.B(n_560),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_706),
.B(n_444),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_714),
.B(n_444),
.Y(n_955)
);

BUFx5_ASAP7_75t_L g956 ( 
.A(n_687),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_767),
.A2(n_438),
.B(n_423),
.Y(n_957)
);

AND2x2_ASAP7_75t_L g958 ( 
.A(n_673),
.B(n_17),
.Y(n_958)
);

NOR2xp33_ASAP7_75t_L g959 ( 
.A(n_661),
.B(n_19),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_714),
.B(n_717),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_769),
.A2(n_438),
.B(n_423),
.Y(n_961)
);

AND2x2_ASAP7_75t_L g962 ( 
.A(n_684),
.B(n_24),
.Y(n_962)
);

OA22x2_ASAP7_75t_L g963 ( 
.A1(n_707),
.A2(n_24),
.B1(n_25),
.B2(n_29),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_813),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_SL g965 ( 
.A(n_797),
.B(n_718),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_818),
.B(n_717),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_905),
.Y(n_967)
);

AOI21xp5_ASAP7_75t_L g968 ( 
.A1(n_782),
.A2(n_740),
.B(n_756),
.Y(n_968)
);

OR2x6_ASAP7_75t_L g969 ( 
.A(n_894),
.B(n_926),
.Y(n_969)
);

AOI21xp5_ASAP7_75t_L g970 ( 
.A1(n_785),
.A2(n_799),
.B(n_775),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_SL g971 ( 
.A(n_791),
.B(n_718),
.Y(n_971)
);

INVx3_ASAP7_75t_L g972 ( 
.A(n_826),
.Y(n_972)
);

O2A1O1Ixp33_ASAP7_75t_L g973 ( 
.A1(n_783),
.A2(n_661),
.B(n_662),
.C(n_723),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_SL g974 ( 
.A(n_792),
.B(n_770),
.Y(n_974)
);

NAND3xp33_ASAP7_75t_SL g975 ( 
.A(n_865),
.B(n_728),
.C(n_676),
.Y(n_975)
);

INVx1_ASAP7_75t_L g976 ( 
.A(n_789),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_795),
.A2(n_740),
.B(n_756),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_L g978 ( 
.A1(n_874),
.A2(n_728),
.B(n_707),
.C(n_662),
.Y(n_978)
);

HB1xp67_ASAP7_75t_L g979 ( 
.A(n_809),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_779),
.A2(n_735),
.B(n_708),
.C(n_709),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_776),
.B(n_720),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_792),
.B(n_884),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_813),
.Y(n_983)
);

OAI22x1_ASAP7_75t_L g984 ( 
.A1(n_885),
.A2(n_633),
.B1(n_752),
.B2(n_747),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_811),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_817),
.Y(n_986)
);

AOI22xp5_ASAP7_75t_L g987 ( 
.A1(n_886),
.A2(n_687),
.B1(n_681),
.B2(n_712),
.Y(n_987)
);

BUFx6f_ASAP7_75t_L g988 ( 
.A(n_813),
.Y(n_988)
);

OAI22xp5_ASAP7_75t_L g989 ( 
.A1(n_796),
.A2(n_740),
.B1(n_713),
.B2(n_739),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_L g990 ( 
.A1(n_889),
.A2(n_879),
.B(n_843),
.C(n_816),
.Y(n_990)
);

INVxp67_ASAP7_75t_L g991 ( 
.A(n_847),
.Y(n_991)
);

AOI21xp5_ASAP7_75t_L g992 ( 
.A1(n_800),
.A2(n_737),
.B(n_746),
.Y(n_992)
);

INVx4_ASAP7_75t_L g993 ( 
.A(n_856),
.Y(n_993)
);

OAI22xp33_ASAP7_75t_L g994 ( 
.A1(n_891),
.A2(n_770),
.B1(n_752),
.B2(n_747),
.Y(n_994)
);

NOR2xp33_ASAP7_75t_L g995 ( 
.A(n_828),
.B(n_743),
.Y(n_995)
);

NOR3xp33_ASAP7_75t_L g996 ( 
.A(n_869),
.B(n_681),
.C(n_741),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_860),
.Y(n_997)
);

INVx2_ASAP7_75t_L g998 ( 
.A(n_917),
.Y(n_998)
);

HB1xp67_ASAP7_75t_L g999 ( 
.A(n_830),
.Y(n_999)
);

OAI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_796),
.A2(n_743),
.B1(n_741),
.B2(n_734),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_856),
.Y(n_1001)
);

BUFx3_ASAP7_75t_L g1002 ( 
.A(n_864),
.Y(n_1002)
);

OAI22x1_ASAP7_75t_L g1003 ( 
.A1(n_824),
.A2(n_633),
.B1(n_721),
.B2(n_734),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_898),
.A2(n_633),
.B1(n_687),
.B2(n_438),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_846),
.B(n_875),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_910),
.B(n_687),
.Y(n_1006)
);

NAND2xp5_ASAP7_75t_L g1007 ( 
.A(n_895),
.B(n_560),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_823),
.B(n_25),
.Y(n_1008)
);

OAI22xp5_ASAP7_75t_L g1009 ( 
.A1(n_924),
.A2(n_881),
.B1(n_835),
.B2(n_892),
.Y(n_1009)
);

NOR2xp33_ASAP7_75t_L g1010 ( 
.A(n_854),
.B(n_31),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_822),
.Y(n_1011)
);

NAND2xp5_ASAP7_75t_L g1012 ( 
.A(n_836),
.B(n_560),
.Y(n_1012)
);

INVx4_ASAP7_75t_SL g1013 ( 
.A(n_856),
.Y(n_1013)
);

HB1xp67_ASAP7_75t_L g1014 ( 
.A(n_852),
.Y(n_1014)
);

OR2x6_ASAP7_75t_L g1015 ( 
.A(n_892),
.B(n_438),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_832),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_866),
.A2(n_438),
.B(n_423),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_831),
.A2(n_438),
.B(n_423),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_852),
.B(n_438),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_838),
.Y(n_1020)
);

NAND2xp5_ASAP7_75t_SL g1021 ( 
.A(n_878),
.B(n_423),
.Y(n_1021)
);

A2O1A1Ixp33_ASAP7_75t_L g1022 ( 
.A1(n_868),
.A2(n_423),
.B(n_421),
.C(n_417),
.Y(n_1022)
);

OR2x2_ASAP7_75t_L g1023 ( 
.A(n_862),
.B(n_31),
.Y(n_1023)
);

OAI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_959),
.A2(n_423),
.B1(n_421),
.B2(n_417),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_819),
.B(n_821),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_798),
.A2(n_423),
.B(n_421),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_SL g1027 ( 
.A(n_777),
.Y(n_1027)
);

AOI21xp5_ASAP7_75t_L g1028 ( 
.A1(n_810),
.A2(n_423),
.B(n_421),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_SL g1029 ( 
.A(n_843),
.B(n_33),
.C(n_35),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_870),
.A2(n_421),
.B(n_417),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_851),
.B(n_421),
.Y(n_1031)
);

BUFx6f_ASAP7_75t_L g1032 ( 
.A(n_896),
.Y(n_1032)
);

CKINVDCx16_ASAP7_75t_R g1033 ( 
.A(n_906),
.Y(n_1033)
);

INVx2_ASAP7_75t_L g1034 ( 
.A(n_919),
.Y(n_1034)
);

OAI22xp5_ASAP7_75t_L g1035 ( 
.A1(n_963),
.A2(n_421),
.B1(n_417),
.B2(n_37),
.Y(n_1035)
);

BUFx6f_ASAP7_75t_L g1036 ( 
.A(n_896),
.Y(n_1036)
);

NOR3xp33_ASAP7_75t_L g1037 ( 
.A(n_842),
.B(n_33),
.C(n_35),
.Y(n_1037)
);

NOR2xp67_ASAP7_75t_L g1038 ( 
.A(n_873),
.B(n_85),
.Y(n_1038)
);

OR2x2_ASAP7_75t_L g1039 ( 
.A(n_825),
.B(n_37),
.Y(n_1039)
);

BUFx10_ASAP7_75t_L g1040 ( 
.A(n_804),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_931),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_787),
.B(n_40),
.Y(n_1042)
);

AOI21xp5_ASAP7_75t_L g1043 ( 
.A1(n_790),
.A2(n_820),
.B(n_913),
.Y(n_1043)
);

BUFx2_ASAP7_75t_L g1044 ( 
.A(n_958),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_935),
.Y(n_1045)
);

AND2x4_ASAP7_75t_L g1046 ( 
.A(n_777),
.B(n_95),
.Y(n_1046)
);

INVx2_ASAP7_75t_L g1047 ( 
.A(n_851),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_876),
.B(n_421),
.Y(n_1048)
);

NAND2xp5_ASAP7_75t_L g1049 ( 
.A(n_803),
.B(n_421),
.Y(n_1049)
);

OAI21xp5_ASAP7_75t_L g1050 ( 
.A1(n_945),
.A2(n_417),
.B(n_68),
.Y(n_1050)
);

AOI21xp5_ASAP7_75t_L g1051 ( 
.A1(n_913),
.A2(n_64),
.B(n_150),
.Y(n_1051)
);

BUFx6f_ASAP7_75t_L g1052 ( 
.A(n_896),
.Y(n_1052)
);

NOR2xp33_ASAP7_75t_L g1053 ( 
.A(n_855),
.B(n_801),
.Y(n_1053)
);

O2A1O1Ixp33_ASAP7_75t_L g1054 ( 
.A1(n_941),
.A2(n_41),
.B(n_44),
.C(n_45),
.Y(n_1054)
);

BUFx2_ASAP7_75t_L g1055 ( 
.A(n_962),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_803),
.B(n_44),
.Y(n_1056)
);

AOI21xp5_ASAP7_75t_L g1057 ( 
.A1(n_897),
.A2(n_97),
.B(n_139),
.Y(n_1057)
);

AOI21xp5_ASAP7_75t_L g1058 ( 
.A1(n_904),
.A2(n_802),
.B(n_882),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_949),
.A2(n_61),
.B(n_137),
.Y(n_1059)
);

INVx2_ASAP7_75t_L g1060 ( 
.A(n_940),
.Y(n_1060)
);

AOI21xp5_ASAP7_75t_L g1061 ( 
.A1(n_949),
.A2(n_152),
.B(n_126),
.Y(n_1061)
);

OR2x2_ASAP7_75t_L g1062 ( 
.A(n_850),
.B(n_45),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_807),
.B(n_125),
.Y(n_1063)
);

OR2x2_ASAP7_75t_L g1064 ( 
.A(n_807),
.B(n_46),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_949),
.A2(n_105),
.B(n_114),
.Y(n_1065)
);

OAI22xp5_ASAP7_75t_L g1066 ( 
.A1(n_963),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1066)
);

AO32x1_ASAP7_75t_L g1067 ( 
.A1(n_911),
.A2(n_49),
.A3(n_51),
.B1(n_880),
.B2(n_827),
.Y(n_1067)
);

BUFx6f_ASAP7_75t_L g1068 ( 
.A(n_907),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_907),
.Y(n_1069)
);

AND2x2_ASAP7_75t_L g1070 ( 
.A(n_786),
.B(n_778),
.Y(n_1070)
);

INVxp67_ASAP7_75t_L g1071 ( 
.A(n_887),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_L g1072 ( 
.A(n_944),
.B(n_786),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_915),
.Y(n_1073)
);

INVxp67_ASAP7_75t_SL g1074 ( 
.A(n_907),
.Y(n_1074)
);

INVxp67_ASAP7_75t_L g1075 ( 
.A(n_780),
.Y(n_1075)
);

NAND2xp5_ASAP7_75t_L g1076 ( 
.A(n_826),
.B(n_839),
.Y(n_1076)
);

AND3x2_ASAP7_75t_L g1077 ( 
.A(n_951),
.B(n_839),
.C(n_780),
.Y(n_1077)
);

AND2x4_ASAP7_75t_SL g1078 ( 
.A(n_848),
.B(n_923),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_923),
.B(n_848),
.Y(n_1079)
);

CKINVDCx5p33_ASAP7_75t_R g1080 ( 
.A(n_863),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_814),
.A2(n_853),
.B(n_805),
.Y(n_1081)
);

INVx2_ASAP7_75t_L g1082 ( 
.A(n_960),
.Y(n_1082)
);

NOR2xp33_ASAP7_75t_L g1083 ( 
.A(n_784),
.B(n_793),
.Y(n_1083)
);

NAND2xp5_ASAP7_75t_L g1084 ( 
.A(n_778),
.B(n_781),
.Y(n_1084)
);

NAND2xp5_ASAP7_75t_SL g1085 ( 
.A(n_784),
.B(n_939),
.Y(n_1085)
);

A2O1A1Ixp33_ASAP7_75t_L g1086 ( 
.A1(n_812),
.A2(n_781),
.B(n_794),
.C(n_899),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_912),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_794),
.B(n_914),
.Y(n_1088)
);

O2A1O1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_827),
.A2(n_900),
.B(n_942),
.C(n_841),
.Y(n_1089)
);

A2O1A1Ixp33_ASAP7_75t_L g1090 ( 
.A1(n_859),
.A2(n_872),
.B(n_861),
.C(n_903),
.Y(n_1090)
);

HB1xp67_ASAP7_75t_L g1091 ( 
.A(n_916),
.Y(n_1091)
);

NOR2xp33_ASAP7_75t_L g1092 ( 
.A(n_841),
.B(n_788),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_927),
.Y(n_1093)
);

AOI22xp33_ASAP7_75t_L g1094 ( 
.A1(n_829),
.A2(n_922),
.B1(n_956),
.B2(n_939),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_SL g1095 ( 
.A1(n_953),
.A2(n_853),
.B1(n_920),
.B2(n_922),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_SL g1096 ( 
.A(n_939),
.B(n_956),
.Y(n_1096)
);

AOI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_805),
.A2(n_806),
.B(n_908),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_929),
.B(n_932),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_934),
.Y(n_1099)
);

OAI22xp33_ASAP7_75t_L g1100 ( 
.A1(n_946),
.A2(n_947),
.B1(n_954),
.B2(n_955),
.Y(n_1100)
);

CKINVDCx5p33_ASAP7_75t_R g1101 ( 
.A(n_939),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_SL g1102 ( 
.A(n_939),
.B(n_956),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_833),
.A2(n_840),
.B(n_845),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_857),
.B(n_858),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_844),
.A2(n_849),
.B(n_871),
.Y(n_1105)
);

INVx2_ASAP7_75t_L g1106 ( 
.A(n_815),
.Y(n_1106)
);

INVx1_ASAP7_75t_SL g1107 ( 
.A(n_938),
.Y(n_1107)
);

NOR2xp33_ASAP7_75t_L g1108 ( 
.A(n_950),
.B(n_952),
.Y(n_1108)
);

AND2x2_ASAP7_75t_L g1109 ( 
.A(n_849),
.B(n_902),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_943),
.Y(n_1110)
);

HB1xp67_ASAP7_75t_L g1111 ( 
.A(n_943),
.Y(n_1111)
);

OAI21x1_ASAP7_75t_L g1112 ( 
.A1(n_970),
.A2(n_808),
.B(n_877),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1097),
.A2(n_867),
.B(n_837),
.Y(n_1113)
);

AOI22xp5_ASAP7_75t_L g1114 ( 
.A1(n_1080),
.A2(n_939),
.B1(n_956),
.B2(n_880),
.Y(n_1114)
);

OAI21x1_ASAP7_75t_L g1115 ( 
.A1(n_1103),
.A2(n_890),
.B(n_883),
.Y(n_1115)
);

CKINVDCx5p33_ASAP7_75t_R g1116 ( 
.A(n_1033),
.Y(n_1116)
);

NOR2xp33_ASAP7_75t_L g1117 ( 
.A(n_982),
.B(n_918),
.Y(n_1117)
);

OAI22xp5_ASAP7_75t_L g1118 ( 
.A1(n_1075),
.A2(n_947),
.B1(n_946),
.B2(n_834),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_1005),
.Y(n_1119)
);

INVx2_ASAP7_75t_SL g1120 ( 
.A(n_979),
.Y(n_1120)
);

BUFx6f_ASAP7_75t_L g1121 ( 
.A(n_964),
.Y(n_1121)
);

AO31x2_ASAP7_75t_L g1122 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_989),
.B(n_1083),
.Y(n_1122)
);

A2O1A1Ixp33_ASAP7_75t_L g1123 ( 
.A1(n_990),
.A2(n_893),
.B(n_901),
.C(n_936),
.Y(n_1123)
);

OAI22xp5_ASAP7_75t_L g1124 ( 
.A1(n_1044),
.A2(n_930),
.B1(n_933),
.B2(n_961),
.Y(n_1124)
);

NAND2xp5_ASAP7_75t_L g1125 ( 
.A(n_995),
.B(n_957),
.Y(n_1125)
);

OR2x6_ASAP7_75t_L g1126 ( 
.A(n_969),
.B(n_888),
.Y(n_1126)
);

INVx2_ASAP7_75t_L g1127 ( 
.A(n_1060),
.Y(n_1127)
);

INVxp67_ASAP7_75t_L g1128 ( 
.A(n_999),
.Y(n_1128)
);

BUFx12f_ASAP7_75t_L g1129 ( 
.A(n_1040),
.Y(n_1129)
);

AND2x2_ASAP7_75t_L g1130 ( 
.A(n_1055),
.B(n_918),
.Y(n_1130)
);

AO32x2_ASAP7_75t_L g1131 ( 
.A1(n_1035),
.A2(n_911),
.A3(n_937),
.B1(n_956),
.B2(n_948),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_1025),
.B(n_956),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_981),
.A2(n_968),
.B(n_1043),
.Y(n_1133)
);

AO21x2_ASAP7_75t_L g1134 ( 
.A1(n_1050),
.A2(n_909),
.B(n_921),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_976),
.Y(n_1135)
);

INVx5_ASAP7_75t_L g1136 ( 
.A(n_964),
.Y(n_1136)
);

AO32x2_ASAP7_75t_L g1137 ( 
.A1(n_1035),
.A2(n_925),
.A3(n_928),
.B1(n_1066),
.B2(n_1004),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_SL g1138 ( 
.A(n_1010),
.B(n_1014),
.Y(n_1138)
);

OAI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1072),
.A2(n_1050),
.B(n_978),
.Y(n_1139)
);

BUFx6f_ASAP7_75t_L g1140 ( 
.A(n_964),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_977),
.A2(n_1105),
.B(n_1081),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_966),
.A2(n_1104),
.B(n_1084),
.Y(n_1142)
);

NOR2xp33_ASAP7_75t_L g1143 ( 
.A(n_991),
.B(n_1053),
.Y(n_1143)
);

AND2x2_ASAP7_75t_L g1144 ( 
.A(n_1023),
.B(n_1039),
.Y(n_1144)
);

NOR2xp33_ASAP7_75t_L g1145 ( 
.A(n_971),
.B(n_1076),
.Y(n_1145)
);

INVx4_ASAP7_75t_L g1146 ( 
.A(n_1069),
.Y(n_1146)
);

AOI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1058),
.A2(n_992),
.B(n_1085),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_1087),
.B(n_1070),
.Y(n_1148)
);

BUFx2_ASAP7_75t_L g1149 ( 
.A(n_997),
.Y(n_1149)
);

OAI21xp33_ASAP7_75t_L g1150 ( 
.A1(n_1008),
.A2(n_1029),
.B(n_1037),
.Y(n_1150)
);

A2O1A1Ixp33_ASAP7_75t_L g1151 ( 
.A1(n_1038),
.A2(n_987),
.B(n_975),
.C(n_973),
.Y(n_1151)
);

A2O1A1Ixp33_ASAP7_75t_L g1152 ( 
.A1(n_1051),
.A2(n_980),
.B(n_1054),
.C(n_1071),
.Y(n_1152)
);

OAI22xp5_ASAP7_75t_L g1153 ( 
.A1(n_1101),
.A2(n_1094),
.B1(n_1086),
.B2(n_972),
.Y(n_1153)
);

AO32x2_ASAP7_75t_L g1154 ( 
.A1(n_1066),
.A2(n_1095),
.A3(n_1009),
.B1(n_1000),
.B2(n_1067),
.Y(n_1154)
);

INVx2_ASAP7_75t_L g1155 ( 
.A(n_967),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_985),
.Y(n_1156)
);

BUFx4f_ASAP7_75t_SL g1157 ( 
.A(n_1002),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_986),
.Y(n_1158)
);

NOR4xp25_ASAP7_75t_L g1159 ( 
.A(n_1042),
.B(n_1089),
.C(n_965),
.D(n_1056),
.Y(n_1159)
);

BUFx6f_ASAP7_75t_L g1160 ( 
.A(n_983),
.Y(n_1160)
);

OAI21x1_ASAP7_75t_L g1161 ( 
.A1(n_1106),
.A2(n_1096),
.B(n_1102),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_1064),
.Y(n_1162)
);

O2A1O1Ixp33_ASAP7_75t_SL g1163 ( 
.A1(n_1073),
.A2(n_1012),
.B(n_1021),
.C(n_1022),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1088),
.A2(n_1098),
.B(n_1108),
.Y(n_1164)
);

O2A1O1Ixp33_ASAP7_75t_L g1165 ( 
.A1(n_1062),
.A2(n_974),
.B(n_996),
.C(n_994),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1011),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_1091),
.B(n_972),
.Y(n_1167)
);

NOR2x1_ASAP7_75t_L g1168 ( 
.A(n_993),
.B(n_969),
.Y(n_1168)
);

OAI21xp5_ASAP7_75t_L g1169 ( 
.A1(n_1092),
.A2(n_1109),
.B(n_1090),
.Y(n_1169)
);

BUFx12f_ASAP7_75t_L g1170 ( 
.A(n_1040),
.Y(n_1170)
);

OAI22x1_ASAP7_75t_L g1171 ( 
.A1(n_1016),
.A2(n_1020),
.B1(n_1063),
.B2(n_1046),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_SL g1172 ( 
.A1(n_1079),
.A2(n_1007),
.B(n_1019),
.C(n_1100),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_1000),
.Y(n_1173)
);

AO31x2_ASAP7_75t_L g1174 ( 
.A1(n_984),
.A2(n_1024),
.A3(n_1018),
.B(n_1030),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1095),
.A2(n_1093),
.B(n_1099),
.Y(n_1175)
);

BUFx10_ASAP7_75t_L g1176 ( 
.A(n_1027),
.Y(n_1176)
);

AO31x2_ASAP7_75t_L g1177 ( 
.A1(n_1024),
.A2(n_1028),
.A3(n_1017),
.B(n_1026),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_998),
.Y(n_1178)
);

INVxp67_ASAP7_75t_L g1179 ( 
.A(n_969),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1048),
.A2(n_1049),
.B(n_1031),
.Y(n_1180)
);

BUFx6f_ASAP7_75t_L g1181 ( 
.A(n_983),
.Y(n_1181)
);

NOR2xp33_ASAP7_75t_SL g1182 ( 
.A(n_1027),
.B(n_993),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1107),
.A2(n_1015),
.B(n_1065),
.Y(n_1183)
);

AOI22xp5_ASAP7_75t_L g1184 ( 
.A1(n_1063),
.A2(n_1046),
.B1(n_1077),
.B2(n_1082),
.Y(n_1184)
);

A2O1A1Ixp33_ASAP7_75t_L g1185 ( 
.A1(n_1059),
.A2(n_1061),
.B(n_1057),
.C(n_1034),
.Y(n_1185)
);

AO31x2_ASAP7_75t_L g1186 ( 
.A1(n_1067),
.A2(n_1047),
.A3(n_1045),
.B(n_1041),
.Y(n_1186)
);

INVx1_ASAP7_75t_SL g1187 ( 
.A(n_983),
.Y(n_1187)
);

O2A1O1Ixp33_ASAP7_75t_L g1188 ( 
.A1(n_1107),
.A2(n_1111),
.B(n_1074),
.C(n_1015),
.Y(n_1188)
);

AOI22xp5_ASAP7_75t_L g1189 ( 
.A1(n_1078),
.A2(n_1110),
.B1(n_1001),
.B2(n_1036),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1013),
.Y(n_1190)
);

INVxp67_ASAP7_75t_SL g1191 ( 
.A(n_988),
.Y(n_1191)
);

AOI22xp33_ASAP7_75t_L g1192 ( 
.A1(n_1006),
.A2(n_1110),
.B1(n_1001),
.B2(n_1052),
.Y(n_1192)
);

INVx2_ASAP7_75t_L g1193 ( 
.A(n_1110),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_1015),
.A2(n_1067),
.B(n_1001),
.Y(n_1194)
);

AOI221xp5_ASAP7_75t_L g1195 ( 
.A1(n_988),
.A2(n_1068),
.B1(n_1032),
.B2(n_1036),
.C(n_1052),
.Y(n_1195)
);

AO32x2_ASAP7_75t_L g1196 ( 
.A1(n_1013),
.A2(n_988),
.A3(n_1032),
.B1(n_1036),
.B2(n_1052),
.Y(n_1196)
);

BUFx2_ASAP7_75t_L g1197 ( 
.A(n_1032),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1068),
.B(n_1013),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_1068),
.Y(n_1199)
);

AOI21xp5_ASAP7_75t_L g1200 ( 
.A1(n_970),
.A2(n_537),
.B(n_1097),
.Y(n_1200)
);

OAI21x1_ASAP7_75t_L g1201 ( 
.A1(n_970),
.A2(n_808),
.B(n_1103),
.Y(n_1201)
);

OAI22xp5_ASAP7_75t_L g1202 ( 
.A1(n_982),
.A2(n_652),
.B1(n_537),
.B2(n_797),
.Y(n_1202)
);

OAI21x1_ASAP7_75t_SL g1203 ( 
.A1(n_1050),
.A2(n_1051),
.B(n_1066),
.Y(n_1203)
);

AO31x2_ASAP7_75t_L g1204 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_989),
.B(n_1083),
.Y(n_1204)
);

O2A1O1Ixp33_ASAP7_75t_SL g1205 ( 
.A1(n_978),
.A2(n_889),
.B(n_1085),
.C(n_1050),
.Y(n_1205)
);

OA21x2_ASAP7_75t_L g1206 ( 
.A1(n_1050),
.A2(n_1081),
.B(n_1097),
.Y(n_1206)
);

NOR2xp33_ASAP7_75t_L g1207 ( 
.A(n_982),
.B(n_652),
.Y(n_1207)
);

O2A1O1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_990),
.A2(n_779),
.B(n_818),
.C(n_630),
.Y(n_1208)
);

NAND2xp5_ASAP7_75t_L g1209 ( 
.A(n_982),
.B(n_630),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1075),
.A2(n_630),
.B(n_644),
.Y(n_1210)
);

AND2x2_ASAP7_75t_L g1211 ( 
.A(n_1044),
.B(n_660),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_982),
.B(n_630),
.Y(n_1212)
);

NOR2xp67_ASAP7_75t_SL g1213 ( 
.A(n_979),
.B(n_613),
.Y(n_1213)
);

AOI21xp5_ASAP7_75t_L g1214 ( 
.A1(n_970),
.A2(n_537),
.B(n_1097),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_1005),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_989),
.B(n_1083),
.Y(n_1216)
);

OAI21x1_ASAP7_75t_L g1217 ( 
.A1(n_970),
.A2(n_808),
.B(n_1103),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_970),
.A2(n_808),
.B(n_1103),
.Y(n_1218)
);

OAI21x1_ASAP7_75t_L g1219 ( 
.A1(n_970),
.A2(n_808),
.B(n_1103),
.Y(n_1219)
);

AOI21xp5_ASAP7_75t_L g1220 ( 
.A1(n_970),
.A2(n_537),
.B(n_1097),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_982),
.B(n_630),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1073),
.Y(n_1222)
);

INVx1_ASAP7_75t_L g1223 ( 
.A(n_1073),
.Y(n_1223)
);

BUFx3_ASAP7_75t_L g1224 ( 
.A(n_997),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1005),
.Y(n_1225)
);

NAND2xp5_ASAP7_75t_L g1226 ( 
.A(n_982),
.B(n_630),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_990),
.A2(n_630),
.B(n_1050),
.C(n_818),
.Y(n_1227)
);

OAI21x1_ASAP7_75t_L g1228 ( 
.A1(n_970),
.A2(n_808),
.B(n_1103),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_SL g1229 ( 
.A1(n_978),
.A2(n_889),
.B(n_1085),
.C(n_1050),
.Y(n_1229)
);

BUFx2_ASAP7_75t_L g1230 ( 
.A(n_1069),
.Y(n_1230)
);

AO31x2_ASAP7_75t_L g1231 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_989),
.B(n_1083),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_1005),
.Y(n_1232)
);

INVx1_ASAP7_75t_L g1233 ( 
.A(n_1005),
.Y(n_1233)
);

NAND2xp5_ASAP7_75t_SL g1234 ( 
.A(n_982),
.B(n_652),
.Y(n_1234)
);

AO31x2_ASAP7_75t_L g1235 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_989),
.B(n_1083),
.Y(n_1235)
);

NAND2x1_ASAP7_75t_L g1236 ( 
.A(n_993),
.B(n_777),
.Y(n_1236)
);

AOI21xp5_ASAP7_75t_L g1237 ( 
.A1(n_970),
.A2(n_537),
.B(n_1097),
.Y(n_1237)
);

NAND2xp5_ASAP7_75t_L g1238 ( 
.A(n_982),
.B(n_630),
.Y(n_1238)
);

NOR2xp33_ASAP7_75t_L g1239 ( 
.A(n_982),
.B(n_652),
.Y(n_1239)
);

AOI22xp33_ASAP7_75t_L g1240 ( 
.A1(n_1010),
.A2(n_865),
.B1(n_874),
.B2(n_818),
.Y(n_1240)
);

NAND2xp5_ASAP7_75t_SL g1241 ( 
.A(n_982),
.B(n_652),
.Y(n_1241)
);

AOI21xp5_ASAP7_75t_L g1242 ( 
.A1(n_970),
.A2(n_537),
.B(n_1097),
.Y(n_1242)
);

INVx2_ASAP7_75t_L g1243 ( 
.A(n_1060),
.Y(n_1243)
);

INVx1_ASAP7_75t_L g1244 ( 
.A(n_1005),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1050),
.A2(n_1081),
.B(n_1097),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_982),
.B(n_630),
.Y(n_1246)
);

AO21x1_ASAP7_75t_L g1247 ( 
.A1(n_1050),
.A2(n_1035),
.B(n_990),
.Y(n_1247)
);

BUFx2_ASAP7_75t_L g1248 ( 
.A(n_1069),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_970),
.A2(n_537),
.B(n_1097),
.Y(n_1249)
);

O2A1O1Ixp5_ASAP7_75t_SL g1250 ( 
.A1(n_1050),
.A2(n_643),
.B(n_783),
.C(n_965),
.Y(n_1250)
);

OR2x2_ASAP7_75t_L g1251 ( 
.A(n_1025),
.B(n_982),
.Y(n_1251)
);

AO31x2_ASAP7_75t_L g1252 ( 
.A1(n_1003),
.A2(n_1004),
.A3(n_989),
.B(n_1083),
.Y(n_1252)
);

O2A1O1Ixp33_ASAP7_75t_SL g1253 ( 
.A1(n_978),
.A2(n_889),
.B(n_1085),
.C(n_1050),
.Y(n_1253)
);

OAI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1075),
.A2(n_630),
.B(n_644),
.Y(n_1254)
);

OAI21x1_ASAP7_75t_L g1255 ( 
.A1(n_970),
.A2(n_808),
.B(n_1103),
.Y(n_1255)
);

CKINVDCx11_ASAP7_75t_R g1256 ( 
.A(n_1040),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1073),
.Y(n_1257)
);

BUFx2_ASAP7_75t_R g1258 ( 
.A(n_997),
.Y(n_1258)
);

AOI221xp5_ASAP7_75t_L g1259 ( 
.A1(n_1010),
.A2(n_874),
.B1(n_545),
.B2(n_518),
.C(n_757),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_1247),
.Y(n_1260)
);

BUFx12f_ASAP7_75t_L g1261 ( 
.A(n_1256),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1210),
.A2(n_1254),
.B1(n_1139),
.B2(n_1203),
.Y(n_1262)
);

BUFx12f_ASAP7_75t_L g1263 ( 
.A(n_1176),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1135),
.Y(n_1264)
);

HB1xp67_ASAP7_75t_L g1265 ( 
.A(n_1169),
.Y(n_1265)
);

CKINVDCx20_ASAP7_75t_R g1266 ( 
.A(n_1157),
.Y(n_1266)
);

AOI22xp33_ASAP7_75t_L g1267 ( 
.A1(n_1209),
.A2(n_1238),
.B1(n_1226),
.B2(n_1221),
.Y(n_1267)
);

OAI22xp33_ASAP7_75t_L g1268 ( 
.A1(n_1212),
.A2(n_1246),
.B1(n_1251),
.B2(n_1225),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_1207),
.B(n_1239),
.Y(n_1269)
);

AOI22xp33_ASAP7_75t_SL g1270 ( 
.A1(n_1206),
.A2(n_1245),
.B1(n_1153),
.B2(n_1202),
.Y(n_1270)
);

AOI22xp33_ASAP7_75t_L g1271 ( 
.A1(n_1144),
.A2(n_1233),
.B1(n_1232),
.B2(n_1244),
.Y(n_1271)
);

INVx3_ASAP7_75t_SL g1272 ( 
.A(n_1199),
.Y(n_1272)
);

CKINVDCx11_ASAP7_75t_R g1273 ( 
.A(n_1176),
.Y(n_1273)
);

BUFx3_ASAP7_75t_L g1274 ( 
.A(n_1224),
.Y(n_1274)
);

AND2x2_ASAP7_75t_L g1275 ( 
.A(n_1211),
.B(n_1162),
.Y(n_1275)
);

OAI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1119),
.A2(n_1215),
.B1(n_1148),
.B2(n_1184),
.Y(n_1276)
);

BUFx12f_ASAP7_75t_L g1277 ( 
.A(n_1116),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1206),
.A2(n_1245),
.B1(n_1143),
.B2(n_1227),
.Y(n_1278)
);

INVx3_ASAP7_75t_L g1279 ( 
.A(n_1121),
.Y(n_1279)
);

OAI22xp33_ASAP7_75t_L g1280 ( 
.A1(n_1222),
.A2(n_1223),
.B1(n_1257),
.B2(n_1175),
.Y(n_1280)
);

AOI22x1_ASAP7_75t_L g1281 ( 
.A1(n_1171),
.A2(n_1164),
.B1(n_1183),
.B2(n_1147),
.Y(n_1281)
);

CKINVDCx11_ASAP7_75t_R g1282 ( 
.A(n_1129),
.Y(n_1282)
);

BUFx2_ASAP7_75t_L g1283 ( 
.A(n_1230),
.Y(n_1283)
);

CKINVDCx16_ASAP7_75t_R g1284 ( 
.A(n_1170),
.Y(n_1284)
);

INVx1_ASAP7_75t_SL g1285 ( 
.A(n_1258),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1138),
.A2(n_1241),
.B1(n_1234),
.B2(n_1145),
.Y(n_1286)
);

BUFx3_ASAP7_75t_L g1287 ( 
.A(n_1149),
.Y(n_1287)
);

OAI22xp5_ASAP7_75t_L g1288 ( 
.A1(n_1114),
.A2(n_1151),
.B1(n_1128),
.B2(n_1152),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1208),
.A2(n_1179),
.B1(n_1120),
.B2(n_1192),
.Y(n_1289)
);

OAI22xp5_ASAP7_75t_L g1290 ( 
.A1(n_1117),
.A2(n_1257),
.B1(n_1222),
.B2(n_1223),
.Y(n_1290)
);

NAND2xp5_ASAP7_75t_L g1291 ( 
.A(n_1167),
.B(n_1213),
.Y(n_1291)
);

OAI22xp33_ASAP7_75t_L g1292 ( 
.A1(n_1156),
.A2(n_1158),
.B1(n_1166),
.B2(n_1125),
.Y(n_1292)
);

OAI22xp5_ASAP7_75t_L g1293 ( 
.A1(n_1188),
.A2(n_1189),
.B1(n_1130),
.B2(n_1168),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1243),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1178),
.Y(n_1295)
);

CKINVDCx20_ASAP7_75t_R g1296 ( 
.A(n_1248),
.Y(n_1296)
);

INVx6_ASAP7_75t_L g1297 ( 
.A(n_1136),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1126),
.A2(n_1132),
.B1(n_1155),
.B2(n_1146),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1142),
.B(n_1159),
.Y(n_1299)
);

AOI22xp33_ASAP7_75t_L g1300 ( 
.A1(n_1126),
.A2(n_1146),
.B1(n_1173),
.B2(n_1124),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1186),
.Y(n_1301)
);

BUFx2_ASAP7_75t_L g1302 ( 
.A(n_1197),
.Y(n_1302)
);

CKINVDCx16_ASAP7_75t_R g1303 ( 
.A(n_1182),
.Y(n_1303)
);

AOI22xp33_ASAP7_75t_L g1304 ( 
.A1(n_1173),
.A2(n_1118),
.B1(n_1134),
.B2(n_1133),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1187),
.B(n_1165),
.Y(n_1305)
);

INVxp67_ASAP7_75t_L g1306 ( 
.A(n_1191),
.Y(n_1306)
);

OAI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1194),
.A2(n_1229),
.B1(n_1205),
.B2(n_1253),
.Y(n_1307)
);

INVx3_ASAP7_75t_L g1308 ( 
.A(n_1121),
.Y(n_1308)
);

BUFx3_ASAP7_75t_L g1309 ( 
.A(n_1198),
.Y(n_1309)
);

CKINVDCx11_ASAP7_75t_R g1310 ( 
.A(n_1140),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1140),
.Y(n_1311)
);

BUFx6f_ASAP7_75t_L g1312 ( 
.A(n_1196),
.Y(n_1312)
);

AOI22xp33_ASAP7_75t_SL g1313 ( 
.A1(n_1154),
.A2(n_1131),
.B1(n_1250),
.B2(n_1220),
.Y(n_1313)
);

AOI22xp33_ASAP7_75t_SL g1314 ( 
.A1(n_1154),
.A2(n_1131),
.B1(n_1214),
.B2(n_1200),
.Y(n_1314)
);

INVx1_ASAP7_75t_SL g1315 ( 
.A(n_1193),
.Y(n_1315)
);

CKINVDCx20_ASAP7_75t_R g1316 ( 
.A(n_1136),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1140),
.Y(n_1317)
);

BUFx3_ASAP7_75t_L g1318 ( 
.A(n_1160),
.Y(n_1318)
);

BUFx12f_ASAP7_75t_L g1319 ( 
.A(n_1160),
.Y(n_1319)
);

NAND2xp5_ASAP7_75t_L g1320 ( 
.A(n_1195),
.B(n_1136),
.Y(n_1320)
);

INVx8_ASAP7_75t_L g1321 ( 
.A(n_1160),
.Y(n_1321)
);

AOI22xp33_ASAP7_75t_L g1322 ( 
.A1(n_1134),
.A2(n_1237),
.B1(n_1249),
.B2(n_1242),
.Y(n_1322)
);

AOI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1141),
.A2(n_1154),
.B1(n_1180),
.B2(n_1113),
.Y(n_1323)
);

AOI22xp33_ASAP7_75t_L g1324 ( 
.A1(n_1190),
.A2(n_1181),
.B1(n_1131),
.B2(n_1161),
.Y(n_1324)
);

BUFx2_ASAP7_75t_L g1325 ( 
.A(n_1181),
.Y(n_1325)
);

AOI22xp33_ASAP7_75t_L g1326 ( 
.A1(n_1190),
.A2(n_1181),
.B1(n_1115),
.B2(n_1137),
.Y(n_1326)
);

INVx4_ASAP7_75t_L g1327 ( 
.A(n_1236),
.Y(n_1327)
);

AND2x2_ASAP7_75t_L g1328 ( 
.A(n_1122),
.B(n_1204),
.Y(n_1328)
);

OAI22xp5_ASAP7_75t_L g1329 ( 
.A1(n_1185),
.A2(n_1123),
.B1(n_1172),
.B2(n_1163),
.Y(n_1329)
);

AOI22xp5_ASAP7_75t_L g1330 ( 
.A1(n_1201),
.A2(n_1217),
.B1(n_1228),
.B2(n_1219),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1137),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1122),
.A2(n_1216),
.B1(n_1231),
.B2(n_1252),
.Y(n_1332)
);

CKINVDCx11_ASAP7_75t_R g1333 ( 
.A(n_1122),
.Y(n_1333)
);

CKINVDCx6p67_ASAP7_75t_R g1334 ( 
.A(n_1174),
.Y(n_1334)
);

BUFx12f_ASAP7_75t_L g1335 ( 
.A(n_1177),
.Y(n_1335)
);

NAND2x1p5_ASAP7_75t_L g1336 ( 
.A(n_1255),
.B(n_1218),
.Y(n_1336)
);

AOI22xp33_ASAP7_75t_L g1337 ( 
.A1(n_1112),
.A2(n_1235),
.B1(n_1252),
.B2(n_1177),
.Y(n_1337)
);

HB1xp67_ASAP7_75t_L g1338 ( 
.A(n_1235),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1252),
.Y(n_1339)
);

OAI22xp33_ASAP7_75t_L g1340 ( 
.A1(n_1177),
.A2(n_1254),
.B1(n_1210),
.B2(n_1259),
.Y(n_1340)
);

INVx3_ASAP7_75t_L g1341 ( 
.A(n_1121),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_1247),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_818),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1135),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1144),
.B(n_1211),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1135),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1196),
.Y(n_1347)
);

BUFx8_ASAP7_75t_L g1348 ( 
.A(n_1149),
.Y(n_1348)
);

INVx1_ASAP7_75t_L g1349 ( 
.A(n_1135),
.Y(n_1349)
);

AOI22xp5_ASAP7_75t_L g1350 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_652),
.B2(n_610),
.Y(n_1350)
);

AOI22xp33_ASAP7_75t_L g1351 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_818),
.Y(n_1351)
);

BUFx3_ASAP7_75t_L g1352 ( 
.A(n_1157),
.Y(n_1352)
);

INVx5_ASAP7_75t_L g1353 ( 
.A(n_1136),
.Y(n_1353)
);

AOI22xp33_ASAP7_75t_L g1354 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_1247),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_1256),
.Y(n_1355)
);

AOI22xp33_ASAP7_75t_SL g1356 ( 
.A1(n_1139),
.A2(n_1066),
.B1(n_1008),
.B2(n_323),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1144),
.B(n_1211),
.Y(n_1357)
);

AOI22xp33_ASAP7_75t_L g1358 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_1247),
.Y(n_1358)
);

CKINVDCx20_ASAP7_75t_R g1359 ( 
.A(n_1157),
.Y(n_1359)
);

CKINVDCx11_ASAP7_75t_R g1360 ( 
.A(n_1256),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_SL g1361 ( 
.A1(n_1139),
.A2(n_1066),
.B1(n_1008),
.B2(n_323),
.Y(n_1361)
);

OAI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1240),
.A2(n_652),
.B1(n_1259),
.B2(n_1227),
.Y(n_1362)
);

INVx4_ASAP7_75t_L g1363 ( 
.A(n_1136),
.Y(n_1363)
);

BUFx3_ASAP7_75t_L g1364 ( 
.A(n_1157),
.Y(n_1364)
);

INVx2_ASAP7_75t_SL g1365 ( 
.A(n_1176),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_818),
.Y(n_1366)
);

CKINVDCx11_ASAP7_75t_R g1367 ( 
.A(n_1256),
.Y(n_1367)
);

CKINVDCx11_ASAP7_75t_R g1368 ( 
.A(n_1256),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_L g1369 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_818),
.Y(n_1369)
);

BUFx6f_ASAP7_75t_L g1370 ( 
.A(n_1196),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_1127),
.Y(n_1371)
);

BUFx8_ASAP7_75t_L g1372 ( 
.A(n_1149),
.Y(n_1372)
);

BUFx5_ASAP7_75t_L g1373 ( 
.A(n_1173),
.Y(n_1373)
);

INVx4_ASAP7_75t_L g1374 ( 
.A(n_1136),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1135),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_L g1376 ( 
.A1(n_1240),
.A2(n_1259),
.B1(n_1150),
.B2(n_1247),
.Y(n_1376)
);

OAI21xp33_ASAP7_75t_L g1377 ( 
.A1(n_1240),
.A2(n_630),
.B(n_818),
.Y(n_1377)
);

INVx4_ASAP7_75t_SL g1378 ( 
.A(n_1190),
.Y(n_1378)
);

OAI22xp5_ASAP7_75t_L g1379 ( 
.A1(n_1240),
.A2(n_652),
.B1(n_1259),
.B2(n_1227),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1135),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1135),
.Y(n_1381)
);

AOI22xp33_ASAP7_75t_SL g1382 ( 
.A1(n_1139),
.A2(n_1066),
.B1(n_1008),
.B2(n_323),
.Y(n_1382)
);

INVx5_ASAP7_75t_L g1383 ( 
.A(n_1136),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1373),
.Y(n_1384)
);

INVx2_ASAP7_75t_L g1385 ( 
.A(n_1373),
.Y(n_1385)
);

HB1xp67_ASAP7_75t_L g1386 ( 
.A(n_1306),
.Y(n_1386)
);

AO21x2_ASAP7_75t_L g1387 ( 
.A1(n_1330),
.A2(n_1340),
.B(n_1307),
.Y(n_1387)
);

BUFx2_ASAP7_75t_L g1388 ( 
.A(n_1312),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1373),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1265),
.B(n_1328),
.Y(n_1390)
);

AOI22xp33_ASAP7_75t_L g1391 ( 
.A1(n_1377),
.A2(n_1379),
.B1(n_1362),
.B2(n_1366),
.Y(n_1391)
);

OR2x2_ASAP7_75t_L g1392 ( 
.A(n_1265),
.B(n_1332),
.Y(n_1392)
);

HB1xp67_ASAP7_75t_L g1393 ( 
.A(n_1306),
.Y(n_1393)
);

OAI22xp33_ASAP7_75t_L g1394 ( 
.A1(n_1350),
.A2(n_1269),
.B1(n_1303),
.B2(n_1288),
.Y(n_1394)
);

A2O1A1Ixp33_ASAP7_75t_L g1395 ( 
.A1(n_1343),
.A2(n_1351),
.B(n_1369),
.C(n_1342),
.Y(n_1395)
);

INVx2_ASAP7_75t_L g1396 ( 
.A(n_1264),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1301),
.Y(n_1397)
);

BUFx6f_ASAP7_75t_L g1398 ( 
.A(n_1335),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1297),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1338),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1275),
.Y(n_1402)
);

INVx2_ASAP7_75t_SL g1403 ( 
.A(n_1297),
.Y(n_1403)
);

CKINVDCx20_ASAP7_75t_R g1404 ( 
.A(n_1266),
.Y(n_1404)
);

AOI22xp33_ASAP7_75t_L g1405 ( 
.A1(n_1356),
.A2(n_1361),
.B1(n_1382),
.B2(n_1354),
.Y(n_1405)
);

INVx2_ASAP7_75t_L g1406 ( 
.A(n_1331),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1356),
.A2(n_1361),
.B1(n_1382),
.B2(n_1354),
.Y(n_1407)
);

INVx2_ASAP7_75t_SL g1408 ( 
.A(n_1297),
.Y(n_1408)
);

OR2x2_ASAP7_75t_L g1409 ( 
.A(n_1339),
.B(n_1299),
.Y(n_1409)
);

INVx2_ASAP7_75t_L g1410 ( 
.A(n_1336),
.Y(n_1410)
);

AOI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1329),
.A2(n_1293),
.B(n_1290),
.Y(n_1411)
);

NOR2xp33_ASAP7_75t_L g1412 ( 
.A(n_1345),
.B(n_1357),
.Y(n_1412)
);

NAND2xp5_ASAP7_75t_L g1413 ( 
.A(n_1267),
.B(n_1271),
.Y(n_1413)
);

OAI22xp33_ASAP7_75t_L g1414 ( 
.A1(n_1305),
.A2(n_1291),
.B1(n_1285),
.B2(n_1276),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1334),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1344),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1360),
.Y(n_1417)
);

INVx2_ASAP7_75t_L g1418 ( 
.A(n_1281),
.Y(n_1418)
);

BUFx6f_ASAP7_75t_L g1419 ( 
.A(n_1347),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1283),
.B(n_1296),
.Y(n_1420)
);

OAI21x1_ASAP7_75t_L g1421 ( 
.A1(n_1322),
.A2(n_1323),
.B(n_1304),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1268),
.B(n_1260),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1367),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1346),
.Y(n_1424)
);

BUFx8_ASAP7_75t_L g1425 ( 
.A(n_1261),
.Y(n_1425)
);

OAI21x1_ASAP7_75t_L g1426 ( 
.A1(n_1323),
.A2(n_1304),
.B(n_1326),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1326),
.A2(n_1337),
.B(n_1324),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1347),
.Y(n_1428)
);

AND2x2_ASAP7_75t_L g1429 ( 
.A(n_1278),
.B(n_1262),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1278),
.B(n_1262),
.Y(n_1430)
);

INVxp67_ASAP7_75t_SL g1431 ( 
.A(n_1268),
.Y(n_1431)
);

OAI21x1_ASAP7_75t_L g1432 ( 
.A1(n_1337),
.A2(n_1324),
.B(n_1300),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1370),
.Y(n_1433)
);

NAND2xp5_ASAP7_75t_L g1434 ( 
.A(n_1260),
.B(n_1358),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1370),
.Y(n_1435)
);

INVx2_ASAP7_75t_L g1436 ( 
.A(n_1349),
.Y(n_1436)
);

AO21x1_ASAP7_75t_L g1437 ( 
.A1(n_1340),
.A2(n_1307),
.B(n_1280),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1280),
.Y(n_1438)
);

OAI21x1_ASAP7_75t_L g1439 ( 
.A1(n_1298),
.A2(n_1375),
.B(n_1381),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1380),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1333),
.B(n_1314),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1292),
.Y(n_1442)
);

HB1xp67_ASAP7_75t_SL g1443 ( 
.A(n_1348),
.Y(n_1443)
);

INVx2_ASAP7_75t_L g1444 ( 
.A(n_1295),
.Y(n_1444)
);

INVx2_ASAP7_75t_L g1445 ( 
.A(n_1294),
.Y(n_1445)
);

BUFx3_ASAP7_75t_L g1446 ( 
.A(n_1353),
.Y(n_1446)
);

AO21x2_ASAP7_75t_L g1447 ( 
.A1(n_1292),
.A2(n_1276),
.B(n_1289),
.Y(n_1447)
);

AND2x2_ASAP7_75t_L g1448 ( 
.A(n_1314),
.B(n_1313),
.Y(n_1448)
);

INVx1_ASAP7_75t_L g1449 ( 
.A(n_1313),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1371),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1270),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1342),
.A2(n_1358),
.B1(n_1376),
.B2(n_1286),
.Y(n_1452)
);

AND2x2_ASAP7_75t_L g1453 ( 
.A(n_1376),
.B(n_1270),
.Y(n_1453)
);

OA21x2_ASAP7_75t_L g1454 ( 
.A1(n_1286),
.A2(n_1320),
.B(n_1315),
.Y(n_1454)
);

INVx8_ASAP7_75t_L g1455 ( 
.A(n_1353),
.Y(n_1455)
);

NAND2x1p5_ASAP7_75t_L g1456 ( 
.A(n_1353),
.B(n_1383),
.Y(n_1456)
);

AOI22xp5_ASAP7_75t_L g1457 ( 
.A1(n_1316),
.A2(n_1284),
.B1(n_1273),
.B2(n_1365),
.Y(n_1457)
);

OA21x2_ASAP7_75t_L g1458 ( 
.A1(n_1325),
.A2(n_1302),
.B(n_1378),
.Y(n_1458)
);

BUFx6f_ASAP7_75t_L g1459 ( 
.A(n_1353),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1383),
.Y(n_1460)
);

OA21x2_ASAP7_75t_L g1461 ( 
.A1(n_1383),
.A2(n_1327),
.B(n_1363),
.Y(n_1461)
);

INVx2_ASAP7_75t_L g1462 ( 
.A(n_1279),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1309),
.B(n_1279),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1287),
.A2(n_1272),
.B1(n_1274),
.B2(n_1363),
.Y(n_1464)
);

INVx1_ASAP7_75t_L g1465 ( 
.A(n_1374),
.Y(n_1465)
);

HB1xp67_ASAP7_75t_L g1466 ( 
.A(n_1308),
.Y(n_1466)
);

NAND2x1_ASAP7_75t_L g1467 ( 
.A(n_1461),
.B(n_1374),
.Y(n_1467)
);

CKINVDCx16_ASAP7_75t_R g1468 ( 
.A(n_1443),
.Y(n_1468)
);

AND2x4_ASAP7_75t_L g1469 ( 
.A(n_1415),
.B(n_1318),
.Y(n_1469)
);

OR2x2_ASAP7_75t_L g1470 ( 
.A(n_1390),
.B(n_1272),
.Y(n_1470)
);

NAND2xp5_ASAP7_75t_L g1471 ( 
.A(n_1431),
.B(n_1442),
.Y(n_1471)
);

BUFx4f_ASAP7_75t_SL g1472 ( 
.A(n_1404),
.Y(n_1472)
);

BUFx2_ASAP7_75t_L g1473 ( 
.A(n_1402),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1442),
.B(n_1341),
.Y(n_1474)
);

OAI22xp5_ASAP7_75t_SL g1475 ( 
.A1(n_1405),
.A2(n_1355),
.B1(n_1359),
.B2(n_1263),
.Y(n_1475)
);

NOR3xp33_ASAP7_75t_SL g1476 ( 
.A(n_1417),
.B(n_1368),
.C(n_1282),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1416),
.Y(n_1477)
);

NAND2xp5_ASAP7_75t_L g1478 ( 
.A(n_1409),
.B(n_1308),
.Y(n_1478)
);

OAI21xp5_ASAP7_75t_L g1479 ( 
.A1(n_1395),
.A2(n_1311),
.B(n_1317),
.Y(n_1479)
);

AOI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1407),
.A2(n_1277),
.B1(n_1372),
.B2(n_1348),
.Y(n_1480)
);

OR2x2_ASAP7_75t_L g1481 ( 
.A(n_1390),
.B(n_1352),
.Y(n_1481)
);

OAI21xp5_ASAP7_75t_L g1482 ( 
.A1(n_1391),
.A2(n_1364),
.B(n_1372),
.Y(n_1482)
);

INVxp67_ASAP7_75t_L g1483 ( 
.A(n_1412),
.Y(n_1483)
);

OAI21xp5_ASAP7_75t_L g1484 ( 
.A1(n_1394),
.A2(n_1319),
.B(n_1310),
.Y(n_1484)
);

OAI22xp5_ASAP7_75t_L g1485 ( 
.A1(n_1452),
.A2(n_1434),
.B1(n_1422),
.B2(n_1413),
.Y(n_1485)
);

AOI221xp5_ASAP7_75t_L g1486 ( 
.A1(n_1414),
.A2(n_1321),
.B1(n_1453),
.B2(n_1437),
.C(n_1451),
.Y(n_1486)
);

AND2x2_ASAP7_75t_L g1487 ( 
.A(n_1441),
.B(n_1321),
.Y(n_1487)
);

INVxp67_ASAP7_75t_L g1488 ( 
.A(n_1466),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1420),
.B(n_1457),
.Y(n_1489)
);

A2O1A1Ixp33_ASAP7_75t_L g1490 ( 
.A1(n_1453),
.A2(n_1430),
.B(n_1429),
.C(n_1401),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1441),
.B(n_1463),
.Y(n_1491)
);

AO32x2_ASAP7_75t_L g1492 ( 
.A1(n_1464),
.A2(n_1403),
.A3(n_1408),
.B1(n_1399),
.B2(n_1449),
.Y(n_1492)
);

AOI21xp5_ASAP7_75t_L g1493 ( 
.A1(n_1437),
.A2(n_1447),
.B(n_1387),
.Y(n_1493)
);

INVxp67_ASAP7_75t_L g1494 ( 
.A(n_1386),
.Y(n_1494)
);

AO21x2_ASAP7_75t_L g1495 ( 
.A1(n_1418),
.A2(n_1447),
.B(n_1387),
.Y(n_1495)
);

OAI22xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1457),
.A2(n_1423),
.B1(n_1454),
.B2(n_1451),
.Y(n_1496)
);

INVxp67_ASAP7_75t_L g1497 ( 
.A(n_1393),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1454),
.B(n_1396),
.Y(n_1498)
);

NAND2xp5_ASAP7_75t_L g1499 ( 
.A(n_1454),
.B(n_1445),
.Y(n_1499)
);

AND2x2_ASAP7_75t_L g1500 ( 
.A(n_1454),
.B(n_1396),
.Y(n_1500)
);

NAND4xp25_ASAP7_75t_L g1501 ( 
.A(n_1449),
.B(n_1430),
.C(n_1429),
.D(n_1438),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1440),
.Y(n_1502)
);

AOI22xp5_ASAP7_75t_L g1503 ( 
.A1(n_1447),
.A2(n_1438),
.B1(n_1387),
.B2(n_1398),
.Y(n_1503)
);

AND2x2_ASAP7_75t_L g1504 ( 
.A(n_1424),
.B(n_1436),
.Y(n_1504)
);

OA21x2_ASAP7_75t_L g1505 ( 
.A1(n_1421),
.A2(n_1426),
.B(n_1418),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1462),
.B(n_1399),
.Y(n_1506)
);

AOI22xp33_ASAP7_75t_L g1507 ( 
.A1(n_1448),
.A2(n_1398),
.B1(n_1392),
.B2(n_1425),
.Y(n_1507)
);

NAND2xp5_ASAP7_75t_L g1508 ( 
.A(n_1444),
.B(n_1440),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1444),
.B(n_1439),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1439),
.B(n_1388),
.Y(n_1510)
);

AO21x2_ASAP7_75t_L g1511 ( 
.A1(n_1411),
.A2(n_1384),
.B(n_1389),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1411),
.A2(n_1432),
.B(n_1427),
.Y(n_1512)
);

BUFx6f_ASAP7_75t_L g1513 ( 
.A(n_1459),
.Y(n_1513)
);

BUFx2_ASAP7_75t_L g1514 ( 
.A(n_1458),
.Y(n_1514)
);

HB1xp67_ASAP7_75t_L g1515 ( 
.A(n_1458),
.Y(n_1515)
);

OR2x6_ASAP7_75t_L g1516 ( 
.A(n_1455),
.B(n_1398),
.Y(n_1516)
);

OAI21xp5_ASAP7_75t_L g1517 ( 
.A1(n_1427),
.A2(n_1460),
.B(n_1450),
.Y(n_1517)
);

NOR2xp33_ASAP7_75t_L g1518 ( 
.A(n_1403),
.B(n_1408),
.Y(n_1518)
);

OR2x2_ASAP7_75t_L g1519 ( 
.A(n_1499),
.B(n_1514),
.Y(n_1519)
);

AND2x4_ASAP7_75t_L g1520 ( 
.A(n_1517),
.B(n_1385),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1505),
.B(n_1512),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1505),
.B(n_1385),
.Y(n_1522)
);

INVx2_ASAP7_75t_L g1523 ( 
.A(n_1509),
.Y(n_1523)
);

AND2x2_ASAP7_75t_L g1524 ( 
.A(n_1517),
.B(n_1448),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1498),
.Y(n_1525)
);

NAND2xp5_ASAP7_75t_L g1526 ( 
.A(n_1500),
.B(n_1397),
.Y(n_1526)
);

HB1xp67_ASAP7_75t_L g1527 ( 
.A(n_1515),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1502),
.Y(n_1528)
);

AND2x2_ASAP7_75t_L g1529 ( 
.A(n_1511),
.B(n_1495),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1511),
.B(n_1406),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1493),
.B(n_1397),
.Y(n_1531)
);

BUFx2_ASAP7_75t_L g1532 ( 
.A(n_1510),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1508),
.Y(n_1533)
);

NOR2xp67_ASAP7_75t_L g1534 ( 
.A(n_1503),
.B(n_1410),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1504),
.Y(n_1535)
);

HB1xp67_ASAP7_75t_L g1536 ( 
.A(n_1477),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1473),
.Y(n_1537)
);

NOR2x1p5_ASAP7_75t_L g1538 ( 
.A(n_1501),
.B(n_1398),
.Y(n_1538)
);

BUFx3_ASAP7_75t_L g1539 ( 
.A(n_1467),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_SL g1540 ( 
.A(n_1496),
.B(n_1398),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1474),
.Y(n_1541)
);

NAND2xp5_ASAP7_75t_L g1542 ( 
.A(n_1494),
.B(n_1400),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1492),
.B(n_1435),
.Y(n_1543)
);

BUFx3_ASAP7_75t_L g1544 ( 
.A(n_1513),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1519),
.B(n_1497),
.Y(n_1545)
);

AND2x2_ASAP7_75t_L g1546 ( 
.A(n_1523),
.B(n_1532),
.Y(n_1546)
);

HB1xp67_ASAP7_75t_L g1547 ( 
.A(n_1527),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1519),
.B(n_1478),
.Y(n_1548)
);

NOR2xp67_ASAP7_75t_L g1549 ( 
.A(n_1519),
.B(n_1501),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1528),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1528),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1528),
.Y(n_1552)
);

AOI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1540),
.A2(n_1484),
.B(n_1482),
.Y(n_1553)
);

INVx2_ASAP7_75t_L g1554 ( 
.A(n_1522),
.Y(n_1554)
);

AND2x2_ASAP7_75t_L g1555 ( 
.A(n_1524),
.B(n_1419),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1528),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1541),
.B(n_1488),
.Y(n_1557)
);

NAND4xp25_ASAP7_75t_L g1558 ( 
.A(n_1540),
.B(n_1480),
.C(n_1490),
.D(n_1486),
.Y(n_1558)
);

OR2x2_ASAP7_75t_L g1559 ( 
.A(n_1519),
.B(n_1478),
.Y(n_1559)
);

NAND2xp33_ASAP7_75t_R g1560 ( 
.A(n_1524),
.B(n_1476),
.Y(n_1560)
);

INVx3_ASAP7_75t_L g1561 ( 
.A(n_1520),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1524),
.B(n_1428),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1524),
.B(n_1525),
.Y(n_1563)
);

HB1xp67_ASAP7_75t_L g1564 ( 
.A(n_1527),
.Y(n_1564)
);

NAND3xp33_ASAP7_75t_L g1565 ( 
.A(n_1534),
.B(n_1484),
.C(n_1485),
.Y(n_1565)
);

INVx4_ASAP7_75t_L g1566 ( 
.A(n_1544),
.Y(n_1566)
);

INVx2_ASAP7_75t_L g1567 ( 
.A(n_1522),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1541),
.B(n_1471),
.Y(n_1568)
);

AOI221xp5_ASAP7_75t_L g1569 ( 
.A1(n_1531),
.A2(n_1485),
.B1(n_1475),
.B2(n_1482),
.C(n_1483),
.Y(n_1569)
);

HB1xp67_ASAP7_75t_L g1570 ( 
.A(n_1530),
.Y(n_1570)
);

OAI21xp5_ASAP7_75t_L g1571 ( 
.A1(n_1534),
.A2(n_1479),
.B(n_1507),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1538),
.A2(n_1489),
.B1(n_1491),
.B2(n_1487),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1543),
.B(n_1433),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1550),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1550),
.Y(n_1575)
);

INVx2_ASAP7_75t_L g1576 ( 
.A(n_1554),
.Y(n_1576)
);

INVxp67_ASAP7_75t_L g1577 ( 
.A(n_1549),
.Y(n_1577)
);

INVx1_ASAP7_75t_SL g1578 ( 
.A(n_1545),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1551),
.Y(n_1579)
);

INVx2_ASAP7_75t_L g1580 ( 
.A(n_1554),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1551),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1568),
.B(n_1536),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1552),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1561),
.B(n_1539),
.Y(n_1586)
);

INVx1_ASAP7_75t_SL g1587 ( 
.A(n_1545),
.Y(n_1587)
);

NAND4xp25_ASAP7_75t_L g1588 ( 
.A(n_1569),
.B(n_1534),
.C(n_1471),
.D(n_1479),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1563),
.B(n_1535),
.Y(n_1589)
);

AND2x4_ASAP7_75t_L g1590 ( 
.A(n_1561),
.B(n_1539),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1568),
.B(n_1536),
.Y(n_1591)
);

OR2x2_ASAP7_75t_L g1592 ( 
.A(n_1548),
.B(n_1526),
.Y(n_1592)
);

INVx2_ASAP7_75t_L g1593 ( 
.A(n_1554),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1556),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1547),
.B(n_1533),
.Y(n_1595)
);

AND2x4_ASAP7_75t_SL g1596 ( 
.A(n_1566),
.B(n_1516),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1556),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1561),
.B(n_1521),
.Y(n_1598)
);

AND2x2_ASAP7_75t_L g1599 ( 
.A(n_1563),
.B(n_1546),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1547),
.B(n_1564),
.Y(n_1600)
);

OR2x2_ASAP7_75t_L g1601 ( 
.A(n_1548),
.B(n_1526),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1567),
.Y(n_1602)
);

INVx1_ASAP7_75t_L g1603 ( 
.A(n_1564),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1548),
.B(n_1531),
.Y(n_1604)
);

AND2x2_ASAP7_75t_L g1605 ( 
.A(n_1546),
.B(n_1521),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1570),
.B(n_1543),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1573),
.Y(n_1607)
);

NAND2xp5_ASAP7_75t_L g1608 ( 
.A(n_1578),
.B(n_1549),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1578),
.B(n_1587),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1603),
.Y(n_1610)
);

INVxp67_ASAP7_75t_L g1611 ( 
.A(n_1583),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1577),
.B(n_1555),
.Y(n_1612)
);

NOR2x1_ASAP7_75t_L g1613 ( 
.A(n_1588),
.B(n_1565),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1587),
.B(n_1537),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1603),
.Y(n_1615)
);

INVx4_ASAP7_75t_L g1616 ( 
.A(n_1596),
.Y(n_1616)
);

INVx2_ASAP7_75t_L g1617 ( 
.A(n_1599),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1600),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1599),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1600),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1574),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1577),
.B(n_1555),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1607),
.B(n_1555),
.Y(n_1623)
);

NOR2xp33_ASAP7_75t_L g1624 ( 
.A(n_1588),
.B(n_1468),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1604),
.B(n_1559),
.Y(n_1625)
);

OAI21xp33_ASAP7_75t_L g1626 ( 
.A1(n_1604),
.A2(n_1558),
.B(n_1565),
.Y(n_1626)
);

NAND2x1p5_ASAP7_75t_L g1627 ( 
.A(n_1586),
.B(n_1538),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1607),
.B(n_1566),
.Y(n_1628)
);

AND2x4_ASAP7_75t_L g1629 ( 
.A(n_1596),
.B(n_1539),
.Y(n_1629)
);

AND2x2_ASAP7_75t_L g1630 ( 
.A(n_1606),
.B(n_1566),
.Y(n_1630)
);

OR2x6_ASAP7_75t_L g1631 ( 
.A(n_1586),
.B(n_1553),
.Y(n_1631)
);

AND2x2_ASAP7_75t_L g1632 ( 
.A(n_1606),
.B(n_1566),
.Y(n_1632)
);

AND2x2_ASAP7_75t_L g1633 ( 
.A(n_1606),
.B(n_1566),
.Y(n_1633)
);

OR2x2_ASAP7_75t_L g1634 ( 
.A(n_1583),
.B(n_1559),
.Y(n_1634)
);

NOR2x1_ASAP7_75t_L g1635 ( 
.A(n_1595),
.B(n_1558),
.Y(n_1635)
);

OAI321xp33_ASAP7_75t_L g1636 ( 
.A1(n_1591),
.A2(n_1571),
.A3(n_1569),
.B1(n_1553),
.B2(n_1572),
.C(n_1557),
.Y(n_1636)
);

OR2x2_ASAP7_75t_L g1637 ( 
.A(n_1591),
.B(n_1559),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1592),
.B(n_1537),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1574),
.Y(n_1639)
);

AOI221x1_ASAP7_75t_L g1640 ( 
.A1(n_1595),
.A2(n_1571),
.B1(n_1557),
.B2(n_1465),
.C(n_1542),
.Y(n_1640)
);

NAND3xp33_ASAP7_75t_L g1641 ( 
.A(n_1575),
.B(n_1560),
.C(n_1529),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1575),
.Y(n_1642)
);

INVx1_ASAP7_75t_SL g1643 ( 
.A(n_1596),
.Y(n_1643)
);

AND2x2_ASAP7_75t_L g1644 ( 
.A(n_1586),
.B(n_1562),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1579),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1592),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1579),
.Y(n_1647)
);

INVx2_ASAP7_75t_SL g1648 ( 
.A(n_1586),
.Y(n_1648)
);

AND2x2_ASAP7_75t_L g1649 ( 
.A(n_1590),
.B(n_1562),
.Y(n_1649)
);

AOI31xp33_ASAP7_75t_L g1650 ( 
.A1(n_1613),
.A2(n_1470),
.A3(n_1425),
.B(n_1481),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1609),
.B(n_1601),
.Y(n_1651)
);

AND2x4_ASAP7_75t_L g1652 ( 
.A(n_1616),
.B(n_1590),
.Y(n_1652)
);

NAND2x1p5_ASAP7_75t_L g1653 ( 
.A(n_1616),
.B(n_1538),
.Y(n_1653)
);

AND2x2_ASAP7_75t_L g1654 ( 
.A(n_1631),
.B(n_1590),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1610),
.Y(n_1655)
);

INVx2_ASAP7_75t_L g1656 ( 
.A(n_1630),
.Y(n_1656)
);

AOI211xp5_ASAP7_75t_SL g1657 ( 
.A1(n_1636),
.A2(n_1590),
.B(n_1585),
.C(n_1598),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1635),
.B(n_1601),
.Y(n_1658)
);

OR2x6_ASAP7_75t_L g1659 ( 
.A(n_1616),
.B(n_1455),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1621),
.Y(n_1660)
);

NAND3xp33_ASAP7_75t_L g1661 ( 
.A(n_1626),
.B(n_1529),
.C(n_1506),
.Y(n_1661)
);

INVx2_ASAP7_75t_SL g1662 ( 
.A(n_1648),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1631),
.B(n_1605),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1621),
.Y(n_1664)
);

INVx1_ASAP7_75t_L g1665 ( 
.A(n_1615),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1639),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1609),
.B(n_1545),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1624),
.B(n_1562),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1639),
.Y(n_1669)
);

INVx1_ASAP7_75t_L g1670 ( 
.A(n_1642),
.Y(n_1670)
);

INVx2_ASAP7_75t_SL g1671 ( 
.A(n_1648),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1630),
.Y(n_1672)
);

INVx1_ASAP7_75t_L g1673 ( 
.A(n_1642),
.Y(n_1673)
);

NAND2xp5_ASAP7_75t_L g1674 ( 
.A(n_1612),
.B(n_1622),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1634),
.B(n_1576),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1632),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1631),
.B(n_1605),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1645),
.Y(n_1678)
);

AO21x2_ASAP7_75t_L g1679 ( 
.A1(n_1641),
.A2(n_1594),
.B(n_1581),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1612),
.B(n_1589),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

INVxp67_ASAP7_75t_SL g1682 ( 
.A(n_1608),
.Y(n_1682)
);

AND2x2_ASAP7_75t_L g1683 ( 
.A(n_1631),
.B(n_1605),
.Y(n_1683)
);

INVx3_ASAP7_75t_SL g1684 ( 
.A(n_1643),
.Y(n_1684)
);

INVx1_ASAP7_75t_L g1685 ( 
.A(n_1660),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1660),
.Y(n_1686)
);

NOR2xp33_ASAP7_75t_L g1687 ( 
.A(n_1684),
.B(n_1425),
.Y(n_1687)
);

OR2x2_ASAP7_75t_L g1688 ( 
.A(n_1674),
.B(n_1638),
.Y(n_1688)
);

INVxp67_ASAP7_75t_SL g1689 ( 
.A(n_1658),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1664),
.Y(n_1690)
);

OAI221xp5_ASAP7_75t_L g1691 ( 
.A1(n_1657),
.A2(n_1661),
.B1(n_1684),
.B2(n_1682),
.C(n_1650),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1656),
.B(n_1622),
.Y(n_1692)
);

INVx1_ASAP7_75t_L g1693 ( 
.A(n_1664),
.Y(n_1693)
);

NAND2xp5_ASAP7_75t_L g1694 ( 
.A(n_1656),
.B(n_1611),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1667),
.B(n_1614),
.Y(n_1695)
);

AOI221xp5_ASAP7_75t_L g1696 ( 
.A1(n_1655),
.A2(n_1620),
.B1(n_1618),
.B2(n_1646),
.C(n_1619),
.Y(n_1696)
);

INVx3_ASAP7_75t_L g1697 ( 
.A(n_1652),
.Y(n_1697)
);

INVx1_ASAP7_75t_SL g1698 ( 
.A(n_1652),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1666),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1652),
.B(n_1644),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1672),
.B(n_1640),
.Y(n_1701)
);

OAI22xp5_ASAP7_75t_L g1702 ( 
.A1(n_1653),
.A2(n_1627),
.B1(n_1629),
.B2(n_1617),
.Y(n_1702)
);

O2A1O1Ixp33_ASAP7_75t_L g1703 ( 
.A1(n_1679),
.A2(n_1627),
.B(n_1640),
.C(n_1628),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1669),
.Y(n_1704)
);

NAND2xp5_ASAP7_75t_L g1705 ( 
.A(n_1672),
.B(n_1617),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1670),
.Y(n_1706)
);

AOI21xp33_ASAP7_75t_L g1707 ( 
.A1(n_1662),
.A2(n_1637),
.B(n_1634),
.Y(n_1707)
);

NAND2xp5_ASAP7_75t_L g1708 ( 
.A(n_1676),
.B(n_1619),
.Y(n_1708)
);

NOR3xp33_ASAP7_75t_L g1709 ( 
.A(n_1662),
.B(n_1628),
.C(n_1632),
.Y(n_1709)
);

OAI21xp5_ASAP7_75t_SL g1710 ( 
.A1(n_1691),
.A2(n_1653),
.B(n_1663),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1685),
.Y(n_1711)
);

AND2x2_ASAP7_75t_L g1712 ( 
.A(n_1700),
.B(n_1687),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1686),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1689),
.B(n_1676),
.Y(n_1714)
);

INVx1_ASAP7_75t_L g1715 ( 
.A(n_1690),
.Y(n_1715)
);

AOI22xp5_ASAP7_75t_L g1716 ( 
.A1(n_1702),
.A2(n_1679),
.B1(n_1659),
.B2(n_1677),
.Y(n_1716)
);

INVx1_ASAP7_75t_L g1717 ( 
.A(n_1693),
.Y(n_1717)
);

OAI22xp5_ASAP7_75t_L g1718 ( 
.A1(n_1698),
.A2(n_1653),
.B1(n_1627),
.B2(n_1659),
.Y(n_1718)
);

NAND2xp5_ASAP7_75t_L g1719 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1697),
.B(n_1671),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1709),
.B(n_1665),
.Y(n_1721)
);

OAI211xp5_ASAP7_75t_SL g1722 ( 
.A1(n_1696),
.A2(n_1668),
.B(n_1651),
.C(n_1681),
.Y(n_1722)
);

INVx1_ASAP7_75t_L g1723 ( 
.A(n_1699),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1709),
.B(n_1654),
.Y(n_1724)
);

AOI22xp33_ASAP7_75t_L g1725 ( 
.A1(n_1688),
.A2(n_1659),
.B1(n_1679),
.B2(n_1663),
.Y(n_1725)
);

AOI22xp5_ASAP7_75t_L g1726 ( 
.A1(n_1692),
.A2(n_1659),
.B1(n_1677),
.B2(n_1683),
.Y(n_1726)
);

AOI221xp5_ASAP7_75t_L g1727 ( 
.A1(n_1696),
.A2(n_1681),
.B1(n_1678),
.B2(n_1673),
.C(n_1683),
.Y(n_1727)
);

OAI21xp5_ASAP7_75t_SL g1728 ( 
.A1(n_1703),
.A2(n_1654),
.B(n_1667),
.Y(n_1728)
);

BUFx2_ASAP7_75t_L g1729 ( 
.A(n_1724),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_L g1730 ( 
.A(n_1724),
.B(n_1704),
.Y(n_1730)
);

NAND2xp5_ASAP7_75t_L g1731 ( 
.A(n_1719),
.B(n_1706),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1720),
.B(n_1694),
.Y(n_1732)
);

CKINVDCx16_ASAP7_75t_R g1733 ( 
.A(n_1712),
.Y(n_1733)
);

OR2x2_ASAP7_75t_L g1734 ( 
.A(n_1714),
.B(n_1695),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1711),
.Y(n_1735)
);

XOR2xp5_ASAP7_75t_L g1736 ( 
.A(n_1726),
.B(n_1705),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1713),
.Y(n_1737)
);

NOR2xp33_ASAP7_75t_L g1738 ( 
.A(n_1710),
.B(n_1707),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1727),
.B(n_1728),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_SL g1740 ( 
.A(n_1733),
.B(n_1703),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1729),
.B(n_1721),
.Y(n_1741)
);

OR2x2_ASAP7_75t_L g1742 ( 
.A(n_1730),
.B(n_1708),
.Y(n_1742)
);

NAND2xp5_ASAP7_75t_L g1743 ( 
.A(n_1738),
.B(n_1723),
.Y(n_1743)
);

NAND4xp75_ASAP7_75t_L g1744 ( 
.A(n_1739),
.B(n_1716),
.C(n_1715),
.D(n_1717),
.Y(n_1744)
);

AOI21xp5_ASAP7_75t_L g1745 ( 
.A1(n_1739),
.A2(n_1725),
.B(n_1722),
.Y(n_1745)
);

INVx1_ASAP7_75t_SL g1746 ( 
.A(n_1734),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1731),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1736),
.B(n_1678),
.Y(n_1748)
);

NOR2xp33_ASAP7_75t_L g1749 ( 
.A(n_1732),
.B(n_1718),
.Y(n_1749)
);

O2A1O1Ixp33_ASAP7_75t_L g1750 ( 
.A1(n_1740),
.A2(n_1735),
.B(n_1737),
.C(n_1701),
.Y(n_1750)
);

OAI211xp5_ASAP7_75t_SL g1751 ( 
.A1(n_1745),
.A2(n_1651),
.B(n_1680),
.C(n_1675),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_SL g1752 ( 
.A(n_1746),
.B(n_1629),
.Y(n_1752)
);

BUFx2_ASAP7_75t_L g1753 ( 
.A(n_1741),
.Y(n_1753)
);

AOI211xp5_ASAP7_75t_L g1754 ( 
.A1(n_1743),
.A2(n_1675),
.B(n_1629),
.C(n_1633),
.Y(n_1754)
);

INVx2_ASAP7_75t_L g1755 ( 
.A(n_1753),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1752),
.B(n_1749),
.Y(n_1756)
);

NAND4xp25_ASAP7_75t_L g1757 ( 
.A(n_1750),
.B(n_1748),
.C(n_1742),
.D(n_1747),
.Y(n_1757)
);

NOR4xp25_ASAP7_75t_L g1758 ( 
.A(n_1751),
.B(n_1744),
.C(n_1633),
.D(n_1637),
.Y(n_1758)
);

AOI222xp33_ASAP7_75t_L g1759 ( 
.A1(n_1754),
.A2(n_1472),
.B1(n_1425),
.B2(n_1623),
.C1(n_1582),
.C2(n_1598),
.Y(n_1759)
);

NAND5xp2_ASAP7_75t_SL g1760 ( 
.A(n_1750),
.B(n_1623),
.C(n_1649),
.D(n_1644),
.E(n_1585),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1755),
.Y(n_1761)
);

NAND4xp75_ASAP7_75t_L g1762 ( 
.A(n_1756),
.B(n_1649),
.C(n_1598),
.D(n_1582),
.Y(n_1762)
);

AOI221xp5_ASAP7_75t_SL g1763 ( 
.A1(n_1757),
.A2(n_1582),
.B1(n_1585),
.B2(n_1625),
.C(n_1576),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1758),
.B(n_1625),
.Y(n_1764)
);

AO22x2_ASAP7_75t_L g1765 ( 
.A1(n_1760),
.A2(n_1580),
.B1(n_1602),
.B2(n_1576),
.Y(n_1765)
);

NOR3xp33_ASAP7_75t_L g1766 ( 
.A(n_1761),
.B(n_1759),
.C(n_1518),
.Y(n_1766)
);

INVx2_ASAP7_75t_SL g1767 ( 
.A(n_1765),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1764),
.B(n_1580),
.Y(n_1768)
);

NAND4xp25_ASAP7_75t_SL g1769 ( 
.A(n_1766),
.B(n_1763),
.C(n_1762),
.D(n_1593),
.Y(n_1769)
);

INVx2_ASAP7_75t_L g1770 ( 
.A(n_1769),
.Y(n_1770)
);

INVx1_ASAP7_75t_SL g1771 ( 
.A(n_1770),
.Y(n_1771)
);

INVx1_ASAP7_75t_L g1772 ( 
.A(n_1770),
.Y(n_1772)
);

AOI22x1_ASAP7_75t_L g1773 ( 
.A1(n_1771),
.A2(n_1767),
.B1(n_1768),
.B2(n_1456),
.Y(n_1773)
);

AOI21xp33_ASAP7_75t_L g1774 ( 
.A1(n_1772),
.A2(n_1469),
.B(n_1465),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1773),
.Y(n_1775)
);

AOI21xp5_ASAP7_75t_L g1776 ( 
.A1(n_1774),
.A2(n_1602),
.B(n_1580),
.Y(n_1776)
);

AOI22xp33_ASAP7_75t_L g1777 ( 
.A1(n_1775),
.A2(n_1539),
.B1(n_1469),
.B2(n_1602),
.Y(n_1777)
);

NAND2x2_ASAP7_75t_L g1778 ( 
.A(n_1777),
.B(n_1776),
.Y(n_1778)
);

BUFx2_ASAP7_75t_L g1779 ( 
.A(n_1778),
.Y(n_1779)
);

AOI221xp5_ASAP7_75t_L g1780 ( 
.A1(n_1779),
.A2(n_1584),
.B1(n_1597),
.B2(n_1594),
.C(n_1581),
.Y(n_1780)
);

AOI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1780),
.A2(n_1459),
.B(n_1460),
.C(n_1446),
.Y(n_1781)
);


endmodule