module fake_netlist_1_2788_n_41 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_41);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_41;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_28;
wire n_23;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_30;
wire n_13;
wire n_26;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_40;
wire n_27;
wire n_39;
NOR2xp33_ASAP7_75t_L g11 ( .A(n_2), .B(n_9), .Y(n_11) );
INVx2_ASAP7_75t_L g12 ( .A(n_8), .Y(n_12) );
CKINVDCx5p33_ASAP7_75t_R g13 ( .A(n_1), .Y(n_13) );
AND2x4_ASAP7_75t_L g14 ( .A(n_5), .B(n_4), .Y(n_14) );
CKINVDCx16_ASAP7_75t_R g15 ( .A(n_0), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_2), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_0), .Y(n_17) );
BUFx3_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NOR3xp33_ASAP7_75t_SL g19 ( .A(n_15), .B(n_1), .C(n_3), .Y(n_19) );
NOR3xp33_ASAP7_75t_SL g20 ( .A(n_15), .B(n_3), .C(n_4), .Y(n_20) );
AND2x2_ASAP7_75t_L g21 ( .A(n_17), .B(n_5), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_17), .B(n_6), .Y(n_22) );
OAI221xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_16), .B1(n_13), .B2(n_11), .C(n_12), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_18), .B(n_12), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_21), .Y(n_25) );
INVx6_ASAP7_75t_L g26 ( .A(n_21), .Y(n_26) );
INVx1_ASAP7_75t_L g27 ( .A(n_24), .Y(n_27) );
INVx1_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
INVx1_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
INVx1_ASAP7_75t_L g30 ( .A(n_28), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_27), .Y(n_31) );
OAI321xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_23), .A3(n_22), .B1(n_27), .B2(n_29), .C(n_20), .Y(n_32) );
AOI22xp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_26), .B1(n_19), .B2(n_14), .Y(n_33) );
INVx2_ASAP7_75t_SL g34 ( .A(n_33), .Y(n_34) );
AOI21xp5_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_14), .B(n_18), .Y(n_35) );
NOR3x1_ASAP7_75t_L g36 ( .A(n_32), .B(n_6), .C(n_7), .Y(n_36) );
OAI211xp5_ASAP7_75t_SL g37 ( .A1(n_34), .A2(n_26), .B(n_14), .C(n_7), .Y(n_37) );
NAND3xp33_ASAP7_75t_L g38 ( .A(n_35), .B(n_14), .C(n_18), .Y(n_38) );
BUFx2_ASAP7_75t_L g39 ( .A(n_38), .Y(n_39) );
INVxp67_ASAP7_75t_SL g40 ( .A(n_37), .Y(n_40) );
AOI22xp5_ASAP7_75t_L g41 ( .A1(n_40), .A2(n_10), .B1(n_36), .B2(n_39), .Y(n_41) );
endmodule