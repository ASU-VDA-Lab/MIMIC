module fake_jpeg_22252_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx3_ASAP7_75t_L g7 ( 
.A(n_6),
.Y(n_7)
);

CKINVDCx20_ASAP7_75t_R g8 ( 
.A(n_6),
.Y(n_8)
);

BUFx12_ASAP7_75t_L g9 ( 
.A(n_4),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_3),
.Y(n_10)
);

NAND2xp5_ASAP7_75t_SL g11 ( 
.A(n_1),
.B(n_2),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

BUFx12f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_0),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_17),
.B(n_18),
.Y(n_28)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_8),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_20),
.B(n_21),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_10),
.B(n_0),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_22),
.Y(n_37)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_27),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_25),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_13),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_5),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_17),
.A2(n_7),
.B1(n_14),
.B2(n_13),
.Y(n_33)
);

XOR2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_7),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g36 ( 
.A1(n_24),
.A2(n_15),
.B(n_14),
.Y(n_36)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_36),
.B(n_18),
.C(n_23),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_32),
.Y(n_43)
);

XOR2xp5_ASAP7_75t_L g45 ( 
.A(n_39),
.B(n_29),
.Y(n_45)
);

OAI21xp5_ASAP7_75t_SL g46 ( 
.A1(n_40),
.A2(n_34),
.B(n_35),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_19),
.Y(n_41)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_41),
.B(n_42),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g42 ( 
.A(n_29),
.B(n_28),
.Y(n_42)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_43),
.A2(n_37),
.B1(n_34),
.B2(n_16),
.Y(n_49)
);

XOR2xp5_ASAP7_75t_L g47 ( 
.A(n_45),
.B(n_46),
.Y(n_47)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_39),
.B1(n_31),
.B2(n_15),
.Y(n_48)
);

INVx1_ASAP7_75t_SL g51 ( 
.A(n_48),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_49),
.B(n_44),
.C(n_16),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_48),
.B(n_47),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_52),
.B(n_47),
.C(n_51),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_48),
.Y(n_54)
);


endmodule