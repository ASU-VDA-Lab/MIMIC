module fake_jpeg_817_n_487 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_487);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_487;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_15;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_292;
wire n_213;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_476;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx5_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx8_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_0),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

BUFx2_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_4),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_11),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_3),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_14),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_3),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_16),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_47),
.Y(n_144)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_48),
.Y(n_146)
);

CKINVDCx14_ASAP7_75t_R g49 ( 
.A(n_28),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_49),
.B(n_52),
.Y(n_104)
);

AND2x2_ASAP7_75t_SL g50 ( 
.A(n_24),
.B(n_7),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_50),
.B(n_85),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

INVx6_ASAP7_75t_L g108 ( 
.A(n_51),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_13),
.Y(n_52)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_24),
.Y(n_53)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g153 ( 
.A(n_54),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_55),
.Y(n_142)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_24),
.Y(n_56)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

HB1xp67_ASAP7_75t_L g57 ( 
.A(n_27),
.Y(n_57)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_57),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g58 ( 
.A(n_34),
.B(n_12),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_58),
.B(n_72),
.Y(n_116)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

INVx5_ASAP7_75t_L g152 ( 
.A(n_59),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_60),
.Y(n_154)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_15),
.Y(n_62)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_62),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_63),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_64),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g145 ( 
.A(n_65),
.Y(n_145)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_66),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx4f_ASAP7_75t_SL g100 ( 
.A(n_67),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_40),
.Y(n_68)
);

BUFx12f_ASAP7_75t_L g112 ( 
.A(n_68),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_69),
.Y(n_136)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_32),
.Y(n_70)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_70),
.Y(n_150)
);

INVx4_ASAP7_75t_L g71 ( 
.A(n_15),
.Y(n_71)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_71),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_41),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g73 ( 
.A1(n_35),
.A2(n_11),
.B1(n_10),
.B2(n_9),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g102 ( 
.A1(n_73),
.A2(n_46),
.B1(n_23),
.B2(n_17),
.Y(n_102)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_35),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_28),
.Y(n_75)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_15),
.Y(n_76)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx12f_ASAP7_75t_L g133 ( 
.A(n_77),
.Y(n_133)
);

INVx6_ASAP7_75t_L g78 ( 
.A(n_30),
.Y(n_78)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_78),
.Y(n_121)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_79),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_30),
.Y(n_80)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_80),
.Y(n_123)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_18),
.Y(n_81)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx5_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_19),
.Y(n_83)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_83),
.Y(n_127)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_84),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_30),
.Y(n_86)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_86),
.Y(n_129)
);

BUFx5_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_89),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g90 ( 
.A(n_29),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_90),
.B(n_95),
.Y(n_124)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_91),
.Y(n_148)
);

INVx8_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_92),
.Y(n_151)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_93),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_20),
.B(n_11),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_94),
.B(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_41),
.Y(n_95)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_34),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_42),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_97),
.B(n_98),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_42),
.Y(n_98)
);

OAI21xp33_ASAP7_75t_L g177 ( 
.A1(n_102),
.A2(n_0),
.B(n_1),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_29),
.B1(n_41),
.B2(n_34),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_106),
.A2(n_109),
.B1(n_140),
.B2(n_73),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_75),
.A2(n_41),
.B1(n_38),
.B2(n_33),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_52),
.B(n_43),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_120),
.B(n_103),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_50),
.B(n_43),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_132),
.B(n_143),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_58),
.A2(n_42),
.B1(n_46),
.B2(n_17),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_134),
.A2(n_135),
.B1(n_156),
.B2(n_39),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_78),
.A2(n_38),
.B1(n_33),
.B2(n_32),
.Y(n_135)
);

AOI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_64),
.A2(n_33),
.B(n_38),
.Y(n_138)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_138),
.B(n_149),
.C(n_39),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g140 ( 
.A1(n_85),
.A2(n_37),
.B1(n_23),
.B2(n_45),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_70),
.B(n_20),
.Y(n_143)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_83),
.B(n_45),
.C(n_44),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_85),
.B(n_31),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_155),
.B(n_125),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g156 ( 
.A1(n_77),
.A2(n_37),
.B1(n_21),
.B2(n_31),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_146),
.Y(n_157)
);

INVx3_ASAP7_75t_L g224 ( 
.A(n_157),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g220 ( 
.A(n_158),
.B(n_193),
.Y(n_220)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_137),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g207 ( 
.A(n_159),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_107),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_160),
.B(n_174),
.Y(n_215)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_121),
.Y(n_161)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_161),
.Y(n_208)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_105),
.B(n_76),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g229 ( 
.A(n_162),
.Y(n_229)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_124),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_163),
.B(n_165),
.Y(n_204)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

INVx3_ASAP7_75t_L g234 ( 
.A(n_164),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_104),
.B(n_22),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_166),
.B(n_191),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g232 ( 
.A(n_167),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_168),
.A2(n_177),
.B1(n_198),
.B2(n_199),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_144),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_171),
.Y(n_213)
);

INVx3_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_172),
.Y(n_218)
);

INVx6_ASAP7_75t_L g173 ( 
.A(n_144),
.Y(n_173)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_173),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_145),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_123),
.Y(n_175)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_175),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_116),
.B(n_149),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_176),
.B(n_178),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_105),
.B(n_36),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_134),
.B(n_36),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_179),
.B(n_183),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_180),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_196),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_138),
.A2(n_98),
.B1(n_97),
.B2(n_91),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_44),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g184 ( 
.A(n_153),
.B(n_84),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_184),
.B(n_189),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_55),
.B1(n_51),
.B2(n_47),
.Y(n_185)
);

INVx3_ASAP7_75t_SL g186 ( 
.A(n_150),
.Y(n_186)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_186),
.Y(n_211)
);

BUFx2_ASAP7_75t_L g187 ( 
.A(n_119),
.Y(n_187)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_187),
.Y(n_221)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_152),
.Y(n_188)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_188),
.Y(n_227)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_129),
.Y(n_190)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_190),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_122),
.B(n_48),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_110),
.B(n_22),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_192),
.B(n_21),
.Y(n_216)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_151),
.Y(n_193)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_147),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_194),
.Y(n_205)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_148),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_195),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_102),
.A2(n_65),
.B1(n_63),
.B2(n_60),
.Y(n_196)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_99),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_197),
.B(n_100),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_119),
.Y(n_198)
);

INVx5_ASAP7_75t_L g199 ( 
.A(n_152),
.Y(n_199)
);

BUFx3_ASAP7_75t_L g200 ( 
.A(n_136),
.Y(n_200)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_200),
.B(n_136),
.Y(n_236)
);

AND2x2_ASAP7_75t_L g201 ( 
.A(n_153),
.B(n_62),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_201),
.B(n_113),
.C(n_126),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_203),
.B(n_71),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_158),
.A2(n_176),
.B1(n_182),
.B2(n_179),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_206),
.A2(n_214),
.B1(n_222),
.B2(n_99),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_162),
.B(n_111),
.C(n_115),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_209),
.B(n_201),
.C(n_113),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_177),
.A2(n_118),
.B1(n_109),
.B2(n_106),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_216),
.B(n_195),
.Y(n_255)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_181),
.A2(n_140),
.B1(n_80),
.B2(n_86),
.Y(n_222)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_236),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_206),
.A2(n_178),
.B(n_162),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g277 ( 
.A1(n_237),
.A2(n_243),
.B(n_246),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_220),
.B(n_183),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_238),
.B(n_251),
.C(n_259),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g239 ( 
.A(n_228),
.B(n_170),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_239),
.B(n_241),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_228),
.B(n_161),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_230),
.Y(n_242)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_242),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_214),
.A2(n_131),
.B1(n_201),
.B2(n_187),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_230),
.Y(n_244)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_244),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_231),
.A2(n_184),
.B1(n_108),
.B2(n_154),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_245),
.A2(n_249),
.B1(n_250),
.B2(n_257),
.Y(n_266)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_222),
.A2(n_157),
.B1(n_188),
.B2(n_172),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_224),
.Y(n_247)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_247),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_215),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_248),
.B(n_255),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_231),
.A2(n_100),
.B1(n_142),
.B2(n_154),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_217),
.A2(n_100),
.B1(n_142),
.B2(n_173),
.Y(n_250)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_253),
.Y(n_286)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_225),
.Y(n_254)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_254),
.Y(n_290)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_229),
.A2(n_135),
.B1(n_199),
.B2(n_200),
.Y(n_256)
);

AND2x2_ASAP7_75t_L g267 ( 
.A(n_256),
.B(n_261),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_220),
.A2(n_145),
.B1(n_141),
.B2(n_130),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_258),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_220),
.B(n_127),
.C(n_130),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_260),
.A2(n_264),
.B1(n_236),
.B2(n_205),
.Y(n_278)
);

OA22x2_ASAP7_75t_L g261 ( 
.A1(n_207),
.A2(n_197),
.B1(n_175),
.B2(n_190),
.Y(n_261)
);

BUFx3_ASAP7_75t_L g262 ( 
.A(n_211),
.Y(n_262)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_262),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_203),
.B(n_114),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_263),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_226),
.A2(n_180),
.B1(n_169),
.B2(n_67),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_167),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_265),
.B(n_218),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_260),
.A2(n_219),
.B1(n_235),
.B2(n_216),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_270),
.A2(n_271),
.B1(n_274),
.B2(n_275),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_249),
.A2(n_207),
.B1(n_227),
.B2(n_224),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_245),
.A2(n_210),
.B1(n_209),
.B2(n_236),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_241),
.B1(n_265),
.B2(n_263),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g303 ( 
.A1(n_278),
.A2(n_285),
.B1(n_272),
.B2(n_280),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_240),
.A2(n_210),
.B1(n_233),
.B2(n_204),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_280),
.A2(n_288),
.B1(n_292),
.B2(n_250),
.Y(n_304)
);

OAI21xp5_ASAP7_75t_L g281 ( 
.A1(n_252),
.A2(n_212),
.B(n_227),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_281),
.A2(n_282),
.B(n_283),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_258),
.A2(n_205),
.B(n_194),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g283 ( 
.A1(n_248),
.A2(n_212),
.B(n_204),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_238),
.B(n_237),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_287),
.B(n_258),
.C(n_255),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_L g288 ( 
.A1(n_246),
.A2(n_233),
.B1(n_223),
.B2(n_202),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g297 ( 
.A(n_289),
.B(n_242),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_238),
.B(n_117),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_291),
.B(n_251),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_243),
.A2(n_223),
.B1(n_218),
.B2(n_202),
.Y(n_292)
);

XNOR2x2_ASAP7_75t_SL g294 ( 
.A(n_258),
.B(n_221),
.Y(n_294)
);

NOR2x1_ASAP7_75t_SL g310 ( 
.A(n_294),
.B(n_295),
.Y(n_310)
);

AND2x4_ASAP7_75t_SL g295 ( 
.A(n_257),
.B(n_128),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_283),
.B(n_239),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_296),
.B(n_313),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_297),
.B(n_298),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_282),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_293),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_300),
.B(n_323),
.Y(n_339)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_273),
.Y(n_301)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_301),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_289),
.Y(n_302)
);

AOI22xp33_ASAP7_75t_L g347 ( 
.A1(n_302),
.A2(n_319),
.B1(n_321),
.B2(n_322),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_303),
.A2(n_304),
.B1(n_314),
.B2(n_266),
.Y(n_334)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_273),
.Y(n_305)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_305),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_287),
.B(n_259),
.Y(n_306)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_306),
.B(n_307),
.Y(n_327)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_263),
.Y(n_307)
);

XNOR2xp5_ASAP7_75t_SL g342 ( 
.A(n_308),
.B(n_291),
.Y(n_342)
);

HB1xp67_ASAP7_75t_L g309 ( 
.A(n_293),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_269),
.B(n_263),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_311),
.B(n_312),
.C(n_221),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_SL g313 ( 
.A(n_276),
.B(n_262),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_278),
.A2(n_267),
.B1(n_270),
.B2(n_274),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_276),
.B(n_232),
.Y(n_315)
);

CKINVDCx16_ASAP7_75t_R g333 ( 
.A(n_315),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_281),
.Y(n_316)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_316),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_267),
.B(n_256),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_317),
.Y(n_329)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_279),
.Y(n_318)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_318),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g319 ( 
.A(n_295),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_268),
.B(n_264),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g350 ( 
.A(n_320),
.Y(n_350)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_279),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_286),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_268),
.B(n_244),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_275),
.B(n_254),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_301),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_299),
.A2(n_267),
.B1(n_266),
.B2(n_292),
.Y(n_326)
);

OAI22xp5_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_330),
.B1(n_332),
.B2(n_334),
.Y(n_356)
);

AOI22x1_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_288),
.B1(n_294),
.B2(n_277),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_314),
.A2(n_324),
.B1(n_302),
.B2(n_317),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_304),
.A2(n_277),
.B1(n_286),
.B2(n_290),
.Y(n_336)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_336),
.A2(n_344),
.B1(n_346),
.B2(n_351),
.Y(n_360)
);

XOR2xp5_ASAP7_75t_L g338 ( 
.A(n_307),
.B(n_306),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g358 ( 
.A(n_338),
.B(n_342),
.Y(n_358)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_297),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_341),
.B(n_321),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_323),
.A2(n_294),
.B1(n_295),
.B2(n_290),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g345 ( 
.A1(n_319),
.A2(n_284),
.B1(n_295),
.B2(n_261),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_345),
.A2(n_234),
.B1(n_186),
.B2(n_164),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_320),
.A2(n_284),
.B1(n_247),
.B2(n_253),
.Y(n_346)
);

XNOR2xp5_ASAP7_75t_SL g348 ( 
.A(n_308),
.B(n_261),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_348),
.B(n_325),
.Y(n_359)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_349),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g351 ( 
.A1(n_298),
.A2(n_261),
.B1(n_262),
.B2(n_202),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_353),
.B(n_355),
.C(n_312),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_325),
.A2(n_310),
.B1(n_300),
.B2(n_318),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_354),
.A2(n_330),
.B1(n_344),
.B2(n_329),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_213),
.C(n_208),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_357),
.B(n_363),
.C(n_378),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_SL g403 ( 
.A(n_359),
.B(n_362),
.Y(n_403)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_327),
.B(n_310),
.Y(n_362)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_362),
.B(n_370),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_327),
.B(n_322),
.C(n_305),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g364 ( 
.A(n_338),
.B(n_353),
.Y(n_364)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_364),
.B(n_367),
.Y(n_394)
);

OAI21xp5_ASAP7_75t_SL g405 ( 
.A1(n_365),
.A2(n_381),
.B(n_26),
.Y(n_405)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_339),
.Y(n_366)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_366),
.Y(n_384)
);

XNOR2xp5_ASAP7_75t_L g367 ( 
.A(n_348),
.B(n_355),
.Y(n_367)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_368),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g369 ( 
.A(n_337),
.B(n_261),
.Y(n_369)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_369),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g370 ( 
.A(n_342),
.B(n_213),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_SL g371 ( 
.A(n_332),
.B(n_208),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_371),
.B(n_380),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_L g372 ( 
.A1(n_350),
.A2(n_223),
.B1(n_234),
.B2(n_211),
.Y(n_372)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_372),
.Y(n_401)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_339),
.Y(n_373)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_373),
.Y(n_402)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_343),
.B(n_139),
.Y(n_374)
);

XOR2xp5_ASAP7_75t_L g385 ( 
.A(n_374),
.B(n_345),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g375 ( 
.A(n_333),
.B(n_341),
.Y(n_375)
);

CKINVDCx16_ASAP7_75t_R g389 ( 
.A(n_375),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_L g376 ( 
.A1(n_326),
.A2(n_347),
.B1(n_351),
.B2(n_330),
.Y(n_376)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_376),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_377),
.A2(n_340),
.B1(n_328),
.B2(n_133),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_343),
.B(n_198),
.C(n_171),
.Y(n_378)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_354),
.A2(n_68),
.B1(n_133),
.B2(n_112),
.Y(n_379)
);

AOI22xp5_ASAP7_75t_L g392 ( 
.A1(n_379),
.A2(n_382),
.B1(n_335),
.B2(n_328),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g380 ( 
.A(n_349),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_331),
.A2(n_37),
.B(n_39),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g382 ( 
.A1(n_331),
.A2(n_346),
.B1(n_352),
.B2(n_335),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_385),
.B(n_397),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_357),
.B(n_340),
.C(n_352),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_387),
.B(n_404),
.Y(n_414)
);

INVx1_ASAP7_75t_SL g388 ( 
.A(n_368),
.Y(n_388)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_388),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g423 ( 
.A1(n_392),
.A2(n_93),
.B1(n_59),
.B2(n_10),
.Y(n_423)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_393),
.A2(n_395),
.B1(n_396),
.B2(n_379),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_361),
.A2(n_112),
.B1(n_90),
.B2(n_26),
.Y(n_395)
);

OAI22xp5_ASAP7_75t_SL g396 ( 
.A1(n_361),
.A2(n_366),
.B1(n_369),
.B2(n_356),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_363),
.B(n_112),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_364),
.B(n_90),
.Y(n_400)
);

XOR2xp5_ASAP7_75t_L g417 ( 
.A(n_400),
.B(n_403),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_367),
.B(n_26),
.Y(n_404)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_405),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_386),
.B(n_358),
.C(n_370),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_406),
.B(n_409),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g407 ( 
.A1(n_387),
.A2(n_359),
.B(n_378),
.Y(n_407)
);

AOI21xp33_ASAP7_75t_L g438 ( 
.A1(n_407),
.A2(n_391),
.B(n_398),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_358),
.C(n_371),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_410),
.Y(n_426)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_401),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_411),
.B(n_413),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_394),
.B(n_360),
.C(n_382),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_394),
.B(n_374),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_415),
.B(n_419),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_389),
.B(n_402),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_SL g436 ( 
.A(n_416),
.B(n_418),
.Y(n_436)
);

CKINVDCx16_ASAP7_75t_R g418 ( 
.A(n_390),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_400),
.C(n_383),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g420 ( 
.A(n_403),
.B(n_377),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_420),
.B(n_392),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_384),
.B(n_381),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_424),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_383),
.B(n_88),
.C(n_92),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_422),
.B(n_388),
.C(n_393),
.Y(n_435)
);

XOR2xp5_ASAP7_75t_L g428 ( 
.A(n_423),
.B(n_405),
.Y(n_428)
);

HB1xp67_ASAP7_75t_L g424 ( 
.A(n_396),
.Y(n_424)
);

HB1xp67_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

XOR2xp5_ASAP7_75t_L g429 ( 
.A(n_417),
.B(n_398),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g444 ( 
.A(n_429),
.B(n_431),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g431 ( 
.A(n_417),
.B(n_385),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g443 ( 
.A(n_434),
.B(n_412),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g456 ( 
.A(n_435),
.B(n_0),
.Y(n_456)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_414),
.A2(n_409),
.B(n_413),
.Y(n_437)
);

OAI21x1_ASAP7_75t_L g454 ( 
.A1(n_437),
.A2(n_441),
.B(n_428),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g446 ( 
.A(n_438),
.B(n_439),
.Y(n_446)
);

NOR2xp33_ASAP7_75t_L g439 ( 
.A(n_408),
.B(n_399),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g440 ( 
.A(n_406),
.B(n_395),
.C(n_1),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g450 ( 
.A(n_440),
.B(n_442),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g441 ( 
.A1(n_425),
.A2(n_8),
.B(n_9),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g442 ( 
.A1(n_410),
.A2(n_9),
.B1(n_8),
.B2(n_2),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g465 ( 
.A(n_443),
.B(n_452),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_433),
.B(n_412),
.C(n_419),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_445),
.B(n_447),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g447 ( 
.A(n_436),
.B(n_415),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_432),
.B(n_420),
.Y(n_449)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_449),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_430),
.B(n_422),
.C(n_9),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_SL g466 ( 
.A(n_451),
.B(n_453),
.Y(n_466)
);

XOR2x2_ASAP7_75t_SL g452 ( 
.A(n_429),
.B(n_431),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g453 ( 
.A1(n_427),
.A2(n_8),
.B(n_1),
.Y(n_453)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_454),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_434),
.B(n_8),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_455),
.B(n_456),
.Y(n_460)
);

OR2x2_ASAP7_75t_L g457 ( 
.A(n_446),
.B(n_426),
.Y(n_457)
);

OAI21x1_ASAP7_75t_L g470 ( 
.A1(n_457),
.A2(n_467),
.B(n_450),
.Y(n_470)
);

NOR2xp67_ASAP7_75t_L g459 ( 
.A(n_444),
.B(n_435),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g474 ( 
.A1(n_459),
.A2(n_5),
.B(n_6),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_448),
.A2(n_426),
.B1(n_440),
.B2(n_4),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g473 ( 
.A(n_461),
.B(n_462),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_445),
.B(n_2),
.C(n_3),
.Y(n_462)
);

NOR2x1_ASAP7_75t_L g467 ( 
.A(n_452),
.B(n_3),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_458),
.B(n_464),
.Y(n_468)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_468),
.B(n_471),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_SL g469 ( 
.A1(n_463),
.A2(n_448),
.B(n_443),
.Y(n_469)
);

OAI21xp5_ASAP7_75t_L g480 ( 
.A1(n_469),
.A2(n_462),
.B(n_5),
.Y(n_480)
);

AO21x1_ASAP7_75t_L g477 ( 
.A1(n_470),
.A2(n_472),
.B(n_466),
.Y(n_477)
);

NOR2x1_ASAP7_75t_L g471 ( 
.A(n_465),
.B(n_4),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g472 ( 
.A(n_465),
.B(n_4),
.Y(n_472)
);

AOI21xp33_ASAP7_75t_L g479 ( 
.A1(n_474),
.A2(n_460),
.B(n_467),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_457),
.B(n_5),
.Y(n_475)
);

CKINVDCx20_ASAP7_75t_R g478 ( 
.A(n_475),
.Y(n_478)
);

CKINVDCx20_ASAP7_75t_R g483 ( 
.A(n_477),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_479),
.B(n_470),
.Y(n_481)
);

NAND3xp33_ASAP7_75t_L g482 ( 
.A(n_480),
.B(n_473),
.C(n_5),
.Y(n_482)
);

AOI21xp5_ASAP7_75t_L g484 ( 
.A1(n_481),
.A2(n_482),
.B(n_476),
.Y(n_484)
);

OAI31xp33_ASAP7_75t_SL g485 ( 
.A1(n_484),
.A2(n_483),
.A3(n_478),
.B(n_6),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_485),
.B(n_5),
.C(n_6),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_486),
.Y(n_487)
);


endmodule