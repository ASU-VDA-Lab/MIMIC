module fake_jpeg_25199_n_337 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_337);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_337;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

CKINVDCx14_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

AND2x4_ASAP7_75t_L g51 ( 
.A(n_35),
.B(n_41),
.Y(n_51)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_34),
.Y(n_37)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_37),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_34),
.Y(n_38)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_34),
.Y(n_39)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_40),
.Y(n_61)
);

BUFx4f_ASAP7_75t_SL g41 ( 
.A(n_17),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_41),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g42 ( 
.A(n_20),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_27),
.Y(n_44)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_16),
.Y(n_45)
);

INVx2_ASAP7_75t_SL g56 ( 
.A(n_45),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_35),
.B(n_18),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_47),
.B(n_53),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_33),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_64),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_45),
.A2(n_27),
.B1(n_19),
.B2(n_31),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_45),
.B1(n_35),
.B2(n_36),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_51),
.B(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_27),
.B1(n_18),
.B2(n_30),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_52),
.A2(n_30),
.B1(n_23),
.B2(n_25),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_41),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_41),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_57),
.B(n_60),
.Y(n_82)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_58),
.Y(n_67)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_67),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_SL g113 ( 
.A(n_68),
.B(n_55),
.C(n_54),
.Y(n_113)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_69),
.B(n_70),
.Y(n_111)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_59),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_71),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_51),
.B(n_37),
.C(n_40),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_83),
.C(n_60),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_50),
.A2(n_35),
.B1(n_36),
.B2(n_43),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_73),
.A2(n_77),
.B1(n_84),
.B2(n_90),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_63),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_74),
.B(n_75),
.Y(n_121)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_59),
.Y(n_76)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_47),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_78),
.A2(n_81),
.B1(n_95),
.B2(n_29),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g80 ( 
.A(n_65),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_58),
.A2(n_36),
.B1(n_43),
.B2(n_28),
.Y(n_81)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_51),
.B(n_38),
.C(n_40),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_58),
.A2(n_19),
.B1(n_31),
.B2(n_16),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_85),
.B(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_52),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_86),
.B(n_89),
.Y(n_98)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_87),
.Y(n_112)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_66),
.Y(n_88)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_63),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g90 ( 
.A1(n_54),
.A2(n_43),
.B1(n_23),
.B2(n_22),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_66),
.Y(n_91)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_91),
.Y(n_125)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_61),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_66),
.Y(n_94)
);

HB1xp67_ASAP7_75t_L g103 ( 
.A(n_94),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_53),
.A2(n_25),
.B1(n_29),
.B2(n_33),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g96 ( 
.A(n_62),
.Y(n_96)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_96),
.Y(n_120)
);

AO21x1_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_85),
.B(n_79),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_75),
.A2(n_28),
.B(n_22),
.Y(n_101)
);

AOI21xp5_ASAP7_75t_L g134 ( 
.A1(n_101),
.A2(n_104),
.B(n_77),
.Y(n_134)
);

OA22x2_ASAP7_75t_L g102 ( 
.A1(n_97),
.A2(n_54),
.B1(n_56),
.B2(n_61),
.Y(n_102)
);

AO22x1_ASAP7_75t_L g142 ( 
.A1(n_102),
.A2(n_56),
.B1(n_55),
.B2(n_48),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g149 ( 
.A1(n_105),
.A2(n_94),
.B1(n_71),
.B2(n_20),
.Y(n_149)
);

BUFx8_ASAP7_75t_L g107 ( 
.A(n_96),
.Y(n_107)
);

INVxp67_ASAP7_75t_L g131 ( 
.A(n_107),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_110),
.B(n_118),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_113),
.A2(n_73),
.B1(n_68),
.B2(n_90),
.Y(n_138)
);

NAND2xp33_ASAP7_75t_SL g114 ( 
.A(n_97),
.B(n_42),
.Y(n_114)
);

NAND2x1p5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_81),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g116 ( 
.A(n_69),
.B(n_64),
.Y(n_116)
);

A2O1A1O1Ixp25_ASAP7_75t_L g135 ( 
.A1(n_116),
.A2(n_124),
.B(n_126),
.C(n_83),
.D(n_72),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_74),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_117),
.B(n_123),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_79),
.B(n_57),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_82),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_67),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_86),
.A2(n_56),
.B1(n_55),
.B2(n_19),
.Y(n_124)
);

AOI32xp33_ASAP7_75t_L g126 ( 
.A1(n_92),
.A2(n_42),
.A3(n_46),
.B1(n_40),
.B2(n_39),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_103),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_127),
.B(n_128),
.Y(n_159)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_98),
.Y(n_128)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_130),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_132),
.B(n_144),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_139),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g166 ( 
.A1(n_134),
.A2(n_135),
.B(n_136),
.Y(n_166)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_117),
.Y(n_137)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_137),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_138),
.A2(n_143),
.B1(n_152),
.B2(n_136),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_119),
.B(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_108),
.Y(n_140)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_141),
.Y(n_171)
);

O2A1O1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_142),
.A2(n_113),
.B(n_106),
.C(n_123),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_115),
.A2(n_82),
.B1(n_76),
.B2(n_70),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_98),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_111),
.B(n_89),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_154),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_118),
.A2(n_87),
.B1(n_91),
.B2(n_88),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_147),
.A2(n_151),
.B1(n_155),
.B2(n_122),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_104),
.B(n_80),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_148),
.B(n_150),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_149),
.A2(n_120),
.B1(n_106),
.B2(n_125),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_116),
.B(n_67),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_71),
.B1(n_40),
.B2(n_39),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_115),
.A2(n_44),
.B1(n_39),
.B2(n_31),
.Y(n_152)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_99),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_153),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_105),
.B(n_19),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_124),
.A2(n_44),
.B1(n_31),
.B2(n_16),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_93),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_156),
.B(n_46),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_121),
.C(n_114),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_158),
.B(n_185),
.C(n_188),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_162),
.A2(n_164),
.B1(n_168),
.B2(n_174),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_145),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g200 ( 
.A(n_165),
.B(n_180),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_150),
.B(n_101),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_167),
.B(n_183),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_148),
.A2(n_102),
.B1(n_126),
.B2(n_109),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_136),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_170),
.B(n_181),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_138),
.A2(n_102),
.B1(n_109),
.B2(n_112),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_176),
.B(n_177),
.Y(n_222)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_151),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_129),
.B(n_102),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_178),
.B(n_62),
.Y(n_205)
);

NAND3xp33_ASAP7_75t_L g180 ( 
.A(n_139),
.B(n_15),
.C(n_13),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_102),
.B1(n_112),
.B2(n_122),
.Y(n_182)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_182),
.A2(n_184),
.B1(n_190),
.B2(n_152),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_134),
.B(n_133),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_147),
.A2(n_125),
.B1(n_120),
.B2(n_44),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_132),
.B(n_48),
.C(n_42),
.Y(n_185)
);

AO22x1_ASAP7_75t_L g186 ( 
.A1(n_142),
.A2(n_48),
.B1(n_107),
.B2(n_16),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_189),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_137),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_187),
.B(n_32),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_143),
.B(n_62),
.C(n_63),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_155),
.A2(n_107),
.B1(n_46),
.B2(n_21),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_142),
.B(n_21),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_191),
.B(n_26),
.Y(n_218)
);

NAND2x1_ASAP7_75t_L g194 ( 
.A(n_170),
.B(n_131),
.Y(n_194)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_194),
.A2(n_186),
.B(n_171),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_196),
.A2(n_202),
.B1(n_207),
.B2(n_221),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_178),
.B(n_127),
.C(n_130),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_197),
.B(n_185),
.C(n_168),
.Y(n_231)
);

INVx2_ASAP7_75t_L g199 ( 
.A(n_160),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_199),
.B(n_209),
.Y(n_244)
);

XOR2x2_ASAP7_75t_SL g201 ( 
.A(n_166),
.B(n_131),
.Y(n_201)
);

XNOR2xp5_ASAP7_75t_SL g223 ( 
.A(n_201),
.B(n_205),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_153),
.B1(n_141),
.B2(n_140),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_166),
.A2(n_107),
.B(n_32),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_212),
.B(n_172),
.Y(n_234)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_206),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_21),
.B1(n_26),
.B2(n_24),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx5_ASAP7_75t_L g210 ( 
.A(n_179),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_210),
.A2(n_220),
.B1(n_171),
.B2(n_186),
.Y(n_232)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_159),
.Y(n_211)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_211),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g212 ( 
.A1(n_173),
.A2(n_32),
.B(n_1),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_163),
.Y(n_213)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_213),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_157),
.B(n_32),
.Y(n_214)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_214),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_21),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g229 ( 
.A(n_215),
.B(n_219),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_161),
.B(n_26),
.Y(n_216)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_216),
.Y(n_237)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_169),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_167),
.B(n_24),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_184),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_162),
.A2(n_24),
.B1(n_1),
.B2(n_2),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_203),
.A2(n_173),
.B1(n_181),
.B2(n_191),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_224),
.A2(n_225),
.B1(n_248),
.B2(n_207),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_203),
.A2(n_176),
.B1(n_188),
.B2(n_164),
.Y(n_225)
);

XNOR2x1_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_158),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_SL g251 ( 
.A(n_230),
.B(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_246),
.C(n_195),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_232),
.B(n_202),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_234),
.B(n_221),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g235 ( 
.A(n_208),
.B(n_157),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g257 ( 
.A1(n_239),
.A2(n_243),
.B(n_245),
.Y(n_257)
);

HB1xp67_ASAP7_75t_L g240 ( 
.A(n_222),
.Y(n_240)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_240),
.Y(n_249)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_208),
.B(n_190),
.Y(n_242)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_242),
.B(n_247),
.Y(n_250)
);

A2O1A1Ixp33_ASAP7_75t_SL g243 ( 
.A1(n_194),
.A2(n_0),
.B(n_1),
.C(n_2),
.Y(n_243)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_194),
.A2(n_0),
.B(n_2),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_195),
.B(n_15),
.C(n_13),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g247 ( 
.A(n_205),
.B(n_13),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_198),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_244),
.Y(n_252)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_252),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_223),
.B(n_197),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_253),
.B(n_262),
.Y(n_276)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_254),
.B(n_263),
.C(n_255),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_215),
.C(n_219),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_255),
.B(n_259),
.C(n_260),
.Y(n_273)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_256),
.B(n_265),
.Y(n_271)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_233),
.Y(n_258)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_258),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g259 ( 
.A(n_229),
.B(n_222),
.C(n_204),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_193),
.C(n_196),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_233),
.Y(n_261)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_261),
.Y(n_285)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_223),
.B(n_212),
.Y(n_262)
);

XOR2xp5_ASAP7_75t_L g263 ( 
.A(n_230),
.B(n_192),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_SL g264 ( 
.A(n_235),
.B(n_192),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_SL g275 ( 
.A(n_264),
.B(n_234),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_266),
.A2(n_269),
.B1(n_225),
.B2(n_224),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_238),
.B(n_199),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g279 ( 
.A(n_267),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_218),
.C(n_210),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_268),
.B(n_246),
.C(n_247),
.Y(n_274)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_274),
.C(n_273),
.Y(n_298)
);

CKINVDCx14_ASAP7_75t_R g299 ( 
.A(n_272),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_SL g289 ( 
.A(n_275),
.B(n_262),
.Y(n_289)
);

AOI22xp5_ASAP7_75t_L g278 ( 
.A1(n_249),
.A2(n_227),
.B1(n_228),
.B2(n_241),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_278),
.B(n_282),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g280 ( 
.A(n_254),
.B(n_236),
.C(n_226),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_280),
.B(n_283),
.Y(n_287)
);

HB1xp67_ASAP7_75t_L g281 ( 
.A(n_268),
.Y(n_281)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_281),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_237),
.B1(n_200),
.B2(n_245),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_253),
.B(n_243),
.C(n_15),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_250),
.B(n_243),
.C(n_4),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_286),
.B(n_3),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_273),
.B(n_250),
.C(n_259),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_289),
.C(n_290),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g303 ( 
.A(n_289),
.B(n_290),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_263),
.Y(n_290)
);

NAND3xp33_ASAP7_75t_L g291 ( 
.A(n_277),
.B(n_257),
.C(n_265),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_291),
.B(n_294),
.Y(n_305)
);

A2O1A1Ixp33_ASAP7_75t_L g292 ( 
.A1(n_271),
.A2(n_264),
.B(n_251),
.C(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_292),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_271),
.A2(n_251),
.B1(n_4),
.B2(n_5),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g308 ( 
.A1(n_293),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_SL g294 ( 
.A(n_274),
.B(n_3),
.Y(n_294)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_295),
.Y(n_313)
);

INVxp33_ASAP7_75t_SL g297 ( 
.A(n_279),
.Y(n_297)
);

AOI22xp33_ASAP7_75t_SL g307 ( 
.A1(n_297),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_298),
.B(n_301),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_281),
.B(n_4),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_SL g302 ( 
.A1(n_287),
.A2(n_285),
.B(n_284),
.Y(n_302)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_302),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_291),
.A2(n_276),
.B(n_279),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g317 ( 
.A1(n_304),
.A2(n_307),
.B1(n_310),
.B2(n_292),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_308),
.B(n_312),
.Y(n_314)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_6),
.B(n_7),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_296),
.B(n_7),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_12),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_SL g316 ( 
.A1(n_305),
.A2(n_300),
.B(n_299),
.Y(n_316)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_316),
.A2(n_303),
.B(n_307),
.Y(n_326)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_317),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_306),
.A2(n_288),
.B1(n_9),
.B2(n_10),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_318),
.B(n_319),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_309),
.B(n_8),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_312),
.B(n_9),
.C(n_10),
.Y(n_320)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_320),
.B(n_321),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_304),
.B(n_11),
.C(n_12),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_322),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_SL g324 ( 
.A1(n_315),
.A2(n_313),
.B(n_310),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_324),
.B(n_326),
.Y(n_331)
);

INVxp67_ASAP7_75t_L g329 ( 
.A(n_328),
.Y(n_329)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_329),
.A2(n_330),
.B(n_314),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_327),
.B(n_318),
.Y(n_330)
);

NOR3xp33_ASAP7_75t_L g333 ( 
.A(n_332),
.B(n_331),
.C(n_323),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_333),
.A2(n_325),
.B(n_320),
.Y(n_334)
);

AOI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_334),
.A2(n_317),
.B(n_321),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_335),
.B(n_303),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g337 ( 
.A1(n_336),
.A2(n_12),
.B(n_334),
.Y(n_337)
);


endmodule