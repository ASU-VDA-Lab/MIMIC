module fake_jpeg_25636_n_38 (n_3, n_2, n_1, n_0, n_4, n_5, n_38);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_38;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_34;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx4_ASAP7_75t_SL g6 ( 
.A(n_4),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_2),
.B(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

AND2x2_ASAP7_75t_SL g10 ( 
.A(n_0),
.B(n_1),
.Y(n_10)
);

INVx1_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_0),
.Y(n_12)
);

AND2x2_ASAP7_75t_L g13 ( 
.A(n_7),
.B(n_10),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g22 ( 
.A(n_13),
.B(n_14),
.Y(n_22)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_L g24 ( 
.A1(n_15),
.A2(n_17),
.B1(n_19),
.B2(n_6),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g21 ( 
.A1(n_16),
.A2(n_18),
.B1(n_11),
.B2(n_12),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_10),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_9),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g20 ( 
.A1(n_14),
.A2(n_10),
.B1(n_8),
.B2(n_6),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_20),
.A2(n_23),
.B1(n_13),
.B2(n_18),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_21),
.A2(n_24),
.B1(n_3),
.B2(n_5),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_16),
.A2(n_6),
.B1(n_12),
.B2(n_9),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g31 ( 
.A1(n_25),
.A2(n_27),
.B1(n_28),
.B2(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_22),
.B(n_13),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_26),
.B(n_20),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_23),
.A2(n_15),
.B1(n_9),
.B2(n_5),
.Y(n_27)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_26),
.A2(n_22),
.B(n_21),
.Y(n_29)
);

OAI21xp33_ASAP7_75t_L g32 ( 
.A1(n_29),
.A2(n_30),
.B(n_31),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_29),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_25),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_34),
.B(n_35),
.Y(n_36)
);

AND2x2_ASAP7_75t_L g35 ( 
.A(n_32),
.B(n_28),
.Y(n_35)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_36),
.B(n_35),
.C(n_27),
.Y(n_37)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_37),
.A2(n_21),
.B1(n_3),
.B2(n_5),
.Y(n_38)
);


endmodule