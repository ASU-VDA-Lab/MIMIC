module fake_jpeg_26770_n_173 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_173);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_173;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx3_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_8),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_6),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_13),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_20),
.B(n_0),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_33),
.B(n_34),
.Y(n_49)
);

HAxp5_ASAP7_75t_SL g34 ( 
.A(n_32),
.B(n_1),
.CON(n_34),
.SN(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_21),
.Y(n_35)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_21),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_21),
.B(n_1),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_38),
.B(n_30),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_16),
.Y(n_39)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

HAxp5_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_1),
.CON(n_41),
.SN(n_41)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_41),
.B(n_2),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g42 ( 
.A(n_30),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_42),
.B(n_26),
.Y(n_52)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_43),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g44 ( 
.A(n_36),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_40),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

HB1xp67_ASAP7_75t_L g46 ( 
.A(n_38),
.Y(n_46)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_55),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_23),
.Y(n_67)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_57),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_43),
.B(n_19),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_58),
.B(n_59),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_39),
.B(n_30),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_17),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_60),
.B(n_23),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_40),
.A2(n_16),
.B1(n_25),
.B2(n_20),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_61),
.A2(n_25),
.B1(n_19),
.B2(n_29),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_39),
.B(n_29),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_22),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_67),
.Y(n_86)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_76),
.B1(n_77),
.B2(n_50),
.Y(n_89)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

OAI21xp33_ASAP7_75t_L g92 ( 
.A1(n_72),
.A2(n_73),
.B(n_82),
.Y(n_92)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_55),
.A2(n_28),
.B(n_27),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g87 ( 
.A(n_74),
.B(n_58),
.Y(n_87)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_63),
.Y(n_75)
);

INVx11_ASAP7_75t_L g95 ( 
.A(n_75),
.Y(n_95)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_51),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g77 ( 
.A1(n_56),
.A2(n_18),
.B1(n_22),
.B2(n_27),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_78),
.B(n_83),
.Y(n_103)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_44),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_79),
.B(n_80),
.Y(n_85)
);

INVxp33_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_62),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_49),
.B(n_17),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_84),
.B(n_49),
.Y(n_90)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_87),
.Y(n_112)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_88),
.B(n_91),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_97),
.B1(n_86),
.B2(n_94),
.Y(n_107)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_81),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_96),
.Y(n_113)
);

OAI32xp33_ASAP7_75t_L g94 ( 
.A1(n_66),
.A2(n_50),
.A3(n_28),
.B1(n_57),
.B2(n_47),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g114 ( 
.A(n_94),
.B(n_99),
.Y(n_114)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_83),
.Y(n_96)
);

AOI22x1_ASAP7_75t_SL g97 ( 
.A1(n_66),
.A2(n_35),
.B1(n_37),
.B2(n_26),
.Y(n_97)
);

OA21x2_ASAP7_75t_SL g111 ( 
.A1(n_97),
.A2(n_102),
.B(n_99),
.Y(n_111)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_81),
.Y(n_98)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_72),
.B(n_36),
.C(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_69),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_102),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_70),
.A2(n_37),
.B(n_36),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_82),
.B(n_18),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_104),
.B(n_81),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_96),
.A2(n_70),
.B1(n_65),
.B2(n_47),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_105),
.A2(n_108),
.B1(n_118),
.B2(n_4),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_95),
.B1(n_100),
.B2(n_53),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_103),
.A2(n_65),
.B1(n_73),
.B2(n_69),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g109 ( 
.A(n_95),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_109),
.B(n_54),
.Y(n_128)
);

AOI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_111),
.A2(n_100),
.B1(n_53),
.B2(n_24),
.Y(n_130)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_85),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_116),
.B(n_120),
.Y(n_137)
);

XOR2xp5_ASAP7_75t_L g117 ( 
.A(n_87),
.B(n_64),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g124 ( 
.A(n_117),
.B(n_119),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_103),
.A2(n_64),
.B1(n_79),
.B2(n_74),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_104),
.B(n_48),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_88),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_121),
.B(n_122),
.Y(n_123)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_115),
.A2(n_98),
.B1(n_93),
.B2(n_48),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g142 ( 
.A1(n_125),
.A2(n_127),
.B(n_134),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_112),
.B(n_92),
.C(n_90),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_126),
.B(n_119),
.C(n_118),
.Y(n_141)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_91),
.B(n_54),
.Y(n_127)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_128),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_129),
.A2(n_108),
.B1(n_115),
.B2(n_105),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_130),
.B(n_132),
.Y(n_146)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_110),
.Y(n_131)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_131),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_45),
.Y(n_132)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_132),
.Y(n_147)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_113),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g134 ( 
.A1(n_114),
.A2(n_2),
.B(n_3),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_114),
.A2(n_3),
.B(n_4),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_SL g140 ( 
.A(n_135),
.B(n_117),
.Y(n_140)
);

OR2x2_ASAP7_75t_L g144 ( 
.A(n_136),
.B(n_107),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_137),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_139),
.B(n_148),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g150 ( 
.A1(n_140),
.A2(n_146),
.B(n_130),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_141),
.B(n_124),
.C(n_126),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g155 ( 
.A1(n_145),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_123),
.Y(n_148)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_149),
.B(n_152),
.C(n_156),
.Y(n_161)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_150),
.A2(n_142),
.B(n_151),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_141),
.B(n_124),
.C(n_127),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_146),
.A2(n_133),
.B1(n_136),
.B2(n_122),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_153),
.A2(n_154),
.B1(n_155),
.B2(n_145),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g154 ( 
.A1(n_142),
.A2(n_135),
.B1(n_134),
.B2(n_109),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_140),
.B(n_10),
.C(n_14),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g163 ( 
.A(n_157),
.B(n_147),
.Y(n_163)
);

OR2x2_ASAP7_75t_L g165 ( 
.A(n_158),
.B(n_5),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_152),
.B(n_149),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_159),
.B(n_160),
.Y(n_166)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_156),
.A2(n_146),
.B(n_144),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_143),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_162),
.B(n_143),
.C(n_138),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_163),
.B(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_165),
.B(n_11),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g170 ( 
.A(n_168),
.B(n_15),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g169 ( 
.A(n_167),
.B(n_166),
.Y(n_169)
);

OAI21x1_ASAP7_75t_L g171 ( 
.A1(n_169),
.A2(n_170),
.B(n_161),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_171),
.B(n_15),
.Y(n_172)
);

BUFx24_ASAP7_75t_SL g173 ( 
.A(n_172),
.Y(n_173)
);


endmodule