module fake_aes_12448_n_36 (n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_36);
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_36;
wire n_20;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_11;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_33;
wire n_30;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
INVx2_ASAP7_75t_L g11 ( .A(n_5), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_0), .Y(n_12) );
INVx2_ASAP7_75t_L g13 ( .A(n_1), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_7), .B(n_9), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_6), .Y(n_15) );
INVx2_ASAP7_75t_SL g16 ( .A(n_11), .Y(n_16) );
NAND2xp5_ASAP7_75t_L g17 ( .A(n_13), .B(n_0), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_15), .B(n_1), .Y(n_18) );
OR2x6_ASAP7_75t_L g19 ( .A(n_16), .B(n_14), .Y(n_19) );
O2A1O1Ixp5_ASAP7_75t_L g20 ( .A1(n_17), .A2(n_14), .B(n_12), .C(n_10), .Y(n_20) );
INVx2_ASAP7_75t_SL g21 ( .A(n_19), .Y(n_21) );
OR2x2_ASAP7_75t_L g22 ( .A(n_19), .B(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx1_ASAP7_75t_L g24 ( .A(n_22), .Y(n_24) );
INVxp67_ASAP7_75t_SL g25 ( .A(n_24), .Y(n_25) );
NAND2xp5_ASAP7_75t_L g26 ( .A(n_23), .B(n_19), .Y(n_26) );
AOI22xp5_ASAP7_75t_L g27 ( .A1(n_25), .A2(n_23), .B1(n_12), .B2(n_20), .Y(n_27) );
AOI22xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_12), .B1(n_3), .B2(n_4), .Y(n_28) );
INVx2_ASAP7_75t_SL g29 ( .A(n_26), .Y(n_29) );
AND2x4_ASAP7_75t_L g30 ( .A(n_29), .B(n_2), .Y(n_30) );
AND2x2_ASAP7_75t_L g31 ( .A(n_28), .B(n_2), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_27), .B(n_3), .Y(n_32) );
NAND3xp33_ASAP7_75t_L g33 ( .A(n_31), .B(n_4), .C(n_5), .Y(n_33) );
AOI21xp5_ASAP7_75t_L g34 ( .A1(n_32), .A2(n_6), .B(n_7), .Y(n_34) );
OAI22xp5_ASAP7_75t_L g35 ( .A1(n_33), .A2(n_30), .B1(n_31), .B2(n_8), .Y(n_35) );
AOI22x1_ASAP7_75t_L g36 ( .A1(n_35), .A2(n_30), .B1(n_34), .B2(n_8), .Y(n_36) );
endmodule