module fake_netlist_5_520_n_1533 (n_137, n_294, n_318, n_82, n_194, n_316, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_61, n_127, n_75, n_235, n_226, n_74, n_57, n_111, n_155, n_43, n_116, n_22, n_284, n_46, n_245, n_21, n_139, n_38, n_105, n_280, n_4, n_17, n_254, n_33, n_23, n_302, n_265, n_293, n_244, n_47, n_173, n_198, n_247, n_314, n_8, n_321, n_292, n_100, n_212, n_119, n_275, n_252, n_26, n_295, n_133, n_330, n_2, n_6, n_39, n_147, n_67, n_307, n_87, n_150, n_106, n_209, n_259, n_301, n_68, n_93, n_186, n_134, n_191, n_51, n_63, n_171, n_153, n_341, n_204, n_250, n_260, n_298, n_320, n_286, n_122, n_282, n_331, n_10, n_24, n_325, n_132, n_90, n_101, n_281, n_240, n_189, n_220, n_291, n_231, n_257, n_31, n_13, n_152, n_317, n_9, n_323, n_195, n_42, n_227, n_45, n_271, n_94, n_335, n_123, n_167, n_234, n_343, n_308, n_267, n_297, n_156, n_5, n_225, n_219, n_157, n_131, n_192, n_223, n_158, n_138, n_264, n_109, n_163, n_276, n_339, n_95, n_183, n_185, n_243, n_347, n_169, n_59, n_255, n_215, n_196, n_211, n_218, n_181, n_3, n_290, n_221, n_178, n_287, n_344, n_72, n_104, n_41, n_56, n_141, n_15, n_336, n_145, n_48, n_50, n_337, n_313, n_88, n_216, n_168, n_164, n_311, n_208, n_142, n_214, n_328, n_140, n_299, n_303, n_296, n_241, n_184, n_65, n_78, n_144, n_114, n_96, n_165, n_213, n_129, n_342, n_98, n_197, n_107, n_69, n_236, n_1, n_249, n_304, n_329, n_203, n_274, n_80, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_333, n_309, n_30, n_14, n_84, n_130, n_322, n_258, n_29, n_79, n_151, n_25, n_306, n_288, n_188, n_190, n_201, n_263, n_44, n_224, n_40, n_34, n_228, n_283, n_112, n_85, n_239, n_55, n_49, n_310, n_54, n_12, n_76, n_170, n_332, n_27, n_77, n_102, n_161, n_273, n_270, n_230, n_81, n_118, n_279, n_70, n_253, n_261, n_174, n_289, n_172, n_206, n_217, n_312, n_345, n_210, n_91, n_176, n_182, n_143, n_83, n_237, n_180, n_340, n_207, n_37, n_346, n_229, n_108, n_66, n_177, n_60, n_16, n_0, n_58, n_18, n_117, n_326, n_233, n_205, n_113, n_246, n_179, n_125, n_269, n_128, n_285, n_120, n_232, n_327, n_135, n_126, n_202, n_266, n_272, n_193, n_251, n_53, n_160, n_154, n_62, n_148, n_71, n_300, n_159, n_334, n_175, n_262, n_238, n_99, n_319, n_20, n_121, n_242, n_36, n_200, n_162, n_64, n_222, n_28, n_89, n_115, n_324, n_199, n_187, n_32, n_103, n_348, n_97, n_166, n_11, n_7, n_256, n_305, n_52, n_278, n_110, n_1533);

input n_137;
input n_294;
input n_318;
input n_82;
input n_194;
input n_316;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_61;
input n_127;
input n_75;
input n_235;
input n_226;
input n_74;
input n_57;
input n_111;
input n_155;
input n_43;
input n_116;
input n_22;
input n_284;
input n_46;
input n_245;
input n_21;
input n_139;
input n_38;
input n_105;
input n_280;
input n_4;
input n_17;
input n_254;
input n_33;
input n_23;
input n_302;
input n_265;
input n_293;
input n_244;
input n_47;
input n_173;
input n_198;
input n_247;
input n_314;
input n_8;
input n_321;
input n_292;
input n_100;
input n_212;
input n_119;
input n_275;
input n_252;
input n_26;
input n_295;
input n_133;
input n_330;
input n_2;
input n_6;
input n_39;
input n_147;
input n_67;
input n_307;
input n_87;
input n_150;
input n_106;
input n_209;
input n_259;
input n_301;
input n_68;
input n_93;
input n_186;
input n_134;
input n_191;
input n_51;
input n_63;
input n_171;
input n_153;
input n_341;
input n_204;
input n_250;
input n_260;
input n_298;
input n_320;
input n_286;
input n_122;
input n_282;
input n_331;
input n_10;
input n_24;
input n_325;
input n_132;
input n_90;
input n_101;
input n_281;
input n_240;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_31;
input n_13;
input n_152;
input n_317;
input n_9;
input n_323;
input n_195;
input n_42;
input n_227;
input n_45;
input n_271;
input n_94;
input n_335;
input n_123;
input n_167;
input n_234;
input n_343;
input n_308;
input n_267;
input n_297;
input n_156;
input n_5;
input n_225;
input n_219;
input n_157;
input n_131;
input n_192;
input n_223;
input n_158;
input n_138;
input n_264;
input n_109;
input n_163;
input n_276;
input n_339;
input n_95;
input n_183;
input n_185;
input n_243;
input n_347;
input n_169;
input n_59;
input n_255;
input n_215;
input n_196;
input n_211;
input n_218;
input n_181;
input n_3;
input n_290;
input n_221;
input n_178;
input n_287;
input n_344;
input n_72;
input n_104;
input n_41;
input n_56;
input n_141;
input n_15;
input n_336;
input n_145;
input n_48;
input n_50;
input n_337;
input n_313;
input n_88;
input n_216;
input n_168;
input n_164;
input n_311;
input n_208;
input n_142;
input n_214;
input n_328;
input n_140;
input n_299;
input n_303;
input n_296;
input n_241;
input n_184;
input n_65;
input n_78;
input n_144;
input n_114;
input n_96;
input n_165;
input n_213;
input n_129;
input n_342;
input n_98;
input n_197;
input n_107;
input n_69;
input n_236;
input n_1;
input n_249;
input n_304;
input n_329;
input n_203;
input n_274;
input n_80;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_333;
input n_309;
input n_30;
input n_14;
input n_84;
input n_130;
input n_322;
input n_258;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_288;
input n_188;
input n_190;
input n_201;
input n_263;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_112;
input n_85;
input n_239;
input n_55;
input n_49;
input n_310;
input n_54;
input n_12;
input n_76;
input n_170;
input n_332;
input n_27;
input n_77;
input n_102;
input n_161;
input n_273;
input n_270;
input n_230;
input n_81;
input n_118;
input n_279;
input n_70;
input n_253;
input n_261;
input n_174;
input n_289;
input n_172;
input n_206;
input n_217;
input n_312;
input n_345;
input n_210;
input n_91;
input n_176;
input n_182;
input n_143;
input n_83;
input n_237;
input n_180;
input n_340;
input n_207;
input n_37;
input n_346;
input n_229;
input n_108;
input n_66;
input n_177;
input n_60;
input n_16;
input n_0;
input n_58;
input n_18;
input n_117;
input n_326;
input n_233;
input n_205;
input n_113;
input n_246;
input n_179;
input n_125;
input n_269;
input n_128;
input n_285;
input n_120;
input n_232;
input n_327;
input n_135;
input n_126;
input n_202;
input n_266;
input n_272;
input n_193;
input n_251;
input n_53;
input n_160;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_159;
input n_334;
input n_175;
input n_262;
input n_238;
input n_99;
input n_319;
input n_20;
input n_121;
input n_242;
input n_36;
input n_200;
input n_162;
input n_64;
input n_222;
input n_28;
input n_89;
input n_115;
input n_324;
input n_199;
input n_187;
input n_32;
input n_103;
input n_348;
input n_97;
input n_166;
input n_11;
input n_7;
input n_256;
input n_305;
input n_52;
input n_278;
input n_110;

output n_1533;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1166;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1150;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1021;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1353;
wire n_800;
wire n_1347;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_864;
wire n_859;
wire n_951;
wire n_1264;
wire n_447;
wire n_1494;
wire n_625;
wire n_854;
wire n_1462;
wire n_674;
wire n_417;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_606;
wire n_877;
wire n_755;
wire n_1118;
wire n_947;
wire n_1285;
wire n_373;
wire n_1359;
wire n_530;
wire n_1107;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_929;
wire n_1124;
wire n_902;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1261;
wire n_938;
wire n_1098;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_1236;
wire n_569;
wire n_920;
wire n_1289;
wire n_1517;
wire n_370;
wire n_976;
wire n_1449;
wire n_1078;
wire n_775;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_955;
wire n_1146;
wire n_882;
wire n_1036;
wire n_1097;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_1040;
wire n_578;
wire n_926;
wire n_1218;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1030;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_496;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_521;
wire n_845;
wire n_663;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_680;
wire n_1473;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_675;
wire n_888;
wire n_1167;
wire n_637;
wire n_1384;
wire n_446;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_468;
wire n_464;
wire n_363;
wire n_1069;
wire n_1075;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_477;
wire n_571;
wire n_461;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_907;
wire n_1447;
wire n_1377;
wire n_989;
wire n_1039;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_838;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1248;
wire n_1331;
wire n_953;
wire n_1014;
wire n_1241;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_476;
wire n_1527;
wire n_534;
wire n_884;
wire n_944;
wire n_647;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_561;
wire n_1319;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_728;
wire n_1162;
wire n_1199;
wire n_352;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_887;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1481;
wire n_434;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1293;
wire n_965;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_759;
wire n_806;
wire n_1477;
wire n_1189;
wire n_1259;
wire n_706;
wire n_746;
wire n_747;
wire n_784;
wire n_1244;
wire n_431;
wire n_1194;
wire n_615;
wire n_851;
wire n_843;
wire n_523;
wire n_913;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_776;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1128;
wire n_744;
wire n_590;
wire n_629;
wire n_1308;
wire n_1233;
wire n_1529;
wire n_526;
wire n_372;
wire n_677;
wire n_1333;
wire n_1121;
wire n_368;
wire n_604;
wire n_433;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_689;
wire n_738;
wire n_640;
wire n_1510;
wire n_624;
wire n_1380;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_610;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_448;
wire n_758;
wire n_999;
wire n_1158;
wire n_1509;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1306;
wire n_1068;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_658;
wire n_1362;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_592;
wire n_1169;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1269;
wire n_1095;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_374;
wire n_396;
wire n_1383;
wire n_1073;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_723;
wire n_1065;
wire n_1336;
wire n_473;
wire n_1309;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_614;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_743;
wire n_613;
wire n_1119;
wire n_1240;
wire n_829;
wire n_1416;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1006;
wire n_1270;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_512;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1349;
wire n_1093;
wire n_1031;
wire n_609;
wire n_1041;
wire n_1265;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_630;
wire n_504;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1455;
wire n_767;
wire n_993;
wire n_1407;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_729;
wire n_1131;
wire n_1084;
wire n_970;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_1209;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_572;
wire n_366;
wire n_815;
wire n_1381;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_426;
wire n_1438;
wire n_1082;
wire n_589;
wire n_716;
wire n_562;
wire n_1436;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_531;
wire n_890;
wire n_764;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_1252;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_950;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1060;
wire n_1141;
wire n_389;
wire n_418;
wire n_912;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_983;
wire n_1305;
wire n_873;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_690;
wire n_583;
wire n_1343;
wire n_1203;
wire n_821;
wire n_1179;
wire n_621;
wire n_753;
wire n_455;
wire n_1048;
wire n_1288;
wire n_385;
wire n_507;
wire n_1228;
wire n_972;
wire n_692;
wire n_820;
wire n_1200;
wire n_1301;
wire n_1363;
wire n_1185;
wire n_991;
wire n_828;
wire n_779;
wire n_576;
wire n_1143;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_992;
wire n_543;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_883;
wire n_470;
wire n_449;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_918;
wire n_942;
wire n_1147;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_356;
wire n_894;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1470;
wire n_1096;
wire n_833;
wire n_1307;
wire n_988;
wire n_814;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_387;
wire n_1149;
wire n_398;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_1219;
wire n_1204;
wire n_1035;
wire n_555;
wire n_783;
wire n_1188;
wire n_661;
wire n_849;
wire n_584;
wire n_681;
wire n_430;
wire n_510;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_875;
wire n_357;
wire n_1110;
wire n_445;
wire n_749;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1419;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1389;
wire n_975;
wire n_1256;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1164;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_876;
wire n_1516;
wire n_1190;
wire n_601;
wire n_917;
wire n_966;
wire n_1116;
wire n_1212;
wire n_726;
wire n_982;
wire n_1453;
wire n_818;
wire n_861;
wire n_1183;
wire n_899;
wire n_1253;
wire n_774;
wire n_1335;
wire n_1514;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_665;
wire n_1440;
wire n_421;
wire n_1356;
wire n_910;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_735;
wire n_1109;
wire n_895;
wire n_1310;
wire n_427;
wire n_1399;
wire n_791;
wire n_732;
wire n_808;
wire n_797;
wire n_1025;
wire n_500;
wire n_1067;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1155;
wire n_1418;
wire n_1524;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1352;
wire n_626;
wire n_1144;
wire n_1137;
wire n_1170;
wire n_676;
wire n_653;
wire n_642;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_664;
wire n_503;
wire n_1372;
wire n_605;
wire n_1273;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_501;
wire n_823;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_581;
wire n_382;
wire n_554;
wire n_898;
wire n_1013;
wire n_1452;
wire n_718;
wire n_1120;
wire n_719;
wire n_443;
wire n_714;
wire n_909;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_508;
wire n_506;
wire n_1320;
wire n_737;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1281;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_733;
wire n_1489;
wire n_1376;
wire n_941;
wire n_981;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_518;
wire n_505;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_381;
wire n_390;
wire n_1330;
wire n_481;
wire n_769;
wire n_1046;
wire n_934;
wire n_826;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1361;
wire n_853;
wire n_377;
wire n_751;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_961;
wire n_771;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1411;
wire n_622;
wire n_1087;
wire n_386;
wire n_994;
wire n_848;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1247;
wire n_922;
wire n_816;
wire n_591;
wire n_1344;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_432;
wire n_839;
wire n_1210;
wire n_1364;
wire n_1250;
wire n_369;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1460;
wire n_772;
wire n_499;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_740;
wire n_384;
wire n_1404;
wire n_1315;
wire n_1061;
wire n_1298;
wire n_462;
wire n_1193;
wire n_1255;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1028;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1245;
wire n_846;
wire n_465;
wire n_362;
wire n_1321;
wire n_585;
wire n_616;
wire n_745;
wire n_1103;
wire n_648;
wire n_1379;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_641;
wire n_730;
wire n_1325;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1220;
wire n_437;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1526;
wire n_863;
wire n_805;
wire n_1275;
wire n_712;
wire n_1042;
wire n_1402;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1196;
wire n_651;
wire n_1340;
wire n_811;
wire n_807;
wire n_835;
wire n_666;
wire n_1433;
wire n_1254;
wire n_1026;
wire n_1234;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_1018;
wire n_438;
wire n_713;
wire n_904;
wire n_1180;
wire n_1271;
wire n_533;
wire n_1251;

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_186),
.Y(n_349)
);

INVx1_ASAP7_75t_SL g350 ( 
.A(n_19),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_325),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_160),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_85),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_196),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_40),
.Y(n_355)
);

INVx2_ASAP7_75t_SL g356 ( 
.A(n_73),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_246),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g358 ( 
.A(n_179),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_312),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_69),
.Y(n_360)
);

INVx1_ASAP7_75t_SL g361 ( 
.A(n_25),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_209),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_151),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_155),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_0),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_210),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_139),
.Y(n_367)
);

BUFx3_ASAP7_75t_L g368 ( 
.A(n_300),
.Y(n_368)
);

BUFx6f_ASAP7_75t_L g369 ( 
.A(n_22),
.Y(n_369)
);

CKINVDCx16_ASAP7_75t_R g370 ( 
.A(n_41),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_324),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_335),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_157),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_338),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_131),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_268),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_328),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_175),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_7),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_296),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_235),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_316),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_119),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_323),
.Y(n_384)
);

CKINVDCx5p33_ASAP7_75t_R g385 ( 
.A(n_244),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_285),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_337),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_19),
.Y(n_388)
);

INVx2_ASAP7_75t_L g389 ( 
.A(n_140),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_346),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_24),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_293),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_91),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_78),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_219),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_322),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_279),
.Y(n_397)
);

BUFx10_ASAP7_75t_L g398 ( 
.A(n_340),
.Y(n_398)
);

CKINVDCx14_ASAP7_75t_R g399 ( 
.A(n_149),
.Y(n_399)
);

INVxp67_ASAP7_75t_L g400 ( 
.A(n_256),
.Y(n_400)
);

CKINVDCx5p33_ASAP7_75t_R g401 ( 
.A(n_329),
.Y(n_401)
);

BUFx3_ASAP7_75t_L g402 ( 
.A(n_261),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_166),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_92),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_313),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_286),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_17),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_14),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_64),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_36),
.Y(n_410)
);

INVxp33_ASAP7_75t_L g411 ( 
.A(n_39),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_199),
.Y(n_412)
);

CKINVDCx5p33_ASAP7_75t_R g413 ( 
.A(n_259),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_105),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_35),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_333),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_242),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_318),
.Y(n_418)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_288),
.Y(n_419)
);

CKINVDCx5p33_ASAP7_75t_R g420 ( 
.A(n_233),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_320),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_113),
.Y(n_422)
);

INVx2_ASAP7_75t_SL g423 ( 
.A(n_330),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g424 ( 
.A(n_75),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_311),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_205),
.Y(n_426)
);

CKINVDCx5p33_ASAP7_75t_R g427 ( 
.A(n_240),
.Y(n_427)
);

BUFx6f_ASAP7_75t_L g428 ( 
.A(n_277),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_306),
.Y(n_429)
);

CKINVDCx16_ASAP7_75t_R g430 ( 
.A(n_295),
.Y(n_430)
);

BUFx2_ASAP7_75t_L g431 ( 
.A(n_61),
.Y(n_431)
);

CKINVDCx5p33_ASAP7_75t_R g432 ( 
.A(n_32),
.Y(n_432)
);

CKINVDCx5p33_ASAP7_75t_R g433 ( 
.A(n_211),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_227),
.Y(n_434)
);

BUFx3_ASAP7_75t_L g435 ( 
.A(n_45),
.Y(n_435)
);

CKINVDCx20_ASAP7_75t_R g436 ( 
.A(n_265),
.Y(n_436)
);

BUFx2_ASAP7_75t_L g437 ( 
.A(n_249),
.Y(n_437)
);

CKINVDCx5p33_ASAP7_75t_R g438 ( 
.A(n_224),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_184),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_291),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_228),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_117),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_342),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_189),
.Y(n_444)
);

CKINVDCx5p33_ASAP7_75t_R g445 ( 
.A(n_141),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_308),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_216),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_43),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_331),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_292),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_302),
.Y(n_451)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_185),
.Y(n_452)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_336),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_3),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_182),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_14),
.Y(n_456)
);

INVx2_ASAP7_75t_L g457 ( 
.A(n_226),
.Y(n_457)
);

INVx2_ASAP7_75t_SL g458 ( 
.A(n_75),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_64),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_150),
.Y(n_460)
);

BUFx10_ASAP7_75t_L g461 ( 
.A(n_190),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_13),
.Y(n_462)
);

BUFx6f_ASAP7_75t_L g463 ( 
.A(n_321),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_197),
.Y(n_464)
);

CKINVDCx5p33_ASAP7_75t_R g465 ( 
.A(n_153),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_314),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_238),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_147),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_193),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_125),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_172),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_169),
.Y(n_472)
);

INVx2_ASAP7_75t_SL g473 ( 
.A(n_158),
.Y(n_473)
);

BUFx10_ASAP7_75t_L g474 ( 
.A(n_232),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_101),
.Y(n_475)
);

BUFx3_ASAP7_75t_L g476 ( 
.A(n_317),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_217),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_146),
.Y(n_478)
);

BUFx6f_ASAP7_75t_L g479 ( 
.A(n_38),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_319),
.Y(n_480)
);

CKINVDCx5p33_ASAP7_75t_R g481 ( 
.A(n_8),
.Y(n_481)
);

CKINVDCx5p33_ASAP7_75t_R g482 ( 
.A(n_110),
.Y(n_482)
);

CKINVDCx5p33_ASAP7_75t_R g483 ( 
.A(n_74),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_176),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_123),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_126),
.Y(n_486)
);

BUFx6f_ASAP7_75t_L g487 ( 
.A(n_47),
.Y(n_487)
);

CKINVDCx5p33_ASAP7_75t_R g488 ( 
.A(n_27),
.Y(n_488)
);

HB1xp67_ASAP7_75t_L g489 ( 
.A(n_138),
.Y(n_489)
);

INVx2_ASAP7_75t_SL g490 ( 
.A(n_43),
.Y(n_490)
);

BUFx5_ASAP7_75t_L g491 ( 
.A(n_121),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_128),
.Y(n_492)
);

HB1xp67_ASAP7_75t_L g493 ( 
.A(n_220),
.Y(n_493)
);

CKINVDCx5p33_ASAP7_75t_R g494 ( 
.A(n_252),
.Y(n_494)
);

CKINVDCx20_ASAP7_75t_R g495 ( 
.A(n_208),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_109),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_212),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_257),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_56),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_99),
.Y(n_500)
);

CKINVDCx20_ASAP7_75t_R g501 ( 
.A(n_327),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_326),
.Y(n_502)
);

BUFx3_ASAP7_75t_L g503 ( 
.A(n_301),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_44),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_156),
.Y(n_505)
);

CKINVDCx5p33_ASAP7_75t_R g506 ( 
.A(n_309),
.Y(n_506)
);

CKINVDCx5p33_ASAP7_75t_R g507 ( 
.A(n_274),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_144),
.Y(n_508)
);

CKINVDCx5p33_ASAP7_75t_R g509 ( 
.A(n_69),
.Y(n_509)
);

CKINVDCx5p33_ASAP7_75t_R g510 ( 
.A(n_30),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_263),
.Y(n_511)
);

BUFx6f_ASAP7_75t_L g512 ( 
.A(n_88),
.Y(n_512)
);

INVx3_ASAP7_75t_L g513 ( 
.A(n_315),
.Y(n_513)
);

CKINVDCx5p33_ASAP7_75t_R g514 ( 
.A(n_86),
.Y(n_514)
);

INVx1_ASAP7_75t_SL g515 ( 
.A(n_5),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_310),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_168),
.Y(n_517)
);

CKINVDCx16_ASAP7_75t_R g518 ( 
.A(n_98),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_23),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_127),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_94),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_34),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_72),
.Y(n_523)
);

CKINVDCx5p33_ASAP7_75t_R g524 ( 
.A(n_183),
.Y(n_524)
);

CKINVDCx5p33_ASAP7_75t_R g525 ( 
.A(n_303),
.Y(n_525)
);

CKINVDCx20_ASAP7_75t_R g526 ( 
.A(n_9),
.Y(n_526)
);

CKINVDCx5p33_ASAP7_75t_R g527 ( 
.A(n_53),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_57),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_41),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_272),
.Y(n_530)
);

INVx1_ASAP7_75t_SL g531 ( 
.A(n_136),
.Y(n_531)
);

INVx1_ASAP7_75t_SL g532 ( 
.A(n_254),
.Y(n_532)
);

CKINVDCx5p33_ASAP7_75t_R g533 ( 
.A(n_40),
.Y(n_533)
);

INVx2_ASAP7_75t_SL g534 ( 
.A(n_180),
.Y(n_534)
);

INVx2_ASAP7_75t_L g535 ( 
.A(n_115),
.Y(n_535)
);

CKINVDCx5p33_ASAP7_75t_R g536 ( 
.A(n_148),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_215),
.Y(n_537)
);

CKINVDCx5p33_ASAP7_75t_R g538 ( 
.A(n_178),
.Y(n_538)
);

BUFx5_ASAP7_75t_L g539 ( 
.A(n_248),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_188),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_489),
.B(n_0),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_369),
.Y(n_542)
);

CKINVDCx5p33_ASAP7_75t_R g543 ( 
.A(n_349),
.Y(n_543)
);

INVxp33_ASAP7_75t_SL g544 ( 
.A(n_489),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_369),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_369),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_351),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g548 ( 
.A(n_526),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_353),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_369),
.Y(n_550)
);

CKINVDCx5p33_ASAP7_75t_R g551 ( 
.A(n_354),
.Y(n_551)
);

HB1xp67_ASAP7_75t_L g552 ( 
.A(n_370),
.Y(n_552)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_479),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_357),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_431),
.B(n_1),
.Y(n_555)
);

CKINVDCx5p33_ASAP7_75t_R g556 ( 
.A(n_362),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_364),
.Y(n_557)
);

CKINVDCx20_ASAP7_75t_R g558 ( 
.A(n_373),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_479),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_479),
.Y(n_560)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_419),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_372),
.Y(n_562)
);

CKINVDCx20_ASAP7_75t_R g563 ( 
.A(n_424),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_375),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_479),
.Y(n_565)
);

BUFx2_ASAP7_75t_L g566 ( 
.A(n_435),
.Y(n_566)
);

CKINVDCx20_ASAP7_75t_R g567 ( 
.A(n_355),
.Y(n_567)
);

INVxp67_ASAP7_75t_SL g568 ( 
.A(n_493),
.Y(n_568)
);

BUFx3_ASAP7_75t_L g569 ( 
.A(n_368),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_365),
.Y(n_570)
);

CKINVDCx20_ASAP7_75t_R g571 ( 
.A(n_436),
.Y(n_571)
);

INVx2_ASAP7_75t_L g572 ( 
.A(n_491),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

INVxp67_ASAP7_75t_SL g574 ( 
.A(n_493),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_484),
.B(n_1),
.Y(n_575)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_437),
.B(n_2),
.Y(n_576)
);

CKINVDCx5p33_ASAP7_75t_R g577 ( 
.A(n_376),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_487),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_487),
.Y(n_579)
);

CKINVDCx20_ASAP7_75t_R g580 ( 
.A(n_495),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_487),
.Y(n_581)
);

CKINVDCx20_ASAP7_75t_R g582 ( 
.A(n_496),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_501),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_388),
.Y(n_584)
);

CKINVDCx5p33_ASAP7_75t_R g585 ( 
.A(n_377),
.Y(n_585)
);

INVxp67_ASAP7_75t_SL g586 ( 
.A(n_402),
.Y(n_586)
);

CKINVDCx5p33_ASAP7_75t_R g587 ( 
.A(n_380),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_391),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_407),
.Y(n_589)
);

HB1xp67_ASAP7_75t_L g590 ( 
.A(n_360),
.Y(n_590)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_409),
.Y(n_591)
);

BUFx3_ASAP7_75t_L g592 ( 
.A(n_503),
.Y(n_592)
);

CKINVDCx5p33_ASAP7_75t_R g593 ( 
.A(n_382),
.Y(n_593)
);

CKINVDCx20_ASAP7_75t_R g594 ( 
.A(n_379),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_448),
.Y(n_595)
);

CKINVDCx20_ASAP7_75t_R g596 ( 
.A(n_408),
.Y(n_596)
);

INVx1_ASAP7_75t_SL g597 ( 
.A(n_350),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_459),
.Y(n_598)
);

CKINVDCx5p33_ASAP7_75t_R g599 ( 
.A(n_385),
.Y(n_599)
);

INVx1_ASAP7_75t_L g600 ( 
.A(n_504),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_522),
.Y(n_601)
);

CKINVDCx5p33_ASAP7_75t_R g602 ( 
.A(n_387),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_523),
.Y(n_603)
);

INVxp33_ASAP7_75t_SL g604 ( 
.A(n_410),
.Y(n_604)
);

CKINVDCx20_ASAP7_75t_R g605 ( 
.A(n_415),
.Y(n_605)
);

INVx1_ASAP7_75t_SL g606 ( 
.A(n_361),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_529),
.Y(n_607)
);

CKINVDCx5p33_ASAP7_75t_R g608 ( 
.A(n_390),
.Y(n_608)
);

CKINVDCx5p33_ASAP7_75t_R g609 ( 
.A(n_394),
.Y(n_609)
);

NOR2xp67_ASAP7_75t_L g610 ( 
.A(n_484),
.B(n_2),
.Y(n_610)
);

CKINVDCx20_ASAP7_75t_R g611 ( 
.A(n_432),
.Y(n_611)
);

CKINVDCx20_ASAP7_75t_R g612 ( 
.A(n_454),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_402),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_400),
.B(n_3),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_456),
.Y(n_615)
);

NOR2xp33_ASAP7_75t_L g616 ( 
.A(n_400),
.B(n_4),
.Y(n_616)
);

CKINVDCx5p33_ASAP7_75t_R g617 ( 
.A(n_395),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_476),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_396),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_476),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_352),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_513),
.B(n_4),
.Y(n_622)
);

BUFx3_ASAP7_75t_L g623 ( 
.A(n_398),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_359),
.Y(n_624)
);

CKINVDCx5p33_ASAP7_75t_R g625 ( 
.A(n_401),
.Y(n_625)
);

INVx2_ASAP7_75t_L g626 ( 
.A(n_491),
.Y(n_626)
);

CKINVDCx5p33_ASAP7_75t_R g627 ( 
.A(n_403),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_363),
.Y(n_628)
);

INVx1_ASAP7_75t_L g629 ( 
.A(n_366),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_367),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_371),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_374),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_381),
.Y(n_633)
);

INVxp67_ASAP7_75t_SL g634 ( 
.A(n_513),
.Y(n_634)
);

CKINVDCx5p33_ASAP7_75t_R g635 ( 
.A(n_404),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_383),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_384),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_386),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_392),
.Y(n_639)
);

INVx3_ASAP7_75t_L g640 ( 
.A(n_378),
.Y(n_640)
);

INVxp67_ASAP7_75t_SL g641 ( 
.A(n_393),
.Y(n_641)
);

CKINVDCx20_ASAP7_75t_R g642 ( 
.A(n_462),
.Y(n_642)
);

INVx1_ASAP7_75t_L g643 ( 
.A(n_397),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_405),
.Y(n_644)
);

CKINVDCx5p33_ASAP7_75t_R g645 ( 
.A(n_412),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_414),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_418),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_421),
.Y(n_648)
);

CKINVDCx20_ASAP7_75t_R g649 ( 
.A(n_481),
.Y(n_649)
);

CKINVDCx20_ASAP7_75t_R g650 ( 
.A(n_483),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_440),
.Y(n_651)
);

CKINVDCx20_ASAP7_75t_R g652 ( 
.A(n_488),
.Y(n_652)
);

INVx1_ASAP7_75t_L g653 ( 
.A(n_441),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_413),
.Y(n_654)
);

INVx2_ASAP7_75t_L g655 ( 
.A(n_491),
.Y(n_655)
);

CKINVDCx20_ASAP7_75t_R g656 ( 
.A(n_502),
.Y(n_656)
);

BUFx3_ASAP7_75t_L g657 ( 
.A(n_398),
.Y(n_657)
);

AND2x4_ASAP7_75t_L g658 ( 
.A(n_634),
.B(n_423),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_542),
.Y(n_659)
);

HB1xp67_ASAP7_75t_L g660 ( 
.A(n_597),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_640),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_640),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_545),
.Y(n_663)
);

AND2x4_ASAP7_75t_L g664 ( 
.A(n_641),
.B(n_473),
.Y(n_664)
);

INVx3_ASAP7_75t_L g665 ( 
.A(n_640),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_550),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_553),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_559),
.Y(n_669)
);

BUFx6f_ASAP7_75t_L g670 ( 
.A(n_560),
.Y(n_670)
);

NAND2xp5_ASAP7_75t_L g671 ( 
.A(n_543),
.B(n_534),
.Y(n_671)
);

BUFx6f_ASAP7_75t_L g672 ( 
.A(n_565),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_573),
.Y(n_673)
);

BUFx3_ASAP7_75t_L g674 ( 
.A(n_569),
.Y(n_674)
);

AND2x2_ASAP7_75t_L g675 ( 
.A(n_590),
.B(n_399),
.Y(n_675)
);

INVx6_ASAP7_75t_L g676 ( 
.A(n_569),
.Y(n_676)
);

NAND2xp5_ASAP7_75t_L g677 ( 
.A(n_547),
.B(n_399),
.Y(n_677)
);

BUFx6f_ASAP7_75t_L g678 ( 
.A(n_578),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_579),
.Y(n_679)
);

AND2x2_ASAP7_75t_L g680 ( 
.A(n_586),
.B(n_358),
.Y(n_680)
);

INVxp67_ASAP7_75t_L g681 ( 
.A(n_552),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_581),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_572),
.Y(n_683)
);

AND2x4_ASAP7_75t_L g684 ( 
.A(n_610),
.B(n_389),
.Y(n_684)
);

AND2x2_ASAP7_75t_SL g685 ( 
.A(n_541),
.B(n_430),
.Y(n_685)
);

AND2x6_ASAP7_75t_L g686 ( 
.A(n_622),
.B(n_378),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_621),
.Y(n_687)
);

AND2x4_ASAP7_75t_L g688 ( 
.A(n_613),
.B(n_406),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_624),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_SL g690 ( 
.A(n_544),
.B(n_518),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_SL g691 ( 
.A(n_576),
.B(n_461),
.Y(n_691)
);

NOR2xp33_ASAP7_75t_L g692 ( 
.A(n_575),
.B(n_411),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_628),
.Y(n_693)
);

INVx2_ASAP7_75t_L g694 ( 
.A(n_572),
.Y(n_694)
);

NAND2xp5_ASAP7_75t_L g695 ( 
.A(n_549),
.B(n_457),
.Y(n_695)
);

AND2x4_ASAP7_75t_L g696 ( 
.A(n_618),
.B(n_478),
.Y(n_696)
);

CKINVDCx20_ASAP7_75t_R g697 ( 
.A(n_548),
.Y(n_697)
);

INVx1_ASAP7_75t_L g698 ( 
.A(n_629),
.Y(n_698)
);

BUFx2_ASAP7_75t_L g699 ( 
.A(n_567),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_584),
.Y(n_700)
);

INVx3_ASAP7_75t_L g701 ( 
.A(n_592),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_620),
.B(n_500),
.Y(n_702)
);

INVx1_ASAP7_75t_L g703 ( 
.A(n_630),
.Y(n_703)
);

INVx4_ASAP7_75t_L g704 ( 
.A(n_551),
.Y(n_704)
);

AND2x4_ASAP7_75t_L g705 ( 
.A(n_592),
.B(n_535),
.Y(n_705)
);

INVx3_ASAP7_75t_L g706 ( 
.A(n_588),
.Y(n_706)
);

INVx3_ASAP7_75t_L g707 ( 
.A(n_589),
.Y(n_707)
);

INVx1_ASAP7_75t_L g708 ( 
.A(n_631),
.Y(n_708)
);

OAI21x1_ASAP7_75t_L g709 ( 
.A1(n_626),
.A2(n_444),
.B(n_442),
.Y(n_709)
);

BUFx2_ASAP7_75t_L g710 ( 
.A(n_567),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_626),
.Y(n_711)
);

AND2x4_ASAP7_75t_L g712 ( 
.A(n_632),
.B(n_447),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_554),
.B(n_450),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_655),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_655),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_556),
.Y(n_716)
);

INVx1_ASAP7_75t_L g717 ( 
.A(n_633),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_636),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_637),
.Y(n_719)
);

AND2x2_ASAP7_75t_L g720 ( 
.A(n_566),
.B(n_411),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_638),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_557),
.B(n_453),
.Y(n_722)
);

BUFx6f_ASAP7_75t_L g723 ( 
.A(n_591),
.Y(n_723)
);

INVx2_ASAP7_75t_L g724 ( 
.A(n_639),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_SL g725 ( 
.A(n_606),
.B(n_461),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_643),
.Y(n_726)
);

INVx2_ASAP7_75t_L g727 ( 
.A(n_644),
.Y(n_727)
);

INVx4_ASAP7_75t_L g728 ( 
.A(n_562),
.Y(n_728)
);

BUFx6f_ASAP7_75t_L g729 ( 
.A(n_595),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_646),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_647),
.Y(n_731)
);

AND2x4_ASAP7_75t_L g732 ( 
.A(n_648),
.B(n_455),
.Y(n_732)
);

OA21x2_ASAP7_75t_L g733 ( 
.A1(n_651),
.A2(n_464),
.B(n_460),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_653),
.Y(n_734)
);

INVx3_ASAP7_75t_L g735 ( 
.A(n_598),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_600),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_L g737 ( 
.A(n_564),
.B(n_467),
.Y(n_737)
);

INVx3_ASAP7_75t_L g738 ( 
.A(n_601),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_603),
.Y(n_739)
);

OA21x2_ASAP7_75t_L g740 ( 
.A1(n_607),
.A2(n_470),
.B(n_469),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_570),
.Y(n_741)
);

INVx1_ASAP7_75t_L g742 ( 
.A(n_614),
.Y(n_742)
);

INVx3_ASAP7_75t_L g743 ( 
.A(n_623),
.Y(n_743)
);

BUFx2_ASAP7_75t_L g744 ( 
.A(n_594),
.Y(n_744)
);

BUFx6f_ASAP7_75t_L g745 ( 
.A(n_616),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_568),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_574),
.B(n_531),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_623),
.Y(n_748)
);

INVx4_ASAP7_75t_L g749 ( 
.A(n_577),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_683),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_SL g751 ( 
.A(n_745),
.B(n_378),
.Y(n_751)
);

OAI22xp33_ASAP7_75t_L g752 ( 
.A1(n_725),
.A2(n_515),
.B1(n_458),
.B2(n_490),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_736),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_660),
.Y(n_754)
);

INVx8_ASAP7_75t_L g755 ( 
.A(n_716),
.Y(n_755)
);

NAND2xp33_ASAP7_75t_SL g756 ( 
.A(n_691),
.B(n_356),
.Y(n_756)
);

AOI22xp33_ASAP7_75t_L g757 ( 
.A1(n_692),
.A2(n_475),
.B1(n_480),
.B2(n_471),
.Y(n_757)
);

INVx2_ASAP7_75t_SL g758 ( 
.A(n_660),
.Y(n_758)
);

INVx2_ASAP7_75t_SL g759 ( 
.A(n_720),
.Y(n_759)
);

OR2x6_ASAP7_75t_L g760 ( 
.A(n_699),
.B(n_657),
.Y(n_760)
);

INVx1_ASAP7_75t_L g761 ( 
.A(n_687),
.Y(n_761)
);

INVx2_ASAP7_75t_L g762 ( 
.A(n_661),
.Y(n_762)
);

BUFx2_ASAP7_75t_L g763 ( 
.A(n_674),
.Y(n_763)
);

INVx1_ASAP7_75t_L g764 ( 
.A(n_689),
.Y(n_764)
);

NAND3xp33_ASAP7_75t_L g765 ( 
.A(n_692),
.B(n_555),
.C(n_585),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_SL g766 ( 
.A(n_745),
.B(n_378),
.Y(n_766)
);

AOI22xp33_ASAP7_75t_L g767 ( 
.A1(n_742),
.A2(n_492),
.B1(n_497),
.B2(n_486),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_693),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_SL g769 ( 
.A(n_745),
.B(n_428),
.Y(n_769)
);

AOI22xp33_ASAP7_75t_L g770 ( 
.A1(n_686),
.A2(n_505),
.B1(n_511),
.B2(n_498),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_698),
.Y(n_771)
);

NAND2xp33_ASAP7_75t_L g772 ( 
.A(n_686),
.B(n_745),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_703),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_708),
.Y(n_774)
);

OAI22xp33_ASAP7_75t_L g775 ( 
.A1(n_691),
.A2(n_747),
.B1(n_690),
.B2(n_746),
.Y(n_775)
);

BUFx2_ASAP7_75t_L g776 ( 
.A(n_674),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_717),
.Y(n_777)
);

NAND2xp33_ASAP7_75t_SL g778 ( 
.A(n_690),
.B(n_521),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_718),
.Y(n_779)
);

INVxp67_ASAP7_75t_L g780 ( 
.A(n_747),
.Y(n_780)
);

AND2x6_ASAP7_75t_L g781 ( 
.A(n_675),
.B(n_428),
.Y(n_781)
);

INVx2_ASAP7_75t_L g782 ( 
.A(n_661),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_721),
.Y(n_783)
);

NAND2xp33_ASAP7_75t_L g784 ( 
.A(n_686),
.B(n_587),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_661),
.Y(n_785)
);

BUFx6f_ASAP7_75t_L g786 ( 
.A(n_661),
.Y(n_786)
);

INVx2_ASAP7_75t_L g787 ( 
.A(n_666),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_700),
.Y(n_788)
);

AOI22xp33_ASAP7_75t_L g789 ( 
.A1(n_686),
.A2(n_530),
.B1(n_452),
.B2(n_463),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_726),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_730),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_SL g792 ( 
.A(n_685),
.B(n_428),
.Y(n_792)
);

AOI22xp5_ASAP7_75t_L g793 ( 
.A1(n_685),
.A2(n_604),
.B1(n_593),
.B2(n_602),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_683),
.Y(n_794)
);

AND2x2_ASAP7_75t_L g795 ( 
.A(n_680),
.B(n_599),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_SL g796 ( 
.A(n_664),
.B(n_428),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_731),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_734),
.Y(n_798)
);

XOR2xp5_ASAP7_75t_L g799 ( 
.A(n_697),
.B(n_558),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_665),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_665),
.Y(n_801)
);

NAND2xp5_ASAP7_75t_L g802 ( 
.A(n_658),
.B(n_608),
.Y(n_802)
);

AOI22xp33_ASAP7_75t_L g803 ( 
.A1(n_686),
.A2(n_463),
.B1(n_512),
.B2(n_452),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_658),
.B(n_609),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_666),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_700),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_700),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_695),
.B(n_617),
.Y(n_808)
);

BUFx3_ASAP7_75t_L g809 ( 
.A(n_676),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_700),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_723),
.Y(n_811)
);

INVx2_ASAP7_75t_L g812 ( 
.A(n_666),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_666),
.Y(n_813)
);

INVx2_ASAP7_75t_SL g814 ( 
.A(n_676),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_723),
.Y(n_815)
);

NAND3xp33_ASAP7_75t_L g816 ( 
.A(n_741),
.B(n_625),
.C(n_619),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_723),
.Y(n_817)
);

INVx2_ASAP7_75t_L g818 ( 
.A(n_694),
.Y(n_818)
);

AOI22xp33_ASAP7_75t_L g819 ( 
.A1(n_684),
.A2(n_740),
.B1(n_664),
.B2(n_733),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_723),
.Y(n_820)
);

INVx3_ASAP7_75t_L g821 ( 
.A(n_669),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_729),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_729),
.Y(n_823)
);

INVx3_ASAP7_75t_L g824 ( 
.A(n_669),
.Y(n_824)
);

INVx8_ASAP7_75t_L g825 ( 
.A(n_716),
.Y(n_825)
);

AOI22xp33_ASAP7_75t_SL g826 ( 
.A1(n_664),
.A2(n_563),
.B1(n_571),
.B2(n_561),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_676),
.Y(n_827)
);

NAND2xp33_ASAP7_75t_L g828 ( 
.A(n_677),
.B(n_627),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_729),
.Y(n_829)
);

INVx1_ASAP7_75t_SL g830 ( 
.A(n_697),
.Y(n_830)
);

AND2x2_ASAP7_75t_L g831 ( 
.A(n_743),
.B(n_635),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_743),
.B(n_645),
.Y(n_832)
);

BUFx6f_ASAP7_75t_L g833 ( 
.A(n_729),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_669),
.Y(n_834)
);

AND2x2_ASAP7_75t_L g835 ( 
.A(n_701),
.B(n_654),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_719),
.Y(n_836)
);

NAND2xp5_ASAP7_75t_SL g837 ( 
.A(n_658),
.B(n_452),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_669),
.Y(n_838)
);

INVx3_ASAP7_75t_L g839 ( 
.A(n_670),
.Y(n_839)
);

NOR2x1p5_ASAP7_75t_L g840 ( 
.A(n_704),
.B(n_657),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_808),
.B(n_713),
.Y(n_841)
);

OAI22xp5_ASAP7_75t_L g842 ( 
.A1(n_757),
.A2(n_722),
.B1(n_737),
.B2(n_684),
.Y(n_842)
);

INVx2_ASAP7_75t_L g843 ( 
.A(n_750),
.Y(n_843)
);

NAND2xp5_ASAP7_75t_L g844 ( 
.A(n_819),
.B(n_733),
.Y(n_844)
);

OAI22xp5_ASAP7_75t_L g845 ( 
.A1(n_757),
.A2(n_684),
.B1(n_582),
.B2(n_583),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_819),
.B(n_733),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_780),
.B(n_740),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_753),
.Y(n_848)
);

INVx1_ASAP7_75t_L g849 ( 
.A(n_761),
.Y(n_849)
);

NAND2xp5_ASAP7_75t_L g850 ( 
.A(n_808),
.B(n_671),
.Y(n_850)
);

NAND2x1_ASAP7_75t_L g851 ( 
.A(n_750),
.B(n_694),
.Y(n_851)
);

INVxp67_ASAP7_75t_SL g852 ( 
.A(n_786),
.Y(n_852)
);

AND2x2_ASAP7_75t_L g853 ( 
.A(n_754),
.B(n_701),
.Y(n_853)
);

INVxp67_ASAP7_75t_L g854 ( 
.A(n_758),
.Y(n_854)
);

BUFx2_ASAP7_75t_L g855 ( 
.A(n_760),
.Y(n_855)
);

NAND2xp5_ASAP7_75t_SL g856 ( 
.A(n_775),
.B(n_704),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_775),
.B(n_704),
.Y(n_857)
);

INVx2_ASAP7_75t_L g858 ( 
.A(n_794),
.Y(n_858)
);

AOI22xp33_ASAP7_75t_L g859 ( 
.A1(n_792),
.A2(n_740),
.B1(n_732),
.B2(n_712),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_L g860 ( 
.A(n_780),
.B(n_728),
.Y(n_860)
);

BUFx6f_ASAP7_75t_SL g861 ( 
.A(n_760),
.Y(n_861)
);

AND2x6_ASAP7_75t_SL g862 ( 
.A(n_760),
.B(n_748),
.Y(n_862)
);

A2O1A1Ixp33_ASAP7_75t_L g863 ( 
.A1(n_792),
.A2(n_756),
.B(n_778),
.C(n_767),
.Y(n_863)
);

A2O1A1Ixp33_ASAP7_75t_L g864 ( 
.A1(n_756),
.A2(n_709),
.B(n_732),
.C(n_712),
.Y(n_864)
);

OR2x6_ASAP7_75t_L g865 ( 
.A(n_755),
.B(n_710),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_835),
.B(n_831),
.Y(n_866)
);

NOR2xp33_ASAP7_75t_L g867 ( 
.A(n_765),
.B(n_728),
.Y(n_867)
);

NAND2x1_ASAP7_75t_L g868 ( 
.A(n_794),
.B(n_711),
.Y(n_868)
);

INVx2_ASAP7_75t_L g869 ( 
.A(n_818),
.Y(n_869)
);

OR2x2_ASAP7_75t_L g870 ( 
.A(n_759),
.B(n_681),
.Y(n_870)
);

AND2x2_ASAP7_75t_L g871 ( 
.A(n_795),
.B(n_728),
.Y(n_871)
);

OR2x2_ASAP7_75t_L g872 ( 
.A(n_830),
.B(n_744),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_802),
.B(n_749),
.Y(n_873)
);

NAND2xp5_ASAP7_75t_L g874 ( 
.A(n_832),
.B(n_749),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_796),
.B(n_749),
.Y(n_875)
);

INVx2_ASAP7_75t_SL g876 ( 
.A(n_763),
.Y(n_876)
);

BUFx6f_ASAP7_75t_SL g877 ( 
.A(n_764),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_768),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_L g879 ( 
.A(n_796),
.B(n_712),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_837),
.B(n_732),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_837),
.B(n_705),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_L g882 ( 
.A(n_771),
.B(n_705),
.Y(n_882)
);

INVx2_ASAP7_75t_SL g883 ( 
.A(n_776),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_773),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_SL g885 ( 
.A(n_804),
.B(n_705),
.Y(n_885)
);

INVx1_ASAP7_75t_SL g886 ( 
.A(n_799),
.Y(n_886)
);

A2O1A1Ixp33_ASAP7_75t_L g887 ( 
.A1(n_778),
.A2(n_709),
.B(n_696),
.C(n_702),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_774),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_SL g889 ( 
.A(n_793),
.B(n_594),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_L g890 ( 
.A(n_777),
.B(n_711),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_818),
.Y(n_891)
);

NOR2xp33_ASAP7_75t_L g892 ( 
.A(n_816),
.B(n_596),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_779),
.B(n_783),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_790),
.B(n_714),
.Y(n_894)
);

BUFx5_ASAP7_75t_L g895 ( 
.A(n_806),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_836),
.Y(n_896)
);

NOR2xp33_ASAP7_75t_R g897 ( 
.A(n_784),
.B(n_580),
.Y(n_897)
);

AND2x2_ASAP7_75t_L g898 ( 
.A(n_840),
.B(n_656),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_752),
.B(n_596),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_SL g900 ( 
.A(n_752),
.B(n_605),
.Y(n_900)
);

OAI221xp5_ASAP7_75t_L g901 ( 
.A1(n_767),
.A2(n_532),
.B1(n_738),
.B2(n_724),
.C(n_727),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_791),
.B(n_714),
.Y(n_902)
);

OR2x2_ASAP7_75t_L g903 ( 
.A(n_814),
.B(n_688),
.Y(n_903)
);

A2O1A1Ixp33_ASAP7_75t_L g904 ( 
.A1(n_797),
.A2(n_696),
.B(n_702),
.C(n_688),
.Y(n_904)
);

AOI22xp33_ASAP7_75t_L g905 ( 
.A1(n_770),
.A2(n_696),
.B1(n_702),
.B2(n_688),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_798),
.Y(n_906)
);

NOR2xp33_ASAP7_75t_L g907 ( 
.A(n_809),
.B(n_605),
.Y(n_907)
);

BUFx2_ASAP7_75t_L g908 ( 
.A(n_809),
.Y(n_908)
);

NOR2xp33_ASAP7_75t_L g909 ( 
.A(n_827),
.B(n_611),
.Y(n_909)
);

AOI22xp5_ASAP7_75t_L g910 ( 
.A1(n_828),
.A2(n_611),
.B1(n_615),
.B2(n_612),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_L g911 ( 
.A(n_800),
.B(n_715),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_801),
.B(n_715),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_786),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_751),
.B(n_738),
.Y(n_914)
);

BUFx6f_ASAP7_75t_L g915 ( 
.A(n_827),
.Y(n_915)
);

NAND2xp5_ASAP7_75t_SL g916 ( 
.A(n_803),
.B(n_612),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_762),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_L g918 ( 
.A(n_751),
.B(n_738),
.Y(n_918)
);

INVx1_ASAP7_75t_L g919 ( 
.A(n_782),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_786),
.Y(n_920)
);

NAND3xp33_ASAP7_75t_SL g921 ( 
.A(n_826),
.B(n_563),
.C(n_615),
.Y(n_921)
);

INVxp67_ASAP7_75t_L g922 ( 
.A(n_826),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_786),
.Y(n_923)
);

OR2x6_ASAP7_75t_L g924 ( 
.A(n_755),
.B(n_739),
.Y(n_924)
);

AOI22xp5_ASAP7_75t_L g925 ( 
.A1(n_772),
.A2(n_649),
.B1(n_650),
.B2(n_642),
.Y(n_925)
);

NAND2xp33_ASAP7_75t_L g926 ( 
.A(n_789),
.B(n_491),
.Y(n_926)
);

NAND2xp5_ASAP7_75t_SL g927 ( 
.A(n_803),
.B(n_642),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_785),
.Y(n_928)
);

AOI22xp33_ASAP7_75t_L g929 ( 
.A1(n_770),
.A2(n_539),
.B1(n_491),
.B2(n_719),
.Y(n_929)
);

NOR2x1_ASAP7_75t_L g930 ( 
.A(n_766),
.B(n_649),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_766),
.B(n_662),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_769),
.B(n_662),
.Y(n_932)
);

INVx2_ASAP7_75t_L g933 ( 
.A(n_821),
.Y(n_933)
);

NOR2xp67_ASAP7_75t_SL g934 ( 
.A(n_769),
.B(n_452),
.Y(n_934)
);

NAND2xp33_ASAP7_75t_L g935 ( 
.A(n_789),
.B(n_491),
.Y(n_935)
);

OAI21xp5_ASAP7_75t_L g936 ( 
.A1(n_807),
.A2(n_727),
.B(n_724),
.Y(n_936)
);

INVx2_ASAP7_75t_L g937 ( 
.A(n_821),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_824),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_810),
.B(n_706),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_841),
.B(n_815),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_848),
.Y(n_941)
);

NAND2x1_ASAP7_75t_L g942 ( 
.A(n_843),
.B(n_824),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_913),
.Y(n_943)
);

NOR2xp33_ASAP7_75t_L g944 ( 
.A(n_850),
.B(n_548),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_844),
.A2(n_811),
.B(n_788),
.Y(n_945)
);

AO21x1_ASAP7_75t_L g946 ( 
.A1(n_856),
.A2(n_820),
.B(n_817),
.Y(n_946)
);

AND2x2_ASAP7_75t_SL g947 ( 
.A(n_892),
.B(n_755),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_L g948 ( 
.A(n_866),
.B(n_822),
.Y(n_948)
);

A2O1A1Ixp33_ASAP7_75t_L g949 ( 
.A1(n_863),
.A2(n_829),
.B(n_823),
.C(n_825),
.Y(n_949)
);

OR2x2_ASAP7_75t_L g950 ( 
.A(n_872),
.B(n_870),
.Y(n_950)
);

AOI21xp5_ASAP7_75t_L g951 ( 
.A1(n_844),
.A2(n_846),
.B(n_879),
.Y(n_951)
);

AOI21xp5_ASAP7_75t_L g952 ( 
.A1(n_846),
.A2(n_811),
.B(n_788),
.Y(n_952)
);

INVx2_ASAP7_75t_L g953 ( 
.A(n_858),
.Y(n_953)
);

AOI21xp5_ASAP7_75t_L g954 ( 
.A1(n_880),
.A2(n_811),
.B(n_788),
.Y(n_954)
);

OAI21xp5_ASAP7_75t_L g955 ( 
.A1(n_847),
.A2(n_781),
.B(n_787),
.Y(n_955)
);

INVx2_ASAP7_75t_L g956 ( 
.A(n_869),
.Y(n_956)
);

AOI22xp5_ASAP7_75t_L g957 ( 
.A1(n_857),
.A2(n_922),
.B1(n_842),
.B2(n_847),
.Y(n_957)
);

AOI22xp33_ASAP7_75t_L g958 ( 
.A1(n_842),
.A2(n_781),
.B1(n_812),
.B2(n_805),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_874),
.B(n_781),
.Y(n_959)
);

O2A1O1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_887),
.A2(n_707),
.B(n_735),
.C(n_706),
.Y(n_960)
);

AOI21xp5_ASAP7_75t_L g961 ( 
.A1(n_885),
.A2(n_811),
.B(n_788),
.Y(n_961)
);

BUFx2_ASAP7_75t_L g962 ( 
.A(n_854),
.Y(n_962)
);

OAI21xp5_ASAP7_75t_L g963 ( 
.A1(n_936),
.A2(n_781),
.B(n_813),
.Y(n_963)
);

AOI21xp5_ASAP7_75t_L g964 ( 
.A1(n_852),
.A2(n_833),
.B(n_834),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_860),
.B(n_781),
.Y(n_965)
);

BUFx4f_ASAP7_75t_L g966 ( 
.A(n_865),
.Y(n_966)
);

NAND2xp5_ASAP7_75t_L g967 ( 
.A(n_875),
.B(n_833),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_L g968 ( 
.A(n_849),
.B(n_833),
.Y(n_968)
);

NAND2xp5_ASAP7_75t_SL g969 ( 
.A(n_871),
.B(n_825),
.Y(n_969)
);

INVx4_ASAP7_75t_L g970 ( 
.A(n_915),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_926),
.A2(n_935),
.B1(n_859),
.B2(n_867),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_878),
.B(n_833),
.Y(n_972)
);

NAND2xp5_ASAP7_75t_L g973 ( 
.A(n_884),
.B(n_838),
.Y(n_973)
);

AOI21xp5_ASAP7_75t_L g974 ( 
.A1(n_881),
.A2(n_839),
.B(n_838),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_853),
.Y(n_975)
);

O2A1O1Ixp33_ASAP7_75t_L g976 ( 
.A1(n_916),
.A2(n_735),
.B(n_707),
.C(n_739),
.Y(n_976)
);

BUFx6f_ASAP7_75t_L g977 ( 
.A(n_915),
.Y(n_977)
);

NAND2xp5_ASAP7_75t_L g978 ( 
.A(n_888),
.B(n_839),
.Y(n_978)
);

AOI21xp5_ASAP7_75t_L g979 ( 
.A1(n_893),
.A2(n_512),
.B(n_463),
.Y(n_979)
);

O2A1O1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_927),
.A2(n_901),
.B(n_864),
.C(n_904),
.Y(n_980)
);

NOR2xp33_ASAP7_75t_L g981 ( 
.A(n_899),
.B(n_650),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_SL g982 ( 
.A(n_845),
.B(n_825),
.Y(n_982)
);

NAND2xp5_ASAP7_75t_L g983 ( 
.A(n_906),
.B(n_652),
.Y(n_983)
);

INVx3_ASAP7_75t_L g984 ( 
.A(n_920),
.Y(n_984)
);

O2A1O1Ixp33_ASAP7_75t_L g985 ( 
.A1(n_900),
.A2(n_659),
.B(n_667),
.C(n_663),
.Y(n_985)
);

AND2x2_ASAP7_75t_L g986 ( 
.A(n_876),
.B(n_652),
.Y(n_986)
);

BUFx4f_ASAP7_75t_L g987 ( 
.A(n_865),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_936),
.A2(n_882),
.B(n_914),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_883),
.B(n_673),
.Y(n_989)
);

BUFx2_ASAP7_75t_L g990 ( 
.A(n_897),
.Y(n_990)
);

OAI21xp5_ASAP7_75t_L g991 ( 
.A1(n_918),
.A2(n_682),
.B(n_679),
.Y(n_991)
);

INVx11_ASAP7_75t_L g992 ( 
.A(n_861),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_845),
.B(n_499),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_896),
.B(n_668),
.Y(n_994)
);

OR2x2_ASAP7_75t_SL g995 ( 
.A(n_921),
.B(n_463),
.Y(n_995)
);

OR2x2_ASAP7_75t_L g996 ( 
.A(n_886),
.B(n_509),
.Y(n_996)
);

NAND2x1p5_ASAP7_75t_L g997 ( 
.A(n_915),
.B(n_908),
.Y(n_997)
);

BUFx4f_ASAP7_75t_L g998 ( 
.A(n_865),
.Y(n_998)
);

INVx1_ASAP7_75t_L g999 ( 
.A(n_911),
.Y(n_999)
);

AOI22xp5_ASAP7_75t_L g1000 ( 
.A1(n_889),
.A2(n_417),
.B1(n_420),
.B2(n_416),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_939),
.A2(n_512),
.B(n_668),
.Y(n_1001)
);

A2O1A1Ixp33_ASAP7_75t_L g1002 ( 
.A1(n_890),
.A2(n_425),
.B(n_426),
.C(n_422),
.Y(n_1002)
);

AOI21xp5_ASAP7_75t_L g1003 ( 
.A1(n_939),
.A2(n_512),
.B(n_429),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_SL g1004 ( 
.A(n_925),
.B(n_427),
.Y(n_1004)
);

OAI22xp5_ASAP7_75t_L g1005 ( 
.A1(n_905),
.A2(n_873),
.B1(n_930),
.B2(n_903),
.Y(n_1005)
);

OR2x2_ASAP7_75t_L g1006 ( 
.A(n_886),
.B(n_510),
.Y(n_1006)
);

BUFx2_ASAP7_75t_L g1007 ( 
.A(n_855),
.Y(n_1007)
);

AOI21xp5_ASAP7_75t_L g1008 ( 
.A1(n_912),
.A2(n_434),
.B(n_433),
.Y(n_1008)
);

AOI21xp5_ASAP7_75t_L g1009 ( 
.A1(n_894),
.A2(n_439),
.B(n_438),
.Y(n_1009)
);

AOI22xp5_ASAP7_75t_L g1010 ( 
.A1(n_902),
.A2(n_445),
.B1(n_446),
.B2(n_443),
.Y(n_1010)
);

NOR3xp33_ASAP7_75t_L g1011 ( 
.A(n_907),
.B(n_527),
.C(n_519),
.Y(n_1011)
);

AOI21xp5_ASAP7_75t_L g1012 ( 
.A1(n_931),
.A2(n_451),
.B(n_449),
.Y(n_1012)
);

NAND2xp5_ASAP7_75t_L g1013 ( 
.A(n_891),
.B(n_465),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_895),
.B(n_466),
.Y(n_1014)
);

OAI21xp5_ASAP7_75t_L g1015 ( 
.A1(n_932),
.A2(n_472),
.B(n_468),
.Y(n_1015)
);

NAND2xp5_ASAP7_75t_L g1016 ( 
.A(n_895),
.B(n_477),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_910),
.B(n_482),
.Y(n_1017)
);

AND2x2_ASAP7_75t_L g1018 ( 
.A(n_909),
.B(n_528),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_944),
.B(n_898),
.Y(n_1019)
);

CKINVDCx5p33_ASAP7_75t_R g1020 ( 
.A(n_990),
.Y(n_1020)
);

AOI21xp5_ASAP7_75t_L g1021 ( 
.A1(n_951),
.A2(n_923),
.B(n_933),
.Y(n_1021)
);

CKINVDCx8_ASAP7_75t_R g1022 ( 
.A(n_1007),
.Y(n_1022)
);

OAI22xp5_ASAP7_75t_L g1023 ( 
.A1(n_957),
.A2(n_924),
.B1(n_937),
.B2(n_938),
.Y(n_1023)
);

AOI22xp33_ASAP7_75t_L g1024 ( 
.A1(n_993),
.A2(n_917),
.B1(n_928),
.B2(n_919),
.Y(n_1024)
);

CKINVDCx6p67_ASAP7_75t_R g1025 ( 
.A(n_986),
.Y(n_1025)
);

OAI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_971),
.A2(n_868),
.B(n_851),
.Y(n_1026)
);

AND2x6_ASAP7_75t_L g1027 ( 
.A(n_971),
.B(n_924),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_L g1028 ( 
.A(n_981),
.B(n_877),
.Y(n_1028)
);

AND2x6_ASAP7_75t_L g1029 ( 
.A(n_957),
.B(n_999),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_941),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_982),
.A2(n_924),
.B(n_929),
.C(n_877),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_947),
.B(n_895),
.Y(n_1032)
);

BUFx8_ASAP7_75t_L g1033 ( 
.A(n_962),
.Y(n_1033)
);

AOI21x1_ASAP7_75t_L g1034 ( 
.A1(n_945),
.A2(n_934),
.B(n_895),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_L g1035 ( 
.A(n_950),
.B(n_861),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_940),
.B(n_895),
.Y(n_1036)
);

AO32x2_ASAP7_75t_L g1037 ( 
.A1(n_1005),
.A2(n_862),
.A3(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_1037)
);

AOI21xp5_ASAP7_75t_L g1038 ( 
.A1(n_967),
.A2(n_494),
.B(n_485),
.Y(n_1038)
);

BUFx2_ASAP7_75t_L g1039 ( 
.A(n_977),
.Y(n_1039)
);

AOI22xp33_ASAP7_75t_L g1040 ( 
.A1(n_1011),
.A2(n_539),
.B1(n_474),
.B2(n_507),
.Y(n_1040)
);

AOI21xp5_ASAP7_75t_L g1041 ( 
.A1(n_988),
.A2(n_508),
.B(n_506),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_SL g1042 ( 
.A(n_977),
.B(n_474),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_994),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_SL g1044 ( 
.A(n_977),
.B(n_514),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_953),
.Y(n_1045)
);

AOI22xp5_ASAP7_75t_L g1046 ( 
.A1(n_1018),
.A2(n_969),
.B1(n_975),
.B2(n_983),
.Y(n_1046)
);

NOR2xp33_ASAP7_75t_L g1047 ( 
.A(n_996),
.B(n_533),
.Y(n_1047)
);

AND2x4_ASAP7_75t_L g1048 ( 
.A(n_970),
.B(n_77),
.Y(n_1048)
);

BUFx2_ASAP7_75t_L g1049 ( 
.A(n_997),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_1006),
.B(n_516),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_956),
.Y(n_1051)
);

NAND3xp33_ASAP7_75t_L g1052 ( 
.A(n_1000),
.B(n_1017),
.C(n_1004),
.Y(n_1052)
);

AOI22xp5_ASAP7_75t_L g1053 ( 
.A1(n_948),
.A2(n_520),
.B1(n_524),
.B2(n_517),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_980),
.B(n_968),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_L g1055 ( 
.A(n_972),
.B(n_525),
.Y(n_1055)
);

A2O1A1Ixp33_ASAP7_75t_L g1056 ( 
.A1(n_949),
.A2(n_537),
.B(n_538),
.C(n_536),
.Y(n_1056)
);

INVx2_ASAP7_75t_L g1057 ( 
.A(n_943),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_SL g1058 ( 
.A(n_970),
.B(n_540),
.Y(n_1058)
);

INVx2_ASAP7_75t_L g1059 ( 
.A(n_943),
.Y(n_1059)
);

CKINVDCx20_ASAP7_75t_R g1060 ( 
.A(n_995),
.Y(n_1060)
);

NOR2xp33_ASAP7_75t_L g1061 ( 
.A(n_1000),
.B(n_5),
.Y(n_1061)
);

INVx4_ASAP7_75t_L g1062 ( 
.A(n_992),
.Y(n_1062)
);

INVx4_ASAP7_75t_L g1063 ( 
.A(n_966),
.Y(n_1063)
);

O2A1O1Ixp33_ASAP7_75t_L g1064 ( 
.A1(n_976),
.A2(n_10),
.B(n_6),
.C(n_9),
.Y(n_1064)
);

INVxp67_ASAP7_75t_L g1065 ( 
.A(n_989),
.Y(n_1065)
);

OAI21xp33_ASAP7_75t_L g1066 ( 
.A1(n_1010),
.A2(n_672),
.B(n_670),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_973),
.B(n_670),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_978),
.B(n_670),
.Y(n_1068)
);

NOR3xp33_ASAP7_75t_SL g1069 ( 
.A(n_1002),
.B(n_10),
.C(n_11),
.Y(n_1069)
);

INVxp67_ASAP7_75t_SL g1070 ( 
.A(n_984),
.Y(n_1070)
);

O2A1O1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_985),
.A2(n_13),
.B(n_11),
.C(n_12),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_952),
.A2(n_678),
.B(n_672),
.Y(n_1072)
);

AND2x2_ASAP7_75t_L g1073 ( 
.A(n_966),
.B(n_672),
.Y(n_1073)
);

OR2x2_ASAP7_75t_L g1074 ( 
.A(n_1013),
.B(n_672),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_984),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1014),
.A2(n_678),
.B(n_80),
.Y(n_1076)
);

NAND2xp5_ASAP7_75t_L g1077 ( 
.A(n_1016),
.B(n_678),
.Y(n_1077)
);

NAND2xp5_ASAP7_75t_L g1078 ( 
.A(n_1015),
.B(n_678),
.Y(n_1078)
);

BUFx6f_ASAP7_75t_L g1079 ( 
.A(n_987),
.Y(n_1079)
);

OAI22xp5_ASAP7_75t_L g1080 ( 
.A1(n_958),
.A2(n_539),
.B1(n_81),
.B2(n_82),
.Y(n_1080)
);

AOI21xp5_ASAP7_75t_L g1081 ( 
.A1(n_954),
.A2(n_83),
.B(n_79),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_959),
.A2(n_87),
.B(n_84),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_965),
.B(n_539),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_1030),
.Y(n_1084)
);

AOI21xp5_ASAP7_75t_L g1085 ( 
.A1(n_1054),
.A2(n_955),
.B(n_960),
.Y(n_1085)
);

INVx2_ASAP7_75t_L g1086 ( 
.A(n_1045),
.Y(n_1086)
);

O2A1O1Ixp5_ASAP7_75t_SL g1087 ( 
.A1(n_1083),
.A2(n_1023),
.B(n_1042),
.C(n_1032),
.Y(n_1087)
);

OAI22xp5_ASAP7_75t_L g1088 ( 
.A1(n_1046),
.A2(n_987),
.B1(n_998),
.B2(n_963),
.Y(n_1088)
);

BUFx5_ASAP7_75t_L g1089 ( 
.A(n_1027),
.Y(n_1089)
);

NOR2xp33_ASAP7_75t_L g1090 ( 
.A(n_1019),
.B(n_998),
.Y(n_1090)
);

AND2x6_ASAP7_75t_L g1091 ( 
.A(n_1048),
.B(n_946),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_1029),
.B(n_1009),
.Y(n_1092)
);

AOI31xp67_ASAP7_75t_L g1093 ( 
.A1(n_1078),
.A2(n_1001),
.A3(n_979),
.B(n_991),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_1036),
.A2(n_961),
.B(n_974),
.Y(n_1094)
);

NAND2xp5_ASAP7_75t_L g1095 ( 
.A(n_1029),
.B(n_1008),
.Y(n_1095)
);

AOI21xp5_ASAP7_75t_L g1096 ( 
.A1(n_1077),
.A2(n_964),
.B(n_942),
.Y(n_1096)
);

OAI21xp5_ASAP7_75t_L g1097 ( 
.A1(n_1052),
.A2(n_1003),
.B(n_1012),
.Y(n_1097)
);

A2O1A1Ixp33_ASAP7_75t_L g1098 ( 
.A1(n_1061),
.A2(n_539),
.B(n_16),
.C(n_12),
.Y(n_1098)
);

AOI22xp5_ASAP7_75t_L g1099 ( 
.A1(n_1028),
.A2(n_539),
.B1(n_17),
.B2(n_15),
.Y(n_1099)
);

INVx5_ASAP7_75t_L g1100 ( 
.A(n_1079),
.Y(n_1100)
);

AOI21xp5_ASAP7_75t_L g1101 ( 
.A1(n_1066),
.A2(n_90),
.B(n_89),
.Y(n_1101)
);

AOI221x1_ASAP7_75t_L g1102 ( 
.A1(n_1056),
.A2(n_15),
.B1(n_16),
.B2(n_18),
.C(n_20),
.Y(n_1102)
);

O2A1O1Ixp33_ASAP7_75t_L g1103 ( 
.A1(n_1071),
.A2(n_18),
.B(n_20),
.C(n_21),
.Y(n_1103)
);

NAND3xp33_ASAP7_75t_L g1104 ( 
.A(n_1047),
.B(n_21),
.C(n_22),
.Y(n_1104)
);

AND2x2_ASAP7_75t_L g1105 ( 
.A(n_1065),
.B(n_23),
.Y(n_1105)
);

NOR2xp33_ASAP7_75t_L g1106 ( 
.A(n_1050),
.B(n_1060),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_1021),
.A2(n_1026),
.B(n_1076),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1067),
.A2(n_95),
.B(n_93),
.Y(n_1108)
);

AOI221xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1064),
.A2(n_1040),
.B1(n_1031),
.B2(n_1080),
.C(n_1043),
.Y(n_1109)
);

A2O1A1Ixp33_ASAP7_75t_L g1110 ( 
.A1(n_1041),
.A2(n_24),
.B(n_25),
.C(n_26),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1068),
.A2(n_1074),
.B(n_1055),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1029),
.B(n_26),
.Y(n_1112)
);

AO22x2_ASAP7_75t_L g1113 ( 
.A1(n_1037),
.A2(n_27),
.B1(n_28),
.B2(n_29),
.Y(n_1113)
);

AO31x2_ASAP7_75t_L g1114 ( 
.A1(n_1072),
.A2(n_1082),
.A3(n_1081),
.B(n_1038),
.Y(n_1114)
);

OR2x2_ASAP7_75t_L g1115 ( 
.A(n_1025),
.B(n_28),
.Y(n_1115)
);

OAI21x1_ASAP7_75t_L g1116 ( 
.A1(n_1034),
.A2(n_97),
.B(n_96),
.Y(n_1116)
);

OAI21x1_ASAP7_75t_L g1117 ( 
.A1(n_1024),
.A2(n_102),
.B(n_100),
.Y(n_1117)
);

NOR2xp33_ASAP7_75t_L g1118 ( 
.A(n_1020),
.B(n_29),
.Y(n_1118)
);

OA21x2_ASAP7_75t_L g1119 ( 
.A1(n_1051),
.A2(n_104),
.B(n_103),
.Y(n_1119)
);

OR2x2_ASAP7_75t_L g1120 ( 
.A(n_1049),
.B(n_30),
.Y(n_1120)
);

NAND2xp5_ASAP7_75t_L g1121 ( 
.A(n_1029),
.B(n_31),
.Y(n_1121)
);

INVx2_ASAP7_75t_L g1122 ( 
.A(n_1057),
.Y(n_1122)
);

INVx5_ASAP7_75t_L g1123 ( 
.A(n_1079),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_1027),
.B(n_31),
.Y(n_1124)
);

OAI22xp5_ASAP7_75t_L g1125 ( 
.A1(n_1070),
.A2(n_32),
.B1(n_33),
.B2(n_34),
.Y(n_1125)
);

AOI21xp5_ASAP7_75t_L g1126 ( 
.A1(n_1058),
.A2(n_107),
.B(n_106),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_1044),
.A2(n_111),
.B(n_108),
.Y(n_1127)
);

INVx4_ASAP7_75t_L g1128 ( 
.A(n_1079),
.Y(n_1128)
);

NOR2xp33_ASAP7_75t_L g1129 ( 
.A(n_1022),
.B(n_33),
.Y(n_1129)
);

AO31x2_ASAP7_75t_L g1130 ( 
.A1(n_1059),
.A2(n_213),
.A3(n_347),
.B(n_345),
.Y(n_1130)
);

OAI21x1_ASAP7_75t_L g1131 ( 
.A1(n_1075),
.A2(n_114),
.B(n_112),
.Y(n_1131)
);

AOI221xp5_ASAP7_75t_SL g1132 ( 
.A1(n_1035),
.A2(n_1073),
.B1(n_1039),
.B2(n_1037),
.C(n_1069),
.Y(n_1132)
);

AOI21xp5_ASAP7_75t_L g1133 ( 
.A1(n_1048),
.A2(n_118),
.B(n_116),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1063),
.B(n_35),
.Y(n_1134)
);

INVxp67_ASAP7_75t_SL g1135 ( 
.A(n_1033),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_1037),
.Y(n_1136)
);

CKINVDCx6p67_ASAP7_75t_R g1137 ( 
.A(n_1062),
.Y(n_1137)
);

NAND2xp5_ASAP7_75t_L g1138 ( 
.A(n_1027),
.B(n_36),
.Y(n_1138)
);

OAI21x1_ASAP7_75t_L g1139 ( 
.A1(n_1053),
.A2(n_122),
.B(n_120),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_1062),
.B(n_1027),
.Y(n_1140)
);

A2O1A1Ixp33_ASAP7_75t_L g1141 ( 
.A1(n_1033),
.A2(n_37),
.B(n_38),
.C(n_39),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1054),
.A2(n_129),
.B(n_124),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1021),
.A2(n_132),
.B(n_130),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1054),
.A2(n_134),
.B(n_133),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_1020),
.Y(n_1145)
);

O2A1O1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1061),
.A2(n_37),
.B(n_42),
.C(n_44),
.Y(n_1146)
);

OAI21xp5_ASAP7_75t_L g1147 ( 
.A1(n_1054),
.A2(n_137),
.B(n_135),
.Y(n_1147)
);

NAND3xp33_ASAP7_75t_SL g1148 ( 
.A(n_1061),
.B(n_42),
.C(n_45),
.Y(n_1148)
);

AO21x2_ASAP7_75t_L g1149 ( 
.A1(n_1078),
.A2(n_143),
.B(n_142),
.Y(n_1149)
);

BUFx4_ASAP7_75t_SL g1150 ( 
.A(n_1020),
.Y(n_1150)
);

OAI21x1_ASAP7_75t_L g1151 ( 
.A1(n_1021),
.A2(n_152),
.B(n_145),
.Y(n_1151)
);

OAI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1021),
.A2(n_159),
.B(n_154),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1054),
.A2(n_162),
.B(n_161),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_1150),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_1137),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_1084),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_SL g1157 ( 
.A1(n_1113),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_1086),
.Y(n_1158)
);

INVx2_ASAP7_75t_SL g1159 ( 
.A(n_1100),
.Y(n_1159)
);

AOI22xp33_ASAP7_75t_L g1160 ( 
.A1(n_1148),
.A2(n_46),
.B1(n_48),
.B2(n_49),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_1122),
.Y(n_1161)
);

INVx4_ASAP7_75t_L g1162 ( 
.A(n_1100),
.Y(n_1162)
);

AOI22xp33_ASAP7_75t_L g1163 ( 
.A1(n_1104),
.A2(n_49),
.B1(n_50),
.B2(n_51),
.Y(n_1163)
);

AOI22xp33_ASAP7_75t_L g1164 ( 
.A1(n_1124),
.A2(n_50),
.B1(n_51),
.B2(n_52),
.Y(n_1164)
);

OAI22xp5_ASAP7_75t_L g1165 ( 
.A1(n_1090),
.A2(n_52),
.B1(n_53),
.B2(n_54),
.Y(n_1165)
);

INVx1_ASAP7_75t_L g1166 ( 
.A(n_1112),
.Y(n_1166)
);

NAND2xp5_ASAP7_75t_L g1167 ( 
.A(n_1106),
.B(n_54),
.Y(n_1167)
);

AOI22xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1113),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_1168)
);

OAI22xp5_ASAP7_75t_L g1169 ( 
.A1(n_1136),
.A2(n_1098),
.B1(n_1121),
.B2(n_1099),
.Y(n_1169)
);

INVx2_ASAP7_75t_L g1170 ( 
.A(n_1131),
.Y(n_1170)
);

BUFx3_ASAP7_75t_L g1171 ( 
.A(n_1145),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_1100),
.Y(n_1172)
);

INVx1_ASAP7_75t_SL g1173 ( 
.A(n_1120),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_1105),
.B(n_55),
.Y(n_1174)
);

INVx1_ASAP7_75t_SL g1175 ( 
.A(n_1123),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_1138),
.Y(n_1176)
);

AOI22xp33_ASAP7_75t_L g1177 ( 
.A1(n_1088),
.A2(n_1147),
.B1(n_1091),
.B2(n_1089),
.Y(n_1177)
);

INVx1_ASAP7_75t_SL g1178 ( 
.A(n_1123),
.Y(n_1178)
);

BUFx6f_ASAP7_75t_L g1179 ( 
.A(n_1123),
.Y(n_1179)
);

INVx4_ASAP7_75t_L g1180 ( 
.A(n_1128),
.Y(n_1180)
);

OAI22x1_ASAP7_75t_L g1181 ( 
.A1(n_1134),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_1140),
.Y(n_1182)
);

INVx2_ASAP7_75t_L g1183 ( 
.A(n_1130),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_1115),
.Y(n_1184)
);

OAI22xp5_ASAP7_75t_L g1185 ( 
.A1(n_1141),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_1185)
);

INVx6_ASAP7_75t_L g1186 ( 
.A(n_1089),
.Y(n_1186)
);

BUFx3_ASAP7_75t_L g1187 ( 
.A(n_1129),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_1139),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1130),
.Y(n_1189)
);

AOI22xp33_ASAP7_75t_SL g1190 ( 
.A1(n_1089),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_1190)
);

INVx1_ASAP7_75t_L g1191 ( 
.A(n_1110),
.Y(n_1191)
);

INVx6_ASAP7_75t_L g1192 ( 
.A(n_1089),
.Y(n_1192)
);

BUFx12f_ASAP7_75t_L g1193 ( 
.A(n_1091),
.Y(n_1193)
);

INVx2_ASAP7_75t_L g1194 ( 
.A(n_1116),
.Y(n_1194)
);

AOI22xp33_ASAP7_75t_SL g1195 ( 
.A1(n_1118),
.A2(n_62),
.B1(n_63),
.B2(n_65),
.Y(n_1195)
);

INVx2_ASAP7_75t_L g1196 ( 
.A(n_1149),
.Y(n_1196)
);

BUFx6f_ASAP7_75t_L g1197 ( 
.A(n_1091),
.Y(n_1197)
);

AOI22xp33_ASAP7_75t_L g1198 ( 
.A1(n_1092),
.A2(n_65),
.B1(n_66),
.B2(n_67),
.Y(n_1198)
);

AOI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1095),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_1199)
);

INVx1_ASAP7_75t_L g1200 ( 
.A(n_1125),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_L g1201 ( 
.A1(n_1101),
.A2(n_1097),
.B1(n_1111),
.B2(n_1133),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1102),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_L g1203 ( 
.A(n_1119),
.Y(n_1203)
);

AOI22xp33_ASAP7_75t_SL g1204 ( 
.A1(n_1135),
.A2(n_68),
.B1(n_70),
.B2(n_71),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_SL g1205 ( 
.A1(n_1117),
.A2(n_70),
.B1(n_71),
.B2(n_72),
.Y(n_1205)
);

AOI22xp33_ASAP7_75t_SL g1206 ( 
.A1(n_1142),
.A2(n_73),
.B1(n_74),
.B2(n_76),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1132),
.B(n_76),
.Y(n_1207)
);

AOI22xp5_ASAP7_75t_L g1208 ( 
.A1(n_1109),
.A2(n_163),
.B1(n_164),
.B2(n_165),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_1146),
.Y(n_1209)
);

AOI22xp33_ASAP7_75t_L g1210 ( 
.A1(n_1127),
.A2(n_167),
.B1(n_170),
.B2(n_171),
.Y(n_1210)
);

NAND2x1p5_ASAP7_75t_L g1211 ( 
.A(n_1143),
.B(n_173),
.Y(n_1211)
);

AOI22xp33_ASAP7_75t_L g1212 ( 
.A1(n_1126),
.A2(n_174),
.B1(n_177),
.B2(n_181),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1151),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1152),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1103),
.B(n_348),
.Y(n_1215)
);

INVx6_ASAP7_75t_L g1216 ( 
.A(n_1087),
.Y(n_1216)
);

BUFx8_ASAP7_75t_L g1217 ( 
.A(n_1108),
.Y(n_1217)
);

AND2x2_ASAP7_75t_L g1218 ( 
.A(n_1144),
.B(n_187),
.Y(n_1218)
);

OAI21xp33_ASAP7_75t_L g1219 ( 
.A1(n_1085),
.A2(n_191),
.B(n_192),
.Y(n_1219)
);

AOI22xp33_ASAP7_75t_L g1220 ( 
.A1(n_1153),
.A2(n_194),
.B1(n_195),
.B2(n_198),
.Y(n_1220)
);

NAND2xp5_ASAP7_75t_L g1221 ( 
.A(n_1107),
.B(n_200),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_L g1222 ( 
.A(n_1094),
.B(n_344),
.Y(n_1222)
);

AOI22xp5_ASAP7_75t_L g1223 ( 
.A1(n_1096),
.A2(n_201),
.B1(n_202),
.B2(n_203),
.Y(n_1223)
);

INVx3_ASAP7_75t_L g1224 ( 
.A(n_1114),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1114),
.Y(n_1225)
);

NAND2x1p5_ASAP7_75t_L g1226 ( 
.A(n_1093),
.B(n_204),
.Y(n_1226)
);

CKINVDCx6p67_ASAP7_75t_R g1227 ( 
.A(n_1100),
.Y(n_1227)
);

BUFx4f_ASAP7_75t_SL g1228 ( 
.A(n_1137),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_1166),
.B(n_206),
.Y(n_1229)
);

AND2x2_ASAP7_75t_L g1230 ( 
.A(n_1176),
.B(n_343),
.Y(n_1230)
);

INVx3_ASAP7_75t_L g1231 ( 
.A(n_1186),
.Y(n_1231)
);

OAI21x1_ASAP7_75t_L g1232 ( 
.A1(n_1224),
.A2(n_207),
.B(n_214),
.Y(n_1232)
);

AND2x2_ASAP7_75t_SL g1233 ( 
.A(n_1177),
.B(n_218),
.Y(n_1233)
);

INVx1_ASAP7_75t_L g1234 ( 
.A(n_1156),
.Y(n_1234)
);

INVxp67_ASAP7_75t_L g1235 ( 
.A(n_1173),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_1207),
.B(n_341),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1158),
.Y(n_1237)
);

BUFx2_ASAP7_75t_L g1238 ( 
.A(n_1225),
.Y(n_1238)
);

INVxp67_ASAP7_75t_L g1239 ( 
.A(n_1173),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_1161),
.Y(n_1240)
);

CKINVDCx8_ASAP7_75t_R g1241 ( 
.A(n_1154),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_1183),
.Y(n_1242)
);

AND2x2_ASAP7_75t_L g1243 ( 
.A(n_1182),
.B(n_221),
.Y(n_1243)
);

BUFx2_ASAP7_75t_L g1244 ( 
.A(n_1182),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1202),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1184),
.B(n_222),
.Y(n_1246)
);

INVxp67_ASAP7_75t_L g1247 ( 
.A(n_1187),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1189),
.Y(n_1248)
);

INVx2_ASAP7_75t_SL g1249 ( 
.A(n_1186),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1170),
.Y(n_1250)
);

INVxp67_ASAP7_75t_L g1251 ( 
.A(n_1184),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_1209),
.B(n_223),
.Y(n_1252)
);

OA21x2_ASAP7_75t_L g1253 ( 
.A1(n_1196),
.A2(n_225),
.B(n_229),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1226),
.Y(n_1254)
);

OR2x6_ASAP7_75t_L g1255 ( 
.A(n_1188),
.B(n_230),
.Y(n_1255)
);

AOI21xp5_ASAP7_75t_L g1256 ( 
.A1(n_1201),
.A2(n_1219),
.B(n_1221),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1197),
.Y(n_1257)
);

AND2x2_ASAP7_75t_L g1258 ( 
.A(n_1197),
.B(n_231),
.Y(n_1258)
);

INVx3_ASAP7_75t_L g1259 ( 
.A(n_1192),
.Y(n_1259)
);

INVx2_ASAP7_75t_L g1260 ( 
.A(n_1226),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1197),
.Y(n_1261)
);

INVx2_ASAP7_75t_L g1262 ( 
.A(n_1194),
.Y(n_1262)
);

INVx1_ASAP7_75t_L g1263 ( 
.A(n_1169),
.Y(n_1263)
);

INVx2_ASAP7_75t_SL g1264 ( 
.A(n_1192),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_1213),
.A2(n_234),
.B(n_236),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1169),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1214),
.Y(n_1267)
);

CKINVDCx5p33_ASAP7_75t_R g1268 ( 
.A(n_1171),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1191),
.Y(n_1269)
);

INVx2_ASAP7_75t_L g1270 ( 
.A(n_1203),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1188),
.Y(n_1271)
);

INVx1_ASAP7_75t_SL g1272 ( 
.A(n_1175),
.Y(n_1272)
);

INVx3_ASAP7_75t_L g1273 ( 
.A(n_1188),
.Y(n_1273)
);

INVx1_ASAP7_75t_L g1274 ( 
.A(n_1172),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1200),
.Y(n_1275)
);

INVx3_ASAP7_75t_L g1276 ( 
.A(n_1203),
.Y(n_1276)
);

INVx1_ASAP7_75t_L g1277 ( 
.A(n_1216),
.Y(n_1277)
);

INVx1_ASAP7_75t_L g1278 ( 
.A(n_1216),
.Y(n_1278)
);

INVx1_ASAP7_75t_L g1279 ( 
.A(n_1175),
.Y(n_1279)
);

INVx4_ASAP7_75t_L g1280 ( 
.A(n_1179),
.Y(n_1280)
);

AOI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1222),
.A2(n_237),
.B(n_239),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1179),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1211),
.Y(n_1283)
);

INVx2_ASAP7_75t_L g1284 ( 
.A(n_1211),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1219),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1208),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1223),
.A2(n_1208),
.B(n_1218),
.Y(n_1287)
);

BUFx3_ASAP7_75t_L g1288 ( 
.A(n_1179),
.Y(n_1288)
);

INVx2_ASAP7_75t_L g1289 ( 
.A(n_1193),
.Y(n_1289)
);

INVx3_ASAP7_75t_L g1290 ( 
.A(n_1217),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1217),
.Y(n_1291)
);

INVx1_ASAP7_75t_L g1292 ( 
.A(n_1178),
.Y(n_1292)
);

HB1xp67_ASAP7_75t_L g1293 ( 
.A(n_1178),
.Y(n_1293)
);

OAI22xp5_ASAP7_75t_L g1294 ( 
.A1(n_1160),
.A2(n_241),
.B1(n_243),
.B2(n_245),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1159),
.Y(n_1295)
);

AO21x1_ASAP7_75t_L g1296 ( 
.A1(n_1185),
.A2(n_247),
.B(n_250),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1163),
.B(n_1164),
.Y(n_1297)
);

OR2x2_ASAP7_75t_L g1298 ( 
.A(n_1244),
.B(n_1235),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1244),
.B(n_1174),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1267),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1239),
.B(n_1167),
.Y(n_1301)
);

OR2x2_ASAP7_75t_L g1302 ( 
.A(n_1251),
.B(n_1215),
.Y(n_1302)
);

INVx3_ASAP7_75t_L g1303 ( 
.A(n_1290),
.Y(n_1303)
);

AOI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1256),
.A2(n_1223),
.B(n_1220),
.Y(n_1304)
);

AND2x2_ASAP7_75t_L g1305 ( 
.A(n_1234),
.B(n_1181),
.Y(n_1305)
);

AO32x2_ASAP7_75t_L g1306 ( 
.A1(n_1249),
.A2(n_1185),
.A3(n_1165),
.B1(n_1168),
.B2(n_1157),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1279),
.B(n_1205),
.Y(n_1307)
);

NOR2x1_ASAP7_75t_SL g1308 ( 
.A(n_1255),
.B(n_1270),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1292),
.B(n_1190),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1245),
.B(n_1198),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1270),
.B(n_1206),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1237),
.B(n_1195),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_1241),
.Y(n_1313)
);

BUFx2_ASAP7_75t_L g1314 ( 
.A(n_1293),
.Y(n_1314)
);

AOI221xp5_ASAP7_75t_L g1315 ( 
.A1(n_1263),
.A2(n_1199),
.B1(n_1204),
.B2(n_1212),
.C(n_1210),
.Y(n_1315)
);

OAI22xp5_ASAP7_75t_L g1316 ( 
.A1(n_1233),
.A2(n_1227),
.B1(n_1155),
.B2(n_1162),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1247),
.B(n_1268),
.Y(n_1317)
);

CKINVDCx5p33_ASAP7_75t_R g1318 ( 
.A(n_1241),
.Y(n_1318)
);

AND2x4_ASAP7_75t_L g1319 ( 
.A(n_1276),
.B(n_1162),
.Y(n_1319)
);

NAND3xp33_ASAP7_75t_L g1320 ( 
.A(n_1266),
.B(n_1180),
.C(n_1228),
.Y(n_1320)
);

AND2x2_ASAP7_75t_L g1321 ( 
.A(n_1236),
.B(n_1180),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1238),
.B(n_251),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1275),
.Y(n_1323)
);

HB1xp67_ASAP7_75t_L g1324 ( 
.A(n_1238),
.Y(n_1324)
);

AND2x2_ASAP7_75t_L g1325 ( 
.A(n_1236),
.B(n_339),
.Y(n_1325)
);

A2O1A1Ixp33_ASAP7_75t_L g1326 ( 
.A1(n_1287),
.A2(n_253),
.B(n_255),
.C(n_258),
.Y(n_1326)
);

AND2x2_ASAP7_75t_L g1327 ( 
.A(n_1274),
.B(n_1240),
.Y(n_1327)
);

AND2x2_ASAP7_75t_SL g1328 ( 
.A(n_1233),
.B(n_260),
.Y(n_1328)
);

AND2x2_ASAP7_75t_L g1329 ( 
.A(n_1243),
.B(n_1289),
.Y(n_1329)
);

AND2x4_ASAP7_75t_L g1330 ( 
.A(n_1276),
.B(n_262),
.Y(n_1330)
);

OR2x6_ASAP7_75t_L g1331 ( 
.A(n_1290),
.B(n_264),
.Y(n_1331)
);

BUFx3_ASAP7_75t_L g1332 ( 
.A(n_1268),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1269),
.B(n_266),
.Y(n_1333)
);

AND2x4_ASAP7_75t_L g1334 ( 
.A(n_1276),
.B(n_334),
.Y(n_1334)
);

AND2x4_ASAP7_75t_L g1335 ( 
.A(n_1290),
.B(n_267),
.Y(n_1335)
);

HB1xp67_ASAP7_75t_L g1336 ( 
.A(n_1272),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1291),
.B(n_332),
.Y(n_1337)
);

AND2x2_ASAP7_75t_L g1338 ( 
.A(n_1243),
.B(n_269),
.Y(n_1338)
);

INVxp67_ASAP7_75t_L g1339 ( 
.A(n_1295),
.Y(n_1339)
);

NOR2x1_ASAP7_75t_L g1340 ( 
.A(n_1291),
.B(n_270),
.Y(n_1340)
);

AOI21xp5_ASAP7_75t_L g1341 ( 
.A1(n_1287),
.A2(n_271),
.B(n_273),
.Y(n_1341)
);

BUFx5_ASAP7_75t_L g1342 ( 
.A(n_1242),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1285),
.B(n_275),
.Y(n_1343)
);

OAI21x1_ASAP7_75t_SL g1344 ( 
.A1(n_1296),
.A2(n_276),
.B(n_278),
.Y(n_1344)
);

O2A1O1Ixp33_ASAP7_75t_SL g1345 ( 
.A1(n_1291),
.A2(n_280),
.B(n_281),
.C(n_282),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1242),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1248),
.Y(n_1347)
);

NOR2xp33_ASAP7_75t_SL g1348 ( 
.A(n_1289),
.B(n_283),
.Y(n_1348)
);

NAND2x1_ASAP7_75t_L g1349 ( 
.A(n_1283),
.B(n_284),
.Y(n_1349)
);

NAND2xp33_ASAP7_75t_R g1350 ( 
.A(n_1258),
.B(n_1231),
.Y(n_1350)
);

INVx1_ASAP7_75t_L g1351 ( 
.A(n_1300),
.Y(n_1351)
);

CKINVDCx20_ASAP7_75t_R g1352 ( 
.A(n_1313),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1300),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1328),
.A2(n_1286),
.B1(n_1297),
.B2(n_1285),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1346),
.Y(n_1355)
);

INVx1_ASAP7_75t_L g1356 ( 
.A(n_1346),
.Y(n_1356)
);

AND2x4_ASAP7_75t_SL g1357 ( 
.A(n_1324),
.B(n_1255),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1314),
.B(n_1286),
.Y(n_1358)
);

NAND2x1p5_ASAP7_75t_L g1359 ( 
.A(n_1341),
.B(n_1253),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1347),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1323),
.Y(n_1361)
);

AOI22xp33_ASAP7_75t_L g1362 ( 
.A1(n_1304),
.A2(n_1296),
.B1(n_1294),
.B2(n_1283),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1327),
.Y(n_1363)
);

NAND3xp33_ASAP7_75t_L g1364 ( 
.A(n_1315),
.B(n_1252),
.C(n_1246),
.Y(n_1364)
);

NAND2xp5_ASAP7_75t_L g1365 ( 
.A(n_1298),
.B(n_1250),
.Y(n_1365)
);

INVx3_ASAP7_75t_L g1366 ( 
.A(n_1342),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1342),
.Y(n_1367)
);

INVx2_ASAP7_75t_L g1368 ( 
.A(n_1342),
.Y(n_1368)
);

INVx2_ASAP7_75t_L g1369 ( 
.A(n_1339),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1303),
.Y(n_1370)
);

AND2x4_ASAP7_75t_L g1371 ( 
.A(n_1303),
.B(n_1271),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1305),
.Y(n_1372)
);

NAND2xp5_ASAP7_75t_L g1373 ( 
.A(n_1336),
.B(n_1250),
.Y(n_1373)
);

BUFx2_ASAP7_75t_L g1374 ( 
.A(n_1319),
.Y(n_1374)
);

INVx2_ASAP7_75t_SL g1375 ( 
.A(n_1319),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1302),
.Y(n_1376)
);

INVx4_ASAP7_75t_L g1377 ( 
.A(n_1331),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1329),
.B(n_1262),
.Y(n_1378)
);

INVx2_ASAP7_75t_L g1379 ( 
.A(n_1308),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1353),
.Y(n_1380)
);

OAI21xp33_ASAP7_75t_L g1381 ( 
.A1(n_1364),
.A2(n_1307),
.B(n_1326),
.Y(n_1381)
);

AND2x2_ASAP7_75t_L g1382 ( 
.A(n_1372),
.B(n_1299),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1351),
.Y(n_1383)
);

NAND2xp5_ASAP7_75t_L g1384 ( 
.A(n_1376),
.B(n_1301),
.Y(n_1384)
);

AND2x2_ASAP7_75t_L g1385 ( 
.A(n_1372),
.B(n_1321),
.Y(n_1385)
);

AOI22xp5_ASAP7_75t_L g1386 ( 
.A1(n_1364),
.A2(n_1316),
.B1(n_1348),
.B2(n_1320),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1376),
.B(n_1317),
.Y(n_1387)
);

AND2x2_ASAP7_75t_L g1388 ( 
.A(n_1374),
.B(n_1332),
.Y(n_1388)
);

OR2x2_ASAP7_75t_L g1389 ( 
.A(n_1369),
.B(n_1310),
.Y(n_1389)
);

AO21x2_ASAP7_75t_L g1390 ( 
.A1(n_1367),
.A2(n_1344),
.B(n_1262),
.Y(n_1390)
);

NAND4xp25_ASAP7_75t_L g1391 ( 
.A(n_1362),
.B(n_1312),
.C(n_1309),
.D(n_1311),
.Y(n_1391)
);

NAND4xp25_ASAP7_75t_SL g1392 ( 
.A(n_1379),
.B(n_1340),
.C(n_1306),
.D(n_1257),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1353),
.Y(n_1393)
);

AND2x2_ASAP7_75t_L g1394 ( 
.A(n_1374),
.B(n_1363),
.Y(n_1394)
);

NOR3xp33_ASAP7_75t_L g1395 ( 
.A(n_1354),
.B(n_1343),
.C(n_1229),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1369),
.Y(n_1396)
);

OA21x2_ASAP7_75t_L g1397 ( 
.A1(n_1367),
.A2(n_1277),
.B(n_1278),
.Y(n_1397)
);

INVx2_ASAP7_75t_L g1398 ( 
.A(n_1353),
.Y(n_1398)
);

OR2x2_ASAP7_75t_SL g1399 ( 
.A(n_1379),
.B(n_1322),
.Y(n_1399)
);

INVx4_ASAP7_75t_L g1400 ( 
.A(n_1377),
.Y(n_1400)
);

OR2x2_ASAP7_75t_L g1401 ( 
.A(n_1369),
.B(n_1271),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1352),
.Y(n_1402)
);

OA21x2_ASAP7_75t_L g1403 ( 
.A1(n_1368),
.A2(n_1254),
.B(n_1260),
.Y(n_1403)
);

AND2x2_ASAP7_75t_L g1404 ( 
.A(n_1394),
.B(n_1375),
.Y(n_1404)
);

AND2x4_ASAP7_75t_SL g1405 ( 
.A(n_1388),
.B(n_1377),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1389),
.B(n_1363),
.Y(n_1406)
);

BUFx3_ASAP7_75t_L g1407 ( 
.A(n_1402),
.Y(n_1407)
);

OR2x2_ASAP7_75t_L g1408 ( 
.A(n_1389),
.B(n_1358),
.Y(n_1408)
);

AND2x4_ASAP7_75t_SL g1409 ( 
.A(n_1388),
.B(n_1377),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1387),
.B(n_1378),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1394),
.B(n_1385),
.Y(n_1411)
);

AND2x2_ASAP7_75t_L g1412 ( 
.A(n_1385),
.B(n_1375),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1383),
.Y(n_1413)
);

BUFx2_ASAP7_75t_L g1414 ( 
.A(n_1400),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1396),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1401),
.Y(n_1416)
);

INVx1_ASAP7_75t_L g1417 ( 
.A(n_1380),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1413),
.Y(n_1418)
);

NAND2xp5_ASAP7_75t_L g1419 ( 
.A(n_1410),
.B(n_1387),
.Y(n_1419)
);

OAI22xp33_ASAP7_75t_L g1420 ( 
.A1(n_1407),
.A2(n_1391),
.B1(n_1386),
.B2(n_1350),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1406),
.Y(n_1421)
);

INVx1_ASAP7_75t_SL g1422 ( 
.A(n_1407),
.Y(n_1422)
);

OAI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1408),
.A2(n_1377),
.B1(n_1400),
.B2(n_1392),
.Y(n_1423)
);

AND2x2_ASAP7_75t_L g1424 ( 
.A(n_1405),
.B(n_1382),
.Y(n_1424)
);

OR2x2_ASAP7_75t_L g1425 ( 
.A(n_1408),
.B(n_1399),
.Y(n_1425)
);

AND2x2_ASAP7_75t_L g1426 ( 
.A(n_1405),
.B(n_1382),
.Y(n_1426)
);

INVx2_ASAP7_75t_L g1427 ( 
.A(n_1411),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1417),
.Y(n_1428)
);

OR2x2_ASAP7_75t_L g1429 ( 
.A(n_1415),
.B(n_1399),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1409),
.B(n_1381),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1411),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1416),
.B(n_1384),
.Y(n_1432)
);

INVxp67_ASAP7_75t_L g1433 ( 
.A(n_1414),
.Y(n_1433)
);

INVx2_ASAP7_75t_L g1434 ( 
.A(n_1422),
.Y(n_1434)
);

AO21x2_ASAP7_75t_L g1435 ( 
.A1(n_1433),
.A2(n_1423),
.B(n_1420),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1427),
.B(n_1414),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1430),
.B(n_1416),
.Y(n_1437)
);

AND2x2_ASAP7_75t_L g1438 ( 
.A(n_1424),
.B(n_1409),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1419),
.B(n_1401),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1418),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_1426),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1431),
.B(n_1404),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1430),
.B(n_1412),
.Y(n_1443)
);

AOI22xp33_ASAP7_75t_L g1444 ( 
.A1(n_1435),
.A2(n_1420),
.B1(n_1395),
.B2(n_1423),
.Y(n_1444)
);

AOI21xp5_ASAP7_75t_L g1445 ( 
.A1(n_1435),
.A2(n_1437),
.B(n_1443),
.Y(n_1445)
);

OAI222xp33_ASAP7_75t_L g1446 ( 
.A1(n_1441),
.A2(n_1425),
.B1(n_1429),
.B2(n_1434),
.C1(n_1433),
.C2(n_1436),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1440),
.Y(n_1447)
);

O2A1O1Ixp33_ASAP7_75t_SL g1448 ( 
.A1(n_1441),
.A2(n_1434),
.B(n_1432),
.C(n_1428),
.Y(n_1448)
);

INVxp67_ASAP7_75t_SL g1449 ( 
.A(n_1436),
.Y(n_1449)
);

INVx2_ASAP7_75t_L g1450 ( 
.A(n_1442),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1442),
.Y(n_1451)
);

INVx1_ASAP7_75t_L g1452 ( 
.A(n_1439),
.Y(n_1452)
);

AOI22xp33_ASAP7_75t_L g1453 ( 
.A1(n_1444),
.A2(n_1445),
.B1(n_1452),
.B2(n_1451),
.Y(n_1453)
);

AND2x4_ASAP7_75t_L g1454 ( 
.A(n_1449),
.B(n_1450),
.Y(n_1454)
);

INVx1_ASAP7_75t_SL g1455 ( 
.A(n_1450),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1447),
.Y(n_1456)
);

O2A1O1Ixp33_ASAP7_75t_L g1457 ( 
.A1(n_1446),
.A2(n_1345),
.B(n_1421),
.C(n_1438),
.Y(n_1457)
);

NOR2xp67_ASAP7_75t_L g1458 ( 
.A(n_1444),
.B(n_1400),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1448),
.B(n_1402),
.Y(n_1459)
);

OAI22xp5_ASAP7_75t_L g1460 ( 
.A1(n_1453),
.A2(n_1318),
.B1(n_1404),
.B2(n_1412),
.Y(n_1460)
);

XNOR2xp5_ASAP7_75t_L g1461 ( 
.A(n_1458),
.B(n_1335),
.Y(n_1461)
);

OAI211xp5_ASAP7_75t_L g1462 ( 
.A1(n_1457),
.A2(n_1258),
.B(n_1349),
.C(n_1325),
.Y(n_1462)
);

NOR3xp33_ASAP7_75t_L g1463 ( 
.A(n_1459),
.B(n_1338),
.C(n_1333),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1455),
.A2(n_1454),
.B1(n_1456),
.B2(n_1359),
.Y(n_1464)
);

OAI31xp33_ASAP7_75t_L g1465 ( 
.A1(n_1454),
.A2(n_1359),
.A3(n_1357),
.B(n_1337),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1454),
.Y(n_1466)
);

INVx1_ASAP7_75t_SL g1467 ( 
.A(n_1459),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1454),
.Y(n_1468)
);

INVx1_ASAP7_75t_L g1469 ( 
.A(n_1466),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1468),
.Y(n_1470)
);

NAND4xp25_ASAP7_75t_L g1471 ( 
.A(n_1467),
.B(n_1462),
.C(n_1463),
.D(n_1464),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1461),
.Y(n_1472)
);

AND2x2_ASAP7_75t_L g1473 ( 
.A(n_1460),
.B(n_1378),
.Y(n_1473)
);

NOR4xp25_ASAP7_75t_L g1474 ( 
.A(n_1465),
.B(n_1230),
.C(n_1261),
.D(n_1361),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1466),
.Y(n_1475)
);

NAND4xp25_ASAP7_75t_L g1476 ( 
.A(n_1467),
.B(n_1337),
.C(n_1335),
.D(n_1334),
.Y(n_1476)
);

NAND3xp33_ASAP7_75t_SL g1477 ( 
.A(n_1469),
.B(n_1230),
.C(n_1280),
.Y(n_1477)
);

NAND4xp25_ASAP7_75t_L g1478 ( 
.A(n_1471),
.B(n_1330),
.C(n_1334),
.D(n_1288),
.Y(n_1478)
);

O2A1O1Ixp33_ASAP7_75t_L g1479 ( 
.A1(n_1470),
.A2(n_1475),
.B(n_1472),
.C(n_1476),
.Y(n_1479)
);

AOI221x1_ASAP7_75t_L g1480 ( 
.A1(n_1473),
.A2(n_1330),
.B1(n_1282),
.B2(n_1280),
.C(n_1380),
.Y(n_1480)
);

AOI321xp33_ASAP7_75t_L g1481 ( 
.A1(n_1474),
.A2(n_1306),
.A3(n_1288),
.B1(n_1373),
.B2(n_1284),
.C(n_1365),
.Y(n_1481)
);

AOI22xp5_ASAP7_75t_L g1482 ( 
.A1(n_1471),
.A2(n_1331),
.B1(n_1357),
.B2(n_1390),
.Y(n_1482)
);

OAI222xp33_ASAP7_75t_L g1483 ( 
.A1(n_1469),
.A2(n_1255),
.B1(n_1359),
.B2(n_1280),
.C1(n_1282),
.C2(n_1249),
.Y(n_1483)
);

AOI221xp5_ASAP7_75t_L g1484 ( 
.A1(n_1479),
.A2(n_1478),
.B1(n_1482),
.B2(n_1477),
.C(n_1483),
.Y(n_1484)
);

AOI211xp5_ASAP7_75t_L g1485 ( 
.A1(n_1481),
.A2(n_1265),
.B(n_1232),
.C(n_1361),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1480),
.B(n_1393),
.Y(n_1486)
);

NAND2x1_ASAP7_75t_L g1487 ( 
.A(n_1482),
.B(n_1397),
.Y(n_1487)
);

AOI221xp5_ASAP7_75t_L g1488 ( 
.A1(n_1479),
.A2(n_1393),
.B1(n_1264),
.B2(n_1390),
.C(n_1357),
.Y(n_1488)
);

OR2x2_ASAP7_75t_L g1489 ( 
.A(n_1478),
.B(n_1398),
.Y(n_1489)
);

HB1xp67_ASAP7_75t_L g1490 ( 
.A(n_1478),
.Y(n_1490)
);

AOI221xp5_ASAP7_75t_L g1491 ( 
.A1(n_1479),
.A2(n_1264),
.B1(n_1390),
.B2(n_1259),
.C(n_1231),
.Y(n_1491)
);

NAND2xp5_ASAP7_75t_L g1492 ( 
.A(n_1479),
.B(n_1398),
.Y(n_1492)
);

NOR2x1_ASAP7_75t_L g1493 ( 
.A(n_1492),
.B(n_1255),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1490),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1489),
.B(n_1486),
.Y(n_1495)
);

NAND2xp5_ASAP7_75t_L g1496 ( 
.A(n_1484),
.B(n_1397),
.Y(n_1496)
);

XNOR2xp5_ASAP7_75t_L g1497 ( 
.A(n_1491),
.B(n_1488),
.Y(n_1497)
);

NOR2xp33_ASAP7_75t_L g1498 ( 
.A(n_1487),
.B(n_1282),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1485),
.B(n_1231),
.Y(n_1499)
);

AND2x2_ASAP7_75t_SL g1500 ( 
.A(n_1490),
.B(n_1253),
.Y(n_1500)
);

OAI22xp5_ASAP7_75t_L g1501 ( 
.A1(n_1485),
.A2(n_1370),
.B1(n_1368),
.B2(n_1371),
.Y(n_1501)
);

XNOR2xp5_ASAP7_75t_L g1502 ( 
.A(n_1490),
.B(n_1281),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1492),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1492),
.Y(n_1504)
);

NOR2xp33_ASAP7_75t_SL g1505 ( 
.A(n_1490),
.B(n_1371),
.Y(n_1505)
);

INVx2_ASAP7_75t_SL g1506 ( 
.A(n_1489),
.Y(n_1506)
);

NAND4xp25_ASAP7_75t_L g1507 ( 
.A(n_1505),
.B(n_1259),
.C(n_1371),
.D(n_1284),
.Y(n_1507)
);

NAND3xp33_ASAP7_75t_L g1508 ( 
.A(n_1494),
.B(n_1253),
.C(n_1259),
.Y(n_1508)
);

INVx2_ASAP7_75t_L g1509 ( 
.A(n_1495),
.Y(n_1509)
);

NAND2x1p5_ASAP7_75t_L g1510 ( 
.A(n_1506),
.B(n_1265),
.Y(n_1510)
);

AOI22xp33_ASAP7_75t_L g1511 ( 
.A1(n_1496),
.A2(n_1371),
.B1(n_1397),
.B2(n_1366),
.Y(n_1511)
);

OAI21xp5_ASAP7_75t_L g1512 ( 
.A1(n_1497),
.A2(n_1232),
.B(n_1281),
.Y(n_1512)
);

OAI21xp5_ASAP7_75t_L g1513 ( 
.A1(n_1502),
.A2(n_1370),
.B(n_1351),
.Y(n_1513)
);

AO22x2_ASAP7_75t_L g1514 ( 
.A1(n_1509),
.A2(n_1504),
.B1(n_1503),
.B2(n_1501),
.Y(n_1514)
);

AOI22xp5_ASAP7_75t_L g1515 ( 
.A1(n_1507),
.A2(n_1499),
.B1(n_1498),
.B2(n_1493),
.Y(n_1515)
);

NAND2xp5_ASAP7_75t_L g1516 ( 
.A(n_1511),
.B(n_1500),
.Y(n_1516)
);

NAND2xp5_ASAP7_75t_SL g1517 ( 
.A(n_1512),
.B(n_1366),
.Y(n_1517)
);

OAI22x1_ASAP7_75t_L g1518 ( 
.A1(n_1515),
.A2(n_1508),
.B1(n_1510),
.B2(n_1513),
.Y(n_1518)
);

HB1xp67_ASAP7_75t_L g1519 ( 
.A(n_1516),
.Y(n_1519)
);

AOI22xp5_ASAP7_75t_L g1520 ( 
.A1(n_1514),
.A2(n_1397),
.B1(n_1366),
.B2(n_1355),
.Y(n_1520)
);

INVx1_ASAP7_75t_L g1521 ( 
.A(n_1517),
.Y(n_1521)
);

OAI22xp5_ASAP7_75t_SL g1522 ( 
.A1(n_1519),
.A2(n_1403),
.B1(n_1366),
.B2(n_1355),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1521),
.Y(n_1523)
);

OAI22x1_ASAP7_75t_L g1524 ( 
.A1(n_1520),
.A2(n_1403),
.B1(n_1356),
.B2(n_1360),
.Y(n_1524)
);

BUFx2_ASAP7_75t_L g1525 ( 
.A(n_1523),
.Y(n_1525)
);

AOI21xp5_ASAP7_75t_L g1526 ( 
.A1(n_1524),
.A2(n_1518),
.B(n_1403),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1522),
.Y(n_1527)
);

INVx2_ASAP7_75t_L g1528 ( 
.A(n_1525),
.Y(n_1528)
);

AOI22xp33_ASAP7_75t_L g1529 ( 
.A1(n_1528),
.A2(n_1527),
.B1(n_1526),
.B2(n_1356),
.Y(n_1529)
);

OAI22x1_ASAP7_75t_L g1530 ( 
.A1(n_1529),
.A2(n_1403),
.B1(n_1273),
.B2(n_1271),
.Y(n_1530)
);

AOI22x1_ASAP7_75t_L g1531 ( 
.A1(n_1530),
.A2(n_287),
.B1(n_289),
.B2(n_290),
.Y(n_1531)
);

OAI221xp5_ASAP7_75t_R g1532 ( 
.A1(n_1531),
.A2(n_294),
.B1(n_297),
.B2(n_298),
.C(n_299),
.Y(n_1532)
);

AOI211xp5_ASAP7_75t_L g1533 ( 
.A1(n_1532),
.A2(n_304),
.B(n_305),
.C(n_307),
.Y(n_1533)
);


endmodule