module fake_netlist_5_7_n_162 (n_16, n_0, n_12, n_9, n_25, n_18, n_27, n_22, n_1, n_8, n_10, n_24, n_21, n_4, n_11, n_17, n_19, n_7, n_15, n_26, n_20, n_5, n_14, n_2, n_23, n_13, n_3, n_6, n_162);

input n_16;
input n_0;
input n_12;
input n_9;
input n_25;
input n_18;
input n_27;
input n_22;
input n_1;
input n_8;
input n_10;
input n_24;
input n_21;
input n_4;
input n_11;
input n_17;
input n_19;
input n_7;
input n_15;
input n_26;
input n_20;
input n_5;
input n_14;
input n_2;
input n_23;
input n_13;
input n_3;
input n_6;

output n_162;

wire n_137;
wire n_91;
wire n_82;
wire n_122;
wire n_142;
wire n_140;
wire n_136;
wire n_86;
wire n_124;
wire n_146;
wire n_143;
wire n_83;
wire n_132;
wire n_61;
wire n_90;
wire n_127;
wire n_75;
wire n_101;
wire n_65;
wire n_78;
wire n_74;
wire n_144;
wire n_114;
wire n_96;
wire n_57;
wire n_37;
wire n_111;
wire n_108;
wire n_129;
wire n_31;
wire n_66;
wire n_98;
wire n_60;
wire n_155;
wire n_152;
wire n_43;
wire n_107;
wire n_69;
wire n_58;
wire n_116;
wire n_42;
wire n_45;
wire n_117;
wire n_46;
wire n_94;
wire n_113;
wire n_38;
wire n_123;
wire n_139;
wire n_105;
wire n_80;
wire n_125;
wire n_35;
wire n_128;
wire n_73;
wire n_92;
wire n_149;
wire n_120;
wire n_135;
wire n_30;
wire n_156;
wire n_33;
wire n_126;
wire n_84;
wire n_130;
wire n_157;
wire n_29;
wire n_79;
wire n_131;
wire n_151;
wire n_47;
wire n_53;
wire n_160;
wire n_158;
wire n_44;
wire n_40;
wire n_34;
wire n_100;
wire n_62;
wire n_138;
wire n_148;
wire n_71;
wire n_154;
wire n_109;
wire n_112;
wire n_85;
wire n_159;
wire n_95;
wire n_119;
wire n_59;
wire n_133;
wire n_55;
wire n_99;
wire n_49;
wire n_39;
wire n_54;
wire n_147;
wire n_67;
wire n_121;
wire n_36;
wire n_76;
wire n_87;
wire n_150;
wire n_77;
wire n_64;
wire n_106;
wire n_102;
wire n_161;
wire n_81;
wire n_118;
wire n_28;
wire n_89;
wire n_115;
wire n_70;
wire n_68;
wire n_93;
wire n_72;
wire n_134;
wire n_32;
wire n_41;
wire n_104;
wire n_103;
wire n_141;
wire n_51;
wire n_63;
wire n_97;
wire n_56;
wire n_153;
wire n_145;
wire n_48;
wire n_50;
wire n_52;
wire n_88;
wire n_110;

INVx1_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

CKINVDCx5p33_ASAP7_75t_R g29 ( 
.A(n_21),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

CKINVDCx5p33_ASAP7_75t_R g31 ( 
.A(n_15),
.Y(n_31)
);

CKINVDCx5p33_ASAP7_75t_R g32 ( 
.A(n_1),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_5),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_9),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

CKINVDCx5p33_ASAP7_75t_R g36 ( 
.A(n_14),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_9),
.Y(n_41)
);

INVxp67_ASAP7_75t_SL g42 ( 
.A(n_27),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_8),
.Y(n_43)
);

CKINVDCx5p33_ASAP7_75t_R g44 ( 
.A(n_25),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

INVxp33_ASAP7_75t_SL g46 ( 
.A(n_24),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_3),
.Y(n_47)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_40),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g50 ( 
.A(n_28),
.Y(n_50)
);

NAND2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_0),
.Y(n_51)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_0),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

BUFx6f_ASAP7_75t_SL g55 ( 
.A(n_40),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_40),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_30),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_46),
.B(n_1),
.Y(n_61)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_31),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_39),
.Y(n_65)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_33),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g68 ( 
.A(n_34),
.B(n_45),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_61),
.B(n_32),
.Y(n_69)
);

NAND2x1p5_ASAP7_75t_L g70 ( 
.A(n_59),
.B(n_47),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_68),
.B(n_29),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_49),
.Y(n_72)
);

NAND2x1p5_ASAP7_75t_L g73 ( 
.A(n_53),
.B(n_47),
.Y(n_73)
);

AO22x2_ASAP7_75t_L g74 ( 
.A1(n_60),
.A2(n_45),
.B1(n_43),
.B2(n_37),
.Y(n_74)
);

OA22x2_ASAP7_75t_L g75 ( 
.A1(n_50),
.A2(n_43),
.B1(n_37),
.B2(n_35),
.Y(n_75)
);

AO22x2_ASAP7_75t_L g76 ( 
.A1(n_60),
.A2(n_34),
.B1(n_35),
.B2(n_42),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_51),
.B(n_36),
.Y(n_77)
);

BUFx8_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

NAND2x1p5_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_44),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_52),
.Y(n_80)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_49),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_54),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_2),
.Y(n_83)
);

NAND2x1p5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_64),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_73),
.A2(n_68),
.B1(n_51),
.B2(n_65),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_72),
.B(n_68),
.Y(n_87)
);

AND2x4_ASAP7_75t_L g88 ( 
.A(n_83),
.B(n_68),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_81),
.B(n_68),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_76),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_76),
.Y(n_93)
);

AND3x1_ASAP7_75t_SL g94 ( 
.A(n_75),
.B(n_63),
.C(n_66),
.Y(n_94)
);

O2A1O1Ixp33_ASAP7_75t_L g95 ( 
.A1(n_92),
.A2(n_93),
.B(n_73),
.C(n_77),
.Y(n_95)
);

OA21x2_ASAP7_75t_L g96 ( 
.A1(n_85),
.A2(n_71),
.B(n_58),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_84),
.B(n_48),
.Y(n_97)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_93),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g99 ( 
.A(n_84),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_92),
.B(n_62),
.Y(n_100)
);

NAND2x1p5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_83),
.Y(n_101)
);

O2A1O1Ixp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_69),
.B(n_64),
.C(n_65),
.Y(n_102)
);

A2O1A1Ixp33_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_92),
.B(n_88),
.C(n_90),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_84),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_98),
.B(n_84),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_99),
.B(n_88),
.Y(n_107)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_98),
.B(n_73),
.Y(n_108)
);

NOR2x1_ASAP7_75t_SL g109 ( 
.A(n_100),
.B(n_89),
.Y(n_109)
);

INVx1_ASAP7_75t_SL g110 ( 
.A(n_106),
.Y(n_110)
);

OAI21x1_ASAP7_75t_SL g111 ( 
.A1(n_109),
.A2(n_95),
.B(n_96),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g112 ( 
.A(n_105),
.B(n_76),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_86),
.Y(n_113)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_107),
.Y(n_114)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_114),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_114),
.Y(n_116)
);

AO21x2_ASAP7_75t_L g117 ( 
.A1(n_111),
.A2(n_103),
.B(n_109),
.Y(n_117)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_112),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_111),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_110),
.Y(n_120)
);

NAND2xp33_ASAP7_75t_SL g121 ( 
.A(n_113),
.B(n_108),
.Y(n_121)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx5_ASAP7_75t_SL g124 ( 
.A(n_114),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_116),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g126 ( 
.A(n_120),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_121),
.A2(n_104),
.B(n_107),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_115),
.B(n_105),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_120),
.B(n_106),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_125),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_130),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_123),
.Y(n_133)
);

AND2x2_ASAP7_75t_L g134 ( 
.A(n_129),
.B(n_118),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_127),
.Y(n_135)
);

OR2x2_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_118),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_131),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_122),
.Y(n_138)
);

NOR3xp33_ASAP7_75t_SL g139 ( 
.A(n_135),
.B(n_119),
.C(n_90),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_136),
.B(n_124),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_134),
.B(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_141),
.B(n_132),
.Y(n_142)
);

NAND4xp75_ASAP7_75t_L g143 ( 
.A(n_139),
.B(n_102),
.C(n_58),
.D(n_57),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g144 ( 
.A(n_140),
.B(n_139),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_137),
.B(n_117),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_138),
.B(n_124),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g147 ( 
.A(n_144),
.B(n_124),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_70),
.B(n_102),
.C(n_6),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_146),
.B(n_124),
.Y(n_149)
);

AOI31xp33_ASAP7_75t_SL g150 ( 
.A1(n_145),
.A2(n_2),
.A3(n_5),
.B(n_7),
.Y(n_150)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_143),
.B(n_11),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_SL g152 ( 
.A1(n_147),
.A2(n_12),
.B(n_13),
.Y(n_152)
);

AOI322xp5_ASAP7_75t_L g153 ( 
.A1(n_150),
.A2(n_12),
.A3(n_13),
.B1(n_15),
.B2(n_16),
.C1(n_56),
.C2(n_74),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_149),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_153),
.A2(n_151),
.B1(n_148),
.B2(n_94),
.Y(n_155)
);

XNOR2x2_ASAP7_75t_L g156 ( 
.A(n_152),
.B(n_17),
.Y(n_156)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_154),
.Y(n_157)
);

AND3x4_ASAP7_75t_L g158 ( 
.A(n_156),
.B(n_18),
.C(n_19),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_155),
.A2(n_96),
.B1(n_78),
.B2(n_91),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_157),
.A2(n_78),
.B1(n_91),
.B2(n_101),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_159),
.B(n_23),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_158),
.B1(n_160),
.B2(n_101),
.Y(n_162)
);


endmodule