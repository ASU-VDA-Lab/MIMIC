module fake_jpeg_4648_n_316 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_316);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_316;

wire n_253;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_11),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_4),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx12_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_12),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_19),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_31),
.B(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_30),
.Y(n_32)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_7),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_19),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_34),
.B(n_35),
.Y(n_56)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_36),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

BUFx3_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_41),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_29),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_40),
.A2(n_27),
.B1(n_22),
.B2(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_21),
.B(n_6),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_44),
.Y(n_77)
);

NOR2x1_ASAP7_75t_R g46 ( 
.A(n_33),
.B(n_15),
.Y(n_46)
);

AND2x2_ASAP7_75t_L g81 ( 
.A(n_46),
.B(n_47),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_33),
.B(n_24),
.Y(n_47)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_49),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_24),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_53),
.B(n_54),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_41),
.B(n_23),
.Y(n_54)
);

OR2x2_ASAP7_75t_SL g55 ( 
.A(n_41),
.B(n_14),
.Y(n_55)
);

AOI21xp33_ASAP7_75t_L g78 ( 
.A1(n_55),
.A2(n_64),
.B(n_21),
.Y(n_78)
);

CKINVDCx12_ASAP7_75t_R g57 ( 
.A(n_35),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_34),
.Y(n_58)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_58),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_60),
.Y(n_72)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_40),
.A2(n_27),
.B1(n_16),
.B2(n_22),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_62),
.A2(n_36),
.B1(n_31),
.B2(n_40),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_35),
.B(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_34),
.B(n_23),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_67),
.A2(n_83),
.B1(n_50),
.B2(n_49),
.Y(n_92)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_68),
.B(n_82),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_46),
.A2(n_43),
.B(n_51),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g99 ( 
.A(n_69),
.B(n_54),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_60),
.A2(n_40),
.B1(n_31),
.B2(n_36),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_70),
.A2(n_74),
.B1(n_80),
.B2(n_62),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_52),
.A2(n_40),
.B1(n_31),
.B2(n_36),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_43),
.A2(n_40),
.B1(n_31),
.B2(n_36),
.Y(n_74)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_78),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g80 ( 
.A1(n_47),
.A2(n_31),
.B1(n_36),
.B2(n_18),
.Y(n_80)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_45),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_52),
.A2(n_18),
.B1(n_28),
.B2(n_34),
.Y(n_83)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_85),
.Y(n_94)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_59),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_86),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_50),
.Y(n_88)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_88),
.Y(n_102)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_75),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_77),
.A2(n_51),
.B1(n_52),
.B2(n_48),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_98),
.B1(n_101),
.B2(n_110),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_75),
.B(n_72),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_104),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_92),
.A2(n_95),
.B1(n_99),
.B2(n_106),
.Y(n_123)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_69),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g138 ( 
.A(n_96),
.B(n_101),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_77),
.A2(n_72),
.B1(n_71),
.B2(n_81),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_56),
.B1(n_61),
.B2(n_50),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_100),
.A2(n_95),
.B1(n_111),
.B2(n_107),
.Y(n_129)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_81),
.Y(n_101)
);

NAND2xp33_ASAP7_75t_SL g103 ( 
.A(n_79),
.B(n_0),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_L g121 ( 
.A1(n_103),
.A2(n_20),
.B(n_55),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_79),
.B(n_64),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_84),
.A2(n_42),
.B1(n_38),
.B2(n_20),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g107 ( 
.A(n_65),
.B(n_53),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_107),
.B(n_112),
.Y(n_130)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_109),
.B(n_76),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_65),
.B(n_56),
.C(n_38),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_111),
.B(n_73),
.C(n_87),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_66),
.B(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_113),
.B(n_119),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g115 ( 
.A1(n_93),
.A2(n_73),
.B(n_87),
.Y(n_115)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_115),
.A2(n_131),
.B(n_136),
.Y(n_163)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_102),
.Y(n_116)
);

CKINVDCx14_ASAP7_75t_R g159 ( 
.A(n_116),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_117),
.A2(n_128),
.B1(n_135),
.B2(n_118),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_118),
.B(n_120),
.C(n_105),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_89),
.B(n_108),
.C(n_98),
.Y(n_120)
);

AOI21xp5_ASAP7_75t_SL g161 ( 
.A1(n_121),
.A2(n_122),
.B(n_15),
.Y(n_161)
);

NOR2x1p5_ASAP7_75t_L g122 ( 
.A(n_100),
.B(n_39),
.Y(n_122)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_109),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_124),
.B(n_125),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_SL g125 ( 
.A(n_108),
.B(n_91),
.Y(n_125)
);

INVx3_ASAP7_75t_L g126 ( 
.A(n_97),
.Y(n_126)
);

INVx6_ASAP7_75t_L g158 ( 
.A(n_126),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_96),
.A2(n_84),
.B1(n_86),
.B2(n_85),
.Y(n_128)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_129),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_104),
.A2(n_57),
.B(n_66),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_97),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_132),
.B(n_133),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_99),
.B(n_66),
.Y(n_133)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_94),
.Y(n_134)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_134),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_90),
.A2(n_82),
.B1(n_68),
.B2(n_37),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_94),
.A2(n_88),
.B1(n_13),
.B2(n_14),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_112),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_137),
.B(n_25),
.Y(n_148)
);

OAI21xp33_ASAP7_75t_L g140 ( 
.A1(n_138),
.A2(n_103),
.B(n_58),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_140),
.B(n_115),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g141 ( 
.A(n_122),
.B(n_105),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_141),
.A2(n_152),
.B(n_161),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_143),
.B(n_157),
.C(n_121),
.Y(n_174)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_128),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_146),
.B(n_147),
.Y(n_188)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_116),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_151),
.Y(n_170)
);

OA22x2_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_39),
.B1(n_37),
.B2(n_32),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_158),
.B1(n_159),
.B2(n_147),
.Y(n_172)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_114),
.B(n_25),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_129),
.B(n_39),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_114),
.B(n_25),
.Y(n_153)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_153),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_130),
.B(n_25),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_154),
.B(n_155),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_135),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_133),
.B(n_39),
.C(n_37),
.Y(n_157)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_130),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g171 ( 
.A(n_160),
.B(n_162),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_SL g162 ( 
.A(n_127),
.B(n_58),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_164),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_120),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_165),
.B(n_166),
.C(n_174),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_131),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_168),
.B(n_152),
.Y(n_215)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_172),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_155),
.A2(n_117),
.B1(n_137),
.B2(n_132),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_173),
.B(n_177),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g175 ( 
.A(n_162),
.Y(n_175)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_145),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_183),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_144),
.B(n_134),
.C(n_126),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_180),
.B(n_181),
.C(n_190),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_124),
.Y(n_181)
);

NOR2xp67_ASAP7_75t_SL g182 ( 
.A(n_163),
.B(n_25),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_182),
.A2(n_149),
.B(n_158),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_144),
.A2(n_39),
.B1(n_37),
.B2(n_32),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_148),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_185),
.B(n_187),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_156),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_156),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_191),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_157),
.B(n_119),
.C(n_37),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_151),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_176),
.A2(n_163),
.B(n_161),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_147),
.B1(n_26),
.B2(n_17),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_171),
.B(n_160),
.Y(n_195)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_195),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_181),
.B(n_154),
.Y(n_202)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_202),
.Y(n_225)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_170),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_205),
.B(n_207),
.Y(n_227)
);

OA21x2_ASAP7_75t_L g206 ( 
.A1(n_182),
.A2(n_149),
.B(n_146),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_209),
.Y(n_234)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_188),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_186),
.B(n_152),
.Y(n_208)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_208),
.Y(n_229)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_172),
.Y(n_209)
);

INVx13_ASAP7_75t_L g210 ( 
.A(n_167),
.Y(n_210)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_210),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_211),
.A2(n_17),
.B1(n_32),
.B2(n_2),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g233 ( 
.A(n_212),
.Y(n_233)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_164),
.C(n_150),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_213),
.B(n_190),
.C(n_168),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_186),
.B(n_175),
.Y(n_214)
);

CKINVDCx14_ASAP7_75t_R g222 ( 
.A(n_214),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g219 ( 
.A(n_215),
.B(n_166),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_169),
.B(n_141),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_216),
.B(n_176),
.Y(n_217)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_217),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g218 ( 
.A1(n_197),
.A2(n_178),
.B1(n_141),
.B2(n_180),
.Y(n_218)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_218),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g242 ( 
.A(n_219),
.B(n_220),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_192),
.B(n_174),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_197),
.A2(n_178),
.B1(n_183),
.B2(n_184),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_221),
.A2(n_209),
.B1(n_203),
.B2(n_211),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_226),
.B(n_235),
.C(n_198),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_228),
.B(n_208),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_26),
.Y(n_230)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_231),
.Y(n_248)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_26),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_215),
.B(n_26),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_232),
.B(n_196),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_32),
.C(n_17),
.Y(n_235)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_236),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_227),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_239),
.B(n_250),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_240),
.B(n_249),
.C(n_256),
.Y(n_260)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g263 ( 
.A(n_244),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_234),
.A2(n_203),
.B1(n_210),
.B2(n_212),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_245),
.A2(n_201),
.B1(n_229),
.B2(n_204),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_224),
.B(n_195),
.Y(n_247)
);

OAI21xp33_ASAP7_75t_L g259 ( 
.A1(n_247),
.A2(n_214),
.B(n_216),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_225),
.B(n_193),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_221),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_233),
.B(n_207),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_251),
.B(n_252),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_223),
.B(n_199),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_253),
.B(n_219),
.Y(n_265)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_217),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_255),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_222),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_202),
.C(n_205),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_231),
.Y(n_258)
);

XNOR2xp5_ASAP7_75t_L g274 ( 
.A(n_258),
.B(n_272),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_259),
.A2(n_261),
.B(n_269),
.Y(n_277)
);

OAI21x1_ASAP7_75t_L g261 ( 
.A1(n_243),
.A2(n_235),
.B(n_237),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_247),
.Y(n_262)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_265),
.B(n_268),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_266),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_242),
.B(n_220),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g269 ( 
.A(n_245),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_242),
.B(n_248),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g279 ( 
.A(n_270),
.B(n_248),
.C(n_230),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_240),
.B(n_232),
.Y(n_272)
);

NOR2x1_ASAP7_75t_L g275 ( 
.A(n_259),
.B(n_201),
.Y(n_275)
);

OA21x2_ASAP7_75t_L g291 ( 
.A1(n_275),
.A2(n_8),
.B(n_13),
.Y(n_291)
);

MAJx2_ASAP7_75t_L g276 ( 
.A(n_267),
.B(n_194),
.C(n_238),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_278),
.B(n_5),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_SL g278 ( 
.A1(n_269),
.A2(n_241),
.B(n_256),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_279),
.B(n_283),
.C(n_286),
.Y(n_295)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_264),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_281),
.B(n_0),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_271),
.B(n_204),
.Y(n_282)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_282),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_268),
.B(n_244),
.C(n_200),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_260),
.B(n_257),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_285),
.B(n_263),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_270),
.B(n_246),
.C(n_206),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_287),
.B(n_289),
.Y(n_301)
);

AOI21x1_ASAP7_75t_L g288 ( 
.A1(n_275),
.A2(n_262),
.B(n_206),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g304 ( 
.A1(n_288),
.A2(n_284),
.B(n_279),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_6),
.Y(n_290)
);

AOI21xp33_ASAP7_75t_L g303 ( 
.A1(n_290),
.A2(n_292),
.B(n_1),
.Y(n_303)
);

FAx1_ASAP7_75t_SL g300 ( 
.A(n_291),
.B(n_296),
.CI(n_0),
.CON(n_300),
.SN(n_300)
);

NOR2xp33_ASAP7_75t_SL g292 ( 
.A(n_277),
.B(n_8),
.Y(n_292)
);

AOI322xp5_ASAP7_75t_L g293 ( 
.A1(n_273),
.A2(n_14),
.A3(n_5),
.B1(n_9),
.B2(n_13),
.C1(n_4),
.C2(n_11),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_293),
.A2(n_297),
.B1(n_276),
.B2(n_10),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_286),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_295),
.B(n_283),
.C(n_284),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g306 ( 
.A(n_298),
.B(n_305),
.C(n_3),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_299),
.B(n_300),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_294),
.B(n_274),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_302),
.A2(n_304),
.B(n_1),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_3),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g305 ( 
.A(n_295),
.B(n_291),
.C(n_293),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_306),
.B(n_307),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g307 ( 
.A(n_298),
.Y(n_307)
);

OAI211xp5_ASAP7_75t_L g313 ( 
.A1(n_309),
.A2(n_310),
.B(n_311),
.C(n_300),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_305),
.A2(n_1),
.B(n_2),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_313),
.A2(n_308),
.B1(n_301),
.B2(n_3),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_314),
.B(n_312),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_315),
.B(n_3),
.Y(n_316)
);


endmodule