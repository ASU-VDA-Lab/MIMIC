module fake_jpeg_13762_n_185 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_185);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_185;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_3),
.Y(n_13)
);

INVxp67_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

INVx8_ASAP7_75t_SL g16 ( 
.A(n_12),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_0),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_5),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_9),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_5),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_15),
.B(n_11),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_33),
.B(n_52),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_22),
.Y(n_34)
);

INVx6_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_35),
.Y(n_72)
);

BUFx2_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_37),
.Y(n_73)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_41),
.Y(n_80)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

AOI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_14),
.A2(n_1),
.B(n_2),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_17),
.C(n_27),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_21),
.Y(n_46)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_46),
.Y(n_77)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_21),
.Y(n_47)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_47),
.Y(n_75)
);

INVx13_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_48),
.Y(n_82)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_49),
.B(n_50),
.Y(n_71)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_32),
.Y(n_50)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_32),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_51),
.B(n_20),
.Y(n_85)
);

INVx11_ASAP7_75t_L g52 ( 
.A(n_32),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_53),
.B(n_54),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_15),
.B(n_11),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_30),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g105 ( 
.A(n_57),
.B(n_85),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_36),
.A2(n_29),
.B1(n_30),
.B2(n_18),
.Y(n_58)
);

AO21x1_ASAP7_75t_L g96 ( 
.A1(n_58),
.A2(n_69),
.B(n_83),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_26),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_65),
.B(n_66),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_17),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_13),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_68),
.B(n_76),
.Y(n_94)
);

A2O1A1Ixp33_ASAP7_75t_L g69 ( 
.A1(n_48),
.A2(n_29),
.B(n_13),
.C(n_18),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_70),
.A2(n_81),
.B1(n_19),
.B2(n_52),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_51),
.B(n_25),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_37),
.B(n_23),
.Y(n_78)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_78),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_40),
.A2(n_34),
.B1(n_43),
.B2(n_45),
.Y(n_81)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_38),
.A2(n_23),
.B1(n_20),
.B2(n_19),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_77),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_87),
.B(n_102),
.Y(n_110)
);

INVx1_ASAP7_75t_SL g88 ( 
.A(n_71),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_88),
.B(n_97),
.Y(n_114)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_82),
.Y(n_91)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_91),
.Y(n_113)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_61),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_93),
.A2(n_74),
.B1(n_79),
.B2(n_56),
.Y(n_119)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_95),
.Y(n_125)
);

INVx1_ASAP7_75t_SL g97 ( 
.A(n_71),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_70),
.A2(n_50),
.B1(n_3),
.B2(n_4),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_98),
.A2(n_79),
.B1(n_64),
.B2(n_74),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_81),
.A2(n_1),
.B1(n_5),
.B2(n_7),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g118 ( 
.A(n_99),
.B(n_84),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_57),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_62),
.Y(n_117)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_84),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_104),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_71),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_75),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_106),
.B(n_107),
.Y(n_123)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_64),
.Y(n_107)
);

AOI21xp5_ASAP7_75t_L g108 ( 
.A1(n_75),
.A2(n_7),
.B(n_8),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g128 ( 
.A1(n_108),
.A2(n_7),
.B(n_8),
.Y(n_128)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_67),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_109),
.B(n_72),
.Y(n_126)
);

NAND2x1_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_56),
.Y(n_112)
);

AOI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_112),
.A2(n_128),
.B(n_108),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_94),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_115),
.B(n_117),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_118),
.A2(n_96),
.B1(n_97),
.B2(n_88),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_119),
.A2(n_122),
.B1(n_90),
.B2(n_102),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_SL g120 ( 
.A(n_100),
.B(n_59),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g142 ( 
.A(n_120),
.B(n_126),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_121),
.B(n_127),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_89),
.B(n_72),
.Y(n_127)
);

OAI21xp5_ASAP7_75t_SL g153 ( 
.A1(n_129),
.A2(n_138),
.B(n_144),
.Y(n_153)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_124),
.Y(n_130)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_130),
.Y(n_155)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_124),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_133),
.Y(n_149)
);

AOI221xp5_ASAP7_75t_L g147 ( 
.A1(n_132),
.A2(n_115),
.B1(n_118),
.B2(n_128),
.C(n_120),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_123),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_111),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_134),
.B(n_137),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_96),
.B1(n_93),
.B2(n_86),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_136),
.A2(n_141),
.B1(n_133),
.B2(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_125),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_110),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_140),
.A2(n_143),
.B1(n_116),
.B2(n_125),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_112),
.A2(n_86),
.B1(n_105),
.B2(n_107),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g143 ( 
.A1(n_122),
.A2(n_105),
.B1(n_95),
.B2(n_92),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_110),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g162 ( 
.A1(n_145),
.A2(n_148),
.B1(n_113),
.B2(n_73),
.Y(n_162)
);

AO22x1_ASAP7_75t_L g146 ( 
.A1(n_129),
.A2(n_112),
.B1(n_116),
.B2(n_114),
.Y(n_146)
);

A2O1A1Ixp33_ASAP7_75t_SL g163 ( 
.A1(n_146),
.A2(n_91),
.B(n_73),
.C(n_111),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g164 ( 
.A(n_147),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_135),
.A2(n_118),
.B1(n_114),
.B2(n_105),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_114),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_151),
.C(n_137),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_144),
.B(n_113),
.C(n_121),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_152),
.A2(n_140),
.B1(n_139),
.B2(n_142),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_157),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_150),
.B(n_153),
.C(n_152),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_158),
.B(n_163),
.C(n_146),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_153),
.A2(n_131),
.B(n_130),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_161),
.C(n_146),
.Y(n_169)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_155),
.Y(n_160)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_160),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_149),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_162),
.A2(n_151),
.B1(n_155),
.B2(n_154),
.Y(n_166)
);

AOI21x1_ASAP7_75t_SL g174 ( 
.A1(n_166),
.A2(n_160),
.B(n_163),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_167),
.A2(n_169),
.B(n_159),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_157),
.B(n_111),
.C(n_10),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_170),
.B(n_156),
.C(n_158),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_171),
.B(n_172),
.C(n_163),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g173 ( 
.A1(n_167),
.A2(n_162),
.B(n_163),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_SL g178 ( 
.A1(n_173),
.A2(n_175),
.B(n_165),
.Y(n_178)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_174),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_168),
.B(n_164),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_178),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_176),
.B(n_164),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_179),
.B(n_9),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_181),
.B(n_182),
.C(n_180),
.Y(n_183)
);

AND2x2_ASAP7_75t_L g182 ( 
.A(n_180),
.B(n_10),
.Y(n_182)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_183),
.A2(n_60),
.B(n_179),
.Y(n_184)
);

BUFx24_ASAP7_75t_SL g185 ( 
.A(n_184),
.Y(n_185)
);


endmodule