module real_aes_1897_n_104 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_104);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_104;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_666;
wire n_320;
wire n_551;
wire n_537;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_815;
wire n_519;
wire n_638;
wire n_564;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_732;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_755;
wire n_284;
wire n_153;
wire n_532;
wire n_316;
wire n_656;
wire n_746;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_142;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_255;
wire n_226;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_569;
wire n_303;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_831;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_804;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_SL g535 ( .A(n_0), .B(n_512), .Y(n_535) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_1), .A2(n_515), .B(n_580), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_2), .B(n_830), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g518 ( .A(n_3), .B(n_222), .Y(n_518) );
INVx1_ASAP7_75t_L g154 ( .A(n_4), .Y(n_154) );
XNOR2xp5_ASAP7_75t_L g123 ( .A(n_5), .B(n_124), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g210 ( .A(n_6), .B(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g588 ( .A(n_7), .B(n_222), .Y(n_588) );
INVx1_ASAP7_75t_L g186 ( .A(n_8), .Y(n_186) );
CKINVDCx16_ASAP7_75t_R g830 ( .A(n_9), .Y(n_830) );
XNOR2xp5_ASAP7_75t_L g124 ( .A(n_10), .B(n_125), .Y(n_124) );
CKINVDCx5p33_ASAP7_75t_R g201 ( .A(n_11), .Y(n_201) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_12), .B(n_219), .Y(n_573) );
INVx2_ASAP7_75t_L g146 ( .A(n_13), .Y(n_146) );
AOI221x1_ASAP7_75t_L g522 ( .A1(n_14), .A2(n_27), .B1(n_512), .B2(n_515), .C(n_523), .Y(n_522) );
CKINVDCx16_ASAP7_75t_R g115 ( .A(n_15), .Y(n_115) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_16), .B(n_512), .Y(n_569) );
INVx1_ASAP7_75t_L g220 ( .A(n_17), .Y(n_220) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_18), .A2(n_183), .B(n_568), .Y(n_567) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_19), .B(n_177), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_20), .B(n_222), .Y(n_562) );
AO21x1_ASAP7_75t_L g511 ( .A1(n_21), .A2(n_512), .B(n_513), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g832 ( .A(n_22), .Y(n_832) );
INVx1_ASAP7_75t_L g119 ( .A(n_23), .Y(n_119) );
NOR2xp33_ASAP7_75t_SL g827 ( .A(n_23), .B(n_120), .Y(n_827) );
INVx1_ASAP7_75t_L g217 ( .A(n_24), .Y(n_217) );
INVx1_ASAP7_75t_SL g271 ( .A(n_25), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_26), .B(n_169), .Y(n_233) );
AOI33xp33_ASAP7_75t_L g257 ( .A1(n_28), .A2(n_56), .A3(n_151), .B1(n_162), .B2(n_258), .B3(n_259), .Y(n_257) );
NAND2x1_ASAP7_75t_L g533 ( .A(n_29), .B(n_222), .Y(n_533) );
AOI22xp5_ASAP7_75t_SL g815 ( .A1(n_30), .A2(n_816), .B1(n_819), .B2(n_820), .Y(n_815) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_30), .Y(n_820) );
NAND2x1_ASAP7_75t_L g587 ( .A(n_31), .B(n_219), .Y(n_587) );
INVx1_ASAP7_75t_L g194 ( .A(n_32), .Y(n_194) );
OA21x2_ASAP7_75t_L g145 ( .A1(n_33), .A2(n_89), .B(n_146), .Y(n_145) );
OR2x2_ASAP7_75t_L g179 ( .A(n_33), .B(n_89), .Y(n_179) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_34), .B(n_149), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g582 ( .A(n_35), .B(n_219), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_36), .B(n_222), .Y(n_572) );
AOI22xp5_ASAP7_75t_L g816 ( .A1(n_37), .A2(n_67), .B1(n_817), .B2(n_818), .Y(n_816) );
CKINVDCx20_ASAP7_75t_R g818 ( .A(n_37), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_38), .B(n_219), .Y(n_517) );
AOI21xp5_ASAP7_75t_L g541 ( .A1(n_39), .A2(n_515), .B(n_542), .Y(n_541) );
AND2x2_ASAP7_75t_L g156 ( .A(n_40), .B(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g161 ( .A(n_40), .Y(n_161) );
AND2x2_ASAP7_75t_L g175 ( .A(n_40), .B(n_154), .Y(n_175) );
OR2x6_ASAP7_75t_L g117 ( .A(n_41), .B(n_118), .Y(n_117) );
NOR3xp33_ASAP7_75t_L g828 ( .A(n_41), .B(n_115), .C(n_829), .Y(n_828) );
CKINVDCx20_ASAP7_75t_R g197 ( .A(n_42), .Y(n_197) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_43), .B(n_512), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g148 ( .A(n_44), .B(n_149), .Y(n_148) );
AOI22xp5_ASAP7_75t_L g226 ( .A1(n_45), .A2(n_144), .B1(n_211), .B2(n_227), .Y(n_226) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_46), .B(n_235), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g272 ( .A(n_47), .B(n_169), .Y(n_272) );
AOI22xp5_ASAP7_75t_L g125 ( .A1(n_48), .A2(n_98), .B1(n_126), .B2(n_127), .Y(n_125) );
CKINVDCx20_ASAP7_75t_R g127 ( .A(n_48), .Y(n_127) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_49), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_50), .B(n_219), .Y(n_543) );
NAND2xp5_ASAP7_75t_SL g188 ( .A(n_51), .B(n_183), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g187 ( .A(n_52), .B(n_169), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g585 ( .A1(n_53), .A2(n_515), .B(n_586), .Y(n_585) );
CKINVDCx5p33_ASAP7_75t_R g230 ( .A(n_54), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g534 ( .A(n_55), .B(n_219), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_57), .B(n_169), .Y(n_168) );
INVx1_ASAP7_75t_L g152 ( .A(n_58), .Y(n_152) );
INVx1_ASAP7_75t_L g171 ( .A(n_58), .Y(n_171) );
AND2x2_ASAP7_75t_L g176 ( .A(n_59), .B(n_177), .Y(n_176) );
AOI221xp5_ASAP7_75t_L g184 ( .A1(n_60), .A2(n_78), .B1(n_149), .B2(n_159), .C(n_185), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_61), .B(n_149), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g111 ( .A(n_62), .B(n_112), .Y(n_111) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_63), .B(n_222), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_64), .B(n_144), .Y(n_203) );
AOI21xp5_ASAP7_75t_SL g241 ( .A1(n_65), .A2(n_159), .B(n_242), .Y(n_241) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_66), .A2(n_515), .B(n_532), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_67), .Y(n_817) );
INVx1_ASAP7_75t_L g214 ( .A(n_68), .Y(n_214) );
AO21x1_ASAP7_75t_L g514 ( .A1(n_69), .A2(n_515), .B(n_516), .Y(n_514) );
NAND2xp5_ASAP7_75t_SL g578 ( .A(n_70), .B(n_512), .Y(n_578) );
INVx1_ASAP7_75t_L g166 ( .A(n_71), .Y(n_166) );
NAND2xp5_ASAP7_75t_SL g589 ( .A(n_72), .B(n_512), .Y(n_589) );
AOI21xp5_ASAP7_75t_L g158 ( .A1(n_73), .A2(n_159), .B(n_165), .Y(n_158) );
AND2x2_ASAP7_75t_L g546 ( .A(n_74), .B(n_178), .Y(n_546) );
INVx1_ASAP7_75t_L g157 ( .A(n_75), .Y(n_157) );
INVx1_ASAP7_75t_L g173 ( .A(n_75), .Y(n_173) );
AND2x2_ASAP7_75t_L g590 ( .A(n_76), .B(n_143), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_77), .B(n_149), .Y(n_260) );
AND2x2_ASAP7_75t_L g273 ( .A(n_79), .B(n_143), .Y(n_273) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_79), .Y(n_821) );
INVx1_ASAP7_75t_L g215 ( .A(n_80), .Y(n_215) );
AOI21xp5_ASAP7_75t_L g269 ( .A1(n_81), .A2(n_159), .B(n_270), .Y(n_269) );
A2O1A1Ixp33_ASAP7_75t_L g231 ( .A1(n_82), .A2(n_159), .B(n_232), .C(n_236), .Y(n_231) );
INVx1_ASAP7_75t_L g120 ( .A(n_83), .Y(n_120) );
NAND2xp5_ASAP7_75t_SL g564 ( .A(n_84), .B(n_512), .Y(n_564) );
AND2x2_ASAP7_75t_SL g239 ( .A(n_85), .B(n_143), .Y(n_239) );
AND2x2_ASAP7_75t_L g576 ( .A(n_86), .B(n_143), .Y(n_576) );
AOI22xp5_ASAP7_75t_L g254 ( .A1(n_87), .A2(n_159), .B1(n_255), .B2(n_256), .Y(n_254) );
AND2x2_ASAP7_75t_L g513 ( .A(n_88), .B(n_211), .Y(n_513) );
AND2x2_ASAP7_75t_L g536 ( .A(n_90), .B(n_143), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_91), .B(n_219), .Y(n_563) );
INVx1_ASAP7_75t_L g243 ( .A(n_92), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g803 ( .A(n_93), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_94), .B(n_222), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_95), .B(n_219), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_96), .A2(n_515), .B(n_561), .Y(n_560) );
AND2x2_ASAP7_75t_L g261 ( .A(n_97), .B(n_143), .Y(n_261) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_98), .Y(n_126) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_99), .B(n_222), .Y(n_581) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_100), .A2(n_192), .B(n_193), .C(n_196), .Y(n_191) );
BUFx2_ASAP7_75t_L g110 ( .A(n_101), .Y(n_110) );
AOI21xp5_ASAP7_75t_L g570 ( .A1(n_102), .A2(n_515), .B(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_103), .B(n_169), .Y(n_244) );
AOI21xp5_ASAP7_75t_SL g104 ( .A1(n_105), .A2(n_824), .B(n_831), .Y(n_104) );
OA22x2_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_121), .B1(n_806), .B2(n_808), .Y(n_105) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_107), .B(n_111), .Y(n_106) );
CKINVDCx11_ASAP7_75t_R g107 ( .A(n_108), .Y(n_107) );
CKINVDCx20_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
HB1xp67_ASAP7_75t_L g109 ( .A(n_110), .Y(n_109) );
CKINVDCx20_ASAP7_75t_R g807 ( .A(n_110), .Y(n_807) );
CKINVDCx20_ASAP7_75t_R g822 ( .A(n_111), .Y(n_822) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
BUFx3_ASAP7_75t_L g813 ( .A(n_114), .Y(n_813) );
NAND2xp5_ASAP7_75t_L g114 ( .A(n_115), .B(n_116), .Y(n_114) );
CKINVDCx16_ASAP7_75t_R g130 ( .A(n_115), .Y(n_130) );
OR2x2_ASAP7_75t_L g805 ( .A(n_115), .B(n_117), .Y(n_805) );
OAI22xp5_ASAP7_75t_SL g121 ( .A1(n_116), .A2(n_122), .B1(n_803), .B2(n_804), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g116 ( .A(n_117), .Y(n_116) );
NAND2xp5_ASAP7_75t_L g118 ( .A(n_119), .B(n_120), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g122 ( .A(n_123), .B(n_128), .Y(n_122) );
OAI22xp5_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_130), .B1(n_131), .B2(n_503), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_130), .Y(n_129) );
INVx2_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
NAND4xp75_ASAP7_75t_L g132 ( .A(n_133), .B(n_375), .C(n_420), .D(n_489), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
NAND2x1_ASAP7_75t_L g134 ( .A(n_135), .B(n_335), .Y(n_134) );
NOR3xp33_ASAP7_75t_L g135 ( .A(n_136), .B(n_291), .C(n_316), .Y(n_135) );
OAI222xp33_ASAP7_75t_L g136 ( .A1(n_137), .A2(n_205), .B1(n_246), .B2(n_262), .C1(n_278), .C2(n_285), .Y(n_136) );
INVxp67_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_139), .B(n_180), .Y(n_138) );
AND2x2_ASAP7_75t_L g500 ( .A(n_139), .B(n_314), .Y(n_500) );
INVx1_ASAP7_75t_L g139 ( .A(n_140), .Y(n_139) );
HB1xp67_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g251 ( .A(n_141), .B(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_141), .B(n_189), .Y(n_290) );
INVx3_ASAP7_75t_L g305 ( .A(n_141), .Y(n_305) );
AND2x2_ASAP7_75t_L g438 ( .A(n_141), .B(n_439), .Y(n_438) );
AO21x2_ASAP7_75t_L g141 ( .A1(n_142), .A2(n_147), .B(n_176), .Y(n_141) );
OAI22xp5_ASAP7_75t_L g190 ( .A1(n_142), .A2(n_143), .B1(n_191), .B2(n_197), .Y(n_190) );
AO21x2_ASAP7_75t_L g323 ( .A1(n_142), .A2(n_147), .B(n_176), .Y(n_323) );
AO21x2_ASAP7_75t_L g529 ( .A1(n_142), .A2(n_530), .B(n_536), .Y(n_529) );
AO21x2_ASAP7_75t_L g539 ( .A1(n_142), .A2(n_540), .B(n_546), .Y(n_539) );
AO21x2_ASAP7_75t_L g551 ( .A1(n_142), .A2(n_530), .B(n_536), .Y(n_551) );
AO21x2_ASAP7_75t_L g553 ( .A1(n_142), .A2(n_540), .B(n_546), .Y(n_553) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx4_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_144), .B(n_200), .Y(n_199) );
INVx3_ASAP7_75t_L g144 ( .A(n_145), .Y(n_144) );
BUFx4f_ASAP7_75t_L g183 ( .A(n_145), .Y(n_183) );
AND2x2_ASAP7_75t_SL g178 ( .A(n_146), .B(n_179), .Y(n_178) );
AND2x4_ASAP7_75t_L g211 ( .A(n_146), .B(n_179), .Y(n_211) );
NAND2xp5_ASAP7_75t_L g147 ( .A(n_148), .B(n_158), .Y(n_147) );
INVx1_ASAP7_75t_L g204 ( .A(n_149), .Y(n_204) );
AND2x4_ASAP7_75t_L g149 ( .A(n_150), .B(n_155), .Y(n_149) );
INVx1_ASAP7_75t_L g228 ( .A(n_150), .Y(n_228) );
AND2x2_ASAP7_75t_L g150 ( .A(n_151), .B(n_153), .Y(n_150) );
OR2x6_ASAP7_75t_L g167 ( .A(n_151), .B(n_163), .Y(n_167) );
INVxp33_ASAP7_75t_L g258 ( .A(n_151), .Y(n_258) );
INVx2_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AND2x2_ASAP7_75t_L g164 ( .A(n_152), .B(n_154), .Y(n_164) );
AND2x4_ASAP7_75t_L g222 ( .A(n_152), .B(n_172), .Y(n_222) );
HB1xp67_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx1_ASAP7_75t_L g229 ( .A(n_155), .Y(n_229) );
BUFx3_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
AND2x6_ASAP7_75t_L g515 ( .A(n_156), .B(n_164), .Y(n_515) );
INVx2_ASAP7_75t_L g163 ( .A(n_157), .Y(n_163) );
AND2x6_ASAP7_75t_L g219 ( .A(n_157), .B(n_170), .Y(n_219) );
INVxp67_ASAP7_75t_L g202 ( .A(n_159), .Y(n_202) );
AND2x4_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
NOR2x1p5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
INVx1_ASAP7_75t_L g259 ( .A(n_162), .Y(n_259) );
INVx3_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
O2A1O1Ixp33_ASAP7_75t_L g165 ( .A1(n_166), .A2(n_167), .B(n_168), .C(n_174), .Y(n_165) );
O2A1O1Ixp33_ASAP7_75t_SL g185 ( .A1(n_167), .A2(n_174), .B(n_186), .C(n_187), .Y(n_185) );
INVxp67_ASAP7_75t_L g192 ( .A(n_167), .Y(n_192) );
OAI22xp5_ASAP7_75t_L g213 ( .A1(n_167), .A2(n_195), .B1(n_214), .B2(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g235 ( .A(n_167), .Y(n_235) );
O2A1O1Ixp33_ASAP7_75t_L g242 ( .A1(n_167), .A2(n_174), .B(n_243), .C(n_244), .Y(n_242) );
O2A1O1Ixp33_ASAP7_75t_SL g270 ( .A1(n_167), .A2(n_174), .B(n_271), .C(n_272), .Y(n_270) );
INVx1_ASAP7_75t_L g195 ( .A(n_169), .Y(n_195) );
AND2x4_ASAP7_75t_L g512 ( .A(n_169), .B(n_175), .Y(n_512) );
AND2x4_ASAP7_75t_L g169 ( .A(n_170), .B(n_172), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_171), .Y(n_170) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_174), .B(n_211), .Y(n_223) );
AOI21xp5_ASAP7_75t_L g232 ( .A1(n_174), .A2(n_233), .B(n_234), .Y(n_232) );
INVx1_ASAP7_75t_L g255 ( .A(n_174), .Y(n_255) );
AOI21xp5_ASAP7_75t_L g516 ( .A1(n_174), .A2(n_517), .B(n_518), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_174), .A2(n_524), .B(n_525), .Y(n_523) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_174), .A2(n_533), .B(n_534), .Y(n_532) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_174), .A2(n_543), .B(n_544), .Y(n_542) );
AOI21xp5_ASAP7_75t_L g561 ( .A1(n_174), .A2(n_562), .B(n_563), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_174), .A2(n_572), .B(n_573), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g580 ( .A1(n_174), .A2(n_581), .B(n_582), .Y(n_580) );
AOI21xp5_ASAP7_75t_L g586 ( .A1(n_174), .A2(n_587), .B(n_588), .Y(n_586) );
INVx5_ASAP7_75t_L g174 ( .A(n_175), .Y(n_174) );
HB1xp67_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
CKINVDCx5p33_ASAP7_75t_R g266 ( .A(n_177), .Y(n_266) );
OA21x2_ASAP7_75t_L g521 ( .A1(n_177), .A2(n_522), .B(n_526), .Y(n_521) );
OA21x2_ASAP7_75t_L g549 ( .A1(n_177), .A2(n_522), .B(n_526), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_177), .A2(n_578), .B(n_579), .Y(n_577) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
AND2x2_ASAP7_75t_L g368 ( .A(n_180), .B(n_321), .Y(n_368) );
AND2x2_ASAP7_75t_L g370 ( .A(n_180), .B(n_371), .Y(n_370) );
INVx3_ASAP7_75t_L g405 ( .A(n_180), .Y(n_405) );
AND2x4_ASAP7_75t_L g180 ( .A(n_181), .B(n_189), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
INVxp67_ASAP7_75t_L g288 ( .A(n_182), .Y(n_288) );
INVx1_ASAP7_75t_L g307 ( .A(n_182), .Y(n_307) );
AND2x4_ASAP7_75t_L g314 ( .A(n_182), .B(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_182), .B(n_252), .Y(n_330) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_182), .Y(n_439) );
INVx1_ASAP7_75t_L g449 ( .A(n_182), .Y(n_449) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_183), .A2(n_184), .B(n_188), .Y(n_182) );
INVx2_ASAP7_75t_SL g236 ( .A(n_183), .Y(n_236) );
INVx1_ASAP7_75t_L g249 ( .A(n_189), .Y(n_249) );
INVx2_ASAP7_75t_L g302 ( .A(n_189), .Y(n_302) );
INVx1_ASAP7_75t_L g383 ( .A(n_189), .Y(n_383) );
OR2x2_ASAP7_75t_L g189 ( .A(n_190), .B(n_198), .Y(n_189) );
NOR2xp33_ASAP7_75t_L g193 ( .A(n_194), .B(n_195), .Y(n_193) );
OAI22xp5_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_202), .B1(n_203), .B2(n_204), .Y(n_198) );
INVx1_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx1_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
AND2x2_ASAP7_75t_SL g206 ( .A(n_207), .B(n_237), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_207), .B(n_264), .Y(n_358) );
INVx2_ASAP7_75t_L g379 ( .A(n_207), .Y(n_379) );
AND2x2_ASAP7_75t_L g387 ( .A(n_207), .B(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g207 ( .A(n_208), .B(n_224), .Y(n_207) );
AND2x4_ASAP7_75t_L g277 ( .A(n_208), .B(n_225), .Y(n_277) );
INVx1_ASAP7_75t_L g284 ( .A(n_208), .Y(n_284) );
AND2x2_ASAP7_75t_L g460 ( .A(n_208), .B(n_265), .Y(n_460) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g298 ( .A(n_209), .B(n_225), .Y(n_298) );
INVx2_ASAP7_75t_L g334 ( .A(n_209), .Y(n_334) );
AND2x2_ASAP7_75t_L g413 ( .A(n_209), .B(n_265), .Y(n_413) );
NOR2x1_ASAP7_75t_SL g456 ( .A(n_209), .B(n_238), .Y(n_456) );
AND2x4_ASAP7_75t_L g209 ( .A(n_210), .B(n_212), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g240 ( .A1(n_211), .A2(n_241), .B(n_245), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g519 ( .A(n_211), .B(n_520), .Y(n_519) );
INVx1_ASAP7_75t_SL g558 ( .A(n_211), .Y(n_558) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_211), .A2(n_569), .B(n_570), .Y(n_568) );
OAI21xp5_ASAP7_75t_L g212 ( .A1(n_213), .A2(n_216), .B(n_223), .Y(n_212) );
OAI22xp5_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B1(n_220), .B2(n_221), .Y(n_216) );
INVxp67_ASAP7_75t_L g218 ( .A(n_219), .Y(n_218) );
INVxp67_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g296 ( .A(n_224), .Y(n_296) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
AND2x2_ASAP7_75t_L g310 ( .A(n_225), .B(n_238), .Y(n_310) );
INVx1_ASAP7_75t_L g326 ( .A(n_225), .Y(n_326) );
HB1xp67_ASAP7_75t_L g434 ( .A(n_225), .Y(n_434) );
AND2x2_ASAP7_75t_L g225 ( .A(n_226), .B(n_231), .Y(n_225) );
NOR3xp33_ASAP7_75t_L g227 ( .A(n_228), .B(n_229), .C(n_230), .Y(n_227) );
AO21x2_ASAP7_75t_L g252 ( .A1(n_236), .A2(n_253), .B(n_261), .Y(n_252) );
AO21x2_ASAP7_75t_L g303 ( .A1(n_236), .A2(n_253), .B(n_261), .Y(n_303) );
AND2x2_ASAP7_75t_L g297 ( .A(n_237), .B(n_298), .Y(n_297) );
OR2x6_ASAP7_75t_L g378 ( .A(n_237), .B(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g416 ( .A(n_237), .B(n_413), .Y(n_416) );
BUFx6f_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
INVx4_ASAP7_75t_L g275 ( .A(n_238), .Y(n_275) );
NAND2xp5_ASAP7_75t_SL g283 ( .A(n_238), .B(n_284), .Y(n_283) );
INVx2_ASAP7_75t_L g345 ( .A(n_238), .Y(n_345) );
OR2x2_ASAP7_75t_L g351 ( .A(n_238), .B(n_265), .Y(n_351) );
AND2x4_ASAP7_75t_L g365 ( .A(n_238), .B(n_326), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_238), .B(n_334), .Y(n_366) );
OR2x6_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
INVx1_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
AND2x2_ASAP7_75t_L g247 ( .A(n_248), .B(n_250), .Y(n_247) );
INVx1_ASAP7_75t_SL g248 ( .A(n_249), .Y(n_248) );
AND2x2_ASAP7_75t_L g410 ( .A(n_249), .B(n_329), .Y(n_410) );
BUFx2_ASAP7_75t_L g462 ( .A(n_249), .Y(n_462) );
INVx1_ASAP7_75t_L g250 ( .A(n_251), .Y(n_250) );
OR2x2_ASAP7_75t_L g493 ( .A(n_251), .B(n_405), .Y(n_493) );
INVx2_ASAP7_75t_L g287 ( .A(n_252), .Y(n_287) );
NAND2xp5_ASAP7_75t_SL g253 ( .A(n_254), .B(n_260), .Y(n_253) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_263), .B(n_274), .Y(n_262) );
AND2x2_ASAP7_75t_L g309 ( .A(n_263), .B(n_310), .Y(n_309) );
HB1xp67_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
AND2x4_ASAP7_75t_SL g294 ( .A(n_264), .B(n_284), .Y(n_294) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
INVx2_ASAP7_75t_L g282 ( .A(n_265), .Y(n_282) );
HB1xp67_ASAP7_75t_L g388 ( .A(n_265), .Y(n_388) );
HB1xp67_ASAP7_75t_L g455 ( .A(n_265), .Y(n_455) );
INVx1_ASAP7_75t_L g495 ( .A(n_265), .Y(n_495) );
AO21x2_ASAP7_75t_L g265 ( .A1(n_266), .A2(n_267), .B(n_273), .Y(n_265) );
AO21x2_ASAP7_75t_L g583 ( .A1(n_266), .A2(n_584), .B(n_590), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_268), .B(n_269), .Y(n_267) );
BUFx2_ASAP7_75t_L g409 ( .A(n_274), .Y(n_409) );
NOR2x1_ASAP7_75t_L g274 ( .A(n_275), .B(n_276), .Y(n_274) );
AND2x4_ASAP7_75t_L g325 ( .A(n_275), .B(n_326), .Y(n_325) );
NOR2xp67_ASAP7_75t_SL g357 ( .A(n_275), .B(n_358), .Y(n_357) );
AND2x2_ASAP7_75t_L g430 ( .A(n_275), .B(n_413), .Y(n_430) );
AND2x4_ASAP7_75t_SL g433 ( .A(n_275), .B(n_434), .Y(n_433) );
OR2x2_ASAP7_75t_L g482 ( .A(n_275), .B(n_483), .Y(n_482) );
INVx2_ASAP7_75t_L g349 ( .A(n_276), .Y(n_349) );
INVx4_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
AND2x2_ASAP7_75t_L g344 ( .A(n_277), .B(n_345), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_277), .B(n_342), .Y(n_362) );
NAND2xp5_ASAP7_75t_L g401 ( .A(n_277), .B(n_402), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_277), .B(n_466), .Y(n_465) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
NOR2x1_ASAP7_75t_L g279 ( .A(n_280), .B(n_283), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
OR2x2_ASAP7_75t_L g427 ( .A(n_281), .B(n_428), .Y(n_427) );
HB1xp67_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
INVx2_ASAP7_75t_L g343 ( .A(n_282), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g285 ( .A(n_286), .B(n_289), .Y(n_285) );
AND2x2_ASAP7_75t_L g461 ( .A(n_286), .B(n_462), .Y(n_461) );
AND2x2_ASAP7_75t_L g469 ( .A(n_286), .B(n_398), .Y(n_469) );
AND2x2_ASAP7_75t_L g286 ( .A(n_287), .B(n_288), .Y(n_286) );
AND2x2_ASAP7_75t_L g338 ( .A(n_287), .B(n_323), .Y(n_338) );
AND2x4_ASAP7_75t_L g371 ( .A(n_287), .B(n_305), .Y(n_371) );
INVx1_ASAP7_75t_L g488 ( .A(n_287), .Y(n_488) );
AND2x2_ASAP7_75t_L g374 ( .A(n_289), .B(n_314), .Y(n_374) );
INVx2_ASAP7_75t_SL g289 ( .A(n_290), .Y(n_289) );
OR2x2_ASAP7_75t_L g395 ( .A(n_290), .B(n_330), .Y(n_395) );
OAI22xp5_ASAP7_75t_L g291 ( .A1(n_292), .A2(n_299), .B1(n_308), .B2(n_311), .Y(n_291) );
AOI21xp5_ASAP7_75t_L g292 ( .A1(n_293), .A2(n_295), .B(n_297), .Y(n_292) );
OAI22xp5_ASAP7_75t_SL g474 ( .A1(n_293), .A2(n_362), .B1(n_470), .B2(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_294), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g363 ( .A(n_294), .B(n_295), .Y(n_363) );
AND2x2_ASAP7_75t_SL g393 ( .A(n_294), .B(n_365), .Y(n_393) );
AOI211xp5_ASAP7_75t_SL g481 ( .A1(n_294), .A2(n_482), .B(n_484), .C(n_485), .Y(n_481) );
AND2x2_ASAP7_75t_SL g412 ( .A(n_295), .B(n_413), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_295), .B(n_341), .Y(n_467) );
INVx2_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g372 ( .A(n_297), .Y(n_372) );
INVx2_ASAP7_75t_L g428 ( .A(n_298), .Y(n_428) );
AND2x2_ASAP7_75t_L g502 ( .A(n_298), .B(n_495), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g450 ( .A1(n_299), .A2(n_451), .B(n_457), .Y(n_450) );
OR2x2_ASAP7_75t_L g299 ( .A(n_300), .B(n_304), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
AND2x4_ASAP7_75t_L g437 ( .A(n_301), .B(n_438), .Y(n_437) );
AND2x2_ASAP7_75t_L g447 ( .A(n_301), .B(n_448), .Y(n_447) );
AND2x2_ASAP7_75t_L g301 ( .A(n_302), .B(n_303), .Y(n_301) );
AND2x2_ASAP7_75t_L g354 ( .A(n_302), .B(n_307), .Y(n_354) );
NOR2xp67_ASAP7_75t_L g356 ( .A(n_302), .B(n_323), .Y(n_356) );
AND2x2_ASAP7_75t_L g398 ( .A(n_302), .B(n_323), .Y(n_398) );
INVx2_ASAP7_75t_L g315 ( .A(n_303), .Y(n_315) );
AND2x4_ASAP7_75t_L g321 ( .A(n_303), .B(n_322), .Y(n_321) );
NAND2x1p5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx3_ASAP7_75t_L g313 ( .A(n_305), .Y(n_313) );
INVx3_ASAP7_75t_L g319 ( .A(n_306), .Y(n_319) );
BUFx3_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
OAI21xp5_ASAP7_75t_L g496 ( .A1(n_310), .A2(n_416), .B(n_492), .Y(n_496) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
AND2x2_ASAP7_75t_L g312 ( .A(n_313), .B(n_314), .Y(n_312) );
INVx1_ASAP7_75t_L g328 ( .A(n_313), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_313), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_313), .B(n_388), .Y(n_403) );
OR2x2_ASAP7_75t_L g418 ( .A(n_313), .B(n_419), .Y(n_418) );
AND2x2_ASAP7_75t_L g425 ( .A(n_313), .B(n_329), .Y(n_425) );
AND2x2_ASAP7_75t_L g381 ( .A(n_314), .B(n_382), .Y(n_381) );
AND2x2_ASAP7_75t_L g397 ( .A(n_314), .B(n_398), .Y(n_397) );
AND2x2_ASAP7_75t_L g414 ( .A(n_314), .B(n_383), .Y(n_414) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_317), .A2(n_324), .B1(n_327), .B2(n_331), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
NOR2xp67_ASAP7_75t_L g391 ( .A(n_319), .B(n_320), .Y(n_391) );
NOR2xp67_ASAP7_75t_SL g429 ( .A(n_319), .B(n_337), .Y(n_429) );
INVxp67_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_L g322 ( .A(n_323), .Y(n_322) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_323), .B(n_449), .Y(n_448) );
AND2x2_ASAP7_75t_L g332 ( .A(n_325), .B(n_333), .Y(n_332) );
AND2x2_ASAP7_75t_L g396 ( .A(n_325), .B(n_342), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_325), .B(n_460), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_328), .B(n_329), .Y(n_327) );
INVx2_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AND2x2_ASAP7_75t_L g499 ( .A(n_333), .B(n_365), .Y(n_499) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
NOR2x1_ASAP7_75t_L g444 ( .A(n_334), .B(n_445), .Y(n_444) );
NOR2xp67_ASAP7_75t_SL g335 ( .A(n_336), .B(n_359), .Y(n_335) );
OAI211xp5_ASAP7_75t_L g336 ( .A1(n_337), .A2(n_339), .B(n_346), .C(n_355), .Y(n_336) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_337), .A2(n_390), .B(n_400), .C(n_404), .Y(n_399) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g479 ( .A(n_338), .B(n_480), .Y(n_479) );
INVx2_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_344), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g390 ( .A(n_342), .B(n_366), .Y(n_390) );
AND2x2_ASAP7_75t_L g477 ( .A(n_342), .B(n_456), .Y(n_477) );
INVx3_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g445 ( .A(n_345), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_352), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2x1_ASAP7_75t_L g348 ( .A(n_349), .B(n_350), .Y(n_348) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_349), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
INVx2_ASAP7_75t_L g419 ( .A(n_354), .Y(n_419) );
NAND2xp33_ASAP7_75t_SL g355 ( .A(n_356), .B(n_357), .Y(n_355) );
OAI221xp5_ASAP7_75t_L g359 ( .A1(n_360), .A2(n_367), .B1(n_369), .B2(n_372), .C(n_373), .Y(n_359) );
NOR4xp25_ASAP7_75t_L g360 ( .A(n_361), .B(n_363), .C(n_364), .D(n_366), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
HB1xp67_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AND2x2_ASAP7_75t_L g478 ( .A(n_365), .B(n_441), .Y(n_478) );
INVx2_ASAP7_75t_L g484 ( .A(n_365), .Y(n_484) );
INVx2_ASAP7_75t_SL g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_368), .B(n_432), .Y(n_431) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
AND2x2_ASAP7_75t_L g471 ( .A(n_371), .B(n_472), .Y(n_471) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
NAND4xp75_ASAP7_75t_L g376 ( .A(n_377), .B(n_399), .C(n_406), .D(n_415), .Y(n_376) );
OA211x2_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_380), .B(n_384), .C(n_392), .Y(n_377) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_378), .B(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g472 ( .A(n_382), .Y(n_472) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g480 ( .A(n_383), .Y(n_480) );
NAND2xp5_ASAP7_75t_SL g384 ( .A(n_385), .B(n_391), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_386), .B(n_389), .Y(n_385) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx2_ASAP7_75t_L g441 ( .A(n_388), .Y(n_441) );
INVx1_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_393), .A2(n_394), .B1(n_396), .B2(n_397), .Y(n_392) );
INVx1_ASAP7_75t_SL g394 ( .A(n_395), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g501 ( .A1(n_396), .A2(n_447), .B(n_502), .Y(n_501) );
INVx1_ASAP7_75t_SL g475 ( .A(n_397), .Y(n_475) );
NAND2x1p5_ASAP7_75t_L g487 ( .A(n_398), .B(n_488), .Y(n_487) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_401), .Y(n_400) );
INVx1_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
NOR2x1_ASAP7_75t_L g406 ( .A(n_407), .B(n_411), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_409), .B(n_410), .Y(n_408) );
INVxp67_ASAP7_75t_L g473 ( .A(n_409), .Y(n_473) );
AND2x2_ASAP7_75t_L g411 ( .A(n_412), .B(n_414), .Y(n_411) );
AND2x2_ASAP7_75t_SL g432 ( .A(n_413), .B(n_433), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g498 ( .A1(n_414), .A2(n_477), .B1(n_499), .B2(n_500), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_416), .B(n_417), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx2_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
NAND3x1_ASAP7_75t_L g421 ( .A(n_422), .B(n_463), .C(n_476), .Y(n_421) );
NOR3x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_435), .C(n_450), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g423 ( .A(n_424), .B(n_431), .Y(n_423) );
AOI22xp5_ASAP7_75t_L g424 ( .A1(n_425), .A2(n_426), .B1(n_429), .B2(n_430), .Y(n_424) );
OAI22xp5_ASAP7_75t_L g435 ( .A1(n_436), .A2(n_440), .B1(n_442), .B2(n_446), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVxp67_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
AND2x2_ASAP7_75t_L g494 ( .A(n_444), .B(n_495), .Y(n_494) );
INVx1_ASAP7_75t_SL g446 ( .A(n_447), .Y(n_446) );
INVx1_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_453), .B(n_456), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_458), .B(n_461), .Y(n_457) );
INVxp67_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_SL g483 ( .A(n_460), .Y(n_483) );
OAI21xp5_ASAP7_75t_SL g491 ( .A1(n_461), .A2(n_492), .B(n_494), .Y(n_491) );
NOR2x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_474), .Y(n_463) );
OAI22xp5_ASAP7_75t_L g464 ( .A1(n_465), .A2(n_468), .B1(n_470), .B2(n_473), .Y(n_464) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
O2A1O1Ixp5_ASAP7_75t_L g476 ( .A1(n_477), .A2(n_478), .B(n_479), .C(n_481), .Y(n_476) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
NOR2x1_ASAP7_75t_SL g489 ( .A(n_490), .B(n_497), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_491), .B(n_496), .Y(n_490) );
INVx1_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g497 ( .A(n_498), .B(n_501), .Y(n_497) );
XOR2x1_ASAP7_75t_SL g814 ( .A(n_503), .B(n_815), .Y(n_814) );
AND2x4_ASAP7_75t_L g503 ( .A(n_504), .B(n_702), .Y(n_503) );
NOR3xp33_ASAP7_75t_L g504 ( .A(n_505), .B(n_639), .C(n_662), .Y(n_504) );
NAND3xp33_ASAP7_75t_SL g505 ( .A(n_506), .B(n_591), .C(n_608), .Y(n_505) );
OAI31xp33_ASAP7_75t_SL g506 ( .A1(n_507), .A2(n_527), .A3(n_547), .B(n_554), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_507), .B(n_666), .Y(n_665) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_521), .Y(n_508) );
AND2x4_ASAP7_75t_L g594 ( .A(n_509), .B(n_521), .Y(n_594) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_509), .B(n_538), .Y(n_623) );
AND2x4_ASAP7_75t_L g625 ( .A(n_509), .B(n_619), .Y(n_625) );
AND2x2_ASAP7_75t_L g756 ( .A(n_509), .B(n_551), .Y(n_756) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
INVx2_ASAP7_75t_L g601 ( .A(n_510), .Y(n_601) );
OAI21x1_ASAP7_75t_SL g510 ( .A1(n_511), .A2(n_514), .B(n_519), .Y(n_510) );
INVx1_ASAP7_75t_L g520 ( .A(n_513), .Y(n_520) );
AND2x2_ASAP7_75t_L g537 ( .A(n_521), .B(n_538), .Y(n_537) );
AND2x2_ASAP7_75t_SL g692 ( .A(n_521), .B(n_600), .Y(n_692) );
AND2x2_ASAP7_75t_L g698 ( .A(n_521), .B(n_539), .Y(n_698) );
AND2x2_ASAP7_75t_L g787 ( .A(n_521), .B(n_788), .Y(n_787) );
INVx1_ASAP7_75t_SL g769 ( .A(n_527), .Y(n_769) );
AND2x2_ASAP7_75t_L g527 ( .A(n_528), .B(n_537), .Y(n_527) );
BUFx2_ASAP7_75t_L g598 ( .A(n_528), .Y(n_598) );
AND2x2_ASAP7_75t_L g632 ( .A(n_528), .B(n_538), .Y(n_632) );
AND2x2_ASAP7_75t_L g681 ( .A(n_528), .B(n_539), .Y(n_681) );
INVx2_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
AND2x2_ASAP7_75t_L g638 ( .A(n_529), .B(n_539), .Y(n_638) );
INVxp67_ASAP7_75t_L g650 ( .A(n_529), .Y(n_650) );
BUFx3_ASAP7_75t_L g695 ( .A(n_529), .Y(n_695) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_531), .B(n_535), .Y(n_530) );
OAI31xp33_ASAP7_75t_L g591 ( .A1(n_537), .A2(n_592), .A3(n_597), .B(n_602), .Y(n_591) );
AND2x2_ASAP7_75t_L g599 ( .A(n_538), .B(n_600), .Y(n_599) );
INVx2_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
AND2x2_ASAP7_75t_L g618 ( .A(n_539), .B(n_619), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_545), .Y(n_540) );
AOI322xp5_ASAP7_75t_L g792 ( .A1(n_547), .A2(n_667), .A3(n_696), .B1(n_701), .B2(n_793), .C1(n_796), .C2(n_797), .Y(n_792) );
AND2x2_ASAP7_75t_L g547 ( .A(n_548), .B(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_548), .B(n_638), .Y(n_643) );
NAND2x1_ASAP7_75t_L g680 ( .A(n_548), .B(n_681), .Y(n_680) );
AND2x4_ASAP7_75t_L g724 ( .A(n_548), .B(n_628), .Y(n_724) );
INVx1_ASAP7_75t_SL g738 ( .A(n_548), .Y(n_738) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g619 ( .A(n_549), .Y(n_619) );
HB1xp67_ASAP7_75t_L g762 ( .A(n_549), .Y(n_762) );
AND2x2_ASAP7_75t_L g691 ( .A(n_550), .B(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_550), .B(n_738), .Y(n_737) );
AND2x4_ASAP7_75t_SL g550 ( .A(n_551), .B(n_552), .Y(n_550) );
BUFx2_ASAP7_75t_L g596 ( .A(n_551), .Y(n_596) );
INVx1_ASAP7_75t_L g788 ( .A(n_551), .Y(n_788) );
OR2x2_ASAP7_75t_L g655 ( .A(n_552), .B(n_600), .Y(n_655) );
NAND2xp5_ASAP7_75t_SL g689 ( .A(n_552), .B(n_625), .Y(n_689) );
INVx2_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g628 ( .A(n_553), .B(n_600), .Y(n_628) );
AND2x2_ASAP7_75t_L g554 ( .A(n_555), .B(n_574), .Y(n_554) );
INVxp67_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g684 ( .A(n_556), .Y(n_684) );
OR2x2_ASAP7_75t_L g711 ( .A(n_556), .B(n_712), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g556 ( .A(n_557), .B(n_567), .Y(n_556) );
NOR2x1_ASAP7_75t_SL g605 ( .A(n_557), .B(n_575), .Y(n_605) );
AND2x2_ASAP7_75t_L g612 ( .A(n_557), .B(n_613), .Y(n_612) );
AND2x2_ASAP7_75t_L g784 ( .A(n_557), .B(n_646), .Y(n_784) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_557) );
NOR2xp33_ASAP7_75t_L g565 ( .A(n_558), .B(n_566), .Y(n_565) );
AO21x2_ASAP7_75t_L g661 ( .A1(n_558), .A2(n_559), .B(n_565), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_560), .B(n_564), .Y(n_559) );
OR2x2_ASAP7_75t_L g606 ( .A(n_567), .B(n_607), .Y(n_606) );
BUFx3_ASAP7_75t_L g615 ( .A(n_567), .Y(n_615) );
INVx2_ASAP7_75t_L g646 ( .A(n_567), .Y(n_646) );
INVx1_ASAP7_75t_L g687 ( .A(n_567), .Y(n_687) );
AND2x2_ASAP7_75t_L g718 ( .A(n_567), .B(n_575), .Y(n_718) );
AND2x2_ASAP7_75t_L g749 ( .A(n_567), .B(n_676), .Y(n_749) );
AND2x2_ASAP7_75t_L g645 ( .A(n_574), .B(n_646), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_574), .B(n_658), .Y(n_657) );
AND2x2_ASAP7_75t_SL g748 ( .A(n_574), .B(n_749), .Y(n_748) );
AND2x2_ASAP7_75t_L g753 ( .A(n_574), .B(n_615), .Y(n_753) );
AND2x2_ASAP7_75t_L g574 ( .A(n_575), .B(n_583), .Y(n_574) );
INVx5_ASAP7_75t_L g613 ( .A(n_575), .Y(n_613) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_575), .B(n_607), .Y(n_685) );
BUFx2_ASAP7_75t_L g745 ( .A(n_575), .Y(n_745) );
OR2x6_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
INVx4_ASAP7_75t_L g607 ( .A(n_583), .Y(n_607) );
AND2x2_ASAP7_75t_L g730 ( .A(n_583), .B(n_613), .Y(n_730) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_585), .B(n_589), .Y(n_584) );
INVx1_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
OAI221xp5_ASAP7_75t_L g719 ( .A1(n_593), .A2(n_720), .B1(n_723), .B2(n_725), .C(n_726), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_594), .B(n_595), .Y(n_593) );
AND2x2_ASAP7_75t_L g741 ( .A(n_594), .B(n_632), .Y(n_741) );
INVx1_ASAP7_75t_SL g767 ( .A(n_594), .Y(n_767) );
AND2x2_ASAP7_75t_L g752 ( .A(n_595), .B(n_724), .Y(n_752) );
INVx2_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g697 ( .A(n_596), .B(n_698), .Y(n_697) );
AND2x2_ASAP7_75t_L g597 ( .A(n_598), .B(n_599), .Y(n_597) );
AND2x2_ASAP7_75t_L g621 ( .A(n_598), .B(n_622), .Y(n_621) );
AND2x2_ASAP7_75t_L g627 ( .A(n_598), .B(n_628), .Y(n_627) );
INVx1_ASAP7_75t_L g651 ( .A(n_599), .Y(n_651) );
AND2x2_ASAP7_75t_L g709 ( .A(n_599), .B(n_637), .Y(n_709) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
BUFx2_ASAP7_75t_L g634 ( .A(n_601), .Y(n_634) );
INVx1_ASAP7_75t_SL g602 ( .A(n_603), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_604), .B(n_606), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVx2_ASAP7_75t_L g630 ( .A(n_606), .Y(n_630) );
OR2x2_ASAP7_75t_L g798 ( .A(n_606), .B(n_799), .Y(n_798) );
INVx2_ASAP7_75t_L g614 ( .A(n_607), .Y(n_614) );
AND2x4_ASAP7_75t_L g670 ( .A(n_607), .B(n_671), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g674 ( .A(n_607), .B(n_675), .Y(n_674) );
NAND2x1p5_ASAP7_75t_L g712 ( .A(n_607), .B(n_613), .Y(n_712) );
AND2x2_ASAP7_75t_L g772 ( .A(n_607), .B(n_675), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_616), .B1(n_629), .B2(n_631), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_609), .B(n_691), .Y(n_690) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
AND3x2_ASAP7_75t_L g611 ( .A(n_612), .B(n_614), .C(n_615), .Y(n_611) );
AND2x4_ASAP7_75t_L g629 ( .A(n_612), .B(n_630), .Y(n_629) );
INVx4_ASAP7_75t_L g669 ( .A(n_613), .Y(n_669) );
AND2x2_ASAP7_75t_SL g802 ( .A(n_613), .B(n_670), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g777 ( .A(n_614), .B(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g714 ( .A(n_615), .Y(n_714) );
AOI322xp5_ASAP7_75t_L g779 ( .A1(n_615), .A2(n_744), .A3(n_780), .B1(n_782), .B2(n_785), .C1(n_789), .C2(n_790), .Y(n_779) );
NAND4xp25_ASAP7_75t_SL g616 ( .A(n_617), .B(n_620), .C(n_624), .D(n_626), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_SL g746 ( .A(n_618), .B(n_634), .Y(n_746) );
BUFx2_ASAP7_75t_L g637 ( .A(n_619), .Y(n_637) );
INVx1_ASAP7_75t_SL g620 ( .A(n_621), .Y(n_620) );
AND2x2_ASAP7_75t_L g761 ( .A(n_622), .B(n_762), .Y(n_761) );
INVx1_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OR2x2_ASAP7_75t_L g775 ( .A(n_623), .B(n_650), .Y(n_775) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g641 ( .A(n_625), .B(n_642), .Y(n_641) );
OAI211xp5_ASAP7_75t_L g693 ( .A1(n_625), .A2(n_694), .B(n_696), .C(n_699), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_625), .B(n_632), .Y(n_751) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_627), .A2(n_709), .B1(n_710), .B2(n_713), .Y(n_708) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_628), .A2(n_664), .B1(n_668), .B2(n_672), .Y(n_663) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_628), .B(n_717), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g764 ( .A(n_628), .B(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_628), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_L g795 ( .A(n_628), .Y(n_795) );
INVx1_ASAP7_75t_L g734 ( .A(n_629), .Y(n_734) );
OAI21xp33_ASAP7_75t_SL g631 ( .A1(n_632), .A2(n_633), .B(n_635), .Y(n_631) );
INVx1_ASAP7_75t_L g642 ( .A(n_632), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_632), .B(n_637), .Y(n_791) );
INVx1_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
AND2x2_ASAP7_75t_L g727 ( .A(n_634), .B(n_638), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_638), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_636), .B(n_654), .Y(n_653) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
OR2x2_ASAP7_75t_L g794 ( .A(n_637), .B(n_795), .Y(n_794) );
INVx1_ASAP7_75t_L g768 ( .A(n_638), .Y(n_768) );
A2O1A1Ixp33_ASAP7_75t_L g639 ( .A1(n_640), .A2(n_643), .B(n_644), .C(n_647), .Y(n_639) );
INVxp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI22xp33_ASAP7_75t_SL g754 ( .A1(n_642), .A2(n_673), .B1(n_720), .B2(n_755), .Y(n_754) );
INVx1_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_646), .B(n_669), .Y(n_677) );
OR2x2_ASAP7_75t_L g706 ( .A(n_646), .B(n_707), .Y(n_706) );
OAI21xp5_ASAP7_75t_SL g647 ( .A1(n_648), .A2(n_652), .B(n_656), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_650), .B(n_651), .Y(n_649) );
INVx1_ASAP7_75t_L g667 ( .A(n_650), .Y(n_667) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
OAI211xp5_ASAP7_75t_SL g705 ( .A1(n_653), .A2(n_706), .B(n_708), .C(n_716), .Y(n_705) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g656 ( .A(n_657), .Y(n_656) );
NOR2xp67_ASAP7_75t_SL g739 ( .A(n_658), .B(n_685), .Y(n_739) );
INVx1_ASAP7_75t_L g742 ( .A(n_658), .Y(n_742) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_660), .B(n_669), .Y(n_799) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g671 ( .A(n_661), .Y(n_671) );
INVx2_ASAP7_75t_L g676 ( .A(n_661), .Y(n_676) );
NAND4xp25_ASAP7_75t_L g662 ( .A(n_663), .B(n_678), .C(n_690), .D(n_693), .Y(n_662) );
INVx1_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
OAI22xp33_ASAP7_75t_L g797 ( .A1(n_666), .A2(n_798), .B1(n_800), .B2(n_801), .Y(n_797) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
AND2x4_ASAP7_75t_L g765 ( .A(n_669), .B(n_695), .Y(n_765) );
AND2x2_ASAP7_75t_L g686 ( .A(n_670), .B(n_687), .Y(n_686) );
INVx2_ASAP7_75t_L g707 ( .A(n_670), .Y(n_707) );
AND2x2_ASAP7_75t_L g717 ( .A(n_670), .B(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
OR2x2_ASAP7_75t_L g673 ( .A(n_674), .B(n_677), .Y(n_673) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_676), .Y(n_731) );
INVx1_ASAP7_75t_L g721 ( .A(n_677), .Y(n_721) );
AOI32xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .A3(n_685), .B1(n_686), .B2(n_688), .Y(n_678) );
OAI21xp33_ASAP7_75t_L g726 ( .A1(n_679), .A2(n_727), .B(n_728), .Y(n_726) );
INVx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI221xp5_ASAP7_75t_L g758 ( .A1(n_682), .A2(n_759), .B1(n_761), .B2(n_763), .C(n_766), .Y(n_758) );
INVx1_ASAP7_75t_SL g682 ( .A(n_683), .Y(n_682) );
INVx1_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AND2x2_ASAP7_75t_L g743 ( .A(n_684), .B(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g701 ( .A(n_685), .Y(n_701) );
AOI22xp5_ASAP7_75t_L g773 ( .A1(n_686), .A2(n_724), .B1(n_774), .B2(n_776), .Y(n_773) );
INVx1_ASAP7_75t_L g700 ( .A(n_687), .Y(n_700) );
AND2x2_ASAP7_75t_L g778 ( .A(n_687), .B(n_731), .Y(n_778) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_SL g781 ( .A(n_694), .B(n_746), .Y(n_781) );
INVx1_ASAP7_75t_L g800 ( .A(n_694), .Y(n_800) );
INVx1_ASAP7_75t_SL g694 ( .A(n_695), .Y(n_694) );
INVx1_ASAP7_75t_L g696 ( .A(n_697), .Y(n_696) );
AND2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_701), .Y(n_699) );
NOR2xp67_ASAP7_75t_L g702 ( .A(n_703), .B(n_757), .Y(n_702) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_704), .B(n_747), .Y(n_703) );
NOR3xp33_ASAP7_75t_SL g704 ( .A(n_705), .B(n_719), .C(n_732), .Y(n_704) );
INVx1_ASAP7_75t_L g722 ( .A(n_707), .Y(n_722) );
INVx1_ASAP7_75t_SL g733 ( .A(n_709), .Y(n_733) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
INVx2_ASAP7_75t_L g715 ( .A(n_712), .Y(n_715) );
INVx2_ASAP7_75t_L g725 ( .A(n_713), .Y(n_725) );
AND2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
AND2x4_ASAP7_75t_L g771 ( .A(n_714), .B(n_772), .Y(n_771) );
AND2x4_ASAP7_75t_L g789 ( .A(n_718), .B(n_772), .Y(n_789) );
NAND2xp5_ASAP7_75t_SL g720 ( .A(n_721), .B(n_722), .Y(n_720) );
INVx1_ASAP7_75t_SL g723 ( .A(n_724), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g728 ( .A(n_729), .B(n_731), .Y(n_728) );
AOI32xp33_ASAP7_75t_L g740 ( .A1(n_729), .A2(n_741), .A3(n_742), .B1(n_743), .B2(n_746), .Y(n_740) );
NOR2xp33_ASAP7_75t_SL g759 ( .A(n_729), .B(n_760), .Y(n_759) );
INVx2_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g760 ( .A(n_731), .Y(n_760) );
OAI211xp5_ASAP7_75t_SL g732 ( .A1(n_733), .A2(n_734), .B(n_735), .C(n_740), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_736), .B(n_739), .Y(n_735) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g796 ( .A(n_744), .B(n_784), .Y(n_796) );
INVx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
NAND2xp5_ASAP7_75t_L g783 ( .A(n_745), .B(n_784), .Y(n_783) );
AOI221xp5_ASAP7_75t_L g747 ( .A1(n_748), .A2(n_750), .B1(n_752), .B2(n_753), .C(n_754), .Y(n_747) );
INVx1_ASAP7_75t_SL g750 ( .A(n_751), .Y(n_750) );
CKINVDCx16_ASAP7_75t_R g755 ( .A(n_756), .Y(n_755) );
NAND4xp25_ASAP7_75t_L g757 ( .A(n_758), .B(n_773), .C(n_779), .D(n_792), .Y(n_757) );
INVxp33_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
O2A1O1Ixp33_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B(n_769), .C(n_770), .Y(n_766) );
INVx2_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
INVx1_ASAP7_75t_L g774 ( .A(n_775), .Y(n_774) );
INVx1_ASAP7_75t_SL g776 ( .A(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g780 ( .A(n_781), .Y(n_780) );
INVx1_ASAP7_75t_L g782 ( .A(n_783), .Y(n_782) );
INVx1_ASAP7_75t_SL g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx2_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx3_ASAP7_75t_SL g801 ( .A(n_802), .Y(n_801) );
BUFx2_ASAP7_75t_L g804 ( .A(n_805), .Y(n_804) );
CKINVDCx5p33_ASAP7_75t_R g806 ( .A(n_807), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_809), .B(n_823), .Y(n_808) );
AOI31xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_814), .A3(n_821), .B(n_822), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_811), .Y(n_810) );
OR3x1_ASAP7_75t_L g823 ( .A(n_811), .B(n_814), .C(n_821), .Y(n_823) );
INVx1_ASAP7_75t_L g811 ( .A(n_812), .Y(n_811) );
HB1xp67_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
INVx1_ASAP7_75t_L g819 ( .A(n_816), .Y(n_819) );
INVx3_ASAP7_75t_L g824 ( .A(n_825), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
NOR2xp33_ASAP7_75t_L g831 ( .A(n_826), .B(n_832), .Y(n_831) );
AND2x2_ASAP7_75t_SL g826 ( .A(n_827), .B(n_828), .Y(n_826) );
endmodule