module fake_jpeg_13965_n_472 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_472);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_472;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_389;
wire n_457;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_15),
.B(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx3_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx24_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

INVx5_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_2),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_13),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

BUFx12_ASAP7_75t_L g37 ( 
.A(n_15),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_13),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_15),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_13),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_12),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_9),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_11),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_0),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g150 ( 
.A(n_49),
.Y(n_150)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_50),
.Y(n_115)
);

INVx4_ASAP7_75t_SL g51 ( 
.A(n_22),
.Y(n_51)
);

INVx5_ASAP7_75t_SL g128 ( 
.A(n_51),
.Y(n_128)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

INVx5_ASAP7_75t_L g121 ( 
.A(n_52),
.Y(n_121)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_53),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_16),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_55),
.Y(n_129)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_31),
.Y(n_56)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_56),
.Y(n_139)
);

BUFx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx5_ASAP7_75t_L g122 ( 
.A(n_57),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_19),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_58),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_17),
.B(n_7),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_59),
.B(n_91),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_17),
.B(n_7),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_60),
.B(n_78),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_61),
.Y(n_102)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_62),
.Y(n_141)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_22),
.Y(n_63)
);

INVx4_ASAP7_75t_L g106 ( 
.A(n_63),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_22),
.Y(n_64)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_64),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g65 ( 
.A(n_26),
.Y(n_65)
);

INVx4_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx4_ASAP7_75t_L g132 ( 
.A(n_66),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_19),
.Y(n_67)
);

INVx6_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_22),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g98 ( 
.A(n_68),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_21),
.A2(n_7),
.B1(n_12),
.B2(n_11),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_69),
.A2(n_43),
.B1(n_41),
.B2(n_24),
.Y(n_100)
);

INVx6_ASAP7_75t_L g70 ( 
.A(n_16),
.Y(n_70)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_70),
.Y(n_114)
);

BUFx2_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx4_ASAP7_75t_L g142 ( 
.A(n_72),
.Y(n_142)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_16),
.Y(n_73)
);

INVx4_ASAP7_75t_L g146 ( 
.A(n_73),
.Y(n_146)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_38),
.Y(n_74)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_26),
.Y(n_76)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_76),
.Y(n_134)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_77),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_37),
.Y(n_78)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_21),
.Y(n_79)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_79),
.Y(n_108)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_16),
.Y(n_80)
);

INVx11_ASAP7_75t_L g138 ( 
.A(n_80),
.Y(n_138)
);

INVx5_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx8_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_83),
.Y(n_147)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_84),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_20),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g99 ( 
.A(n_85),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_86),
.B(n_90),
.Y(n_148)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_20),
.Y(n_87)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_87),
.Y(n_116)
);

INVx5_ASAP7_75t_L g88 ( 
.A(n_21),
.Y(n_88)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_88),
.Y(n_149)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_29),
.Y(n_89)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_89),
.Y(n_152)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_36),
.Y(n_90)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_36),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_18),
.B(n_39),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_92),
.B(n_93),
.Y(n_123)
);

INVx5_ASAP7_75t_L g93 ( 
.A(n_36),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_32),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_94),
.B(n_96),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g95 ( 
.A(n_29),
.Y(n_95)
);

OAI21xp33_ASAP7_75t_L g104 ( 
.A1(n_95),
.A2(n_51),
.B(n_35),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_32),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_97),
.B(n_27),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g154 ( 
.A(n_100),
.B(n_104),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_95),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_103),
.B(n_52),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_59),
.A2(n_40),
.B1(n_28),
.B2(n_46),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_109),
.A2(n_144),
.B1(n_145),
.B2(n_98),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_60),
.A2(n_28),
.B1(n_40),
.B2(n_32),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_111),
.A2(n_118),
.B1(n_119),
.B2(n_25),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_64),
.A2(n_40),
.B1(n_28),
.B2(n_43),
.Y(n_112)
);

OAI22xp33_ASAP7_75t_L g203 ( 
.A1(n_112),
.A2(n_127),
.B1(n_130),
.B2(n_135),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_55),
.A2(n_46),
.B1(n_45),
.B2(n_44),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_70),
.A2(n_39),
.B1(n_45),
.B2(n_44),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_54),
.A2(n_40),
.B1(n_48),
.B2(n_23),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_58),
.A2(n_48),
.B1(n_23),
.B2(n_25),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_64),
.A2(n_43),
.B1(n_24),
.B2(n_41),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_136),
.B(n_153),
.Y(n_190)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_63),
.A2(n_24),
.B1(n_41),
.B2(n_47),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_72),
.A2(n_47),
.B1(n_35),
.B2(n_33),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_73),
.B(n_42),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_155),
.B(n_168),
.Y(n_213)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_156),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_157),
.Y(n_215)
);

INVx3_ASAP7_75t_L g158 ( 
.A(n_146),
.Y(n_158)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_158),
.Y(n_219)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_107),
.Y(n_159)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

INVx6_ASAP7_75t_L g160 ( 
.A(n_117),
.Y(n_160)
);

INVx3_ASAP7_75t_L g205 ( 
.A(n_160),
.Y(n_205)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_128),
.Y(n_161)
);

INVx3_ASAP7_75t_L g236 ( 
.A(n_161),
.Y(n_236)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_146),
.Y(n_162)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_162),
.Y(n_207)
);

INVx4_ASAP7_75t_L g163 ( 
.A(n_99),
.Y(n_163)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_163),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g164 ( 
.A(n_150),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_164),
.Y(n_226)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_152),
.Y(n_165)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_165),
.Y(n_211)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_99),
.Y(n_166)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_166),
.Y(n_220)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_167),
.Y(n_221)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_148),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_169),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_170),
.Y(n_233)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_121),
.Y(n_171)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_171),
.Y(n_227)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_115),
.Y(n_172)
);

INVxp67_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_104),
.Y(n_173)
);

OAI21xp33_ASAP7_75t_L g218 ( 
.A1(n_173),
.A2(n_180),
.B(n_182),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_110),
.B(n_18),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_174),
.B(n_184),
.Y(n_230)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_116),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_175),
.Y(n_242)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_137),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_176),
.B(n_177),
.Y(n_232)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_141),
.Y(n_177)
);

INVx2_ASAP7_75t_SL g178 ( 
.A(n_121),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g210 ( 
.A(n_178),
.Y(n_210)
);

INVx2_ASAP7_75t_SL g179 ( 
.A(n_122),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_179),
.B(n_181),
.Y(n_239)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

CKINVDCx6p67_ASAP7_75t_R g182 ( 
.A(n_138),
.Y(n_182)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_151),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_183),
.B(n_186),
.Y(n_212)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_149),
.Y(n_184)
);

INVx1_ASAP7_75t_SL g185 ( 
.A(n_139),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_185),
.A2(n_187),
.B1(n_189),
.B2(n_200),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_123),
.Y(n_186)
);

INVx1_ASAP7_75t_SL g187 ( 
.A(n_140),
.Y(n_187)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_120),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_191),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_135),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_134),
.Y(n_191)
);

NAND3xp33_ASAP7_75t_SL g192 ( 
.A(n_133),
.B(n_42),
.C(n_33),
.Y(n_192)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_192),
.A2(n_143),
.B1(n_142),
.B2(n_106),
.Y(n_237)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_120),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_193),
.B(n_194),
.Y(n_235)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_113),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_195),
.B(n_196),
.Y(n_240)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_113),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_147),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_197),
.B(n_199),
.Y(n_243)
);

OA22x2_ASAP7_75t_L g217 ( 
.A1(n_198),
.A2(n_137),
.B1(n_83),
.B2(n_96),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_132),
.B(n_125),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g200 ( 
.A(n_138),
.Y(n_200)
);

INVxp33_ASAP7_75t_L g201 ( 
.A(n_127),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g222 ( 
.A1(n_201),
.A2(n_80),
.B1(n_102),
.B2(n_105),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_130),
.B(n_131),
.Y(n_202)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_202),
.B(n_85),
.Y(n_231)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_203),
.A2(n_114),
.B1(n_105),
.B2(n_102),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_206),
.A2(n_229),
.B1(n_217),
.B2(n_161),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_173),
.A2(n_112),
.B1(n_145),
.B2(n_114),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g255 ( 
.A1(n_209),
.A2(n_223),
.B1(n_234),
.B2(n_238),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g274 ( 
.A(n_217),
.B(n_231),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_222),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_189),
.A2(n_144),
.B1(n_67),
.B2(n_97),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_L g224 ( 
.A1(n_154),
.A2(n_27),
.B(n_126),
.Y(n_224)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_224),
.A2(n_179),
.B(n_170),
.Y(n_252)
);

OAI22x1_ASAP7_75t_L g225 ( 
.A1(n_203),
.A2(n_106),
.B1(n_142),
.B2(n_125),
.Y(n_225)
);

OAI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_201),
.B1(n_166),
.B2(n_163),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_190),
.A2(n_87),
.B1(n_61),
.B2(n_75),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_237),
.B(n_185),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g238 ( 
.A1(n_154),
.A2(n_94),
.B1(n_129),
.B2(n_71),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g244 ( 
.A(n_233),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g308 ( 
.A(n_244),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_212),
.B(n_157),
.C(n_187),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_245),
.B(n_241),
.C(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_246),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_215),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_248),
.B(n_253),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_251),
.B1(n_268),
.B2(n_279),
.Y(n_280)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_216),
.Y(n_250)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_250),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g298 ( 
.A(n_252),
.Y(n_298)
);

NOR2xp33_ASAP7_75t_L g253 ( 
.A(n_213),
.B(n_230),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_240),
.Y(n_254)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_254),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_267),
.Y(n_312)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_240),
.Y(n_257)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_257),
.Y(n_313)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_258),
.B(n_259),
.Y(n_287)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_204),
.Y(n_259)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_260),
.A2(n_276),
.B1(n_278),
.B2(n_228),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g299 ( 
.A(n_261),
.B(n_263),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_218),
.B1(n_209),
.B2(n_223),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g300 ( 
.A1(n_262),
.A2(n_255),
.B1(n_252),
.B2(n_274),
.Y(n_300)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

OAI21xp33_ASAP7_75t_L g264 ( 
.A1(n_212),
.A2(n_182),
.B(n_10),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_SL g301 ( 
.A1(n_264),
.A2(n_277),
.B(n_210),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_158),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_266),
.Y(n_285)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_208),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_235),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g268 ( 
.A1(n_206),
.A2(n_217),
.B1(n_231),
.B2(n_224),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_211),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_269),
.B(n_270),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_162),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_236),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_271),
.B(n_275),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_229),
.A2(n_27),
.B(n_194),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_272),
.A2(n_273),
.B(n_220),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_243),
.A2(n_196),
.B(n_181),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_235),
.B(n_160),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_236),
.Y(n_276)
);

OA22x2_ASAP7_75t_L g277 ( 
.A1(n_217),
.A2(n_129),
.B1(n_132),
.B2(n_188),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_211),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_225),
.A2(n_169),
.B1(n_176),
.B2(n_122),
.Y(n_279)
);

XOR2xp5_ASAP7_75t_L g281 ( 
.A(n_245),
.B(n_238),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_281),
.B(n_289),
.C(n_290),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_275),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_282),
.B(n_293),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_268),
.A2(n_234),
.B1(n_221),
.B2(n_230),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g318 ( 
.A1(n_283),
.A2(n_306),
.B1(n_310),
.B2(n_280),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_246),
.B(n_250),
.C(n_254),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_270),
.Y(n_293)
);

MAJx2_ASAP7_75t_L g295 ( 
.A(n_257),
.B(n_265),
.C(n_274),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_L g334 ( 
.A(n_295),
.B(n_302),
.Y(n_334)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_258),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_296),
.B(n_207),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_262),
.A2(n_221),
.B1(n_232),
.B2(n_205),
.Y(n_297)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_297),
.A2(n_300),
.B1(n_277),
.B2(n_266),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_301),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g302 ( 
.A(n_261),
.B(n_241),
.C(n_227),
.Y(n_302)
);

INVxp67_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g304 ( 
.A(n_273),
.B(n_255),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_305),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_274),
.B(n_242),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g306 ( 
.A1(n_247),
.A2(n_205),
.B1(n_210),
.B2(n_227),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_SL g331 ( 
.A1(n_307),
.A2(n_214),
.B(n_233),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_272),
.B(n_226),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g335 ( 
.A(n_309),
.B(n_311),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_247),
.A2(n_207),
.B1(n_219),
.B2(n_226),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g311 ( 
.A(n_259),
.B(n_182),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_329),
.Y(n_345)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_291),
.Y(n_315)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_315),
.Y(n_350)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_299),
.Y(n_316)
);

NOR2xp33_ASAP7_75t_L g368 ( 
.A(n_316),
.B(n_325),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_318),
.A2(n_339),
.B1(n_342),
.B2(n_284),
.Y(n_344)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_291),
.Y(n_319)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_293),
.B(n_278),
.Y(n_320)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_320),
.Y(n_353)
);

NOR2x1_ASAP7_75t_R g321 ( 
.A(n_284),
.B(n_263),
.Y(n_321)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_321),
.Y(n_365)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_322),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_283),
.A2(n_277),
.B1(n_269),
.B2(n_271),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_L g348 ( 
.A1(n_324),
.A2(n_304),
.B1(n_292),
.B2(n_313),
.Y(n_348)
);

NAND3xp33_ASAP7_75t_L g325 ( 
.A(n_286),
.B(n_248),
.C(n_8),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g327 ( 
.A1(n_298),
.A2(n_276),
.B(n_220),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_L g356 ( 
.A1(n_327),
.A2(n_331),
.B(n_340),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g328 ( 
.A1(n_280),
.A2(n_277),
.B1(n_260),
.B2(n_244),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g361 ( 
.A(n_328),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g329 ( 
.A1(n_300),
.A2(n_260),
.B1(n_214),
.B2(n_219),
.Y(n_329)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_330),
.Y(n_360)
);

AND2x6_ASAP7_75t_L g332 ( 
.A(n_295),
.B(n_178),
.Y(n_332)
);

INVx6_ASAP7_75t_L g358 ( 
.A(n_332),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g336 ( 
.A(n_288),
.B(n_0),
.Y(n_336)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_288),
.Y(n_337)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_337),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_312),
.B(n_193),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g347 ( 
.A(n_338),
.Y(n_347)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_285),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_297),
.A2(n_171),
.B1(n_52),
.B2(n_82),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_290),
.B(n_37),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g354 ( 
.A(n_341),
.B(n_298),
.C(n_281),
.Y(n_354)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_344),
.A2(n_348),
.B1(n_362),
.B2(n_370),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_SL g346 ( 
.A(n_334),
.B(n_323),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g383 ( 
.A(n_346),
.B(n_349),
.Y(n_383)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_334),
.B(n_289),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_317),
.B(n_305),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g384 ( 
.A(n_351),
.B(n_326),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_354),
.B(n_355),
.C(n_364),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_317),
.B(n_309),
.C(n_311),
.Y(n_355)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_333),
.A2(n_343),
.B(n_307),
.Y(n_357)
);

AOI21xp5_ASAP7_75t_L g386 ( 
.A1(n_357),
.A2(n_366),
.B(n_327),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_L g359 ( 
.A1(n_333),
.A2(n_301),
.B(n_282),
.Y(n_359)
);

INVxp67_ASAP7_75t_L g371 ( 
.A(n_359),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_324),
.A2(n_342),
.B1(n_339),
.B2(n_337),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_323),
.B(n_313),
.C(n_294),
.Y(n_364)
);

OAI21xp5_ASAP7_75t_L g366 ( 
.A1(n_331),
.A2(n_294),
.B(n_292),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_315),
.A2(n_296),
.B1(n_302),
.B2(n_308),
.Y(n_370)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_353),
.Y(n_372)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_372),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g373 ( 
.A(n_362),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_SL g401 ( 
.A(n_373),
.B(n_376),
.Y(n_401)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_353),
.Y(n_374)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_374),
.Y(n_409)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_347),
.B(n_314),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_351),
.B(n_335),
.C(n_341),
.Y(n_378)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_378),
.B(n_379),
.C(n_350),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g379 ( 
.A(n_349),
.B(n_335),
.C(n_320),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_361),
.A2(n_344),
.B1(n_358),
.B2(n_368),
.Y(n_380)
);

HB1xp67_ASAP7_75t_L g403 ( 
.A(n_380),
.Y(n_403)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_369),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_382),
.Y(n_402)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_369),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g395 ( 
.A(n_384),
.B(n_388),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_308),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_385),
.A2(n_389),
.B1(n_365),
.B2(n_360),
.Y(n_398)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_386),
.A2(n_392),
.B1(n_367),
.B2(n_365),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g387 ( 
.A(n_364),
.B(n_319),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_387),
.B(n_391),
.Y(n_397)
);

XOR2xp5_ASAP7_75t_L g388 ( 
.A(n_346),
.B(n_332),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_352),
.Y(n_389)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_355),
.B(n_322),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_390),
.B(n_359),
.Y(n_396)
);

XNOR2xp5_ASAP7_75t_L g391 ( 
.A(n_354),
.B(n_370),
.Y(n_391)
);

OA22x2_ASAP7_75t_L g392 ( 
.A1(n_348),
.A2(n_329),
.B1(n_321),
.B2(n_306),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_SL g393 ( 
.A(n_358),
.B(n_343),
.C(n_336),
.Y(n_393)
);

FAx1_ASAP7_75t_SL g404 ( 
.A(n_393),
.B(n_356),
.CI(n_366),
.CON(n_404),
.SN(n_404)
);

XNOR2x1_ASAP7_75t_L g412 ( 
.A(n_394),
.B(n_405),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g425 ( 
.A(n_396),
.B(n_399),
.Y(n_425)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_398),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g399 ( 
.A(n_391),
.B(n_357),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_400),
.B(n_410),
.Y(n_416)
);

NOR2xp33_ASAP7_75t_L g424 ( 
.A(n_404),
.B(n_9),
.Y(n_424)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_375),
.A2(n_367),
.B1(n_371),
.B2(n_374),
.Y(n_405)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_405),
.A2(n_411),
.B1(n_340),
.B2(n_310),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_390),
.B(n_352),
.C(n_363),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g414 ( 
.A(n_407),
.B(n_387),
.Y(n_414)
);

OAI22xp5_ASAP7_75t_L g408 ( 
.A1(n_371),
.A2(n_345),
.B1(n_363),
.B2(n_356),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_408),
.B(n_8),
.Y(n_422)
);

XOR2xp5_ASAP7_75t_L g410 ( 
.A(n_378),
.B(n_345),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_388),
.A2(n_392),
.B1(n_384),
.B2(n_393),
.Y(n_411)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_412),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_400),
.B(n_377),
.C(n_379),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_SL g434 ( 
.A(n_413),
.B(n_414),
.Y(n_434)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_401),
.B(n_377),
.Y(n_415)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_415),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_403),
.A2(n_392),
.B1(n_386),
.B2(n_383),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_418),
.B(n_423),
.Y(n_430)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_397),
.B(n_383),
.C(n_392),
.Y(n_419)
);

NOR2xp67_ASAP7_75t_SL g435 ( 
.A(n_419),
.B(n_396),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g429 ( 
.A1(n_420),
.A2(n_421),
.B1(n_406),
.B2(n_409),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g421 ( 
.A1(n_411),
.A2(n_9),
.B1(n_15),
.B2(n_4),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_422),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_394),
.A2(n_8),
.B1(n_12),
.B2(n_4),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_424),
.A2(n_426),
.B(n_402),
.Y(n_428)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_404),
.A2(n_6),
.B(n_12),
.Y(n_426)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_428),
.B(n_433),
.Y(n_443)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_417),
.B(n_402),
.Y(n_432)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_432),
.Y(n_442)
);

CKINVDCx14_ASAP7_75t_R g433 ( 
.A(n_422),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g446 ( 
.A1(n_435),
.A2(n_407),
.B(n_425),
.Y(n_446)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_423),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g445 ( 
.A(n_437),
.B(n_438),
.Y(n_445)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_418),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_R g439 ( 
.A(n_426),
.B(n_404),
.C(n_399),
.Y(n_439)
);

AOI21xp5_ASAP7_75t_L g444 ( 
.A1(n_439),
.A2(n_419),
.B(n_425),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g441 ( 
.A(n_434),
.B(n_413),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g453 ( 
.A(n_441),
.B(n_449),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_444),
.A2(n_446),
.B(n_450),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_427),
.B(n_416),
.C(n_410),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_447),
.B(n_448),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g448 ( 
.A(n_431),
.B(n_416),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_SL g449 ( 
.A(n_432),
.B(n_397),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_439),
.A2(n_412),
.B(n_395),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_447),
.B(n_444),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_455),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_442),
.B(n_428),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_L g456 ( 
.A1(n_443),
.A2(n_430),
.B(n_436),
.C(n_395),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_456),
.B(n_457),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_440),
.A2(n_421),
.B1(n_430),
.B2(n_429),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g458 ( 
.A(n_445),
.Y(n_458)
);

AOI21xp33_ASAP7_75t_L g461 ( 
.A1(n_458),
.A2(n_450),
.B(n_6),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g459 ( 
.A(n_453),
.Y(n_459)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_459),
.A2(n_37),
.B(n_5),
.Y(n_466)
);

AOI21xp5_ASAP7_75t_L g464 ( 
.A1(n_461),
.A2(n_454),
.B(n_10),
.Y(n_464)
);

O2A1O1Ixp33_ASAP7_75t_SL g463 ( 
.A1(n_453),
.A2(n_4),
.B(n_5),
.C(n_10),
.Y(n_463)
);

OAI321xp33_ASAP7_75t_L g465 ( 
.A1(n_463),
.A2(n_452),
.A3(n_10),
.B1(n_4),
.B2(n_5),
.C(n_11),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_464),
.B(n_466),
.C(n_5),
.Y(n_468)
);

NOR3xp33_ASAP7_75t_L g467 ( 
.A(n_465),
.B(n_460),
.C(n_462),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_467),
.B(n_468),
.C(n_1),
.Y(n_469)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_469),
.A2(n_1),
.B(n_2),
.Y(n_470)
);

AOI21xp5_ASAP7_75t_L g471 ( 
.A1(n_470),
.A2(n_1),
.B(n_37),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_471),
.B(n_1),
.C(n_37),
.Y(n_472)
);


endmodule