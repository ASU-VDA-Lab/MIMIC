module real_aes_12034_n_281 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_254, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_258, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_281);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_281;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_761;
wire n_421;
wire n_329;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_330;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_292;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_553;
wire n_744;
wire n_1367;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_1199;
wire n_951;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_343;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_812;
wire n_817;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_323;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1589;
wire n_947;
wire n_970;
wire n_1149;
wire n_368;
wire n_527;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1346;
wire n_1383;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_1600;
wire n_805;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1583;
wire n_360;
wire n_1284;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_488;
wire n_501;
wire n_1380;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_306;
wire n_1003;
wire n_346;
wire n_293;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_290;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_420;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1495;
wire n_1510;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_724;
wire n_440;
wire n_1231;
wire n_1305;
wire n_315;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_1391;
wire n_375;
wire n_597;
wire n_1036;
wire n_687;
wire n_1538;
wire n_652;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_337;
wire n_1572;
wire n_1514;
wire n_480;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_667;
wire n_991;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1370;
wire n_1417;
wire n_979;
wire n_445;
wire n_596;
wire n_1197;
wire n_657;
wire n_328;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_1014;
wire n_742;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_560;
wire n_1094;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_1269;
wire n_677;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_333;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1479;
wire n_1612;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1070;
wire n_1189;
wire n_535;
wire n_882;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_311;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_602;
wire n_402;
wire n_733;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_286;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1620;
wire n_985;
wire n_777;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_296;
wire n_1347;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_334;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_643;
wire n_1403;
wire n_486;
wire n_291;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_282;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_300;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_313;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_325;
wire n_1298;
wire n_442;
wire n_1633;
wire n_740;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_474;
wire n_1159;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_307;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_285;
wire n_1377;
wire n_800;
wire n_1170;
wire n_778;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_299;
wire n_322;
wire n_900;
wire n_841;
wire n_318;
wire n_1218;
wire n_736;
wire n_766;
wire n_852;
wire n_1268;
wire n_1113;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_594;
wire n_856;
wire n_1146;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_332;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_289;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_356;
wire n_584;
wire n_896;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_284;
wire n_316;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_996;
wire n_523;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1263;
wire n_1411;
wire n_1115;
wire n_310;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_324;
wire n_664;
wire n_367;
wire n_1017;
wire n_936;
wire n_581;
wire n_1215;
wire n_582;
wire n_641;
wire n_940;
wire n_745;
wire n_339;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1603;
wire n_1450;
wire n_714;
wire n_1331;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_288;
wire n_303;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1605;
wire n_1592;
wire n_1056;
wire n_663;
wire n_588;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_295;
wire n_845;
wire n_1619;
wire n_1127;
wire n_484;
wire n_326;
wire n_893;
wire n_1068;
wire n_747;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1355;
wire n_309;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_418;
wire n_771;
wire n_524;
wire n_1378;
wire n_1496;
wire n_705;
wire n_1191;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1617;
wire n_1226;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_929;
wire n_1143;
wire n_1190;
wire n_543;
wire n_305;
wire n_585;
wire n_465;
wire n_719;
wire n_1343;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_1396;
wire n_921;
wire n_1176;
wire n_640;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_1480;
wire n_1101;
wire n_1076;
wire n_1251;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1192;
wire n_1292;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_319;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_376;
wire n_308;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_317;
wire n_1595;
wire n_321;
wire n_666;
wire n_320;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1541;
wire n_1272;
wire n_408;
wire n_372;
wire n_578;
wire n_892;
wire n_938;
wire n_327;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_301;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1257;
wire n_1082;
wire n_1360;
wire n_468;
wire n_532;
wire n_1025;
wire n_298;
wire n_924;
wire n_1264;
wire n_1527;
wire n_297;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_304;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1290;
wire n_1318;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_398;
wire n_1100;
wire n_1519;
wire n_425;
wire n_879;
wire n_1640;
wire n_331;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_302;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1132;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_344;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_336;
wire n_1573;
wire n_1130;
wire n_794;
wire n_283;
wire n_314;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_312;
wire n_1183;
wire n_335;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_1300;
wire n_575;
wire n_338;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_340;
wire n_483;
wire n_1630;
wire n_394;
wire n_729;
wire n_1280;
wire n_1323;
wire n_1352;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_342;
wire n_348;
wire n_1528;
wire n_603;
wire n_1288;
wire n_868;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_429;
AO221x1_ASAP7_75t_L g1299 ( .A1(n_0), .A2(n_169), .B1(n_1300), .B2(n_1306), .C(n_1309), .Y(n_1299) );
CKINVDCx5p33_ASAP7_75t_R g1245 ( .A(n_1), .Y(n_1245) );
AOI21xp33_ASAP7_75t_L g905 ( .A1(n_2), .A2(n_490), .B(n_644), .Y(n_905) );
INVx1_ASAP7_75t_L g925 ( .A(n_2), .Y(n_925) );
INVx1_ASAP7_75t_L g675 ( .A(n_3), .Y(n_675) );
OAI221xp5_ASAP7_75t_L g711 ( .A1(n_3), .A2(n_29), .B1(n_712), .B2(n_713), .C(n_714), .Y(n_711) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_4), .Y(n_295) );
AND2x2_ASAP7_75t_L g384 ( .A(n_4), .B(n_385), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_4), .B(n_213), .Y(n_421) );
INVx1_ASAP7_75t_L g439 ( .A(n_4), .Y(n_439) );
AOI22xp33_ASAP7_75t_L g1194 ( .A1(n_5), .A2(n_19), .B1(n_1141), .B2(n_1195), .Y(n_1194) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_5), .A2(n_215), .B1(n_1153), .B2(n_1224), .Y(n_1223) );
OAI211xp5_ASAP7_75t_L g1236 ( .A1(n_6), .A2(n_1237), .B(n_1238), .C(n_1266), .Y(n_1236) );
AOI22xp5_ASAP7_75t_L g1337 ( .A1(n_7), .A2(n_126), .B1(n_1300), .B2(n_1308), .Y(n_1337) );
OAI221xp5_ASAP7_75t_L g948 ( .A1(n_8), .A2(n_417), .B1(n_606), .B2(n_949), .C(n_955), .Y(n_948) );
INVx1_ASAP7_75t_L g974 ( .A(n_8), .Y(n_974) );
XNOR2x2_ASAP7_75t_L g583 ( .A(n_9), .B(n_584), .Y(n_583) );
CKINVDCx5p33_ASAP7_75t_R g1252 ( .A(n_10), .Y(n_1252) );
AOI221xp5_ASAP7_75t_L g1591 ( .A1(n_11), .A2(n_117), .B1(n_1526), .B2(n_1592), .C(n_1594), .Y(n_1591) );
AOI22xp33_ASAP7_75t_SL g1615 ( .A1(n_11), .A2(n_164), .B1(n_1616), .B2(n_1617), .Y(n_1615) );
AOI221xp5_ASAP7_75t_L g945 ( .A1(n_12), .A2(n_61), .B1(n_435), .B2(n_539), .C(n_946), .Y(n_945) );
INVx1_ASAP7_75t_L g979 ( .A(n_12), .Y(n_979) );
INVx1_ASAP7_75t_L g940 ( .A(n_13), .Y(n_940) );
AOI22xp33_ASAP7_75t_L g976 ( .A1(n_13), .A2(n_62), .B1(n_484), .B2(n_798), .Y(n_976) );
INVx1_ASAP7_75t_L g780 ( .A(n_14), .Y(n_780) );
AO22x2_ASAP7_75t_L g984 ( .A1(n_15), .A2(n_985), .B1(n_1041), .B2(n_1042), .Y(n_984) );
CKINVDCx14_ASAP7_75t_R g1041 ( .A(n_15), .Y(n_1041) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_16), .A2(n_92), .B1(n_342), .B2(n_344), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g451 ( .A1(n_16), .A2(n_30), .B1(n_383), .B2(n_419), .Y(n_451) );
AOI22xp33_ASAP7_75t_SL g682 ( .A1(n_17), .A2(n_242), .B1(n_452), .B2(n_683), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_17), .A2(n_76), .B1(n_489), .B2(n_724), .C(n_725), .Y(n_723) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_18), .A2(n_76), .B1(n_686), .B2(n_688), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_18), .A2(n_242), .B1(n_493), .B2(n_514), .Y(n_726) );
AOI221xp5_ASAP7_75t_L g1219 ( .A1(n_19), .A2(n_99), .B1(n_1033), .B2(n_1220), .C(n_1221), .Y(n_1219) );
AO221x2_ASAP7_75t_L g1390 ( .A1(n_20), .A2(n_189), .B1(n_1306), .B2(n_1391), .C(n_1393), .Y(n_1390) );
AOI221xp5_ASAP7_75t_L g487 ( .A1(n_21), .A2(n_239), .B1(n_488), .B2(n_489), .C(n_490), .Y(n_487) );
INVx1_ASAP7_75t_L g541 ( .A(n_21), .Y(n_541) );
OAI221xp5_ASAP7_75t_L g884 ( .A1(n_22), .A2(n_830), .B1(n_885), .B2(n_890), .C(n_896), .Y(n_884) );
AOI22xp33_ASAP7_75t_L g919 ( .A1(n_22), .A2(n_191), .B1(n_431), .B2(n_920), .Y(n_919) );
CKINVDCx5p33_ASAP7_75t_R g956 ( .A(n_23), .Y(n_956) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_24), .A2(n_162), .B1(n_429), .B2(n_431), .C(n_435), .Y(n_428) );
OAI22xp5_ASAP7_75t_L g470 ( .A1(n_24), .A2(n_238), .B1(n_471), .B2(n_472), .Y(n_470) );
INVx2_ASAP7_75t_L g320 ( .A(n_25), .Y(n_320) );
OR2x2_ASAP7_75t_L g466 ( .A(n_25), .B(n_365), .Y(n_466) );
AO22x1_ASAP7_75t_L g935 ( .A1(n_26), .A2(n_936), .B1(n_982), .B2(n_983), .Y(n_935) );
INVx1_ASAP7_75t_L g983 ( .A(n_26), .Y(n_983) );
AOI22xp33_ASAP7_75t_L g321 ( .A1(n_27), .A2(n_66), .B1(n_322), .B2(n_327), .Y(n_321) );
INVx1_ASAP7_75t_L g416 ( .A(n_27), .Y(n_416) );
OAI22xp5_ASAP7_75t_L g841 ( .A1(n_28), .A2(n_250), .B1(n_713), .B2(n_842), .Y(n_841) );
OAI221xp5_ASAP7_75t_L g857 ( .A1(n_28), .A2(n_250), .B1(n_551), .B2(n_858), .C(n_859), .Y(n_857) );
INVx1_ASAP7_75t_L g671 ( .A(n_29), .Y(n_671) );
OAI222xp33_ASAP7_75t_L g455 ( .A1(n_30), .A2(n_162), .B1(n_167), .B2(n_456), .C1(n_459), .C2(n_467), .Y(n_455) );
BUFx2_ASAP7_75t_L g316 ( .A(n_31), .Y(n_316) );
BUFx2_ASAP7_75t_L g352 ( .A(n_31), .Y(n_352) );
INVx1_ASAP7_75t_L g367 ( .A(n_31), .Y(n_367) );
OR2x2_ASAP7_75t_L g529 ( .A(n_31), .B(n_421), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g1198 ( .A1(n_32), .A2(n_163), .B1(n_1197), .B2(n_1199), .Y(n_1198) );
INVxp33_ASAP7_75t_SL g1228 ( .A(n_32), .Y(n_1228) );
OAI221xp5_ASAP7_75t_L g1246 ( .A1(n_33), .A2(n_228), .B1(n_756), .B2(n_757), .C(n_858), .Y(n_1246) );
INVx1_ASAP7_75t_L g1279 ( .A(n_33), .Y(n_1279) );
AOI221xp5_ASAP7_75t_L g1525 ( .A1(n_34), .A2(n_111), .B1(n_719), .B2(n_1526), .C(n_1527), .Y(n_1525) );
INVx1_ASAP7_75t_L g1552 ( .A(n_34), .Y(n_1552) );
OAI22xp33_ASAP7_75t_L g1072 ( .A1(n_35), .A2(n_180), .B1(n_653), .B2(n_655), .Y(n_1072) );
INVx1_ASAP7_75t_L g1104 ( .A(n_35), .Y(n_1104) );
INVx1_ASAP7_75t_L g988 ( .A(n_36), .Y(n_988) );
AOI21xp33_ASAP7_75t_L g1032 ( .A1(n_36), .A2(n_484), .B(n_1033), .Y(n_1032) );
INVxp33_ASAP7_75t_SL g1190 ( .A(n_37), .Y(n_1190) );
AOI221xp5_ASAP7_75t_L g1210 ( .A1(n_37), .A2(n_225), .B1(n_1211), .B2(n_1212), .C(n_1213), .Y(n_1210) );
CKINVDCx5p33_ASAP7_75t_R g1000 ( .A(n_38), .Y(n_1000) );
AOI221xp5_ASAP7_75t_L g1535 ( .A1(n_39), .A2(n_170), .B1(n_511), .B2(n_1536), .C(n_1538), .Y(n_1535) );
INVx1_ASAP7_75t_L g1561 ( .A(n_39), .Y(n_1561) );
OAI22xp5_ASAP7_75t_L g497 ( .A1(n_40), .A2(n_75), .B1(n_498), .B2(n_500), .Y(n_497) );
OAI221xp5_ASAP7_75t_L g547 ( .A1(n_40), .A2(n_75), .B1(n_548), .B2(n_551), .C(n_554), .Y(n_547) );
AOI22xp33_ASAP7_75t_L g904 ( .A1(n_41), .A2(n_150), .B1(n_484), .B2(n_798), .Y(n_904) );
INVx1_ASAP7_75t_L g926 ( .A(n_41), .Y(n_926) );
INVx1_ASAP7_75t_L g783 ( .A(n_42), .Y(n_783) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_43), .A2(n_221), .B1(n_342), .B2(n_834), .Y(n_833) );
INVx1_ASAP7_75t_L g864 ( .A(n_43), .Y(n_864) );
OAI221xp5_ASAP7_75t_L g1034 ( .A1(n_44), .A2(n_233), .B1(n_794), .B2(n_1035), .C(n_1036), .Y(n_1034) );
INVx1_ASAP7_75t_L g1039 ( .A(n_44), .Y(n_1039) );
AOI22xp33_ASAP7_75t_SL g1134 ( .A1(n_45), .A2(n_112), .B1(n_1135), .B2(n_1136), .Y(n_1134) );
AOI221xp5_ASAP7_75t_L g1157 ( .A1(n_45), .A2(n_74), .B1(n_811), .B2(n_1158), .C(n_1160), .Y(n_1157) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_46), .A2(n_57), .B1(n_692), .B2(n_694), .Y(n_691) );
INVx1_ASAP7_75t_L g728 ( .A(n_46), .Y(n_728) );
INVx1_ASAP7_75t_L g954 ( .A(n_47), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g969 ( .A1(n_47), .A2(n_155), .B1(n_798), .B2(n_895), .Y(n_969) );
OAI22xp5_ASAP7_75t_L g947 ( .A1(n_48), .A2(n_171), .B1(n_443), .B2(n_448), .Y(n_947) );
OAI22xp5_ASAP7_75t_SL g966 ( .A1(n_48), .A2(n_171), .B1(n_357), .B2(n_370), .Y(n_966) );
AOI22xp33_ASAP7_75t_L g589 ( .A1(n_49), .A2(n_54), .B1(n_590), .B2(n_592), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g664 ( .A1(n_49), .A2(n_73), .B1(n_471), .B2(n_472), .Y(n_664) );
CKINVDCx5p33_ASAP7_75t_R g1531 ( .A(n_50), .Y(n_1531) );
INVx1_ASAP7_75t_L g374 ( .A(n_51), .Y(n_374) );
OAI221xp5_ASAP7_75t_L g442 ( .A1(n_51), .A2(n_93), .B1(n_443), .B2(n_448), .C(n_450), .Y(n_442) );
OAI22xp5_ASAP7_75t_L g1235 ( .A1(n_52), .A2(n_1236), .B1(n_1290), .B2(n_1291), .Y(n_1235) );
INVx1_ASAP7_75t_L g1291 ( .A(n_52), .Y(n_1291) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_53), .A2(n_83), .B1(n_349), .B2(n_1070), .Y(n_1069) );
OAI22xp5_ASAP7_75t_L g1074 ( .A1(n_53), .A2(n_83), .B1(n_1075), .B2(n_1076), .Y(n_1074) );
INVxp67_ASAP7_75t_SL g661 ( .A(n_54), .Y(n_661) );
INVxp67_ASAP7_75t_SL g1600 ( .A(n_55), .Y(n_1600) );
AOI221xp5_ASAP7_75t_L g1628 ( .A1(n_55), .A2(n_108), .B1(n_1136), .B2(n_1629), .C(n_1630), .Y(n_1628) );
INVxp67_ASAP7_75t_SL g1604 ( .A(n_56), .Y(n_1604) );
OAI211xp5_ASAP7_75t_SL g1620 ( .A1(n_56), .A2(n_562), .B(n_1621), .C(n_1622), .Y(n_1620) );
INVx1_ASAP7_75t_L g722 ( .A(n_57), .Y(n_722) );
INVx1_ASAP7_75t_L g1607 ( .A(n_58), .Y(n_1607) );
OAI22xp33_ASAP7_75t_L g906 ( .A1(n_59), .A2(n_191), .B1(n_521), .B2(n_524), .Y(n_906) );
AOI22xp33_ASAP7_75t_L g917 ( .A1(n_59), .A2(n_274), .B1(n_914), .B2(n_918), .Y(n_917) );
INVx1_ASAP7_75t_L g614 ( .A(n_60), .Y(n_614) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_61), .A2(n_118), .B1(n_472), .B2(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g941 ( .A(n_62), .Y(n_941) );
AOI221xp5_ASAP7_75t_L g832 ( .A1(n_63), .A2(n_77), .B1(n_489), .B2(n_511), .C(n_724), .Y(n_832) );
INVxp67_ASAP7_75t_SL g867 ( .A(n_63), .Y(n_867) );
INVx1_ASAP7_75t_L g750 ( .A(n_64), .Y(n_750) );
AOI22xp33_ASAP7_75t_L g1058 ( .A1(n_65), .A2(n_151), .B1(n_1059), .B2(n_1060), .Y(n_1058) );
INVxp67_ASAP7_75t_SL g1084 ( .A(n_65), .Y(n_1084) );
INVx1_ASAP7_75t_L g414 ( .A(n_66), .Y(n_414) );
OAI221xp5_ASAP7_75t_L g753 ( .A1(n_67), .A2(n_229), .B1(n_754), .B2(n_756), .C(n_757), .Y(n_753) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_67), .A2(n_229), .B1(n_792), .B2(n_794), .Y(n_791) );
INVxp67_ASAP7_75t_L g771 ( .A(n_68), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_68), .A2(n_128), .B1(n_813), .B2(n_814), .Y(n_812) );
INVx1_ASAP7_75t_L g1244 ( .A(n_69), .Y(n_1244) );
AOI221xp5_ASAP7_75t_L g1285 ( .A1(n_69), .A2(n_142), .B1(n_1162), .B2(n_1286), .C(n_1288), .Y(n_1285) );
AOI22xp33_ASAP7_75t_SL g1589 ( .A1(n_70), .A2(n_164), .B1(n_1527), .B2(n_1590), .Y(n_1589) );
AOI22xp33_ASAP7_75t_L g1618 ( .A1(n_70), .A2(n_117), .B1(n_452), .B2(n_1619), .Y(n_1618) );
INVx1_ASAP7_75t_L g1315 ( .A(n_71), .Y(n_1315) );
AOI22xp33_ASAP7_75t_L g1528 ( .A1(n_72), .A2(n_195), .B1(n_1212), .B2(n_1529), .Y(n_1528) );
INVx1_ASAP7_75t_L g1550 ( .A(n_72), .Y(n_1550) );
AOI221xp5_ASAP7_75t_L g595 ( .A1(n_73), .A2(n_201), .B1(n_435), .B2(n_596), .C(n_598), .Y(n_595) );
AOI22xp33_ASAP7_75t_L g1131 ( .A1(n_74), .A2(n_138), .B1(n_1132), .B2(n_1133), .Y(n_1131) );
INVxp67_ASAP7_75t_SL g871 ( .A(n_77), .Y(n_871) );
AOI22xp33_ASAP7_75t_L g513 ( .A1(n_78), .A2(n_267), .B1(n_514), .B2(n_515), .Y(n_513) );
INVx1_ASAP7_75t_L g561 ( .A(n_78), .Y(n_561) );
AOI22xp33_ASAP7_75t_L g1595 ( .A1(n_79), .A2(n_103), .B1(n_1212), .B2(n_1590), .Y(n_1595) );
INVxp67_ASAP7_75t_SL g1634 ( .A(n_79), .Y(n_1634) );
INVx1_ASAP7_75t_L g1261 ( .A(n_80), .Y(n_1261) );
OAI22xp5_ASAP7_75t_L g1289 ( .A1(n_80), .A2(n_251), .B1(n_521), .B2(n_524), .Y(n_1289) );
AOI22xp33_ASAP7_75t_SL g1140 ( .A1(n_81), .A2(n_95), .B1(n_1094), .B2(n_1141), .Y(n_1140) );
INVx1_ASAP7_75t_L g1156 ( .A(n_81), .Y(n_1156) );
AOI221xp5_ASAP7_75t_L g1596 ( .A1(n_82), .A2(n_165), .B1(n_719), .B2(n_1527), .C(n_1597), .Y(n_1596) );
INVxp33_ASAP7_75t_SL g1625 ( .A(n_82), .Y(n_1625) );
AO221x1_ASAP7_75t_L g1344 ( .A1(n_84), .A2(n_137), .B1(n_1300), .B2(n_1308), .C(n_1345), .Y(n_1344) );
INVx1_ASAP7_75t_L g1395 ( .A(n_85), .Y(n_1395) );
INVx1_ASAP7_75t_L g1126 ( .A(n_86), .Y(n_1126) );
AOI221xp5_ASAP7_75t_L g1151 ( .A1(n_86), .A2(n_106), .B1(n_1152), .B2(n_1153), .C(n_1154), .Y(n_1151) );
CKINVDCx5p33_ASAP7_75t_R g1541 ( .A(n_87), .Y(n_1541) );
AO221x1_ASAP7_75t_L g1340 ( .A1(n_88), .A2(n_185), .B1(n_1300), .B2(n_1308), .C(n_1341), .Y(n_1340) );
AOI22xp33_ASAP7_75t_L g1138 ( .A1(n_89), .A2(n_226), .B1(n_1136), .B2(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1168 ( .A(n_89), .Y(n_1168) );
INVx1_ASAP7_75t_L g319 ( .A(n_90), .Y(n_319) );
INVx1_ASAP7_75t_L g365 ( .A(n_90), .Y(n_365) );
INVx1_ASAP7_75t_L g827 ( .A(n_91), .Y(n_827) );
INVx1_ASAP7_75t_L g441 ( .A(n_92), .Y(n_441) );
INVx1_ASAP7_75t_L g368 ( .A(n_93), .Y(n_368) );
INVx1_ASAP7_75t_L g1065 ( .A(n_94), .Y(n_1065) );
OAI221xp5_ASAP7_75t_L g1077 ( .A1(n_94), .A2(n_606), .B1(n_619), .B2(n_1078), .C(n_1081), .Y(n_1077) );
INVx1_ASAP7_75t_L g1167 ( .A(n_95), .Y(n_1167) );
INVx1_ASAP7_75t_L g1342 ( .A(n_96), .Y(n_1342) );
INVx1_ASAP7_75t_L g891 ( .A(n_97), .Y(n_891) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_97), .A2(n_168), .B1(n_431), .B2(n_912), .Y(n_911) );
INVx1_ASAP7_75t_L g1092 ( .A(n_98), .Y(n_1092) );
OAI22xp5_ASAP7_75t_L g1106 ( .A1(n_98), .A2(n_123), .B1(n_472), .B2(n_981), .Y(n_1106) );
AOI22xp33_ASAP7_75t_SL g1196 ( .A1(n_99), .A2(n_215), .B1(n_1132), .B2(n_1197), .Y(n_1196) );
INVx1_ASAP7_75t_L g1111 ( .A(n_100), .Y(n_1111) );
INVx1_ASAP7_75t_L g617 ( .A(n_101), .Y(n_617) );
AOI221xp5_ASAP7_75t_L g629 ( .A1(n_101), .A2(n_270), .B1(n_630), .B2(n_633), .C(n_635), .Y(n_629) );
INVxp67_ASAP7_75t_L g765 ( .A(n_102), .Y(n_765) );
AOI221xp5_ASAP7_75t_L g806 ( .A1(n_102), .A2(n_125), .B1(n_807), .B2(n_809), .C(n_811), .Y(n_806) );
INVxp33_ASAP7_75t_L g1626 ( .A(n_103), .Y(n_1626) );
OAI22xp5_ASAP7_75t_L g880 ( .A1(n_104), .A2(n_881), .B1(n_930), .B2(n_931), .Y(n_880) );
INVxp67_ASAP7_75t_SL g930 ( .A(n_104), .Y(n_930) );
OAI22xp5_ASAP7_75t_L g1175 ( .A1(n_105), .A2(n_1176), .B1(n_1177), .B2(n_1230), .Y(n_1175) );
INVx1_ASAP7_75t_L g1230 ( .A(n_105), .Y(n_1230) );
INVx1_ASAP7_75t_L g1121 ( .A(n_106), .Y(n_1121) );
AOI22xp33_ASAP7_75t_SL g332 ( .A1(n_107), .A2(n_174), .B1(n_333), .B2(n_338), .Y(n_332) );
AOI21xp33_ASAP7_75t_L g404 ( .A1(n_107), .A2(n_405), .B(n_408), .Y(n_404) );
OAI211xp5_ASAP7_75t_SL g1587 ( .A1(n_108), .A2(n_524), .B(n_1588), .C(n_1598), .Y(n_1587) );
CKINVDCx5p33_ASAP7_75t_R g1204 ( .A(n_109), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_110), .A2(n_232), .B1(n_1300), .B2(n_1308), .Y(n_1355) );
INVx1_ASAP7_75t_L g1554 ( .A(n_111), .Y(n_1554) );
AOI22xp33_ASAP7_75t_L g1161 ( .A1(n_112), .A2(n_138), .B1(n_1162), .B2(n_1165), .Y(n_1161) );
INVx1_ASAP7_75t_L g1265 ( .A(n_113), .Y(n_1265) );
OAI211xp5_ASAP7_75t_SL g1267 ( .A1(n_113), .A2(n_1268), .B(n_1269), .C(n_1275), .Y(n_1267) );
INVx1_ASAP7_75t_L g1189 ( .A(n_114), .Y(n_1189) );
AOI221xp5_ASAP7_75t_L g1093 ( .A1(n_115), .A2(n_123), .B1(n_1094), .B2(n_1096), .C(n_1098), .Y(n_1093) );
OAI22xp5_ASAP7_75t_L g1107 ( .A1(n_115), .A2(n_208), .B1(n_459), .B2(n_467), .Y(n_1107) );
AOI22xp33_ASAP7_75t_L g838 ( .A1(n_116), .A2(n_243), .B1(n_839), .B2(n_840), .Y(n_838) );
INVx1_ASAP7_75t_L g855 ( .A(n_116), .Y(n_855) );
AOI22xp33_ASAP7_75t_L g943 ( .A1(n_118), .A2(n_134), .B1(n_425), .B2(n_944), .Y(n_943) );
AOI22xp33_ASAP7_75t_SL g1201 ( .A1(n_119), .A2(n_139), .B1(n_683), .B2(n_1141), .Y(n_1201) );
INVxp33_ASAP7_75t_L g1227 ( .A(n_119), .Y(n_1227) );
INVxp33_ASAP7_75t_L g746 ( .A(n_120), .Y(n_746) );
AOI221xp5_ASAP7_75t_L g796 ( .A1(n_120), .A2(n_154), .B1(n_797), .B2(n_799), .C(n_801), .Y(n_796) );
AOI221xp5_ASAP7_75t_L g837 ( .A1(n_121), .A2(n_227), .B1(n_489), .B2(n_490), .C(n_644), .Y(n_837) );
INVx1_ASAP7_75t_L g854 ( .A(n_121), .Y(n_854) );
INVx1_ASAP7_75t_L g1347 ( .A(n_122), .Y(n_1347) );
INVx1_ASAP7_75t_L g287 ( .A(n_124), .Y(n_287) );
INVxp67_ASAP7_75t_L g768 ( .A(n_125), .Y(n_768) );
CKINVDCx5p33_ASAP7_75t_R g522 ( .A(n_127), .Y(n_522) );
INVx1_ASAP7_75t_L g762 ( .A(n_128), .Y(n_762) );
INVx1_ASAP7_75t_L g580 ( .A(n_129), .Y(n_580) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_130), .A2(n_202), .B1(n_590), .B2(n_690), .Y(n_689) );
INVx1_ASAP7_75t_L g729 ( .A(n_130), .Y(n_729) );
CKINVDCx5p33_ASAP7_75t_R g997 ( .A(n_131), .Y(n_997) );
INVxp67_ASAP7_75t_SL g1182 ( .A(n_132), .Y(n_1182) );
OAI22xp5_ASAP7_75t_L g1208 ( .A1(n_132), .A2(n_280), .B1(n_1148), .B2(n_1209), .Y(n_1208) );
AOI22xp33_ASAP7_75t_L g491 ( .A1(n_133), .A2(n_204), .B1(n_492), .B2(n_493), .Y(n_491) );
INVx1_ASAP7_75t_L g533 ( .A(n_133), .Y(n_533) );
INVx1_ASAP7_75t_L g978 ( .A(n_134), .Y(n_978) );
AOI22xp5_ASAP7_75t_L g1332 ( .A1(n_135), .A2(n_216), .B1(n_1324), .B2(n_1327), .Y(n_1332) );
INVx1_ASAP7_75t_L g748 ( .A(n_136), .Y(n_748) );
INVxp67_ASAP7_75t_SL g1225 ( .A(n_139), .Y(n_1225) );
AOI22xp5_ASAP7_75t_L g1333 ( .A1(n_140), .A2(n_192), .B1(n_1300), .B2(n_1308), .Y(n_1333) );
AOI22xp5_ASAP7_75t_L g1356 ( .A1(n_141), .A2(n_279), .B1(n_1324), .B2(n_1327), .Y(n_1356) );
INVx1_ASAP7_75t_L g1242 ( .A(n_142), .Y(n_1242) );
INVx1_ASAP7_75t_L g622 ( .A(n_143), .Y(n_622) );
INVx1_ASAP7_75t_L g1187 ( .A(n_144), .Y(n_1187) );
CKINVDCx5p33_ASAP7_75t_R g699 ( .A(n_145), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g1003 ( .A(n_146), .Y(n_1003) );
INVx1_ASAP7_75t_L g731 ( .A(n_147), .Y(n_731) );
XNOR2xp5_ASAP7_75t_L g309 ( .A(n_148), .B(n_310), .Y(n_309) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_149), .Y(n_900) );
OAI22xp5_ASAP7_75t_L g927 ( .A1(n_150), .A2(n_260), .B1(n_928), .B2(n_929), .Y(n_927) );
INVxp67_ASAP7_75t_SL g1088 ( .A(n_151), .Y(n_1088) );
INVx1_ASAP7_75t_L g1143 ( .A(n_152), .Y(n_1143) );
CKINVDCx5p33_ASAP7_75t_R g519 ( .A(n_153), .Y(n_519) );
INVxp33_ASAP7_75t_L g751 ( .A(n_154), .Y(n_751) );
INVx1_ASAP7_75t_L g952 ( .A(n_155), .Y(n_952) );
INVx1_ASAP7_75t_L g697 ( .A(n_156), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g716 ( .A1(n_156), .A2(n_240), .B1(n_324), .B2(n_328), .Y(n_716) );
INVx1_ASAP7_75t_L g1068 ( .A(n_157), .Y(n_1068) );
OAI211xp5_ASAP7_75t_SL g1089 ( .A1(n_157), .A2(n_587), .B(n_1090), .C(n_1099), .Y(n_1089) );
INVx1_ASAP7_75t_L g989 ( .A(n_158), .Y(n_989) );
AOI22xp33_ASAP7_75t_SL g1030 ( .A1(n_158), .A2(n_206), .B1(n_798), .B2(n_1031), .Y(n_1030) );
CKINVDCx5p33_ASAP7_75t_R g1125 ( .A(n_159), .Y(n_1125) );
OAI22xp5_ASAP7_75t_L g601 ( .A1(n_160), .A2(n_186), .B1(n_443), .B2(n_448), .Y(n_601) );
OAI221xp5_ASAP7_75t_L g652 ( .A1(n_160), .A2(n_186), .B1(n_653), .B2(n_655), .C(n_656), .Y(n_652) );
CKINVDCx5p33_ASAP7_75t_R g506 ( .A(n_161), .Y(n_506) );
INVxp67_ASAP7_75t_SL g1207 ( .A(n_163), .Y(n_1207) );
OAI21xp33_ASAP7_75t_SL g1612 ( .A1(n_165), .A2(n_1613), .B(n_1614), .Y(n_1612) );
INVx1_ASAP7_75t_L g831 ( .A(n_166), .Y(n_831) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_167), .A2(n_238), .B1(n_424), .B2(n_425), .Y(n_423) );
INVx1_ASAP7_75t_L g887 ( .A(n_168), .Y(n_887) );
INVx1_ASAP7_75t_L g1563 ( .A(n_170), .Y(n_1563) );
AOI22xp33_ASAP7_75t_SL g347 ( .A1(n_172), .A2(n_181), .B1(n_348), .B2(n_349), .Y(n_347) );
INVx1_ASAP7_75t_L g390 ( .A(n_172), .Y(n_390) );
INVxp67_ASAP7_75t_SL g1256 ( .A(n_173), .Y(n_1256) );
AOI221xp5_ASAP7_75t_L g1273 ( .A1(n_173), .A2(n_205), .B1(n_1220), .B2(n_1221), .C(n_1274), .Y(n_1273) );
INVx1_ASAP7_75t_L g403 ( .A(n_174), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g1012 ( .A1(n_175), .A2(n_231), .B1(n_528), .B2(n_928), .Y(n_1012) );
AOI22xp33_ASAP7_75t_SL g1025 ( .A1(n_175), .A2(n_200), .B1(n_484), .B2(n_798), .Y(n_1025) );
AOI221xp5_ASAP7_75t_L g507 ( .A1(n_176), .A2(n_241), .B1(n_508), .B2(n_510), .C(n_511), .Y(n_507) );
INVx1_ASAP7_75t_L g570 ( .A(n_176), .Y(n_570) );
AOI21xp33_ASAP7_75t_L g894 ( .A1(n_177), .A2(n_811), .B(n_895), .Y(n_894) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_177), .A2(n_259), .B1(n_914), .B2(n_915), .Y(n_913) );
OAI22xp5_ASAP7_75t_L g1009 ( .A1(n_178), .A2(n_200), .B1(n_1010), .B2(n_1011), .Y(n_1009) );
INVx1_ASAP7_75t_L g1021 ( .A(n_178), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g1047 ( .A(n_179), .Y(n_1047) );
INVx1_ASAP7_75t_L g1102 ( .A(n_180), .Y(n_1102) );
INVx1_ASAP7_75t_L g396 ( .A(n_181), .Y(n_396) );
HB1xp67_ASAP7_75t_L g289 ( .A(n_182), .Y(n_289) );
AND3x2_ASAP7_75t_L g1304 ( .A(n_182), .B(n_287), .C(n_1305), .Y(n_1304) );
NAND2xp5_ASAP7_75t_L g1312 ( .A(n_182), .B(n_287), .Y(n_1312) );
CKINVDCx5p33_ASAP7_75t_R g998 ( .A(n_183), .Y(n_998) );
OA332x1_ASAP7_75t_L g986 ( .A1(n_184), .A2(n_556), .A3(n_987), .B1(n_992), .B2(n_996), .B3(n_999), .C1(n_1005), .C2(n_1006), .Y(n_986) );
AOI21xp5_ASAP7_75t_L g1026 ( .A1(n_184), .A2(n_490), .B(n_1027), .Y(n_1026) );
INVx2_ASAP7_75t_L g300 ( .A(n_187), .Y(n_300) );
INVx1_ASAP7_75t_L g844 ( .A(n_188), .Y(n_844) );
INVx1_ASAP7_75t_L g776 ( .A(n_190), .Y(n_776) );
OAI211xp5_ASAP7_75t_L g938 ( .A1(n_193), .A2(n_587), .B(n_939), .C(n_942), .Y(n_938) );
INVx1_ASAP7_75t_L g975 ( .A(n_193), .Y(n_975) );
AOI22xp33_ASAP7_75t_L g1540 ( .A1(n_194), .A2(n_236), .B1(n_327), .B2(n_813), .Y(n_1540) );
INVx1_ASAP7_75t_L g1559 ( .A(n_194), .Y(n_1559) );
INVx1_ASAP7_75t_L g1555 ( .A(n_195), .Y(n_1555) );
INVx1_ASAP7_75t_L g1346 ( .A(n_196), .Y(n_1346) );
CKINVDCx5p33_ASAP7_75t_R g899 ( .A(n_197), .Y(n_899) );
INVx1_ASAP7_75t_L g612 ( .A(n_198), .Y(n_612) );
INVx1_ASAP7_75t_L g1305 ( .A(n_199), .Y(n_1305) );
INVxp67_ASAP7_75t_SL g663 ( .A(n_201), .Y(n_663) );
INVx1_ASAP7_75t_L g710 ( .A(n_202), .Y(n_710) );
OAI211xp5_ASAP7_75t_SL g1601 ( .A1(n_203), .A2(n_1602), .B(n_1603), .C(n_1609), .Y(n_1601) );
INVx1_ASAP7_75t_L g1632 ( .A(n_203), .Y(n_1632) );
INVx1_ASAP7_75t_L g544 ( .A(n_204), .Y(n_544) );
INVxp67_ASAP7_75t_SL g1251 ( .A(n_205), .Y(n_1251) );
INVx1_ASAP7_75t_L g993 ( .A(n_206), .Y(n_993) );
CKINVDCx5p33_ASAP7_75t_R g730 ( .A(n_207), .Y(n_730) );
INVx1_ASAP7_75t_L g1091 ( .A(n_208), .Y(n_1091) );
OAI211xp5_ASAP7_75t_L g586 ( .A1(n_209), .A2(n_587), .B(n_588), .C(n_602), .Y(n_586) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_209), .A2(n_219), .B1(n_641), .B2(n_643), .C(n_646), .Y(n_640) );
OAI22xp33_ASAP7_75t_L g1532 ( .A1(n_210), .A2(n_212), .B1(n_794), .B2(n_1533), .Y(n_1532) );
OAI221xp5_ASAP7_75t_L g1556 ( .A1(n_210), .A2(n_212), .B1(n_754), .B2(n_756), .C(n_757), .Y(n_1556) );
CKINVDCx5p33_ASAP7_75t_R g486 ( .A(n_211), .Y(n_486) );
INVx1_ASAP7_75t_L g302 ( .A(n_213), .Y(n_302) );
INVx2_ASAP7_75t_L g385 ( .A(n_213), .Y(n_385) );
INVx1_ASAP7_75t_L g603 ( .A(n_214), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g1336 ( .A1(n_217), .A2(n_235), .B1(n_1324), .B2(n_1327), .Y(n_1336) );
INVx1_ASAP7_75t_L g774 ( .A(n_218), .Y(n_774) );
OAI221xp5_ASAP7_75t_L g605 ( .A1(n_219), .A2(n_606), .B1(n_608), .B2(n_615), .C(n_619), .Y(n_605) );
OR2x2_ASAP7_75t_L g882 ( .A(n_220), .B(n_527), .Y(n_882) );
INVx1_ASAP7_75t_L g872 ( .A(n_221), .Y(n_872) );
INVx1_ASAP7_75t_L g964 ( .A(n_222), .Y(n_964) );
OAI22xp5_ASAP7_75t_L g821 ( .A1(n_223), .A2(n_822), .B1(n_878), .B2(n_879), .Y(n_821) );
INVx1_ASAP7_75t_L g879 ( .A(n_223), .Y(n_879) );
INVx1_ASAP7_75t_L g701 ( .A(n_224), .Y(n_701) );
AOI21xp33_ASAP7_75t_L g717 ( .A1(n_224), .A2(n_718), .B(n_719), .Y(n_717) );
INVxp33_ASAP7_75t_SL g1186 ( .A(n_225), .Y(n_1186) );
INVx1_ASAP7_75t_L g1146 ( .A(n_226), .Y(n_1146) );
INVx1_ASAP7_75t_L g851 ( .A(n_227), .Y(n_851) );
INVx1_ASAP7_75t_L g1281 ( .A(n_228), .Y(n_1281) );
XNOR2xp5_ASAP7_75t_L g1518 ( .A(n_230), .B(n_1519), .Y(n_1518) );
INVx1_ASAP7_75t_L g1037 ( .A(n_231), .Y(n_1037) );
INVx1_ASAP7_75t_L g1040 ( .A(n_233), .Y(n_1040) );
INVx1_ASAP7_75t_L g1254 ( .A(n_234), .Y(n_1254) );
INVx1_ASAP7_75t_L g1564 ( .A(n_236), .Y(n_1564) );
INVx1_ASAP7_75t_L g1545 ( .A(n_237), .Y(n_1545) );
INVx1_ASAP7_75t_L g537 ( .A(n_239), .Y(n_537) );
INVx1_ASAP7_75t_L g702 ( .A(n_240), .Y(n_702) );
INVx1_ASAP7_75t_L g566 ( .A(n_241), .Y(n_566) );
INVx1_ASAP7_75t_L g849 ( .A(n_243), .Y(n_849) );
INVx1_ASAP7_75t_L g1258 ( .A(n_244), .Y(n_1258) );
OAI211xp5_ASAP7_75t_L g1276 ( .A1(n_244), .A2(n_1277), .B(n_1278), .C(n_1282), .Y(n_1276) );
INVx1_ASAP7_75t_L g1303 ( .A(n_245), .Y(n_1303) );
NAND2xp5_ASAP7_75t_L g1318 ( .A(n_245), .B(n_1314), .Y(n_1318) );
INVx1_ASAP7_75t_L g836 ( .A(n_246), .Y(n_836) );
INVx1_ASAP7_75t_L g1044 ( .A(n_247), .Y(n_1044) );
CKINVDCx5p33_ASAP7_75t_R g788 ( .A(n_248), .Y(n_788) );
INVx1_ASAP7_75t_L g1119 ( .A(n_249), .Y(n_1119) );
OAI22xp5_ASAP7_75t_L g1147 ( .A1(n_249), .A2(n_262), .B1(n_1148), .B2(n_1149), .Y(n_1147) );
INVx1_ASAP7_75t_L g1263 ( .A(n_251), .Y(n_1263) );
INVx1_ASAP7_75t_L g1608 ( .A(n_252), .Y(n_1608) );
INVx1_ASAP7_75t_L g819 ( .A(n_253), .Y(n_819) );
AO22x1_ASAP7_75t_L g1321 ( .A1(n_254), .A2(n_266), .B1(n_1308), .B2(n_1322), .Y(n_1321) );
AOI22xp33_ASAP7_75t_L g1577 ( .A1(n_254), .A2(n_1578), .B1(n_1583), .B2(n_1637), .Y(n_1577) );
AOI22x1_ASAP7_75t_L g1584 ( .A1(n_254), .A2(n_1585), .B1(n_1635), .B2(n_1636), .Y(n_1584) );
INVxp67_ASAP7_75t_L g1635 ( .A(n_254), .Y(n_1635) );
CKINVDCx5p33_ASAP7_75t_R g1544 ( .A(n_255), .Y(n_1544) );
CKINVDCx5p33_ASAP7_75t_R g959 ( .A(n_256), .Y(n_959) );
INVx2_ASAP7_75t_L g299 ( .A(n_257), .Y(n_299) );
AO22x1_ASAP7_75t_L g1323 ( .A1(n_258), .A2(n_272), .B1(n_1324), .B2(n_1327), .Y(n_1323) );
INVx1_ASAP7_75t_L g889 ( .A(n_259), .Y(n_889) );
INVx1_ASAP7_75t_L g902 ( .A(n_260), .Y(n_902) );
CKINVDCx5p33_ASAP7_75t_R g994 ( .A(n_261), .Y(n_994) );
INVx1_ASAP7_75t_L g1116 ( .A(n_262), .Y(n_1116) );
CKINVDCx5p33_ASAP7_75t_R g1241 ( .A(n_263), .Y(n_1241) );
INVx1_ASAP7_75t_L g604 ( .A(n_264), .Y(n_604) );
INVx1_ASAP7_75t_L g1053 ( .A(n_265), .Y(n_1053) );
INVx1_ASAP7_75t_L g573 ( .A(n_267), .Y(n_573) );
INVx1_ASAP7_75t_L g525 ( .A(n_268), .Y(n_525) );
CKINVDCx5p33_ASAP7_75t_R g1543 ( .A(n_269), .Y(n_1543) );
AOI21xp33_ASAP7_75t_L g618 ( .A1(n_270), .A2(n_408), .B(n_596), .Y(n_618) );
CKINVDCx5p33_ASAP7_75t_R g1123 ( .A(n_271), .Y(n_1123) );
INVx1_ASAP7_75t_L g1057 ( .A(n_273), .Y(n_1057) );
OAI211xp5_ASAP7_75t_SL g897 ( .A1(n_274), .A2(n_708), .B(n_898), .C(n_901), .Y(n_897) );
BUFx3_ASAP7_75t_L g326 ( .A(n_275), .Y(n_326) );
INVx1_ASAP7_75t_L g331 ( .A(n_275), .Y(n_331) );
INVx1_ASAP7_75t_L g325 ( .A(n_276), .Y(n_325) );
BUFx3_ASAP7_75t_L g330 ( .A(n_276), .Y(n_330) );
INVx1_ASAP7_75t_L g826 ( .A(n_277), .Y(n_826) );
INVx1_ASAP7_75t_L g1599 ( .A(n_278), .Y(n_1599) );
INVxp67_ASAP7_75t_SL g1183 ( .A(n_280), .Y(n_1183) );
AOI21xp5_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_303), .B(n_1293), .Y(n_281) );
HB1xp67_ASAP7_75t_L g282 ( .A(n_283), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g284 ( .A(n_285), .B(n_290), .Y(n_284) );
AND2x4_ASAP7_75t_L g1582 ( .A(n_285), .B(n_291), .Y(n_1582) );
NOR2xp33_ASAP7_75t_SL g285 ( .A(n_286), .B(n_288), .Y(n_285) );
INVx1_ASAP7_75t_SL g1576 ( .A(n_286), .Y(n_1576) );
NAND2xp5_ASAP7_75t_L g1644 ( .A(n_286), .B(n_288), .Y(n_1644) );
HB1xp67_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
AND2x2_ASAP7_75t_L g1575 ( .A(n_288), .B(n_1576), .Y(n_1575) );
INVx1_ASAP7_75t_L g288 ( .A(n_289), .Y(n_288) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_296), .Y(n_291) );
INVxp67_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
HB1xp67_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AND2x2_ASAP7_75t_L g681 ( .A(n_294), .B(n_302), .Y(n_681) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
OR2x2_ASAP7_75t_L g408 ( .A(n_295), .B(n_409), .Y(n_408) );
OR2x6_ASAP7_75t_L g296 ( .A(n_297), .B(n_301), .Y(n_296) );
OR2x2_ASAP7_75t_L g528 ( .A(n_297), .B(n_529), .Y(n_528) );
BUFx2_ASAP7_75t_L g560 ( .A(n_297), .Y(n_560) );
BUFx6f_ASAP7_75t_L g761 ( .A(n_297), .Y(n_761) );
INVx1_ASAP7_75t_L g779 ( .A(n_297), .Y(n_779) );
INVx2_ASAP7_75t_SL g863 ( .A(n_297), .Y(n_863) );
INVx2_ASAP7_75t_SL g958 ( .A(n_297), .Y(n_958) );
BUFx6f_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_299), .B(n_300), .Y(n_298) );
AND2x4_ASAP7_75t_L g388 ( .A(n_299), .B(n_389), .Y(n_388) );
INVx2_ASAP7_75t_L g393 ( .A(n_299), .Y(n_393) );
INVx1_ASAP7_75t_L g402 ( .A(n_299), .Y(n_402) );
AND2x2_ASAP7_75t_L g407 ( .A(n_299), .B(n_300), .Y(n_407) );
INVx1_ASAP7_75t_L g434 ( .A(n_299), .Y(n_434) );
INVx2_ASAP7_75t_L g389 ( .A(n_300), .Y(n_389) );
INVx1_ASAP7_75t_L g395 ( .A(n_300), .Y(n_395) );
INVx1_ASAP7_75t_L g401 ( .A(n_300), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_300), .B(n_393), .Y(n_413) );
INVx1_ASAP7_75t_L g446 ( .A(n_300), .Y(n_446) );
INVx2_ASAP7_75t_SL g301 ( .A(n_302), .Y(n_301) );
XNOR2xp5_ASAP7_75t_L g303 ( .A(n_304), .B(n_734), .Y(n_303) );
HB1xp67_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
XNOR2xp5_ASAP7_75t_L g306 ( .A(n_307), .B(n_582), .Y(n_306) );
AO22x2_ASAP7_75t_L g307 ( .A1(n_308), .A2(n_475), .B1(n_476), .B2(n_581), .Y(n_307) );
INVxp67_ASAP7_75t_SL g581 ( .A(n_308), .Y(n_581) );
INVxp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
NOR4xp75_ASAP7_75t_L g310 ( .A(n_311), .B(n_379), .C(n_455), .D(n_470), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_355), .Y(n_311) );
AOI33xp33_ASAP7_75t_L g312 ( .A1(n_313), .A2(n_321), .A3(n_332), .B1(n_341), .B2(n_347), .B3(n_351), .Y(n_312) );
INVx3_ASAP7_75t_L g313 ( .A(n_314), .Y(n_313) );
OAI22xp5_ASAP7_75t_SL g967 ( .A1(n_314), .A2(n_968), .B1(n_970), .B2(n_971), .Y(n_967) );
OR2x2_ASAP7_75t_L g314 ( .A(n_315), .B(n_317), .Y(n_314) );
BUFx2_ASAP7_75t_L g620 ( .A(n_315), .Y(n_620) );
INVx2_ASAP7_75t_L g625 ( .A(n_315), .Y(n_625) );
OR2x6_ASAP7_75t_L g638 ( .A(n_315), .B(n_639), .Y(n_638) );
AND2x4_ASAP7_75t_L g680 ( .A(n_315), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g922 ( .A(n_315), .B(n_436), .Y(n_922) );
AND2x4_ASAP7_75t_L g1130 ( .A(n_315), .B(n_681), .Y(n_1130) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
BUFx2_ASAP7_75t_L g454 ( .A(n_316), .Y(n_454) );
OR2x6_ASAP7_75t_L g556 ( .A(n_316), .B(n_408), .Y(n_556) );
INVx1_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
BUFx3_ASAP7_75t_L g512 ( .A(n_318), .Y(n_512) );
INVx2_ASAP7_75t_L g639 ( .A(n_318), .Y(n_639) );
INVx2_ASAP7_75t_SL g811 ( .A(n_318), .Y(n_811) );
INVx1_ASAP7_75t_L g1033 ( .A(n_318), .Y(n_1033) );
AND2x2_ASAP7_75t_L g318 ( .A(n_319), .B(n_320), .Y(n_318) );
AND2x4_ASAP7_75t_L g353 ( .A(n_319), .B(n_354), .Y(n_353) );
INVx2_ASAP7_75t_L g354 ( .A(n_320), .Y(n_354) );
INVx2_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
OAI22xp5_ASAP7_75t_L g635 ( .A1(n_323), .A2(n_612), .B1(n_614), .B2(n_636), .Y(n_635) );
INVx2_ASAP7_75t_L g659 ( .A(n_323), .Y(n_659) );
INVx1_ASAP7_75t_L g1220 ( .A(n_323), .Y(n_1220) );
INVx2_ASAP7_75t_SL g323 ( .A(n_324), .Y(n_323) );
BUFx3_ASAP7_75t_L g348 ( .A(n_324), .Y(n_348) );
BUFx6f_ASAP7_75t_L g469 ( .A(n_324), .Y(n_469) );
BUFx6f_ASAP7_75t_L g484 ( .A(n_324), .Y(n_484) );
BUFx2_ASAP7_75t_L g492 ( .A(n_324), .Y(n_492) );
BUFx6f_ASAP7_75t_L g724 ( .A(n_324), .Y(n_724) );
HB1xp67_ASAP7_75t_L g839 ( .A(n_324), .Y(n_839) );
BUFx6f_ASAP7_75t_L g895 ( .A(n_324), .Y(n_895) );
HB1xp67_ASAP7_75t_L g1284 ( .A(n_324), .Y(n_1284) );
AND2x4_ASAP7_75t_L g324 ( .A(n_325), .B(n_326), .Y(n_324) );
INVx1_ASAP7_75t_L g464 ( .A(n_325), .Y(n_464) );
INVx2_ASAP7_75t_L g336 ( .A(n_326), .Y(n_336) );
AND2x2_ASAP7_75t_L g340 ( .A(n_326), .B(n_330), .Y(n_340) );
AOI22xp33_ASAP7_75t_L g1015 ( .A1(n_327), .A2(n_634), .B1(n_997), .B2(n_1003), .Y(n_1015) );
INVx2_ASAP7_75t_SL g1272 ( .A(n_327), .Y(n_1272) );
BUFx6f_ASAP7_75t_L g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g636 ( .A(n_328), .Y(n_636) );
INVx1_ASAP7_75t_L g650 ( .A(n_328), .Y(n_650) );
HB1xp67_ASAP7_75t_L g834 ( .A(n_328), .Y(n_834) );
BUFx6f_ASAP7_75t_L g1062 ( .A(n_328), .Y(n_1062) );
INVx2_ASAP7_75t_L g1530 ( .A(n_328), .Y(n_1530) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g350 ( .A(n_329), .Y(n_350) );
INVx2_ASAP7_75t_L g496 ( .A(n_329), .Y(n_496) );
BUFx6f_ASAP7_75t_L g798 ( .A(n_329), .Y(n_798) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_331), .Y(n_329) );
INVx2_ASAP7_75t_L g337 ( .A(n_330), .Y(n_337) );
INVx1_ASAP7_75t_L g463 ( .A(n_331), .Y(n_463) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
BUFx6f_ASAP7_75t_L g343 ( .A(n_334), .Y(n_343) );
INVx2_ASAP7_75t_L g634 ( .A(n_334), .Y(n_634) );
INVx2_ASAP7_75t_SL g718 ( .A(n_334), .Y(n_718) );
INVx1_ASAP7_75t_L g1031 ( .A(n_334), .Y(n_1031) );
INVx2_ASAP7_75t_L g1164 ( .A(n_334), .Y(n_1164) );
INVx6_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g458 ( .A(n_335), .B(n_363), .Y(n_458) );
BUFx2_ASAP7_75t_L g514 ( .A(n_335), .Y(n_514) );
INVx2_ASAP7_75t_L g645 ( .A(n_335), .Y(n_645) );
AND2x4_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
INVx1_ASAP7_75t_L g373 ( .A(n_336), .Y(n_373) );
INVx1_ASAP7_75t_L g360 ( .A(n_337), .Y(n_360) );
INVx1_ASAP7_75t_L g642 ( .A(n_338), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_338), .B(n_378), .Y(n_656) );
BUFx2_ASAP7_75t_SL g1160 ( .A(n_338), .Y(n_1160) );
INVx1_ASAP7_75t_L g1287 ( .A(n_338), .Y(n_1287) );
BUFx6f_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
AND2x4_ASAP7_75t_L g505 ( .A(n_339), .B(n_485), .Y(n_505) );
INVx1_ASAP7_75t_L g509 ( .A(n_339), .Y(n_509) );
AND2x4_ASAP7_75t_L g516 ( .A(n_339), .B(n_517), .Y(n_516) );
BUFx4f_ASAP7_75t_L g1017 ( .A(n_339), .Y(n_1017) );
INVx1_ASAP7_75t_L g1222 ( .A(n_339), .Y(n_1222) );
BUFx3_ASAP7_75t_L g1526 ( .A(n_339), .Y(n_1526) );
INVx2_ASAP7_75t_SL g1539 ( .A(n_339), .Y(n_1539) );
BUFx6f_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
BUFx6f_ASAP7_75t_L g346 ( .A(n_340), .Y(n_346) );
INVx2_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVx1_ASAP7_75t_L g488 ( .A(n_343), .Y(n_488) );
INVx4_ASAP7_75t_L g1527 ( .A(n_343), .Y(n_1527) );
INVx2_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
INVx3_ASAP7_75t_L g489 ( .A(n_345), .Y(n_489) );
INVx2_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
INVx1_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
BUFx6f_ASAP7_75t_L g632 ( .A(n_346), .Y(n_632) );
BUFx6f_ASAP7_75t_L g810 ( .A(n_346), .Y(n_810) );
BUFx3_ASAP7_75t_L g1070 ( .A(n_348), .Y(n_1070) );
BUFx2_ASAP7_75t_L g1211 ( .A(n_349), .Y(n_1211) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g471 ( .A(n_350), .B(n_465), .Y(n_471) );
OR2x6_ASAP7_75t_L g981 ( .A(n_350), .B(n_465), .Y(n_981) );
AND2x4_ASAP7_75t_L g351 ( .A(n_352), .B(n_353), .Y(n_351) );
AND2x4_ASAP7_75t_L g457 ( .A(n_352), .B(n_458), .Y(n_457) );
AND2x4_ASAP7_75t_L g651 ( .A(n_352), .B(n_353), .Y(n_651) );
INVx2_ASAP7_75t_SL g490 ( .A(n_353), .Y(n_490) );
CKINVDCx5p33_ASAP7_75t_R g719 ( .A(n_353), .Y(n_719) );
HB1xp67_ASAP7_75t_L g803 ( .A(n_353), .Y(n_803) );
INVx2_ASAP7_75t_L g1217 ( .A(n_353), .Y(n_1217) );
AND2x4_ASAP7_75t_L g363 ( .A(n_354), .B(n_364), .Y(n_363) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_356), .A2(n_368), .B1(n_369), .B2(n_374), .C(n_375), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
INVx2_ASAP7_75t_L g654 ( .A(n_357), .Y(n_654) );
NAND2x1p5_ASAP7_75t_L g357 ( .A(n_358), .B(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx2_ASAP7_75t_L g502 ( .A(n_359), .Y(n_502) );
INVx1_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx2_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
OR2x6_ASAP7_75t_L g370 ( .A(n_362), .B(n_371), .Y(n_370) );
INVx1_ASAP7_75t_L g378 ( .A(n_362), .Y(n_378) );
OR2x2_ASAP7_75t_L g655 ( .A(n_362), .B(n_371), .Y(n_655) );
NAND2x1p5_ASAP7_75t_L g362 ( .A(n_363), .B(n_366), .Y(n_362) );
AND2x4_ASAP7_75t_L g499 ( .A(n_363), .B(n_372), .Y(n_499) );
AND2x4_ASAP7_75t_L g501 ( .A(n_363), .B(n_502), .Y(n_501) );
BUFx2_ASAP7_75t_L g517 ( .A(n_363), .Y(n_517) );
AND2x4_ASAP7_75t_L g793 ( .A(n_363), .B(n_502), .Y(n_793) );
AND2x2_ASAP7_75t_L g795 ( .A(n_363), .B(n_372), .Y(n_795) );
INVx1_ASAP7_75t_L g817 ( .A(n_363), .Y(n_817) );
AND2x2_ASAP7_75t_L g1150 ( .A(n_363), .B(n_372), .Y(n_1150) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
OR2x6_ASAP7_75t_L g579 ( .A(n_366), .B(n_437), .Y(n_579) );
INVx1_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
OR2x2_ASAP7_75t_L g465 ( .A(n_367), .B(n_466), .Y(n_465) );
AND2x4_ASAP7_75t_L g536 ( .A(n_367), .B(n_384), .Y(n_536) );
INVx2_ASAP7_75t_L g369 ( .A(n_370), .Y(n_369) );
OR2x2_ASAP7_75t_L g1209 ( .A(n_371), .B(n_817), .Y(n_1209) );
INVx2_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NOR3xp33_ASAP7_75t_L g965 ( .A(n_375), .B(n_966), .C(n_967), .Y(n_965) );
BUFx2_ASAP7_75t_L g1071 ( .A(n_375), .Y(n_1071) );
AND2x2_ASAP7_75t_L g375 ( .A(n_376), .B(n_378), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
AOI21x1_ASAP7_75t_L g379 ( .A1(n_380), .A2(n_422), .B(n_453), .Y(n_379) );
AOI221x1_ASAP7_75t_L g380 ( .A1(n_381), .A2(n_390), .B1(n_391), .B2(n_396), .C(n_397), .Y(n_380) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_381), .A2(n_391), .B1(n_603), .B2(n_604), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g939 ( .A1(n_381), .A2(n_391), .B1(n_940), .B2(n_941), .Y(n_939) );
INVx3_ASAP7_75t_L g1076 ( .A(n_381), .Y(n_1076) );
AND2x4_ASAP7_75t_L g381 ( .A(n_382), .B(n_386), .Y(n_381) );
AND2x4_ASAP7_75t_L g440 ( .A(n_382), .B(n_432), .Y(n_440) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g391 ( .A(n_384), .B(n_392), .Y(n_391) );
AND2x4_ASAP7_75t_L g607 ( .A(n_384), .B(n_430), .Y(n_607) );
INVx1_ASAP7_75t_L g409 ( .A(n_385), .Y(n_409) );
INVx1_ASAP7_75t_L g438 ( .A(n_385), .Y(n_438) );
INVx1_ASAP7_75t_L g415 ( .A(n_386), .Y(n_415) );
INVx2_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
INVx1_ASAP7_75t_L g572 ( .A(n_387), .Y(n_572) );
INVx1_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
INVx3_ASAP7_75t_L g427 ( .A(n_388), .Y(n_427) );
BUFx6f_ASAP7_75t_L g782 ( .A(n_388), .Y(n_782) );
AND2x4_ASAP7_75t_L g433 ( .A(n_389), .B(n_434), .Y(n_433) );
INVx3_ASAP7_75t_L g1075 ( .A(n_391), .Y(n_1075) );
BUFx6f_ASAP7_75t_L g424 ( .A(n_392), .Y(n_424) );
BUFx6f_ASAP7_75t_L g546 ( .A(n_392), .Y(n_546) );
INVx1_ASAP7_75t_L g591 ( .A(n_392), .Y(n_591) );
INVx1_ASAP7_75t_L g687 ( .A(n_392), .Y(n_687) );
BUFx6f_ASAP7_75t_L g944 ( .A(n_392), .Y(n_944) );
BUFx2_ASAP7_75t_L g1616 ( .A(n_392), .Y(n_1616) );
AND2x4_ASAP7_75t_L g392 ( .A(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g449 ( .A(n_393), .Y(n_449) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
OAI21xp5_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_410), .B(n_417), .Y(n_397) );
OAI21xp5_ASAP7_75t_SL g398 ( .A1(n_399), .A2(n_403), .B(n_404), .Y(n_398) );
INVx1_ASAP7_75t_L g764 ( .A(n_399), .Y(n_764) );
BUFx2_ASAP7_75t_L g775 ( .A(n_399), .Y(n_775) );
OAI221xp5_ASAP7_75t_L g955 ( .A1(n_399), .A2(n_956), .B1(n_957), .B2(n_959), .C(n_960), .Y(n_955) );
INVx3_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
INVx2_ASAP7_75t_L g418 ( .A(n_400), .Y(n_418) );
INVx2_ASAP7_75t_L g616 ( .A(n_400), .Y(n_616) );
AND2x2_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_401), .B(n_402), .Y(n_565) );
INVx1_ASAP7_75t_L g674 ( .A(n_402), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g626 ( .A(n_405), .B(n_627), .Y(n_626) );
AND2x2_ASAP7_75t_L g1007 ( .A(n_405), .B(n_536), .Y(n_1007) );
INVx2_ASAP7_75t_SL g405 ( .A(n_406), .Y(n_405) );
INVx2_ASAP7_75t_L g452 ( .A(n_406), .Y(n_452) );
INVx2_ASAP7_75t_SL g543 ( .A(n_406), .Y(n_543) );
INVx3_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
BUFx6f_ASAP7_75t_L g430 ( .A(n_407), .Y(n_430) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B1(n_415), .B2(n_416), .Y(n_410) );
INVx2_ASAP7_75t_L g569 ( .A(n_411), .Y(n_569) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx3_ASAP7_75t_L g870 ( .A(n_412), .Y(n_870) );
INVx1_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g611 ( .A(n_413), .Y(n_611) );
BUFx2_ASAP7_75t_L g951 ( .A(n_413), .Y(n_951) );
INVx1_ASAP7_75t_L g918 ( .A(n_415), .Y(n_918) );
OR2x6_ASAP7_75t_L g417 ( .A(n_418), .B(n_419), .Y(n_417) );
OAI22xp33_ASAP7_75t_L g578 ( .A1(n_418), .A2(n_506), .B1(n_519), .B2(n_558), .Y(n_578) );
OR2x2_ASAP7_75t_L g619 ( .A(n_418), .B(n_419), .Y(n_619) );
INVx1_ASAP7_75t_L g866 ( .A(n_418), .Y(n_866) );
INVx1_ASAP7_75t_L g447 ( .A(n_419), .Y(n_447) );
OR2x6_ASAP7_75t_L g448 ( .A(n_419), .B(n_449), .Y(n_448) );
INVx1_ASAP7_75t_L g627 ( .A(n_419), .Y(n_627) );
INVx2_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
INVx1_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
AOI221xp5_ASAP7_75t_SL g422 ( .A1(n_423), .A2(n_428), .B1(n_440), .B2(n_441), .C(n_442), .Y(n_422) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_425), .Y(n_770) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx3_ASAP7_75t_L g1260 ( .A(n_426), .Y(n_1260) );
INVx2_ASAP7_75t_L g1629 ( .A(n_426), .Y(n_1629) );
BUFx6f_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx3_ASAP7_75t_L g535 ( .A(n_427), .Y(n_535) );
INVx3_ASAP7_75t_L g594 ( .A(n_427), .Y(n_594) );
BUFx2_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
INVx3_ASAP7_75t_L g921 ( .A(n_430), .Y(n_921) );
BUFx6f_ASAP7_75t_L g946 ( .A(n_430), .Y(n_946) );
HB1xp67_ASAP7_75t_L g1195 ( .A(n_431), .Y(n_1195) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
BUFx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
BUFx3_ASAP7_75t_L g539 ( .A(n_433), .Y(n_539) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_433), .Y(n_600) );
BUFx2_ASAP7_75t_L g677 ( .A(n_433), .Y(n_677) );
BUFx6f_ASAP7_75t_L g684 ( .A(n_433), .Y(n_684) );
INVx2_ASAP7_75t_SL g435 ( .A(n_436), .Y(n_435) );
INVx1_ASAP7_75t_L g1098 ( .A(n_436), .Y(n_1098) );
INVx2_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2x1p5_ASAP7_75t_L g437 ( .A(n_438), .B(n_439), .Y(n_437) );
INVx8_ASAP7_75t_L g587 ( .A(n_440), .Y(n_587) );
NAND2x1p5_ASAP7_75t_L g443 ( .A(n_444), .B(n_447), .Y(n_443) );
NAND2x1_ASAP7_75t_SL g549 ( .A(n_444), .B(n_550), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g1622 ( .A1(n_444), .A2(n_553), .B1(n_1607), .B2(n_1608), .Y(n_1622) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
HB1xp67_ASAP7_75t_L g670 ( .A(n_446), .Y(n_670) );
CKINVDCx11_ASAP7_75t_R g1103 ( .A(n_448), .Y(n_1103) );
INVx1_ASAP7_75t_L g553 ( .A(n_449), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
INVx2_ASAP7_75t_L g480 ( .A(n_453), .Y(n_480) );
OAI31xp33_ASAP7_75t_L g1013 ( .A1(n_453), .A2(n_1014), .A3(n_1019), .B(n_1034), .Y(n_1013) );
BUFx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g962 ( .A(n_454), .Y(n_962) );
AND2x4_ASAP7_75t_L g527 ( .A(n_456), .B(n_528), .Y(n_527) );
INVx2_ASAP7_75t_L g456 ( .A(n_457), .Y(n_456) );
OR2x6_ASAP7_75t_L g623 ( .A(n_457), .B(n_624), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g1036 ( .A(n_458), .B(n_1037), .Y(n_1036) );
INVx2_ASAP7_75t_L g1606 ( .A(n_458), .Y(n_1606) );
OR2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_465), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx2_ASAP7_75t_L g802 ( .A(n_461), .Y(n_802) );
INVx2_ASAP7_75t_L g886 ( .A(n_461), .Y(n_886) );
INVx2_ASAP7_75t_L g1064 ( .A(n_461), .Y(n_1064) );
HB1xp67_ASAP7_75t_L g1271 ( .A(n_461), .Y(n_1271) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
OR2x2_ASAP7_75t_L g521 ( .A(n_462), .B(n_466), .Y(n_521) );
INVx1_ASAP7_75t_L g973 ( .A(n_462), .Y(n_973) );
BUFx2_ASAP7_75t_L g1052 ( .A(n_462), .Y(n_1052) );
OR2x2_ASAP7_75t_L g462 ( .A(n_463), .B(n_464), .Y(n_462) );
AND2x2_ASAP7_75t_L g474 ( .A(n_463), .B(n_464), .Y(n_474) );
OR2x2_ASAP7_75t_L g467 ( .A(n_465), .B(n_468), .Y(n_467) );
OR2x6_ASAP7_75t_L g472 ( .A(n_465), .B(n_473), .Y(n_472) );
INVx1_ASAP7_75t_L g660 ( .A(n_465), .Y(n_660) );
INVx2_ASAP7_75t_L g485 ( .A(n_466), .Y(n_485) );
OR2x2_ASAP7_75t_L g524 ( .A(n_466), .B(n_496), .Y(n_524) );
A2O1A1Ixp33_ASAP7_75t_L g1014 ( .A1(n_466), .A2(n_1015), .B(n_1016), .C(n_1018), .Y(n_1014) );
INVx1_ASAP7_75t_L g1152 ( .A(n_468), .Y(n_1152) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
BUFx4f_ASAP7_75t_L g510 ( .A(n_469), .Y(n_510) );
AND2x2_ASAP7_75t_L g709 ( .A(n_469), .B(n_485), .Y(n_709) );
INVx1_ASAP7_75t_L g1159 ( .A(n_469), .Y(n_1159) );
INVx1_ASAP7_75t_L g1067 ( .A(n_473), .Y(n_1067) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g715 ( .A(n_474), .Y(n_715) );
BUFx4f_ASAP7_75t_L g893 ( .A(n_474), .Y(n_893) );
INVx1_ASAP7_75t_L g1024 ( .A(n_474), .Y(n_1024) );
INVx1_ASAP7_75t_L g1056 ( .A(n_474), .Y(n_1056) );
BUFx2_ASAP7_75t_L g1215 ( .A(n_474), .Y(n_1215) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
XOR2x2_ASAP7_75t_L g476 ( .A(n_477), .B(n_580), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_478), .B(n_530), .Y(n_477) );
AOI22xp33_ASAP7_75t_L g478 ( .A1(n_479), .A2(n_481), .B1(n_525), .B2(n_526), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g704 ( .A1(n_479), .A2(n_526), .B1(n_705), .B2(n_730), .Y(n_704) );
INVx1_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AOI31xp33_ASAP7_75t_L g789 ( .A1(n_480), .A2(n_790), .A3(n_804), .B(n_818), .Y(n_789) );
AOI31xp33_ASAP7_75t_L g1144 ( .A1(n_480), .A2(n_1145), .A3(n_1155), .B(n_1166), .Y(n_1144) );
NAND3xp33_ASAP7_75t_L g481 ( .A(n_482), .B(n_503), .C(n_518), .Y(n_481) );
AOI221xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_486), .B1(n_487), .B2(n_491), .C(n_497), .Y(n_482) );
AOI211xp5_ASAP7_75t_L g790 ( .A1(n_483), .A2(n_774), .B(n_791), .C(n_796), .Y(n_790) );
AOI211xp5_ASAP7_75t_SL g1145 ( .A1(n_483), .A2(n_1146), .B(n_1147), .C(n_1151), .Y(n_1145) );
AOI211xp5_ASAP7_75t_L g1206 ( .A1(n_483), .A2(n_1207), .B(n_1208), .C(n_1210), .Y(n_1206) );
INVx1_ASAP7_75t_L g1277 ( .A(n_483), .Y(n_1277) );
AOI221xp5_ASAP7_75t_L g1524 ( .A1(n_483), .A2(n_1525), .B1(n_1528), .B2(n_1531), .C(n_1532), .Y(n_1524) );
AOI22xp33_ASAP7_75t_L g1598 ( .A1(n_483), .A2(n_520), .B1(n_1599), .B2(n_1600), .Y(n_1598) );
AND2x4_ASAP7_75t_L g483 ( .A(n_484), .B(n_485), .Y(n_483) );
INVx2_ASAP7_75t_SL g808 ( .A(n_484), .Y(n_808) );
OAI22xp5_ASAP7_75t_L g574 ( .A1(n_486), .A2(n_522), .B1(n_575), .B2(n_576), .Y(n_574) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g814 ( .A(n_495), .Y(n_814) );
INVx2_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g515 ( .A(n_496), .Y(n_515) );
INVx2_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx2_ASAP7_75t_SL g713 ( .A(n_499), .Y(n_713) );
AOI22xp5_ASAP7_75t_L g898 ( .A1(n_499), .A2(n_501), .B1(n_899), .B2(n_900), .Y(n_898) );
INVx2_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
INVx4_ASAP7_75t_L g712 ( .A(n_501), .Y(n_712) );
INVx1_ASAP7_75t_SL g842 ( .A(n_501), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_506), .B1(n_507), .B2(n_513), .C(n_516), .Y(n_503) );
HB1xp67_ASAP7_75t_L g504 ( .A(n_505), .Y(n_504) );
HB1xp67_ASAP7_75t_L g721 ( .A(n_505), .Y(n_721) );
BUFx6f_ASAP7_75t_L g805 ( .A(n_505), .Y(n_805) );
INVx2_ASAP7_75t_SL g830 ( .A(n_505), .Y(n_830) );
INVx1_ASAP7_75t_L g1602 ( .A(n_505), .Y(n_1602) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
INVx1_ASAP7_75t_L g647 ( .A(n_510), .Y(n_647) );
INVx3_ASAP7_75t_L g511 ( .A(n_512), .Y(n_511) );
INVxp67_ASAP7_75t_L g725 ( .A(n_512), .Y(n_725) );
INVx1_ASAP7_75t_L g1594 ( .A(n_512), .Y(n_1594) );
AOI221xp5_ASAP7_75t_L g720 ( .A1(n_516), .A2(n_721), .B1(n_722), .B2(n_723), .C(n_726), .Y(n_720) );
AOI221xp5_ASAP7_75t_L g828 ( .A1(n_516), .A2(n_829), .B1(n_831), .B2(n_832), .C(n_833), .Y(n_828) );
INVx1_ASAP7_75t_L g896 ( .A(n_516), .Y(n_896) );
INVx1_ASAP7_75t_L g1018 ( .A(n_516), .Y(n_1018) );
AOI221xp5_ASAP7_75t_L g1534 ( .A1(n_516), .A2(n_805), .B1(n_1535), .B2(n_1540), .C(n_1541), .Y(n_1534) );
AOI22xp33_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B1(n_522), .B2(n_523), .Y(n_518) );
AOI22xp33_ASAP7_75t_L g727 ( .A1(n_520), .A2(n_523), .B1(n_728), .B2(n_729), .Y(n_727) );
AOI22xp33_ASAP7_75t_L g818 ( .A1(n_520), .A2(n_523), .B1(n_780), .B2(n_783), .Y(n_818) );
AOI22xp5_ASAP7_75t_L g825 ( .A1(n_520), .A2(n_523), .B1(n_826), .B2(n_827), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g1166 ( .A1(n_520), .A2(n_523), .B1(n_1167), .B2(n_1168), .Y(n_1166) );
AOI22xp33_ASAP7_75t_L g1226 ( .A1(n_520), .A2(n_523), .B1(n_1227), .B2(n_1228), .Y(n_1226) );
AOI22xp33_ASAP7_75t_L g1542 ( .A1(n_520), .A2(n_523), .B1(n_1543), .B2(n_1544), .Y(n_1542) );
INVx6_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
INVx4_ASAP7_75t_L g523 ( .A(n_524), .Y(n_523) );
INVx2_ASAP7_75t_L g526 ( .A(n_527), .Y(n_526) );
INVx5_ASAP7_75t_L g787 ( .A(n_527), .Y(n_787) );
INVx2_ASAP7_75t_SL g845 ( .A(n_527), .Y(n_845) );
INVx1_ASAP7_75t_L g1203 ( .A(n_527), .Y(n_1203) );
INVx1_ASAP7_75t_L g1546 ( .A(n_527), .Y(n_1546) );
INVx3_ASAP7_75t_L g550 ( .A(n_529), .Y(n_550) );
NOR3xp33_ASAP7_75t_L g530 ( .A(n_531), .B(n_547), .C(n_555), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_532), .B(n_540), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_533), .A2(n_534), .B1(n_537), .B2(n_538), .Y(n_532) );
BUFx2_ASAP7_75t_L g698 ( .A(n_534), .Y(n_698) );
BUFx2_ASAP7_75t_L g747 ( .A(n_534), .Y(n_747) );
BUFx2_ASAP7_75t_L g1122 ( .A(n_534), .Y(n_1122) );
BUFx2_ASAP7_75t_L g1551 ( .A(n_534), .Y(n_1551) );
AND2x4_ASAP7_75t_L g534 ( .A(n_535), .B(n_536), .Y(n_534) );
BUFx3_ASAP7_75t_L g577 ( .A(n_535), .Y(n_577) );
INVx2_ASAP7_75t_L g613 ( .A(n_535), .Y(n_613) );
INVx1_ASAP7_75t_L g953 ( .A(n_535), .Y(n_953) );
AND2x6_ASAP7_75t_L g538 ( .A(n_536), .B(n_539), .Y(n_538) );
AND2x4_ASAP7_75t_L g542 ( .A(n_536), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g545 ( .A(n_536), .B(n_546), .Y(n_545) );
AND2x2_ASAP7_75t_L g703 ( .A(n_536), .B(n_546), .Y(n_703) );
AND2x2_ASAP7_75t_L g752 ( .A(n_536), .B(n_546), .Y(n_752) );
AND2x2_ASAP7_75t_L g850 ( .A(n_536), .B(n_594), .Y(n_850) );
AND2x2_ASAP7_75t_L g852 ( .A(n_536), .B(n_684), .Y(n_852) );
AND2x2_ASAP7_75t_L g856 ( .A(n_536), .B(n_546), .Y(n_856) );
AND2x2_ASAP7_75t_L g1127 ( .A(n_536), .B(n_546), .Y(n_1127) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_538), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
AOI22xp33_ASAP7_75t_L g745 ( .A1(n_538), .A2(n_746), .B1(n_747), .B2(n_748), .Y(n_745) );
AOI22xp33_ASAP7_75t_L g1120 ( .A1(n_538), .A2(n_1121), .B1(n_1122), .B2(n_1123), .Y(n_1120) );
AOI22xp33_ASAP7_75t_L g1185 ( .A1(n_538), .A2(n_747), .B1(n_1186), .B2(n_1187), .Y(n_1185) );
AOI22xp33_ASAP7_75t_L g1240 ( .A1(n_538), .A2(n_698), .B1(n_1241), .B2(n_1242), .Y(n_1240) );
AOI22xp33_ASAP7_75t_L g1549 ( .A1(n_538), .A2(n_1550), .B1(n_1551), .B2(n_1552), .Y(n_1549) );
INVx1_ASAP7_75t_SL g1613 ( .A(n_538), .Y(n_1613) );
NAND2x1p5_ASAP7_75t_L g554 ( .A(n_539), .B(n_550), .Y(n_554) );
BUFx2_ASAP7_75t_L g1619 ( .A(n_539), .Y(n_1619) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_542), .B1(n_544), .B2(n_545), .Y(n_540) );
AOI22xp33_ASAP7_75t_L g700 ( .A1(n_542), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_542), .A2(n_750), .B1(n_751), .B2(n_752), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g853 ( .A1(n_542), .A2(n_854), .B1(n_855), .B2(n_856), .Y(n_853) );
AOI221xp5_ASAP7_75t_L g924 ( .A1(n_542), .A2(n_752), .B1(n_925), .B2(n_926), .C(n_927), .Y(n_924) );
AOI22xp33_ASAP7_75t_L g1124 ( .A1(n_542), .A2(n_1125), .B1(n_1126), .B2(n_1127), .Y(n_1124) );
AOI22xp33_ASAP7_75t_L g1188 ( .A1(n_542), .A2(n_752), .B1(n_1189), .B2(n_1190), .Y(n_1188) );
AOI22xp33_ASAP7_75t_L g1243 ( .A1(n_542), .A2(n_545), .B1(n_1244), .B2(n_1245), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1553 ( .A1(n_542), .A2(n_703), .B1(n_1554), .B2(n_1555), .Y(n_1553) );
AOI22xp33_ASAP7_75t_L g1624 ( .A1(n_542), .A2(n_1127), .B1(n_1625), .B2(n_1626), .Y(n_1624) );
INVx1_ASAP7_75t_L g597 ( .A(n_543), .Y(n_597) );
INVx1_ASAP7_75t_L g693 ( .A(n_543), .Y(n_693) );
BUFx2_ASAP7_75t_L g912 ( .A(n_543), .Y(n_912) );
BUFx3_ASAP7_75t_L g1141 ( .A(n_543), .Y(n_1141) );
INVx2_ASAP7_75t_SL g1137 ( .A(n_546), .Y(n_1137) );
HB1xp67_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
INVx2_ASAP7_75t_L g755 ( .A(n_549), .Y(n_755) );
NAND2x1p5_ASAP7_75t_L g552 ( .A(n_550), .B(n_553), .Y(n_552) );
AND2x4_ASAP7_75t_L g669 ( .A(n_550), .B(n_670), .Y(n_669) );
AND2x4_ASAP7_75t_L g672 ( .A(n_550), .B(n_673), .Y(n_672) );
AND2x4_ASAP7_75t_L g676 ( .A(n_550), .B(n_677), .Y(n_676) );
AOI32xp33_ASAP7_75t_L g1614 ( .A1(n_550), .A2(n_1130), .A3(n_1615), .B1(n_1618), .B2(n_1620), .Y(n_1614) );
BUFx4f_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
BUFx4f_ASAP7_75t_L g756 ( .A(n_552), .Y(n_756) );
BUFx2_ASAP7_75t_L g757 ( .A(n_554), .Y(n_757) );
BUFx3_ASAP7_75t_L g859 ( .A(n_554), .Y(n_859) );
OAI33xp33_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .A3(n_567), .B1(n_574), .B2(n_578), .B3(n_579), .Y(n_555) );
OAI33xp33_ASAP7_75t_L g758 ( .A1(n_556), .A2(n_759), .A3(n_766), .B1(n_772), .B2(n_777), .B3(n_784), .Y(n_758) );
OAI33xp33_ASAP7_75t_L g860 ( .A1(n_556), .A2(n_861), .A3(n_868), .B1(n_873), .B2(n_875), .B3(n_877), .Y(n_860) );
OAI33xp33_ASAP7_75t_L g1247 ( .A1(n_556), .A2(n_784), .A3(n_1248), .B1(n_1253), .B2(n_1257), .B3(n_1262), .Y(n_1247) );
OAI33xp33_ASAP7_75t_L g1557 ( .A1(n_556), .A2(n_877), .A3(n_1558), .B1(n_1562), .B2(n_1566), .B3(n_1571), .Y(n_1557) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_558), .A2(n_561), .B1(n_562), .B2(n_566), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g1621 ( .A(n_559), .Y(n_1621) );
INVx2_ASAP7_75t_SL g559 ( .A(n_560), .Y(n_559) );
INVx2_ASAP7_75t_L g562 ( .A(n_563), .Y(n_562) );
INVx2_ASAP7_75t_L g1633 ( .A(n_563), .Y(n_1633) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
BUFx3_ASAP7_75t_L g876 ( .A(n_564), .Y(n_876) );
BUFx3_ASAP7_75t_L g995 ( .A(n_564), .Y(n_995) );
OAI22xp33_ASAP7_75t_L g996 ( .A1(n_564), .A2(n_761), .B1(n_997), .B2(n_998), .Y(n_996) );
BUFx6f_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g567 ( .A1(n_568), .A2(n_570), .B1(n_571), .B2(n_573), .Y(n_567) );
INVx2_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx1_ASAP7_75t_L g575 ( .A(n_569), .Y(n_575) );
INVx2_ASAP7_75t_L g767 ( .A(n_569), .Y(n_767) );
INVx2_ASAP7_75t_L g773 ( .A(n_569), .Y(n_773) );
INVx1_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_572), .Y(n_688) );
INVx1_ASAP7_75t_L g874 ( .A(n_572), .Y(n_874) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx6_ASAP7_75t_L g695 ( .A(n_579), .Y(n_695) );
INVx5_ASAP7_75t_L g785 ( .A(n_579), .Y(n_785) );
AO22x1_ASAP7_75t_SL g582 ( .A1(n_583), .A2(n_665), .B1(n_732), .B2(n_733), .Y(n_582) );
INVx1_ASAP7_75t_L g732 ( .A(n_583), .Y(n_732) );
NAND4xp25_ASAP7_75t_L g584 ( .A(n_585), .B(n_621), .C(n_628), .D(n_657), .Y(n_584) );
OAI21xp5_ASAP7_75t_SL g585 ( .A1(n_586), .A2(n_605), .B(n_620), .Y(n_585) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_589), .A2(n_595), .B(n_601), .Y(n_588) );
INVx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_L g592 ( .A(n_593), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
INVx2_ASAP7_75t_L g916 ( .A(n_594), .Y(n_916) );
HB1xp67_ASAP7_75t_L g991 ( .A(n_594), .Y(n_991) );
INVx1_ASAP7_75t_L g1087 ( .A(n_594), .Y(n_1087) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_SL g599 ( .A(n_600), .Y(n_599) );
BUFx2_ASAP7_75t_L g694 ( .A(n_600), .Y(n_694) );
OAI22xp5_ASAP7_75t_L g646 ( .A1(n_603), .A2(n_604), .B1(n_647), .B2(n_648), .Y(n_646) );
CKINVDCx6p67_ASAP7_75t_R g606 ( .A(n_607), .Y(n_606) );
OAI22xp5_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_612), .B1(n_613), .B2(n_614), .Y(n_608) );
OAI22xp5_ASAP7_75t_L g873 ( .A1(n_609), .A2(n_827), .B1(n_836), .B2(n_874), .Y(n_873) );
INVx1_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
HB1xp67_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g1002 ( .A(n_611), .Y(n_1002) );
INVx1_ASAP7_75t_L g1569 ( .A(n_611), .Y(n_1569) );
INVx1_ASAP7_75t_L g690 ( .A(n_613), .Y(n_690) );
OAI22xp5_ASAP7_75t_L g868 ( .A1(n_613), .A2(n_869), .B1(n_871), .B2(n_872), .Y(n_868) );
OAI21xp5_ASAP7_75t_SL g615 ( .A1(n_616), .A2(n_617), .B(n_618), .Y(n_615) );
CKINVDCx8_ASAP7_75t_R g843 ( .A(n_620), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_622), .B(n_623), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g963 ( .A(n_623), .B(n_964), .Y(n_963) );
NAND2xp5_ASAP7_75t_L g1046 ( .A(n_623), .B(n_1047), .Y(n_1046) );
NOR2xp67_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
INVx2_ASAP7_75t_L g908 ( .A(n_625), .Y(n_908) );
AND2x2_ASAP7_75t_L g1101 ( .A(n_627), .B(n_670), .Y(n_1101) );
AOI221xp5_ASAP7_75t_L g628 ( .A1(n_629), .A2(n_637), .B1(n_640), .B2(n_651), .C(n_652), .Y(n_628) );
INVx1_ASAP7_75t_L g630 ( .A(n_631), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x4_ASAP7_75t_L g815 ( .A(n_632), .B(n_816), .Y(n_815) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_634), .Y(n_633) );
BUFx3_ASAP7_75t_L g813 ( .A(n_634), .Y(n_813) );
INVx1_ASAP7_75t_L g840 ( .A(n_636), .Y(n_840) );
INVx1_ASAP7_75t_L g1050 ( .A(n_637), .Y(n_1050) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
BUFx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
AND2x2_ASAP7_75t_L g662 ( .A(n_644), .B(n_660), .Y(n_662) );
INVx2_ASAP7_75t_SL g644 ( .A(n_645), .Y(n_644) );
INVx1_ASAP7_75t_L g1027 ( .A(n_645), .Y(n_1027) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
INVx4_ASAP7_75t_L g970 ( .A(n_651), .Y(n_970) );
INVx1_ASAP7_75t_L g653 ( .A(n_654), .Y(n_653) );
AOI221xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_661), .B1(n_662), .B2(n_663), .C(n_664), .Y(n_657) );
AOI221xp5_ASAP7_75t_L g977 ( .A1(n_658), .A2(n_662), .B1(n_978), .B2(n_979), .C(n_980), .Y(n_977) );
AND2x2_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g1016 ( .A1(n_659), .A2(n_998), .B1(n_1000), .B2(n_1017), .Y(n_1016) );
INVx1_ASAP7_75t_L g733 ( .A(n_665), .Y(n_733) );
XNOR2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_731), .Y(n_665) );
NAND2x1_ASAP7_75t_L g666 ( .A(n_667), .B(n_704), .Y(n_666) );
AND4x1_ASAP7_75t_L g667 ( .A(n_668), .B(n_678), .C(n_696), .D(n_700), .Y(n_667) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_669), .A2(n_671), .B1(n_672), .B2(n_675), .C(n_676), .Y(n_668) );
AOI221xp5_ASAP7_75t_L g923 ( .A1(n_669), .A2(n_672), .B1(n_676), .B2(n_899), .C(n_900), .Y(n_923) );
AOI221xp5_ASAP7_75t_L g1038 ( .A1(n_669), .A2(n_672), .B1(n_676), .B2(n_1039), .C(n_1040), .Y(n_1038) );
INVx1_ASAP7_75t_L g1118 ( .A(n_669), .Y(n_1118) );
AOI221xp5_ASAP7_75t_L g1179 ( .A1(n_669), .A2(n_1180), .B1(n_1182), .B2(n_1183), .C(n_1184), .Y(n_1179) );
HB1xp67_ASAP7_75t_L g1115 ( .A(n_672), .Y(n_1115) );
INVx1_ASAP7_75t_L g1181 ( .A(n_672), .Y(n_1181) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_676), .A2(n_1115), .B1(n_1116), .B2(n_1117), .C(n_1119), .Y(n_1114) );
HB1xp67_ASAP7_75t_L g1184 ( .A(n_676), .Y(n_1184) );
AOI33xp33_ASAP7_75t_L g678 ( .A1(n_679), .A2(n_682), .A3(n_685), .B1(n_689), .B2(n_691), .B3(n_695), .Y(n_678) );
BUFx2_ASAP7_75t_L g679 ( .A(n_680), .Y(n_679) );
AOI33xp33_ASAP7_75t_L g910 ( .A1(n_680), .A2(n_911), .A3(n_913), .B1(n_917), .B2(n_919), .B3(n_922), .Y(n_910) );
BUFx2_ASAP7_75t_SL g960 ( .A(n_681), .Y(n_960) );
INVx1_ASAP7_75t_L g1080 ( .A(n_681), .Y(n_1080) );
BUFx6f_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
INVx2_ASAP7_75t_SL g1095 ( .A(n_684), .Y(n_1095) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g914 ( .A(n_687), .Y(n_914) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
INVx2_ASAP7_75t_L g877 ( .A(n_695), .Y(n_877) );
INVx1_ASAP7_75t_L g1005 ( .A(n_695), .Y(n_1005) );
AOI33xp33_ASAP7_75t_L g1128 ( .A1(n_695), .A2(n_1129), .A3(n_1131), .B1(n_1134), .B2(n_1138), .B3(n_1140), .Y(n_1128) );
AOI33xp33_ASAP7_75t_L g1191 ( .A1(n_695), .A2(n_1192), .A3(n_1194), .B1(n_1196), .B2(n_1198), .B3(n_1201), .Y(n_1191) );
AOI22xp5_ASAP7_75t_L g1627 ( .A1(n_695), .A2(n_1551), .B1(n_1628), .B2(n_1634), .Y(n_1627) );
OAI211xp5_ASAP7_75t_L g714 ( .A1(n_699), .A2(n_715), .B(n_716), .C(n_717), .Y(n_714) );
NAND3xp33_ASAP7_75t_L g705 ( .A(n_706), .B(n_720), .C(n_727), .Y(n_705) );
AOI21xp5_ASAP7_75t_SL g706 ( .A1(n_707), .A2(n_710), .B(n_711), .Y(n_706) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
AOI221xp5_ASAP7_75t_L g835 ( .A1(n_709), .A2(n_836), .B1(n_837), .B2(n_838), .C(n_841), .Y(n_835) );
OAI221xp5_ASAP7_75t_L g801 ( .A1(n_715), .A2(n_748), .B1(n_750), .B2(n_802), .C(n_803), .Y(n_801) );
OAI221xp5_ASAP7_75t_L g1154 ( .A1(n_715), .A2(n_803), .B1(n_972), .B2(n_1123), .C(n_1125), .Y(n_1154) );
INVx2_ASAP7_75t_L g800 ( .A(n_724), .Y(n_800) );
INVx2_ASAP7_75t_SL g1593 ( .A(n_724), .Y(n_1593) );
OAI22xp33_ASAP7_75t_L g1393 ( .A1(n_731), .A2(n_1394), .B1(n_1395), .B2(n_1396), .Y(n_1393) );
AOI22xp5_ASAP7_75t_L g734 ( .A1(n_735), .A2(n_736), .B1(n_1170), .B2(n_1171), .Y(n_734) );
INVx1_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
AO22x2_ASAP7_75t_L g736 ( .A1(n_737), .A2(n_738), .B1(n_1110), .B2(n_1169), .Y(n_736) );
INVx2_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
XNOR2xp5_ASAP7_75t_L g738 ( .A(n_739), .B(n_933), .Y(n_738) );
OAI22xp5_ASAP7_75t_L g739 ( .A1(n_740), .A2(n_741), .B1(n_820), .B2(n_932), .Y(n_739) );
INVx2_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
XNOR2x1_ASAP7_75t_L g741 ( .A(n_742), .B(n_819), .Y(n_741) );
AND2x2_ASAP7_75t_L g742 ( .A(n_743), .B(n_786), .Y(n_742) );
NOR3xp33_ASAP7_75t_L g743 ( .A(n_744), .B(n_753), .C(n_758), .Y(n_743) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_749), .Y(n_744) );
INVx2_ASAP7_75t_SL g754 ( .A(n_755), .Y(n_754) );
INVx2_ASAP7_75t_L g858 ( .A(n_755), .Y(n_858) );
OAI22xp33_ASAP7_75t_L g759 ( .A1(n_760), .A2(n_762), .B1(n_763), .B2(n_765), .Y(n_759) );
OAI22xp33_ASAP7_75t_L g1571 ( .A1(n_760), .A2(n_876), .B1(n_1541), .B2(n_1543), .Y(n_1571) );
BUFx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
OAI22xp33_ASAP7_75t_L g875 ( .A1(n_761), .A2(n_826), .B1(n_831), .B2(n_876), .Y(n_875) );
OAI22xp33_ASAP7_75t_L g1253 ( .A1(n_761), .A2(n_1254), .B1(n_1255), .B2(n_1256), .Y(n_1253) );
OAI22xp33_ASAP7_75t_L g1262 ( .A1(n_761), .A2(n_1263), .B1(n_1264), .B2(n_1265), .Y(n_1262) );
INVx1_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
INVx1_ASAP7_75t_L g1264 ( .A(n_764), .Y(n_1264) );
OAI22xp5_ASAP7_75t_L g766 ( .A1(n_767), .A2(n_768), .B1(n_769), .B2(n_771), .Y(n_766) );
OAI221xp5_ASAP7_75t_L g1090 ( .A1(n_767), .A2(n_1004), .B1(n_1091), .B2(n_1092), .C(n_1093), .Y(n_1090) );
OAI22xp5_ASAP7_75t_SL g1562 ( .A1(n_767), .A2(n_1563), .B1(n_1564), .B2(n_1565), .Y(n_1562) );
INVx1_ASAP7_75t_L g769 ( .A(n_770), .Y(n_769) );
OAI22xp5_ASAP7_75t_L g772 ( .A1(n_773), .A2(n_774), .B1(n_775), .B2(n_776), .Y(n_772) );
OAI221xp5_ASAP7_75t_L g1078 ( .A1(n_775), .A2(n_957), .B1(n_1053), .B2(n_1057), .C(n_1079), .Y(n_1078) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_776), .A2(n_805), .B1(n_806), .B2(n_812), .C(n_815), .Y(n_804) );
OAI22xp5_ASAP7_75t_L g777 ( .A1(n_778), .A2(n_780), .B1(n_781), .B2(n_783), .Y(n_777) );
INVx2_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g1560 ( .A(n_779), .Y(n_1560) );
INVx1_ASAP7_75t_L g1631 ( .A(n_779), .Y(n_1631) );
INVx2_ASAP7_75t_SL g1132 ( .A(n_781), .Y(n_1132) );
INVx2_ASAP7_75t_L g1617 ( .A(n_781), .Y(n_1617) );
INVx4_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx2_ASAP7_75t_SL g1004 ( .A(n_782), .Y(n_1004) );
BUFx3_ASAP7_75t_L g1139 ( .A(n_782), .Y(n_1139) );
INVx2_ASAP7_75t_SL g1200 ( .A(n_782), .Y(n_1200) );
CKINVDCx8_ASAP7_75t_R g784 ( .A(n_785), .Y(n_784) );
AOI21xp33_ASAP7_75t_SL g786 ( .A1(n_787), .A2(n_788), .B(n_789), .Y(n_786) );
AOI21xp5_ASAP7_75t_L g1142 ( .A1(n_787), .A2(n_1143), .B(n_1144), .Y(n_1142) );
INVx1_ASAP7_75t_L g1237 ( .A(n_787), .Y(n_1237) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
INVx2_ASAP7_75t_SL g1035 ( .A(n_793), .Y(n_1035) );
INVx2_ASAP7_75t_L g1148 ( .A(n_793), .Y(n_1148) );
AOI22xp33_ASAP7_75t_L g1278 ( .A1(n_793), .A2(n_1279), .B1(n_1280), .B2(n_1281), .Y(n_1278) );
INVx1_ASAP7_75t_L g1533 ( .A(n_793), .Y(n_1533) );
AOI222xp33_ASAP7_75t_L g1603 ( .A1(n_793), .A2(n_1150), .B1(n_1604), .B2(n_1605), .C1(n_1607), .C2(n_1608), .Y(n_1603) );
INVx3_ASAP7_75t_L g794 ( .A(n_795), .Y(n_794) );
BUFx6f_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g888 ( .A(n_798), .Y(n_888) );
BUFx3_ASAP7_75t_L g1153 ( .A(n_798), .Y(n_1153) );
INVx2_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
OAI221xp5_ASAP7_75t_L g968 ( .A1(n_802), .A2(n_892), .B1(n_956), .B2(n_959), .C(n_969), .Y(n_968) );
AOI221xp5_ASAP7_75t_L g1155 ( .A1(n_805), .A2(n_815), .B1(n_1156), .B2(n_1157), .C(n_1161), .Y(n_1155) );
AOI221xp5_ASAP7_75t_L g1218 ( .A1(n_805), .A2(n_815), .B1(n_1219), .B2(n_1223), .C(n_1225), .Y(n_1218) );
INVx1_ASAP7_75t_L g1268 ( .A(n_805), .Y(n_1268) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g1059 ( .A(n_808), .Y(n_1059) );
HB1xp67_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
BUFx2_ASAP7_75t_L g1274 ( .A(n_811), .Y(n_1274) );
INVx1_ASAP7_75t_L g1275 ( .A(n_815), .Y(n_1275) );
INVx1_ASAP7_75t_L g1609 ( .A(n_815), .Y(n_1609) );
INVx1_ASAP7_75t_SL g816 ( .A(n_817), .Y(n_816) );
INVx2_ASAP7_75t_L g932 ( .A(n_820), .Y(n_932) );
XOR2x2_ASAP7_75t_L g820 ( .A(n_821), .B(n_880), .Y(n_820) );
INVx1_ASAP7_75t_L g878 ( .A(n_822), .Y(n_878) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_846), .Y(n_822) );
AOI22xp5_ASAP7_75t_L g823 ( .A1(n_824), .A2(n_843), .B1(n_844), .B2(n_845), .Y(n_823) );
NAND3xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_828), .C(n_835), .Y(n_824) );
INVx1_ASAP7_75t_L g829 ( .A(n_830), .Y(n_829) );
INVx2_ASAP7_75t_L g1229 ( .A(n_843), .Y(n_1229) );
NOR3xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_857), .C(n_860), .Y(n_846) );
NAND2xp5_ASAP7_75t_SL g847 ( .A(n_848), .B(n_853), .Y(n_847) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_849), .A2(n_850), .B1(n_851), .B2(n_852), .Y(n_848) );
INVx2_ASAP7_75t_L g928 ( .A(n_850), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_852), .Y(n_929) );
INVxp67_ASAP7_75t_L g1011 ( .A(n_852), .Y(n_1011) );
INVx1_ASAP7_75t_L g1010 ( .A(n_856), .Y(n_1010) );
OAI22xp33_ASAP7_75t_L g861 ( .A1(n_862), .A2(n_864), .B1(n_865), .B2(n_867), .Y(n_861) );
INVx2_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx1_ASAP7_75t_L g865 ( .A(n_866), .Y(n_865) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_SL g1083 ( .A(n_870), .Y(n_1083) );
OAI22xp33_ASAP7_75t_L g1558 ( .A1(n_876), .A2(n_1559), .B1(n_1560), .B2(n_1561), .Y(n_1558) );
OAI22xp33_ASAP7_75t_L g1341 ( .A1(n_879), .A2(n_1310), .B1(n_1317), .B2(n_1342), .Y(n_1341) );
INVx1_ASAP7_75t_L g931 ( .A(n_881), .Y(n_931) );
NAND4xp75_ASAP7_75t_L g881 ( .A(n_882), .B(n_883), .C(n_909), .D(n_924), .Y(n_881) );
OAI31xp33_ASAP7_75t_L g883 ( .A1(n_884), .A2(n_897), .A3(n_906), .B(n_907), .Y(n_883) );
OAI22xp5_ASAP7_75t_L g885 ( .A1(n_886), .A2(n_887), .B1(n_888), .B2(n_889), .Y(n_885) );
INVx1_ASAP7_75t_L g1590 ( .A(n_888), .Y(n_1590) );
OAI21xp33_ASAP7_75t_L g890 ( .A1(n_891), .A2(n_892), .B(n_894), .Y(n_890) );
OAI221xp5_ASAP7_75t_L g971 ( .A1(n_892), .A2(n_972), .B1(n_974), .B2(n_975), .C(n_976), .Y(n_971) );
INVx2_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
INVx1_ASAP7_75t_L g903 ( .A(n_893), .Y(n_903) );
INVx1_ASAP7_75t_L g1029 ( .A(n_893), .Y(n_1029) );
BUFx3_ASAP7_75t_L g1212 ( .A(n_895), .Y(n_1212) );
INVx2_ASAP7_75t_L g1537 ( .A(n_895), .Y(n_1537) );
OAI211xp5_ASAP7_75t_L g901 ( .A1(n_902), .A2(n_903), .B(n_904), .C(n_905), .Y(n_901) );
OAI31xp33_ASAP7_75t_L g1266 ( .A1(n_907), .A2(n_1267), .A3(n_1276), .B(n_1289), .Y(n_1266) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
OAI31xp33_ASAP7_75t_SL g1073 ( .A1(n_908), .A2(n_1074), .A3(n_1077), .B(n_1089), .Y(n_1073) );
AND2x2_ASAP7_75t_SL g909 ( .A(n_910), .B(n_923), .Y(n_909) );
INVx1_ASAP7_75t_L g915 ( .A(n_916), .Y(n_915) );
INVx2_ASAP7_75t_L g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_SL g1135 ( .A(n_921), .Y(n_1135) );
AOI22xp33_ASAP7_75t_L g933 ( .A1(n_934), .A2(n_1043), .B1(n_1108), .B2(n_1109), .Y(n_933) );
INVx1_ASAP7_75t_L g1108 ( .A(n_934), .Y(n_1108) );
XNOR2x1_ASAP7_75t_L g934 ( .A(n_935), .B(n_984), .Y(n_934) );
INVx1_ASAP7_75t_L g982 ( .A(n_936), .Y(n_982) );
NAND4xp25_ASAP7_75t_L g936 ( .A(n_937), .B(n_963), .C(n_965), .D(n_977), .Y(n_936) );
OAI21xp5_ASAP7_75t_L g937 ( .A1(n_938), .A2(n_948), .B(n_961), .Y(n_937) );
AOI21xp5_ASAP7_75t_L g942 ( .A1(n_943), .A2(n_945), .B(n_947), .Y(n_942) );
BUFx3_ASAP7_75t_L g1197 ( .A(n_944), .Y(n_1197) );
INVx1_ASAP7_75t_L g1097 ( .A(n_946), .Y(n_1097) );
OAI22xp5_ASAP7_75t_L g949 ( .A1(n_950), .A2(n_952), .B1(n_953), .B2(n_954), .Y(n_949) );
OAI22xp5_ASAP7_75t_L g987 ( .A1(n_950), .A2(n_988), .B1(n_989), .B2(n_990), .Y(n_987) );
BUFx2_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx2_ASAP7_75t_L g1250 ( .A(n_951), .Y(n_1250) );
OAI22xp33_ASAP7_75t_L g992 ( .A1(n_957), .A2(n_993), .B1(n_994), .B2(n_995), .Y(n_992) );
INVx3_ASAP7_75t_L g957 ( .A(n_958), .Y(n_957) );
INVx5_ASAP7_75t_L g1610 ( .A(n_961), .Y(n_1610) );
BUFx8_ASAP7_75t_SL g961 ( .A(n_962), .Y(n_961) );
INVx2_ASAP7_75t_L g1522 ( .A(n_962), .Y(n_1522) );
OAI22xp33_ASAP7_75t_L g1049 ( .A1(n_970), .A2(n_1050), .B1(n_1051), .B2(n_1063), .Y(n_1049) );
OAI221xp5_ASAP7_75t_L g1213 ( .A1(n_972), .A2(n_1187), .B1(n_1189), .B2(n_1214), .C(n_1216), .Y(n_1213) );
INVx2_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
INVx1_ASAP7_75t_SL g1042 ( .A(n_985), .Y(n_1042) );
NAND4xp75_ASAP7_75t_L g985 ( .A(n_986), .B(n_1008), .C(n_1013), .D(n_1038), .Y(n_985) );
INVx1_ASAP7_75t_L g990 ( .A(n_991), .Y(n_990) );
OAI211xp5_ASAP7_75t_L g1028 ( .A1(n_994), .A2(n_1029), .B(n_1030), .C(n_1032), .Y(n_1028) );
BUFx3_ASAP7_75t_L g1255 ( .A(n_995), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g999 ( .A1(n_1000), .A2(n_1001), .B1(n_1003), .B2(n_1004), .Y(n_999) );
BUFx2_ASAP7_75t_L g1001 ( .A(n_1002), .Y(n_1001) );
INVx1_ASAP7_75t_L g1006 ( .A(n_1007), .Y(n_1006) );
NOR2x1_ASAP7_75t_L g1008 ( .A(n_1009), .B(n_1012), .Y(n_1008) );
NAND2xp5_ASAP7_75t_L g1019 ( .A(n_1020), .B(n_1028), .Y(n_1019) );
OAI211xp5_ASAP7_75t_L g1020 ( .A1(n_1021), .A2(n_1022), .B(n_1025), .C(n_1026), .Y(n_1020) );
INVx1_ASAP7_75t_L g1022 ( .A(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g1023 ( .A(n_1024), .Y(n_1023) );
HB1xp67_ASAP7_75t_L g1224 ( .A(n_1031), .Y(n_1224) );
INVxp67_ASAP7_75t_SL g1109 ( .A(n_1043), .Y(n_1109) );
XNOR2xp5_ASAP7_75t_L g1043 ( .A(n_1044), .B(n_1045), .Y(n_1043) );
AND4x1_ASAP7_75t_L g1045 ( .A(n_1046), .B(n_1048), .C(n_1073), .D(n_1105), .Y(n_1045) );
NOR3xp33_ASAP7_75t_L g1048 ( .A(n_1049), .B(n_1071), .C(n_1072), .Y(n_1048) );
OAI221xp5_ASAP7_75t_L g1051 ( .A1(n_1052), .A2(n_1053), .B1(n_1054), .B2(n_1057), .C(n_1058), .Y(n_1051) );
INVx2_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
INVx1_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
INVx1_ASAP7_75t_L g1060 ( .A(n_1061), .Y(n_1060) );
INVx1_ASAP7_75t_L g1061 ( .A(n_1062), .Y(n_1061) );
HB1xp67_ASAP7_75t_L g1165 ( .A(n_1062), .Y(n_1165) );
OAI221xp5_ASAP7_75t_L g1063 ( .A1(n_1064), .A2(n_1065), .B1(n_1066), .B2(n_1068), .C(n_1069), .Y(n_1063) );
INVx2_ASAP7_75t_L g1066 ( .A(n_1067), .Y(n_1066) );
INVx2_ASAP7_75t_L g1079 ( .A(n_1080), .Y(n_1079) );
OAI22xp5_ASAP7_75t_L g1081 ( .A1(n_1082), .A2(n_1084), .B1(n_1085), .B2(n_1088), .Y(n_1081) );
BUFx2_ASAP7_75t_L g1082 ( .A(n_1083), .Y(n_1082) );
OAI22xp5_ASAP7_75t_L g1248 ( .A1(n_1085), .A2(n_1249), .B1(n_1251), .B2(n_1252), .Y(n_1248) );
INVx2_ASAP7_75t_SL g1085 ( .A(n_1086), .Y(n_1085) );
INVx1_ASAP7_75t_L g1086 ( .A(n_1087), .Y(n_1086) );
INVx2_ASAP7_75t_L g1094 ( .A(n_1095), .Y(n_1094) );
INVx2_ASAP7_75t_SL g1133 ( .A(n_1095), .Y(n_1133) );
INVx1_ASAP7_75t_L g1096 ( .A(n_1097), .Y(n_1096) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_1100), .A2(n_1102), .B1(n_1103), .B2(n_1104), .Y(n_1099) );
HB1xp67_ASAP7_75t_L g1100 ( .A(n_1101), .Y(n_1100) );
NOR2xp33_ASAP7_75t_L g1105 ( .A(n_1106), .B(n_1107), .Y(n_1105) );
INVx1_ASAP7_75t_L g1169 ( .A(n_1110), .Y(n_1169) );
XNOR2x1_ASAP7_75t_L g1110 ( .A(n_1111), .B(n_1112), .Y(n_1110) );
AND2x4_ASAP7_75t_L g1112 ( .A(n_1113), .B(n_1142), .Y(n_1112) );
AND4x1_ASAP7_75t_L g1113 ( .A(n_1114), .B(n_1120), .C(n_1124), .D(n_1128), .Y(n_1113) );
INVx1_ASAP7_75t_L g1117 ( .A(n_1118), .Y(n_1117) );
BUFx3_ASAP7_75t_L g1129 ( .A(n_1130), .Y(n_1129) );
INVx2_ASAP7_75t_L g1193 ( .A(n_1130), .Y(n_1193) );
INVx3_ASAP7_75t_L g1136 ( .A(n_1137), .Y(n_1136) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1139), .Y(n_1565) );
INVx2_ASAP7_75t_SL g1149 ( .A(n_1150), .Y(n_1149) );
INVx1_ASAP7_75t_L g1158 ( .A(n_1159), .Y(n_1158) );
INVx2_ASAP7_75t_L g1162 ( .A(n_1163), .Y(n_1162) );
INVx1_ASAP7_75t_L g1163 ( .A(n_1164), .Y(n_1163) );
INVx1_ASAP7_75t_L g1170 ( .A(n_1171), .Y(n_1170) );
AOI22xp5_ASAP7_75t_L g1171 ( .A1(n_1172), .A2(n_1173), .B1(n_1231), .B2(n_1292), .Y(n_1171) );
INVx1_ASAP7_75t_L g1172 ( .A(n_1173), .Y(n_1172) );
INVx1_ASAP7_75t_L g1173 ( .A(n_1174), .Y(n_1173) );
HB1xp67_ASAP7_75t_L g1174 ( .A(n_1175), .Y(n_1174) );
INVx2_ASAP7_75t_L g1176 ( .A(n_1177), .Y(n_1176) );
AND2x2_ASAP7_75t_L g1177 ( .A(n_1178), .B(n_1202), .Y(n_1177) );
AND4x1_ASAP7_75t_L g1178 ( .A(n_1179), .B(n_1185), .C(n_1188), .D(n_1191), .Y(n_1178) );
INVx1_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx2_ASAP7_75t_L g1192 ( .A(n_1193), .Y(n_1192) );
INVx1_ASAP7_75t_L g1199 ( .A(n_1200), .Y(n_1199) );
AOI21xp33_ASAP7_75t_SL g1202 ( .A1(n_1203), .A2(n_1204), .B(n_1205), .Y(n_1202) );
AOI31xp33_ASAP7_75t_L g1205 ( .A1(n_1206), .A2(n_1218), .A3(n_1226), .B(n_1229), .Y(n_1205) );
INVx1_ASAP7_75t_L g1280 ( .A(n_1209), .Y(n_1280) );
INVx1_ASAP7_75t_L g1214 ( .A(n_1215), .Y(n_1214) );
INVx1_ASAP7_75t_L g1216 ( .A(n_1217), .Y(n_1216) );
BUFx2_ASAP7_75t_L g1288 ( .A(n_1217), .Y(n_1288) );
INVx1_ASAP7_75t_L g1221 ( .A(n_1222), .Y(n_1221) );
INVx1_ASAP7_75t_L g1231 ( .A(n_1232), .Y(n_1231) );
INVx1_ASAP7_75t_L g1232 ( .A(n_1233), .Y(n_1232) );
INVx1_ASAP7_75t_L g1292 ( .A(n_1233), .Y(n_1292) );
HB1xp67_ASAP7_75t_L g1233 ( .A(n_1234), .Y(n_1233) );
INVx1_ASAP7_75t_L g1234 ( .A(n_1235), .Y(n_1234) );
INVx1_ASAP7_75t_L g1290 ( .A(n_1236), .Y(n_1290) );
NOR3xp33_ASAP7_75t_L g1238 ( .A(n_1239), .B(n_1246), .C(n_1247), .Y(n_1238) );
NAND2xp5_ASAP7_75t_L g1239 ( .A(n_1240), .B(n_1243), .Y(n_1239) );
OAI221xp5_ASAP7_75t_L g1282 ( .A1(n_1241), .A2(n_1245), .B1(n_1272), .B2(n_1283), .C(n_1285), .Y(n_1282) );
OAI22xp5_ASAP7_75t_L g1257 ( .A1(n_1249), .A2(n_1258), .B1(n_1259), .B2(n_1261), .Y(n_1257) );
INVx2_ASAP7_75t_L g1249 ( .A(n_1250), .Y(n_1249) );
OAI221xp5_ASAP7_75t_L g1269 ( .A1(n_1252), .A2(n_1254), .B1(n_1270), .B2(n_1272), .C(n_1273), .Y(n_1269) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1260), .Y(n_1259) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1260), .Y(n_1570) );
INVx1_ASAP7_75t_L g1270 ( .A(n_1271), .Y(n_1270) );
INVx1_ASAP7_75t_L g1283 ( .A(n_1284), .Y(n_1283) );
INVx1_ASAP7_75t_L g1286 ( .A(n_1287), .Y(n_1286) );
OAI22xp33_ASAP7_75t_L g1309 ( .A1(n_1291), .A2(n_1310), .B1(n_1315), .B2(n_1316), .Y(n_1309) );
OAI221xp5_ASAP7_75t_L g1293 ( .A1(n_1294), .A2(n_1514), .B1(n_1518), .B2(n_1572), .C(n_1577), .Y(n_1293) );
AND4x1_ASAP7_75t_L g1294 ( .A(n_1295), .B(n_1427), .C(n_1462), .D(n_1492), .Y(n_1294) );
A2O1A1Ixp33_ASAP7_75t_L g1295 ( .A1(n_1296), .A2(n_1380), .B(n_1381), .C(n_1411), .Y(n_1295) );
OAI211xp5_ASAP7_75t_SL g1296 ( .A1(n_1297), .A2(n_1329), .B(n_1359), .C(n_1362), .Y(n_1296) );
OR2x2_ASAP7_75t_L g1297 ( .A(n_1298), .B(n_1319), .Y(n_1297) );
NAND2xp5_ASAP7_75t_L g1403 ( .A(n_1298), .B(n_1377), .Y(n_1403) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_1298), .B(n_1320), .Y(n_1408) );
AND2x4_ASAP7_75t_SL g1503 ( .A(n_1298), .B(n_1319), .Y(n_1503) );
INVx2_ASAP7_75t_SL g1298 ( .A(n_1299), .Y(n_1298) );
AND2x2_ASAP7_75t_L g1375 ( .A(n_1299), .B(n_1319), .Y(n_1375) );
INVx2_ASAP7_75t_L g1380 ( .A(n_1299), .Y(n_1380) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1300), .Y(n_1392) );
AND2x4_ASAP7_75t_L g1300 ( .A(n_1301), .B(n_1304), .Y(n_1300) );
AND2x2_ASAP7_75t_L g1322 ( .A(n_1301), .B(n_1304), .Y(n_1322) );
HB1xp67_ASAP7_75t_L g1641 ( .A(n_1301), .Y(n_1641) );
INVx1_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
AND2x4_ASAP7_75t_L g1308 ( .A(n_1302), .B(n_1304), .Y(n_1308) );
INVx1_ASAP7_75t_L g1302 ( .A(n_1303), .Y(n_1302) );
NAND2xp5_ASAP7_75t_L g1313 ( .A(n_1303), .B(n_1314), .Y(n_1313) );
INVx1_ASAP7_75t_L g1314 ( .A(n_1305), .Y(n_1314) );
INVx2_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
INVx1_ASAP7_75t_L g1517 ( .A(n_1307), .Y(n_1517) );
INVx2_ASAP7_75t_L g1307 ( .A(n_1308), .Y(n_1307) );
OAI22xp5_ASAP7_75t_L g1345 ( .A1(n_1310), .A2(n_1317), .B1(n_1346), .B2(n_1347), .Y(n_1345) );
BUFx3_ASAP7_75t_L g1394 ( .A(n_1310), .Y(n_1394) );
BUFx6f_ASAP7_75t_L g1310 ( .A(n_1311), .Y(n_1310) );
OR2x2_ASAP7_75t_L g1311 ( .A(n_1312), .B(n_1313), .Y(n_1311) );
OR2x2_ASAP7_75t_L g1317 ( .A(n_1312), .B(n_1318), .Y(n_1317) );
INVx1_ASAP7_75t_L g1326 ( .A(n_1312), .Y(n_1326) );
INVx1_ASAP7_75t_L g1325 ( .A(n_1313), .Y(n_1325) );
HB1xp67_ASAP7_75t_L g1643 ( .A(n_1314), .Y(n_1643) );
HB1xp67_ASAP7_75t_L g1316 ( .A(n_1317), .Y(n_1316) );
INVx1_ASAP7_75t_L g1397 ( .A(n_1317), .Y(n_1397) );
INVx1_ASAP7_75t_L g1328 ( .A(n_1318), .Y(n_1328) );
AND2x2_ASAP7_75t_L g1365 ( .A(n_1319), .B(n_1354), .Y(n_1365) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_1319), .B(n_1378), .Y(n_1416) );
OAI221xp5_ASAP7_75t_L g1463 ( .A1(n_1319), .A2(n_1445), .B1(n_1464), .B2(n_1466), .C(n_1468), .Y(n_1463) );
AND2x2_ASAP7_75t_L g1471 ( .A(n_1319), .B(n_1429), .Y(n_1471) );
CKINVDCx6p67_ASAP7_75t_R g1319 ( .A(n_1320), .Y(n_1319) );
AND2x2_ASAP7_75t_L g1387 ( .A(n_1320), .B(n_1388), .Y(n_1387) );
AND2x2_ASAP7_75t_L g1400 ( .A(n_1320), .B(n_1354), .Y(n_1400) );
NAND2xp5_ASAP7_75t_L g1432 ( .A(n_1320), .B(n_1433), .Y(n_1432) );
AOI221xp5_ASAP7_75t_L g1479 ( .A1(n_1320), .A2(n_1360), .B1(n_1480), .B2(n_1483), .C(n_1485), .Y(n_1479) );
A2O1A1Ixp33_ASAP7_75t_L g1493 ( .A1(n_1320), .A2(n_1447), .B(n_1494), .C(n_1495), .Y(n_1493) );
AOI221xp5_ASAP7_75t_L g1495 ( .A1(n_1320), .A2(n_1387), .B1(n_1439), .B2(n_1496), .C(n_1497), .Y(n_1495) );
OR2x6_ASAP7_75t_L g1320 ( .A(n_1321), .B(n_1323), .Y(n_1320) );
AND2x4_ASAP7_75t_L g1324 ( .A(n_1325), .B(n_1326), .Y(n_1324) );
AND2x4_ASAP7_75t_L g1327 ( .A(n_1326), .B(n_1328), .Y(n_1327) );
AOI211xp5_ASAP7_75t_L g1329 ( .A1(n_1330), .A2(n_1338), .B(n_1348), .C(n_1352), .Y(n_1329) );
AND2x2_ASAP7_75t_L g1405 ( .A(n_1330), .B(n_1406), .Y(n_1405) );
NAND2xp5_ASAP7_75t_L g1448 ( .A(n_1330), .B(n_1350), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1465 ( .A(n_1330), .B(n_1339), .Y(n_1465) );
AND2x2_ASAP7_75t_L g1330 ( .A(n_1331), .B(n_1334), .Y(n_1330) );
NAND2xp5_ASAP7_75t_L g1349 ( .A(n_1331), .B(n_1350), .Y(n_1349) );
INVx4_ASAP7_75t_L g1357 ( .A(n_1331), .Y(n_1357) );
INVx3_ASAP7_75t_L g1370 ( .A(n_1331), .Y(n_1370) );
NOR2xp67_ASAP7_75t_SL g1421 ( .A(n_1331), .B(n_1422), .Y(n_1421) );
NOR2xp33_ASAP7_75t_L g1455 ( .A(n_1331), .B(n_1456), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1477 ( .A(n_1331), .B(n_1339), .Y(n_1477) );
OR2x2_ASAP7_75t_L g1505 ( .A(n_1331), .B(n_1354), .Y(n_1505) );
AND2x4_ASAP7_75t_L g1331 ( .A(n_1332), .B(n_1333), .Y(n_1331) );
AND2x2_ASAP7_75t_L g1360 ( .A(n_1334), .B(n_1361), .Y(n_1360) );
OR2x2_ASAP7_75t_L g1371 ( .A(n_1334), .B(n_1372), .Y(n_1371) );
NAND2xp5_ASAP7_75t_L g1422 ( .A(n_1334), .B(n_1343), .Y(n_1422) );
NOR2xp33_ASAP7_75t_L g1430 ( .A(n_1334), .B(n_1343), .Y(n_1430) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_1334), .B(n_1477), .Y(n_1476) );
BUFx3_ASAP7_75t_L g1334 ( .A(n_1335), .Y(n_1334) );
INVx2_ASAP7_75t_L g1386 ( .A(n_1335), .Y(n_1386) );
AND2x2_ASAP7_75t_L g1401 ( .A(n_1335), .B(n_1372), .Y(n_1401) );
AND2x2_ASAP7_75t_L g1410 ( .A(n_1335), .B(n_1350), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1335), .B(n_1339), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1443 ( .A(n_1335), .B(n_1406), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1491 ( .A(n_1335), .B(n_1460), .Y(n_1491) );
AND2x2_ASAP7_75t_L g1335 ( .A(n_1336), .B(n_1337), .Y(n_1335) );
AOI21xp33_ASAP7_75t_L g1424 ( .A1(n_1338), .A2(n_1425), .B(n_1426), .Y(n_1424) );
AOI21xp5_ASAP7_75t_L g1490 ( .A1(n_1338), .A2(n_1426), .B(n_1491), .Y(n_1490) );
INVx1_ASAP7_75t_L g1338 ( .A(n_1339), .Y(n_1338) );
NAND2xp5_ASAP7_75t_L g1384 ( .A(n_1339), .B(n_1385), .Y(n_1384) );
NAND2xp5_ASAP7_75t_L g1482 ( .A(n_1339), .B(n_1370), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1339 ( .A(n_1340), .B(n_1343), .Y(n_1339) );
INVx1_ASAP7_75t_L g1351 ( .A(n_1340), .Y(n_1351) );
INVx1_ASAP7_75t_L g1372 ( .A(n_1340), .Y(n_1372) );
AND2x2_ASAP7_75t_L g1406 ( .A(n_1340), .B(n_1344), .Y(n_1406) );
AND2x2_ASAP7_75t_L g1358 ( .A(n_1343), .B(n_1351), .Y(n_1358) );
INVx2_ASAP7_75t_L g1366 ( .A(n_1343), .Y(n_1366) );
AND2x2_ASAP7_75t_L g1489 ( .A(n_1343), .B(n_1386), .Y(n_1489) );
INVx2_ASAP7_75t_L g1343 ( .A(n_1344), .Y(n_1343) );
AND2x2_ASAP7_75t_L g1350 ( .A(n_1344), .B(n_1351), .Y(n_1350) );
INVx1_ASAP7_75t_L g1348 ( .A(n_1349), .Y(n_1348) );
AND2x2_ASAP7_75t_L g1361 ( .A(n_1350), .B(n_1357), .Y(n_1361) );
INVx1_ASAP7_75t_L g1460 ( .A(n_1350), .Y(n_1460) );
AND2x2_ASAP7_75t_L g1467 ( .A(n_1350), .B(n_1385), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1352 ( .A(n_1353), .B(n_1358), .Y(n_1352) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1353), .Y(n_1498) );
AND2x2_ASAP7_75t_L g1353 ( .A(n_1354), .B(n_1357), .Y(n_1353) );
CKINVDCx5p33_ASAP7_75t_R g1378 ( .A(n_1354), .Y(n_1378) );
INVx1_ASAP7_75t_SL g1388 ( .A(n_1354), .Y(n_1388) );
INVx1_ASAP7_75t_L g1423 ( .A(n_1354), .Y(n_1423) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1354), .Y(n_1452) );
AND2x2_ASAP7_75t_L g1354 ( .A(n_1355), .B(n_1356), .Y(n_1354) );
NAND2xp5_ASAP7_75t_L g1364 ( .A(n_1357), .B(n_1365), .Y(n_1364) );
AND2x2_ASAP7_75t_L g1385 ( .A(n_1357), .B(n_1386), .Y(n_1385) );
AND2x2_ASAP7_75t_L g1414 ( .A(n_1357), .B(n_1415), .Y(n_1414) );
INVx1_ASAP7_75t_L g1429 ( .A(n_1357), .Y(n_1429) );
AND2x2_ASAP7_75t_L g1439 ( .A(n_1357), .B(n_1440), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1461 ( .A(n_1357), .B(n_1387), .Y(n_1461) );
AND2x2_ASAP7_75t_L g1500 ( .A(n_1357), .B(n_1400), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1446 ( .A(n_1358), .B(n_1386), .Y(n_1446) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1358), .Y(n_1506) );
NAND2xp5_ASAP7_75t_L g1511 ( .A(n_1358), .B(n_1512), .Y(n_1511) );
INVx1_ASAP7_75t_L g1359 ( .A(n_1360), .Y(n_1359) );
AOI221xp5_ASAP7_75t_L g1413 ( .A1(n_1361), .A2(n_1365), .B1(n_1414), .B2(n_1416), .C(n_1417), .Y(n_1413) );
A2O1A1Ixp33_ASAP7_75t_L g1362 ( .A1(n_1363), .A2(n_1366), .B(n_1367), .C(n_1373), .Y(n_1362) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1418 ( .A(n_1365), .B(n_1405), .Y(n_1418) );
A2O1A1Ixp33_ASAP7_75t_L g1486 ( .A1(n_1365), .A2(n_1389), .B(n_1487), .C(n_1490), .Y(n_1486) );
INVxp67_ASAP7_75t_L g1367 ( .A(n_1368), .Y(n_1367) );
OR2x2_ASAP7_75t_L g1368 ( .A(n_1369), .B(n_1371), .Y(n_1368) );
NAND2xp5_ASAP7_75t_L g1426 ( .A(n_1369), .B(n_1416), .Y(n_1426) );
A2O1A1Ixp33_ASAP7_75t_L g1507 ( .A1(n_1369), .A2(n_1508), .B(n_1509), .C(n_1510), .Y(n_1507) );
INVx2_ASAP7_75t_L g1369 ( .A(n_1370), .Y(n_1369) );
NOR2xp33_ASAP7_75t_L g1436 ( .A(n_1370), .B(n_1437), .Y(n_1436) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1370), .B(n_1446), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1450 ( .A(n_1370), .B(n_1430), .Y(n_1450) );
NAND2xp5_ASAP7_75t_L g1488 ( .A(n_1370), .B(n_1489), .Y(n_1488) );
NOR2x1_ASAP7_75t_L g1415 ( .A(n_1372), .B(n_1386), .Y(n_1415) );
NAND2xp5_ASAP7_75t_L g1425 ( .A(n_1372), .B(n_1386), .Y(n_1425) );
NAND2xp5_ASAP7_75t_L g1373 ( .A(n_1374), .B(n_1376), .Y(n_1373) );
INVx1_ASAP7_75t_L g1374 ( .A(n_1375), .Y(n_1374) );
NAND2xp5_ASAP7_75t_L g1376 ( .A(n_1377), .B(n_1379), .Y(n_1376) );
AOI321xp33_ASAP7_75t_L g1427 ( .A1(n_1377), .A2(n_1387), .A3(n_1428), .B1(n_1431), .B2(n_1434), .C(n_1444), .Y(n_1427) );
OR2x2_ASAP7_75t_L g1447 ( .A(n_1377), .B(n_1448), .Y(n_1447) );
NOR2xp33_ASAP7_75t_L g1466 ( .A(n_1377), .B(n_1467), .Y(n_1466) );
INVx3_ASAP7_75t_L g1377 ( .A(n_1378), .Y(n_1377) );
NOR2xp33_ASAP7_75t_L g1464 ( .A(n_1378), .B(n_1465), .Y(n_1464) );
NAND2xp5_ASAP7_75t_L g1513 ( .A(n_1378), .B(n_1503), .Y(n_1513) );
NAND2xp5_ASAP7_75t_L g1398 ( .A(n_1379), .B(n_1390), .Y(n_1398) );
NOR2xp33_ASAP7_75t_L g1412 ( .A(n_1379), .B(n_1390), .Y(n_1412) );
AOI21xp5_ASAP7_75t_SL g1492 ( .A1(n_1379), .A2(n_1493), .B(n_1501), .Y(n_1492) );
NOR3xp33_ASAP7_75t_L g1504 ( .A(n_1379), .B(n_1505), .C(n_1506), .Y(n_1504) );
INVx2_ASAP7_75t_L g1379 ( .A(n_1380), .Y(n_1379) );
AND2x2_ASAP7_75t_L g1399 ( .A(n_1380), .B(n_1400), .Y(n_1399) );
INVx2_ASAP7_75t_L g1442 ( .A(n_1380), .Y(n_1442) );
INVxp67_ASAP7_75t_SL g1381 ( .A(n_1382), .Y(n_1381) );
OAI211xp5_ASAP7_75t_L g1411 ( .A1(n_1382), .A2(n_1412), .B(n_1413), .C(n_1419), .Y(n_1411) );
AOI221xp5_ASAP7_75t_L g1382 ( .A1(n_1383), .A2(n_1398), .B1(n_1399), .B2(n_1401), .C(n_1402), .Y(n_1382) );
OAI21xp33_ASAP7_75t_SL g1383 ( .A1(n_1384), .A2(n_1387), .B(n_1389), .Y(n_1383) );
AND2x2_ASAP7_75t_L g1440 ( .A(n_1386), .B(n_1406), .Y(n_1440) );
OR2x2_ASAP7_75t_L g1481 ( .A(n_1386), .B(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1473 ( .A(n_1387), .Y(n_1473) );
A2O1A1Ixp33_ASAP7_75t_L g1434 ( .A1(n_1389), .A2(n_1435), .B(n_1438), .C(n_1441), .Y(n_1434) );
INVx2_ASAP7_75t_L g1457 ( .A(n_1389), .Y(n_1457) );
BUFx3_ASAP7_75t_L g1389 ( .A(n_1390), .Y(n_1389) );
INVx1_ASAP7_75t_L g1433 ( .A(n_1390), .Y(n_1433) );
AOI21xp5_ASAP7_75t_L g1449 ( .A1(n_1390), .A2(n_1450), .B(n_1451), .Y(n_1449) );
AOI31xp33_ASAP7_75t_L g1501 ( .A1(n_1390), .A2(n_1502), .A3(n_1507), .B(n_1511), .Y(n_1501) );
INVx1_ASAP7_75t_L g1391 ( .A(n_1392), .Y(n_1391) );
INVx1_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
INVx1_ASAP7_75t_L g1474 ( .A(n_1398), .Y(n_1474) );
INVx1_ASAP7_75t_L g1478 ( .A(n_1399), .Y(n_1478) );
AND2x2_ASAP7_75t_L g1485 ( .A(n_1399), .B(n_1410), .Y(n_1485) );
AOI21xp33_ASAP7_75t_L g1454 ( .A1(n_1400), .A2(n_1455), .B(n_1457), .Y(n_1454) );
NAND2xp5_ASAP7_75t_L g1499 ( .A(n_1401), .B(n_1500), .Y(n_1499) );
OAI22xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1404), .B1(n_1407), .B2(n_1409), .Y(n_1402) );
INVx1_ASAP7_75t_L g1510 ( .A(n_1403), .Y(n_1510) );
INVx1_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVx1_ASAP7_75t_L g1456 ( .A(n_1406), .Y(n_1456) );
NAND2xp5_ASAP7_75t_SL g1483 ( .A(n_1407), .B(n_1484), .Y(n_1483) );
INVx2_ASAP7_75t_L g1407 ( .A(n_1408), .Y(n_1407) );
AOI221xp5_ASAP7_75t_L g1502 ( .A1(n_1408), .A2(n_1420), .B1(n_1421), .B2(n_1503), .C(n_1504), .Y(n_1502) );
INVx1_ASAP7_75t_L g1409 ( .A(n_1410), .Y(n_1409) );
OAI21xp5_ASAP7_75t_L g1453 ( .A1(n_1414), .A2(n_1416), .B(n_1421), .Y(n_1453) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1415), .Y(n_1437) );
INVx1_ASAP7_75t_L g1417 ( .A(n_1418), .Y(n_1417) );
O2A1O1Ixp33_ASAP7_75t_L g1419 ( .A1(n_1420), .A2(n_1421), .B(n_1423), .C(n_1424), .Y(n_1419) );
NAND2xp5_ASAP7_75t_SL g1469 ( .A(n_1422), .B(n_1470), .Y(n_1469) );
INVx1_ASAP7_75t_L g1484 ( .A(n_1423), .Y(n_1484) );
INVx1_ASAP7_75t_L g1508 ( .A(n_1425), .Y(n_1508) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1430), .Y(n_1428) );
AOI331xp33_ASAP7_75t_L g1444 ( .A1(n_1431), .A2(n_1445), .A3(n_1447), .B1(n_1449), .B2(n_1453), .B3(n_1454), .C1(n_1458), .Y(n_1444) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
INVx1_ASAP7_75t_L g1435 ( .A(n_1436), .Y(n_1435) );
INVxp67_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
INVx1_ASAP7_75t_L g1470 ( .A(n_1440), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1441 ( .A(n_1442), .B(n_1443), .Y(n_1441) );
NOR2xp33_ASAP7_75t_L g1472 ( .A(n_1446), .B(n_1473), .Y(n_1472) );
INVx1_ASAP7_75t_L g1451 ( .A(n_1452), .Y(n_1451) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
NOR2xp33_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1461), .Y(n_1459) );
AOI21xp5_ASAP7_75t_L g1462 ( .A1(n_1463), .A2(n_1474), .B(n_1475), .Y(n_1462) );
INVx1_ASAP7_75t_L g1494 ( .A(n_1465), .Y(n_1494) );
AOI21xp5_ASAP7_75t_SL g1468 ( .A1(n_1469), .A2(n_1471), .B(n_1472), .Y(n_1468) );
OAI21xp33_ASAP7_75t_L g1497 ( .A1(n_1470), .A2(n_1498), .B(n_1499), .Y(n_1497) );
OAI211xp5_ASAP7_75t_SL g1475 ( .A1(n_1476), .A2(n_1478), .B(n_1479), .C(n_1486), .Y(n_1475) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1476), .Y(n_1496) );
INVx1_ASAP7_75t_L g1480 ( .A(n_1481), .Y(n_1480) );
INVx1_ASAP7_75t_L g1487 ( .A(n_1488), .Y(n_1487) );
INVx1_ASAP7_75t_L g1509 ( .A(n_1491), .Y(n_1509) );
INVx1_ASAP7_75t_L g1512 ( .A(n_1513), .Y(n_1512) );
CKINVDCx5p33_ASAP7_75t_R g1514 ( .A(n_1515), .Y(n_1514) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1516), .Y(n_1515) );
INVx1_ASAP7_75t_L g1516 ( .A(n_1517), .Y(n_1516) );
BUFx2_ASAP7_75t_L g1519 ( .A(n_1520), .Y(n_1519) );
AND2x2_ASAP7_75t_L g1520 ( .A(n_1521), .B(n_1547), .Y(n_1520) );
AOI22xp5_ASAP7_75t_L g1521 ( .A1(n_1522), .A2(n_1523), .B1(n_1545), .B2(n_1546), .Y(n_1521) );
NAND3xp33_ASAP7_75t_L g1523 ( .A(n_1524), .B(n_1534), .C(n_1542), .Y(n_1523) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
OAI22xp5_ASAP7_75t_L g1566 ( .A1(n_1531), .A2(n_1544), .B1(n_1567), .B2(n_1570), .Y(n_1566) );
INVx1_ASAP7_75t_L g1536 ( .A(n_1537), .Y(n_1536) );
INVx2_ASAP7_75t_L g1538 ( .A(n_1539), .Y(n_1538) );
INVx1_ASAP7_75t_L g1597 ( .A(n_1539), .Y(n_1597) );
NOR3xp33_ASAP7_75t_L g1547 ( .A(n_1548), .B(n_1556), .C(n_1557), .Y(n_1547) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1549), .B(n_1553), .Y(n_1548) );
INVx1_ASAP7_75t_L g1567 ( .A(n_1568), .Y(n_1567) );
INVx1_ASAP7_75t_L g1568 ( .A(n_1569), .Y(n_1568) );
CKINVDCx14_ASAP7_75t_R g1572 ( .A(n_1573), .Y(n_1572) );
INVx2_ASAP7_75t_L g1573 ( .A(n_1574), .Y(n_1573) );
CKINVDCx5p33_ASAP7_75t_R g1574 ( .A(n_1575), .Y(n_1574) );
A2O1A1Ixp33_ASAP7_75t_L g1639 ( .A1(n_1576), .A2(n_1640), .B(n_1642), .C(n_1644), .Y(n_1639) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1579 ( .A(n_1580), .Y(n_1579) );
INVx1_ASAP7_75t_L g1580 ( .A(n_1581), .Y(n_1580) );
INVx1_ASAP7_75t_L g1581 ( .A(n_1582), .Y(n_1581) );
INVx1_ASAP7_75t_L g1583 ( .A(n_1584), .Y(n_1583) );
INVx2_ASAP7_75t_SL g1636 ( .A(n_1585), .Y(n_1636) );
AND2x2_ASAP7_75t_L g1585 ( .A(n_1586), .B(n_1611), .Y(n_1585) );
OAI21xp33_ASAP7_75t_L g1586 ( .A1(n_1587), .A2(n_1601), .B(n_1610), .Y(n_1586) );
AOI22xp5_ASAP7_75t_L g1588 ( .A1(n_1589), .A2(n_1591), .B1(n_1595), .B2(n_1596), .Y(n_1588) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
OAI22xp33_ASAP7_75t_L g1630 ( .A1(n_1599), .A2(n_1631), .B1(n_1632), .B2(n_1633), .Y(n_1630) );
INVx2_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
NOR2xp33_ASAP7_75t_L g1611 ( .A(n_1612), .B(n_1623), .Y(n_1611) );
NAND2xp5_ASAP7_75t_L g1623 ( .A(n_1624), .B(n_1627), .Y(n_1623) );
BUFx2_ASAP7_75t_L g1637 ( .A(n_1638), .Y(n_1637) );
HB1xp67_ASAP7_75t_L g1638 ( .A(n_1639), .Y(n_1638) );
INVx1_ASAP7_75t_L g1640 ( .A(n_1641), .Y(n_1640) );
INVx1_ASAP7_75t_L g1642 ( .A(n_1643), .Y(n_1642) );
endmodule