module real_aes_3835_n_296 (n_17, n_28, n_226, n_76, n_202, n_255, n_149, n_286, n_56, n_1078, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_257, n_261, n_262, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_285, n_134, n_32, n_30, n_263, n_230, n_165, n_51, n_195, n_246, n_248, n_252, n_283, n_176, n_27, n_163, n_222, n_249, n_61, n_29, n_20, n_52, n_221, n_287, n_174, n_156, n_57, n_64, n_66, n_254, n_1077, n_18, n_207, n_104, n_21, n_31, n_8, n_251, n_183, n_266, n_205, n_220, n_211, n_10, n_281, n_177, n_83, n_181, n_197, n_293, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_284, n_75, n_178, n_219, n_256, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_253, n_35, n_42, n_147, n_150, n_288, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_274, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_269, n_152, n_198, n_201, n_122, n_7, n_228, n_272, n_196, n_141, n_1079, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_275, n_69, n_279, n_46, n_109, n_59, n_25, n_203, n_236, n_278, n_73, n_77, n_218, n_81, n_133, n_48, n_267, n_270, n_260, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_273, n_138, n_50, n_114, n_276, n_89, n_295, n_170, n_277, n_26, n_235, n_265, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_271, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_294, n_227, n_67, n_92, n_33, n_206, n_258, n_291, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_250, n_292, n_116, n_94, n_229, n_289, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_280, n_38, n_290, n_259, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_268, n_136, n_87, n_171, n_0, n_157, n_78, n_264, n_282, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_296);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_255;
input n_149;
input n_286;
input n_56;
input n_1078;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_257;
input n_261;
input n_262;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_285;
input n_134;
input n_32;
input n_30;
input n_263;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_252;
input n_283;
input n_176;
input n_27;
input n_163;
input n_222;
input n_249;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_287;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_254;
input n_1077;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_251;
input n_183;
input n_266;
input n_205;
input n_220;
input n_211;
input n_10;
input n_281;
input n_177;
input n_83;
input n_181;
input n_197;
input n_293;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_284;
input n_75;
input n_178;
input n_219;
input n_256;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_253;
input n_35;
input n_42;
input n_147;
input n_150;
input n_288;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_274;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_269;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_272;
input n_196;
input n_141;
input n_1079;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_275;
input n_69;
input n_279;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_278;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_267;
input n_270;
input n_260;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_273;
input n_138;
input n_50;
input n_114;
input n_276;
input n_89;
input n_295;
input n_170;
input n_277;
input n_26;
input n_235;
input n_265;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_271;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_294;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_258;
input n_291;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_250;
input n_292;
input n_116;
input n_94;
input n_229;
input n_289;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_280;
input n_38;
input n_290;
input n_259;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_268;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_264;
input n_282;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_296;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_1066;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_1018;
wire n_980;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_977;
wire n_943;
wire n_357;
wire n_503;
wire n_792;
wire n_673;
wire n_386;
wire n_1067;
wire n_518;
wire n_635;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_991;
wire n_577;
wire n_580;
wire n_1004;
wire n_469;
wire n_987;
wire n_362;
wire n_759;
wire n_979;
wire n_445;
wire n_1065;
wire n_596;
wire n_592;
wire n_540;
wire n_1064;
wire n_1075;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_974;
wire n_857;
wire n_919;
wire n_461;
wire n_1047;
wire n_1016;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_1034;
wire n_952;
wire n_429;
wire n_976;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_989;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_1044;
wire n_321;
wire n_963;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_983;
wire n_767;
wire n_696;
wire n_889;
wire n_955;
wire n_975;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_1046;
wire n_677;
wire n_958;
wire n_1021;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_961;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_815;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_953;
wire n_462;
wire n_615;
wire n_990;
wire n_550;
wire n_966;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_495;
wire n_994;
wire n_892;
wire n_370;
wire n_1072;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_951;
wire n_875;
wire n_327;
wire n_774;
wire n_992;
wire n_813;
wire n_791;
wire n_981;
wire n_1053;
wire n_1049;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_984;
wire n_1019;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_1070;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_962;
wire n_468;
wire n_746;
wire n_656;
wire n_316;
wire n_532;
wire n_755;
wire n_1025;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_996;
wire n_439;
wire n_1062;
wire n_576;
wire n_924;
wire n_956;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_973;
wire n_671;
wire n_960;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_565;
wire n_443;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_1029;
wire n_1020;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_1059;
wire n_950;
wire n_381;
wire n_993;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_1013;
wire n_1017;
wire n_581;
wire n_610;
wire n_936;
wire n_1035;
wire n_620;
wire n_582;
wire n_1063;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_1042;
wire n_879;
wire n_331;
wire n_449;
wire n_363;
wire n_417;
wire n_754;
wire n_607;
wire n_1006;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_970;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_1012;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1054;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_1050;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_658;
wire n_676;
wire n_986;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_1031;
wire n_1037;
wire n_1008;
wire n_807;
wire n_1011;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_999;
wire n_619;
wire n_391;
wire n_360;
wire n_1060;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_361;
wire n_917;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_985;
wire n_501;
wire n_488;
wire n_1041;
wire n_910;
wire n_642;
wire n_613;
wire n_387;
wire n_957;
wire n_995;
wire n_954;
wire n_702;
wire n_969;
wire n_912;
wire n_1009;
wire n_1007;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_604;
wire n_734;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_1022;
wire n_404;
wire n_1073;
wire n_756;
wire n_598;
wire n_713;
wire n_728;
wire n_334;
wire n_735;
wire n_569;
wire n_303;
wire n_997;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_843;
wire n_810;
wire n_306;
wire n_579;
wire n_1033;
wire n_699;
wire n_533;
wire n_1000;
wire n_1003;
wire n_1028;
wire n_366;
wire n_346;
wire n_727;
wire n_1014;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_470;
wire n_851;
wire n_915;
wire n_1002;
wire n_934;
wire n_494;
wire n_1001;
wire n_711;
wire n_864;
wire n_1027;
wire n_377;
wire n_1058;
wire n_927;
wire n_1038;
wire n_965;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_1043;
wire n_354;
wire n_720;
wire n_968;
wire n_972;
wire n_435;
wire n_1026;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_1068;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_1023;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_1057;
wire n_411;
wire n_697;
wire n_978;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_1005;
wire n_487;
wire n_831;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_928;
wire n_899;
wire n_692;
wire n_544;
wire n_789;
wire n_1051;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_922;
wire n_926;
wire n_942;
wire n_1048;
wire n_472;
wire n_971;
wire n_866;
wire n_452;
wire n_1052;
wire n_1071;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_959;
wire n_946;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_741;
wire n_753;
wire n_314;
wire n_623;
wire n_1032;
wire n_446;
wire n_721;
wire n_681;
wire n_982;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_712;
wire n_433;
wire n_516;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_418;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_1010;
wire n_811;
wire n_1015;
wire n_459;
wire n_558;
wire n_863;
wire n_998;
wire n_724;
wire n_440;
wire n_525;
wire n_1074;
wire n_644;
wire n_674;
wire n_836;
wire n_888;
wire n_793;
wire n_1056;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_949;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_967;
wire n_837;
wire n_1045;
wire n_871;
wire n_474;
wire n_829;
wire n_1030;
wire n_988;
wire n_1055;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_1036;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_1040;
wire n_703;
wire n_652;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_1039;
wire n_424;
wire n_802;
wire n_868;
wire n_877;
wire n_574;
wire n_1069;
wire n_337;
wire n_1024;
wire n_842;
wire n_849;
wire n_1061;
wire n_554;
wire n_475;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
AOI22xp5_ASAP7_75t_L g562 ( .A1(n_0), .A2(n_164), .B1(n_534), .B2(n_563), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g770 ( .A1(n_1), .A2(n_159), .B1(n_504), .B2(n_685), .Y(n_770) );
INVx1_ASAP7_75t_L g715 ( .A(n_2), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g729 ( .A1(n_3), .A2(n_6), .B1(n_530), .B2(n_567), .Y(n_729) );
HB1xp67_ASAP7_75t_L g307 ( .A(n_4), .Y(n_307) );
AND2x4_ASAP7_75t_L g816 ( .A(n_4), .B(n_286), .Y(n_816) );
AND2x4_ASAP7_75t_L g825 ( .A(n_4), .B(n_826), .Y(n_825) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_5), .A2(n_157), .B1(n_819), .B2(n_836), .Y(n_848) );
AOI221x1_ASAP7_75t_L g670 ( .A1(n_7), .A2(n_89), .B1(n_671), .B2(n_672), .C(n_673), .Y(n_670) );
AOI22xp33_ASAP7_75t_L g517 ( .A1(n_8), .A2(n_254), .B1(n_518), .B2(n_519), .Y(n_517) );
AOI22xp5_ASAP7_75t_L g429 ( .A1(n_9), .A2(n_195), .B1(n_389), .B2(n_396), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_10), .A2(n_175), .B1(n_404), .B2(n_432), .Y(n_431) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_11), .A2(n_70), .B1(n_428), .B2(n_538), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g425 ( .A1(n_12), .A2(n_154), .B1(n_426), .B2(n_428), .Y(n_425) );
AOI22xp33_ASAP7_75t_SL g413 ( .A1(n_13), .A2(n_253), .B1(n_414), .B2(n_416), .Y(n_413) );
INVx1_ASAP7_75t_L g451 ( .A(n_14), .Y(n_451) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_15), .Y(n_686) );
AOI22xp33_ASAP7_75t_L g466 ( .A1(n_16), .A2(n_115), .B1(n_407), .B2(n_467), .Y(n_466) );
AOI22xp33_ASAP7_75t_L g576 ( .A1(n_17), .A2(n_18), .B1(n_442), .B2(n_577), .Y(n_576) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_19), .A2(n_117), .B1(n_389), .B2(n_540), .Y(n_628) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_20), .A2(n_204), .B1(n_470), .B2(n_471), .Y(n_469) );
AO22x1_ASAP7_75t_L g742 ( .A1(n_21), .A2(n_147), .B1(n_627), .B2(n_743), .Y(n_742) );
CKINVDCx20_ASAP7_75t_R g903 ( .A(n_22), .Y(n_903) );
INVxp33_ASAP7_75t_SL g829 ( .A(n_23), .Y(n_829) );
AO22x2_ASAP7_75t_L g857 ( .A1(n_24), .A2(n_81), .B1(n_819), .B2(n_836), .Y(n_857) );
XNOR2x1_ASAP7_75t_L g1032 ( .A(n_24), .B(n_1033), .Y(n_1032) );
AOI22xp33_ASAP7_75t_L g1051 ( .A1(n_24), .A2(n_1052), .B1(n_1071), .B2(n_1073), .Y(n_1051) );
INVx1_ASAP7_75t_L g480 ( .A(n_25), .Y(n_480) );
INVx1_ASAP7_75t_L g792 ( .A(n_26), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_27), .A2(n_262), .B1(n_563), .B2(n_661), .Y(n_746) );
AO22x1_ASAP7_75t_L g858 ( .A1(n_28), .A2(n_295), .B1(n_841), .B2(n_847), .Y(n_858) );
AOI211x1_ASAP7_75t_L g472 ( .A1(n_29), .A2(n_376), .B(n_473), .C(n_485), .Y(n_472) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_30), .A2(n_95), .B1(n_515), .B2(n_519), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_31), .B(n_354), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g728 ( .A1(n_32), .A2(n_103), .B1(n_410), .B2(n_677), .Y(n_728) );
INVx1_ASAP7_75t_L g548 ( .A(n_33), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g689 ( .A(n_34), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g481 ( .A1(n_35), .A2(n_151), .B1(n_482), .B2(n_483), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g750 ( .A1(n_36), .A2(n_199), .B1(n_446), .B2(n_482), .Y(n_750) );
AOI22xp5_ASAP7_75t_L g786 ( .A1(n_37), .A2(n_104), .B1(n_467), .B2(n_538), .Y(n_786) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_38), .B(n_441), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g433 ( .A1(n_39), .A2(n_289), .B1(n_434), .B2(n_435), .Y(n_433) );
AOI22xp33_ASAP7_75t_SL g676 ( .A1(n_40), .A2(n_73), .B1(n_410), .B2(n_677), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_41), .B(n_643), .Y(n_642) );
AOI22xp33_ASAP7_75t_L g765 ( .A1(n_42), .A2(n_263), .B1(n_512), .B2(n_518), .Y(n_765) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_43), .A2(n_113), .B1(n_502), .B2(n_504), .Y(n_1035) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_44), .A2(n_282), .B1(n_407), .B2(n_409), .Y(n_406) );
AOI22xp33_ASAP7_75t_L g1064 ( .A1(n_45), .A2(n_194), .B1(n_446), .B2(n_618), .Y(n_1064) );
AOI22xp33_ASAP7_75t_L g726 ( .A1(n_46), .A2(n_187), .B1(n_534), .B2(n_608), .Y(n_726) );
AOI22xp33_ASAP7_75t_L g833 ( .A1(n_47), .A2(n_149), .B1(n_813), .B2(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_48), .A2(n_100), .B1(n_530), .B2(n_531), .Y(n_529) );
AOI22xp33_ASAP7_75t_L g542 ( .A1(n_49), .A2(n_292), .B1(n_446), .B2(n_482), .Y(n_542) );
NOR2xp33_ASAP7_75t_L g305 ( .A(n_50), .B(n_230), .Y(n_305) );
INVx1_ASAP7_75t_L g338 ( .A(n_50), .Y(n_338) );
INVxp67_ASAP7_75t_L g351 ( .A(n_50), .Y(n_351) );
AOI22xp33_ASAP7_75t_L g511 ( .A1(n_51), .A2(n_174), .B1(n_512), .B2(n_513), .Y(n_511) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_52), .A2(n_244), .B1(n_819), .B2(n_869), .Y(n_868) );
INVx1_ASAP7_75t_L g718 ( .A(n_53), .Y(n_718) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_54), .A2(n_92), .B1(n_627), .B2(n_661), .Y(n_660) );
INVx1_ASAP7_75t_L g754 ( .A(n_55), .Y(n_754) );
AOI22xp33_ASAP7_75t_SL g400 ( .A1(n_56), .A2(n_76), .B1(n_401), .B2(n_404), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_57), .B(n_592), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g863 ( .A1(n_58), .A2(n_152), .B1(n_841), .B2(n_843), .Y(n_863) );
AOI21xp5_ASAP7_75t_L g1038 ( .A1(n_59), .A2(n_509), .B(n_1039), .Y(n_1038) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_60), .B(n_323), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g1069 ( .A1(n_61), .A2(n_160), .B1(n_512), .B2(n_518), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_62), .A2(n_65), .B1(n_401), .B2(n_404), .Y(n_468) );
INVx1_ASAP7_75t_L g707 ( .A(n_63), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g1068 ( .A1(n_64), .A2(n_179), .B1(n_515), .B2(n_565), .Y(n_1068) );
AOI22xp5_ASAP7_75t_L g566 ( .A1(n_66), .A2(n_197), .B1(n_530), .B2(n_567), .Y(n_566) );
AOI22xp33_ASAP7_75t_SL g655 ( .A1(n_67), .A2(n_183), .B1(n_656), .B2(n_657), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g861 ( .A1(n_68), .A2(n_261), .B1(n_836), .B2(n_862), .Y(n_861) );
AOI22xp5_ASAP7_75t_L g1066 ( .A1(n_69), .A2(n_180), .B1(n_743), .B2(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g574 ( .A(n_71), .Y(n_574) );
INVx2_ASAP7_75t_L g302 ( .A(n_72), .Y(n_302) );
INVxp33_ASAP7_75t_SL g904 ( .A(n_74), .Y(n_904) );
INVx1_ASAP7_75t_L g815 ( .A(n_75), .Y(n_815) );
AND2x4_ASAP7_75t_L g820 ( .A(n_75), .B(n_302), .Y(n_820) );
INVx1_ASAP7_75t_SL g842 ( .A(n_75), .Y(n_842) );
AOI22xp33_ASAP7_75t_L g543 ( .A1(n_77), .A2(n_215), .B1(n_378), .B2(n_544), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g725 ( .A1(n_78), .A2(n_276), .B1(n_389), .B2(n_540), .Y(n_725) );
AOI22xp5_ASAP7_75t_L g783 ( .A1(n_79), .A2(n_226), .B1(n_434), .B2(n_608), .Y(n_783) );
INVx1_ASAP7_75t_L g491 ( .A(n_80), .Y(n_491) );
NAND2xp5_ASAP7_75t_SL g755 ( .A(n_82), .B(n_643), .Y(n_755) );
INVx1_ASAP7_75t_L g1060 ( .A(n_83), .Y(n_1060) );
INVx1_ASAP7_75t_L g712 ( .A(n_84), .Y(n_712) );
AOI21xp5_ASAP7_75t_L g315 ( .A1(n_85), .A2(n_316), .B(n_341), .Y(n_315) );
AOI22xp5_ASAP7_75t_L g787 ( .A1(n_86), .A2(n_258), .B1(n_396), .B2(n_657), .Y(n_787) );
INVx1_ASAP7_75t_L g594 ( .A(n_87), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g606 ( .A1(n_88), .A2(n_257), .B1(n_470), .B2(n_471), .Y(n_606) );
BUFx6f_ASAP7_75t_L g323 ( .A(n_90), .Y(n_323) );
AOI22xp33_ASAP7_75t_L g629 ( .A1(n_91), .A2(n_125), .B1(n_534), .B2(n_563), .Y(n_629) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_93), .B(n_507), .Y(n_771) );
AOI22xp33_ASAP7_75t_L g1045 ( .A1(n_94), .A2(n_238), .B1(n_521), .B2(n_522), .Y(n_1045) );
AOI22xp33_ASAP7_75t_L g1036 ( .A1(n_96), .A2(n_280), .B1(n_501), .B2(n_505), .Y(n_1036) );
AOI22xp33_ASAP7_75t_L g1044 ( .A1(n_97), .A2(n_188), .B1(n_518), .B2(n_519), .Y(n_1044) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_98), .A2(n_170), .B1(n_490), .B2(n_618), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g375 ( .A1(n_99), .A2(n_121), .B1(n_376), .B2(n_381), .Y(n_375) );
AOI21xp5_ASAP7_75t_L g644 ( .A1(n_101), .A2(n_645), .B(n_647), .Y(n_644) );
INVx1_ASAP7_75t_SL g669 ( .A(n_102), .Y(n_669) );
NOR3xp33_ASAP7_75t_L g697 ( .A(n_102), .B(n_698), .C(n_699), .Y(n_697) );
INVx1_ASAP7_75t_L g492 ( .A(n_105), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g649 ( .A1(n_106), .A2(n_207), .B1(n_487), .B2(n_577), .Y(n_649) );
AOI221xp5_ASAP7_75t_L g572 ( .A1(n_107), .A2(n_193), .B1(n_501), .B2(n_509), .C(n_573), .Y(n_572) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_108), .A2(n_287), .B1(n_446), .B2(n_447), .Y(n_575) );
INVx1_ASAP7_75t_L g1040 ( .A(n_109), .Y(n_1040) );
AOI22xp5_ASAP7_75t_L g793 ( .A1(n_110), .A2(n_209), .B1(n_487), .B2(n_577), .Y(n_793) );
AOI22xp33_ASAP7_75t_L g520 ( .A1(n_111), .A2(n_235), .B1(n_521), .B2(n_522), .Y(n_520) );
INVx1_ASAP7_75t_L g324 ( .A(n_112), .Y(n_324) );
NAND2xp5_ASAP7_75t_L g348 ( .A(n_112), .B(n_229), .Y(n_348) );
INVx1_ASAP7_75t_L g709 ( .A(n_114), .Y(n_709) );
AOI22xp5_ASAP7_75t_L g537 ( .A1(n_116), .A2(n_216), .B1(n_428), .B2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_118), .A2(n_163), .B1(n_540), .B2(n_657), .Y(n_741) );
AOI22xp5_ASAP7_75t_L g650 ( .A1(n_119), .A2(n_184), .B1(n_446), .B2(n_447), .Y(n_650) );
AOI21xp5_ASAP7_75t_SL g790 ( .A1(n_120), .A2(n_645), .B(n_791), .Y(n_790) );
CKINVDCx5p33_ASAP7_75t_R g691 ( .A(n_122), .Y(n_691) );
AOI22xp33_ASAP7_75t_L g503 ( .A1(n_123), .A2(n_130), .B1(n_504), .B2(n_505), .Y(n_503) );
INVx1_ASAP7_75t_L g497 ( .A(n_124), .Y(n_497) );
AOI22xp5_ASAP7_75t_L g539 ( .A1(n_126), .A2(n_237), .B1(n_389), .B2(n_540), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g514 ( .A1(n_127), .A2(n_228), .B1(n_515), .B2(n_516), .Y(n_514) );
INVx1_ASAP7_75t_L g559 ( .A(n_128), .Y(n_559) );
CKINVDCx20_ASAP7_75t_R g796 ( .A(n_129), .Y(n_796) );
AO221x2_ASAP7_75t_L g900 ( .A1(n_129), .A2(n_132), .B1(n_869), .B2(n_901), .C(n_902), .Y(n_900) );
AOI22xp5_ASAP7_75t_L g835 ( .A1(n_131), .A2(n_291), .B1(n_824), .B2(n_836), .Y(n_835) );
OAI22xp5_ASAP7_75t_L g1052 ( .A1(n_133), .A2(n_1053), .B1(n_1054), .B2(n_1055), .Y(n_1052) );
CKINVDCx5p33_ASAP7_75t_R g1053 ( .A(n_133), .Y(n_1053) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_134), .A2(n_158), .B1(n_414), .B2(n_465), .Y(n_464) );
AOI21xp33_ASAP7_75t_L g546 ( .A1(n_135), .A2(n_509), .B(n_547), .Y(n_546) );
INVx1_ASAP7_75t_L g775 ( .A(n_136), .Y(n_775) );
INVx1_ASAP7_75t_L g599 ( .A(n_137), .Y(n_599) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_138), .A2(n_239), .B1(n_407), .B2(n_428), .Y(n_605) );
AOI22xp33_ASAP7_75t_L g678 ( .A1(n_139), .A2(n_161), .B1(n_513), .B2(n_516), .Y(n_678) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_140), .A2(n_283), .B1(n_515), .B2(n_516), .Y(n_767) );
AOI22xp33_ASAP7_75t_L g568 ( .A1(n_141), .A2(n_203), .B1(n_569), .B2(n_570), .Y(n_568) );
AOI22xp33_ASAP7_75t_L g653 ( .A1(n_142), .A2(n_246), .B1(n_540), .B2(n_654), .Y(n_653) );
AOI21xp33_ASAP7_75t_L g773 ( .A1(n_143), .A2(n_501), .B(n_774), .Y(n_773) );
AOI22xp33_ASAP7_75t_L g607 ( .A1(n_144), .A2(n_269), .B1(n_434), .B2(n_608), .Y(n_607) );
AOI22xp33_ASAP7_75t_L g500 ( .A1(n_145), .A2(n_176), .B1(n_501), .B2(n_502), .Y(n_500) );
AOI22xp33_ASAP7_75t_L g620 ( .A1(n_146), .A2(n_182), .B1(n_544), .B2(n_621), .Y(n_620) );
AOI22x1_ASAP7_75t_L g583 ( .A1(n_148), .A2(n_584), .B1(n_585), .B2(n_609), .Y(n_583) );
INVx1_ASAP7_75t_L g609 ( .A(n_148), .Y(n_609) );
AOI22xp5_ASAP7_75t_L g768 ( .A1(n_150), .A2(n_214), .B1(n_513), .B2(n_519), .Y(n_768) );
CKINVDCx16_ASAP7_75t_R g455 ( .A(n_153), .Y(n_455) );
INVx1_ASAP7_75t_L g648 ( .A(n_155), .Y(n_648) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_156), .A2(n_173), .B1(n_521), .B2(n_522), .Y(n_766) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_162), .B(n_592), .Y(n_619) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_165), .A2(n_234), .B1(n_841), .B2(n_843), .Y(n_840) );
AOI21xp5_ASAP7_75t_L g588 ( .A1(n_166), .A2(n_438), .B(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g564 ( .A1(n_167), .A2(n_241), .B1(n_389), .B2(n_565), .Y(n_564) );
AOI22xp33_ASAP7_75t_L g445 ( .A1(n_168), .A2(n_248), .B1(n_446), .B2(n_447), .Y(n_445) );
AOI22xp5_ASAP7_75t_L g533 ( .A1(n_169), .A2(n_192), .B1(n_534), .B2(n_536), .Y(n_533) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_171), .A2(n_290), .B1(n_819), .B2(n_836), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g1043 ( .A1(n_172), .A2(n_213), .B1(n_515), .B2(n_516), .Y(n_1043) );
AOI22xp33_ASAP7_75t_L g1070 ( .A1(n_177), .A2(n_211), .B1(n_521), .B2(n_522), .Y(n_1070) );
AOI22xp33_ASAP7_75t_L g784 ( .A1(n_178), .A2(n_288), .B1(n_404), .B2(n_432), .Y(n_784) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_181), .B(n_602), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g440 ( .A1(n_185), .A2(n_270), .B1(n_441), .B2(n_442), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_186), .A2(n_225), .B1(n_623), .B2(n_624), .Y(n_622) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_189), .A2(n_294), .B1(n_366), .B2(n_371), .Y(n_365) );
AOI22xp5_ASAP7_75t_L g659 ( .A1(n_190), .A2(n_255), .B1(n_428), .B2(n_538), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g720 ( .A1(n_191), .A2(n_240), .B1(n_502), .B2(n_721), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g448 ( .A1(n_196), .A2(n_449), .B(n_450), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g1058 ( .A1(n_198), .A2(n_247), .B1(n_501), .B2(n_507), .C(n_1059), .Y(n_1058) );
AOI22x1_ASAP7_75t_L g311 ( .A1(n_200), .A2(n_312), .B1(n_313), .B2(n_419), .Y(n_311) );
INVx1_ASAP7_75t_L g419 ( .A(n_200), .Y(n_419) );
OAI22xp5_ASAP7_75t_L g456 ( .A1(n_200), .A2(n_312), .B1(n_313), .B2(n_419), .Y(n_456) );
AOI22xp33_ASAP7_75t_L g872 ( .A1(n_200), .A2(n_224), .B1(n_813), .B2(n_824), .Y(n_872) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_201), .A2(n_208), .B1(n_544), .B2(n_714), .Y(n_749) );
INVx1_ASAP7_75t_L g342 ( .A(n_202), .Y(n_342) );
INVx1_ASAP7_75t_L g631 ( .A(n_205), .Y(n_631) );
AOI22xp5_ASAP7_75t_L g745 ( .A1(n_206), .A2(n_278), .B1(n_428), .B2(n_538), .Y(n_745) );
OA22x2_ASAP7_75t_L g328 ( .A1(n_210), .A2(n_230), .B1(n_323), .B2(n_327), .Y(n_328) );
INVx1_ASAP7_75t_L g364 ( .A(n_210), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_212), .A2(n_275), .B1(n_453), .B2(n_507), .Y(n_506) );
CKINVDCx5p33_ASAP7_75t_R g683 ( .A(n_217), .Y(n_683) );
AO22x2_ASAP7_75t_L g701 ( .A1(n_218), .A2(n_702), .B1(n_703), .B2(n_704), .Y(n_701) );
INVx1_ASAP7_75t_L g702 ( .A(n_218), .Y(n_702) );
AND2x2_ASAP7_75t_L g673 ( .A(n_219), .B(n_354), .Y(n_673) );
NAND2xp33_ASAP7_75t_L g437 ( .A(n_220), .B(n_438), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_221), .A2(n_273), .B1(n_388), .B2(n_396), .Y(n_387) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_222), .A2(n_260), .B1(n_404), .B2(n_627), .Y(n_626) );
INVx1_ASAP7_75t_L g817 ( .A(n_223), .Y(n_817) );
AOI22xp33_ASAP7_75t_L g846 ( .A1(n_227), .A2(n_243), .B1(n_824), .B2(n_847), .Y(n_846) );
INVx1_ASAP7_75t_L g340 ( .A(n_229), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_229), .B(n_361), .Y(n_360) );
OAI21xp33_ASAP7_75t_L g374 ( .A1(n_230), .A2(n_251), .B(n_352), .Y(n_374) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_231), .A2(n_249), .B1(n_404), .B2(n_530), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g772 ( .A1(n_232), .A2(n_256), .B1(n_505), .B2(n_509), .Y(n_772) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_233), .A2(n_267), .B1(n_518), .B2(n_530), .Y(n_668) );
XNOR2x2_ASAP7_75t_SL g762 ( .A(n_234), .B(n_763), .Y(n_762) );
XNOR2x1_ASAP7_75t_L g798 ( .A(n_234), .B(n_763), .Y(n_798) );
INVx1_ASAP7_75t_L g526 ( .A(n_236), .Y(n_526) );
INVx1_ASAP7_75t_L g474 ( .A(n_242), .Y(n_474) );
OAI21x1_ASAP7_75t_L g737 ( .A1(n_243), .A2(n_738), .B(n_756), .Y(n_737) );
NAND2xp5_ASAP7_75t_L g759 ( .A(n_243), .B(n_741), .Y(n_759) );
INVx1_ASAP7_75t_L g488 ( .A(n_245), .Y(n_488) );
INVx1_ASAP7_75t_SL g821 ( .A(n_250), .Y(n_821) );
NOR2xp33_ASAP7_75t_L g306 ( .A(n_251), .B(n_277), .Y(n_306) );
INVx1_ASAP7_75t_L g326 ( .A(n_251), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_252), .B(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g1061 ( .A1(n_259), .A2(n_272), .B1(n_1062), .B2(n_1063), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g827 ( .A(n_264), .Y(n_827) );
INVx1_ASAP7_75t_L g596 ( .A(n_265), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_266), .B(n_438), .Y(n_789) );
INVx1_ASAP7_75t_L g590 ( .A(n_268), .Y(n_590) );
AOI22xp33_ASAP7_75t_L g1042 ( .A1(n_271), .A2(n_274), .B1(n_512), .B2(n_513), .Y(n_1042) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_277), .B(n_333), .Y(n_332) );
AOI22x1_ASAP7_75t_L g794 ( .A1(n_279), .A2(n_285), .B1(n_446), .B2(n_795), .Y(n_794) );
NAND2xp5_ASAP7_75t_L g1037 ( .A(n_281), .B(n_577), .Y(n_1037) );
AOI21xp33_ASAP7_75t_L g752 ( .A1(n_284), .A2(n_449), .B(n_753), .Y(n_752) );
INVx1_ASAP7_75t_L g826 ( .A(n_286), .Y(n_826) );
INVx1_ASAP7_75t_L g639 ( .A(n_293), .Y(n_639) );
NOR2xp33_ASAP7_75t_L g663 ( .A(n_293), .B(n_658), .Y(n_663) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_297), .A2(n_308), .B(n_803), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
BUFx4_ASAP7_75t_SL g298 ( .A(n_299), .Y(n_298) );
NAND3xp33_ASAP7_75t_L g299 ( .A(n_300), .B(n_303), .C(n_307), .Y(n_299) );
AND2x2_ASAP7_75t_L g1048 ( .A(n_300), .B(n_1049), .Y(n_1048) );
AND2x2_ASAP7_75t_L g1072 ( .A(n_300), .B(n_1050), .Y(n_1072) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
OA21x2_ASAP7_75t_L g1074 ( .A1(n_301), .A2(n_842), .B(n_1075), .Y(n_1074) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g814 ( .A(n_302), .B(n_815), .Y(n_814) );
AND3x4_ASAP7_75t_L g841 ( .A(n_302), .B(n_825), .C(n_842), .Y(n_841) );
NOR2xp33_ASAP7_75t_L g1049 ( .A(n_303), .B(n_1050), .Y(n_1049) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
AO21x2_ASAP7_75t_L g357 ( .A1(n_304), .A2(n_358), .B(n_359), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_305), .B(n_306), .Y(n_304) );
INVx1_ASAP7_75t_L g1050 ( .A(n_307), .Y(n_1050) );
XNOR2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_554), .Y(n_308) );
OAI22xp33_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_458), .B1(n_459), .B2(n_553), .Y(n_309) );
INVx1_ASAP7_75t_L g553 ( .A(n_310), .Y(n_553) );
OAI22xp5_ASAP7_75t_L g310 ( .A1(n_311), .A2(n_420), .B1(n_456), .B2(n_457), .Y(n_310) );
INVx2_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g313 ( .A(n_314), .B(n_386), .Y(n_313) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_315), .B(n_365), .C(n_375), .Y(n_314) );
BUFx3_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
INVx2_ASAP7_75t_L g318 ( .A(n_319), .Y(n_318) );
INVx3_ASAP7_75t_L g439 ( .A(n_319), .Y(n_439) );
BUFx3_ASAP7_75t_L g623 ( .A(n_319), .Y(n_623) );
AND2x2_ASAP7_75t_L g319 ( .A(n_320), .B(n_329), .Y(n_319) );
AND2x2_ASAP7_75t_L g385 ( .A(n_320), .B(n_380), .Y(n_385) );
AND2x4_ASAP7_75t_L g402 ( .A(n_320), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g415 ( .A(n_320), .B(n_393), .Y(n_415) );
AND2x4_ASAP7_75t_L g504 ( .A(n_320), .B(n_380), .Y(n_504) );
AND2x2_ASAP7_75t_L g509 ( .A(n_320), .B(n_329), .Y(n_509) );
AND2x4_ASAP7_75t_L g512 ( .A(n_320), .B(n_398), .Y(n_512) );
AND2x4_ASAP7_75t_L g518 ( .A(n_320), .B(n_393), .Y(n_518) );
AND2x2_ASAP7_75t_L g535 ( .A(n_320), .B(n_393), .Y(n_535) );
AND2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_328), .Y(n_320) );
INVx1_ASAP7_75t_L g370 ( .A(n_321), .Y(n_370) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
NAND2xp33_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
INVx2_ASAP7_75t_L g327 ( .A(n_323), .Y(n_327) );
INVx3_ASAP7_75t_L g333 ( .A(n_323), .Y(n_333) );
NAND2xp33_ASAP7_75t_L g339 ( .A(n_323), .B(n_340), .Y(n_339) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_323), .Y(n_347) );
INVx1_ASAP7_75t_L g352 ( .A(n_323), .Y(n_352) );
NAND2xp5_ASAP7_75t_L g363 ( .A(n_324), .B(n_364), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g325 ( .A(n_326), .B(n_327), .Y(n_325) );
OAI21xp5_ASAP7_75t_L g350 ( .A1(n_326), .A2(n_351), .B(n_352), .Y(n_350) );
AND2x2_ASAP7_75t_L g349 ( .A(n_328), .B(n_350), .Y(n_349) );
AND2x2_ASAP7_75t_L g369 ( .A(n_328), .B(n_370), .Y(n_369) );
INVx1_ASAP7_75t_L g392 ( .A(n_328), .Y(n_392) );
AND2x4_ASAP7_75t_L g368 ( .A(n_329), .B(n_369), .Y(n_368) );
AND2x4_ASAP7_75t_L g372 ( .A(n_329), .B(n_373), .Y(n_372) );
AND2x2_ASAP7_75t_L g412 ( .A(n_329), .B(n_391), .Y(n_412) );
AND2x4_ASAP7_75t_L g505 ( .A(n_329), .B(n_373), .Y(n_505) );
AND2x2_ASAP7_75t_L g507 ( .A(n_329), .B(n_369), .Y(n_507) );
AND2x4_ASAP7_75t_L g522 ( .A(n_329), .B(n_391), .Y(n_522) );
AND2x4_ASAP7_75t_L g329 ( .A(n_330), .B(n_335), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
AND2x2_ASAP7_75t_L g345 ( .A(n_331), .B(n_346), .Y(n_345) );
AND2x4_ASAP7_75t_L g380 ( .A(n_331), .B(n_335), .Y(n_380) );
AND2x4_ASAP7_75t_L g393 ( .A(n_331), .B(n_394), .Y(n_393) );
OR2x2_ASAP7_75t_L g399 ( .A(n_331), .B(n_395), .Y(n_399) );
AND2x4_ASAP7_75t_L g331 ( .A(n_332), .B(n_334), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g337 ( .A(n_333), .B(n_338), .Y(n_337) );
INVxp67_ASAP7_75t_L g361 ( .A(n_333), .Y(n_361) );
NAND3xp33_ASAP7_75t_L g359 ( .A(n_334), .B(n_360), .C(n_362), .Y(n_359) );
INVx1_ASAP7_75t_L g335 ( .A(n_336), .Y(n_335) );
INVx1_ASAP7_75t_L g395 ( .A(n_336), .Y(n_395) );
AND2x2_ASAP7_75t_L g336 ( .A(n_337), .B(n_339), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g341 ( .A1(n_342), .A2(n_343), .B(n_353), .Y(n_341) );
INVx2_ASAP7_75t_L g447 ( .A(n_343), .Y(n_447) );
INVx3_ASAP7_75t_L g602 ( .A(n_343), .Y(n_602) );
INVx4_ASAP7_75t_L g795 ( .A(n_343), .Y(n_795) );
INVx5_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
BUFx4f_ASAP7_75t_L g482 ( .A(n_344), .Y(n_482) );
BUFx2_ASAP7_75t_L g618 ( .A(n_344), .Y(n_618) );
AND2x4_ASAP7_75t_L g344 ( .A(n_345), .B(n_349), .Y(n_344) );
AND2x2_ASAP7_75t_L g502 ( .A(n_345), .B(n_349), .Y(n_502) );
AND2x4_ASAP7_75t_L g685 ( .A(n_345), .B(n_349), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
INVx1_ASAP7_75t_L g358 ( .A(n_347), .Y(n_358) );
INVx4_ASAP7_75t_L g354 ( .A(n_355), .Y(n_354) );
INVx3_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
INVx4_ASAP7_75t_L g484 ( .A(n_356), .Y(n_484) );
INVx3_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
BUFx6f_ASAP7_75t_L g454 ( .A(n_357), .Y(n_454) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_361), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_L g373 ( .A(n_362), .B(n_374), .Y(n_373) );
INVx2_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
INVx3_ASAP7_75t_L g592 ( .A(n_367), .Y(n_592) );
INVx2_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
BUFx3_ASAP7_75t_L g441 ( .A(n_368), .Y(n_441) );
INVx2_ASAP7_75t_L g479 ( .A(n_368), .Y(n_479) );
BUFx6f_ASAP7_75t_L g577 ( .A(n_368), .Y(n_577) );
BUFx8_ASAP7_75t_SL g671 ( .A(n_368), .Y(n_671) );
BUFx6f_ASAP7_75t_L g714 ( .A(n_368), .Y(n_714) );
AND2x4_ASAP7_75t_L g379 ( .A(n_369), .B(n_380), .Y(n_379) );
AND2x4_ASAP7_75t_L g501 ( .A(n_369), .B(n_380), .Y(n_501) );
AND2x4_ASAP7_75t_L g391 ( .A(n_370), .B(n_392), .Y(n_391) );
BUFx6f_ASAP7_75t_L g371 ( .A(n_372), .Y(n_371) );
INVx3_ASAP7_75t_L g443 ( .A(n_372), .Y(n_443) );
BUFx6f_ASAP7_75t_L g544 ( .A(n_372), .Y(n_544) );
AND2x4_ASAP7_75t_L g405 ( .A(n_373), .B(n_398), .Y(n_405) );
AND2x4_ASAP7_75t_L g418 ( .A(n_373), .B(n_393), .Y(n_418) );
AND2x4_ASAP7_75t_L g513 ( .A(n_373), .B(n_398), .Y(n_513) );
AND2x4_ASAP7_75t_L g519 ( .A(n_373), .B(n_393), .Y(n_519) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
BUFx6f_ASAP7_75t_L g449 ( .A(n_379), .Y(n_449) );
BUFx3_ASAP7_75t_L g621 ( .A(n_379), .Y(n_621) );
INVx1_ASAP7_75t_L g646 ( .A(n_379), .Y(n_646) );
AND2x4_ASAP7_75t_L g408 ( .A(n_380), .B(n_391), .Y(n_408) );
AND2x4_ASAP7_75t_L g521 ( .A(n_380), .B(n_391), .Y(n_521) );
INVx1_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx6f_ASAP7_75t_L g600 ( .A(n_384), .Y(n_600) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
BUFx6f_ASAP7_75t_L g446 ( .A(n_385), .Y(n_446) );
BUFx3_ASAP7_75t_L g490 ( .A(n_385), .Y(n_490) );
NAND4xp25_ASAP7_75t_SL g386 ( .A(n_387), .B(n_400), .C(n_406), .D(n_413), .Y(n_386) );
BUFx12f_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
BUFx12f_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_390), .Y(n_470) );
BUFx6f_ASAP7_75t_L g657 ( .A(n_390), .Y(n_657) );
AND2x4_ASAP7_75t_L g390 ( .A(n_391), .B(n_393), .Y(n_390) );
AND2x4_ASAP7_75t_L g397 ( .A(n_391), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g515 ( .A(n_391), .B(n_393), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_391), .B(n_403), .Y(n_516) );
INVx1_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
BUFx6f_ASAP7_75t_L g471 ( .A(n_397), .Y(n_471) );
BUFx6f_ASAP7_75t_L g540 ( .A(n_397), .Y(n_540) );
BUFx6f_ASAP7_75t_L g565 ( .A(n_397), .Y(n_565) );
INVx2_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
INVx2_ASAP7_75t_L g403 ( .A(n_399), .Y(n_403) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
BUFx12f_ASAP7_75t_L g432 ( .A(n_402), .Y(n_432) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_402), .Y(n_530) );
BUFx6f_ASAP7_75t_L g627 ( .A(n_402), .Y(n_627) );
BUFx12f_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx6_ASAP7_75t_L g532 ( .A(n_405), .Y(n_532) );
BUFx6f_ASAP7_75t_L g407 ( .A(n_408), .Y(n_407) );
INVx3_ASAP7_75t_L g427 ( .A(n_408), .Y(n_427) );
BUFx12f_ASAP7_75t_L g538 ( .A(n_408), .Y(n_538) );
BUFx6f_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
INVx2_ASAP7_75t_L g410 ( .A(n_411), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
BUFx6f_ASAP7_75t_L g428 ( .A(n_412), .Y(n_428) );
BUFx5_ASAP7_75t_L g467 ( .A(n_412), .Y(n_467) );
BUFx3_ASAP7_75t_L g570 ( .A(n_412), .Y(n_570) );
BUFx8_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
BUFx6f_ASAP7_75t_L g434 ( .A(n_415), .Y(n_434) );
INVx4_ASAP7_75t_L g416 ( .A(n_417), .Y(n_416) );
INVx2_ASAP7_75t_L g435 ( .A(n_417), .Y(n_435) );
INVx1_ASAP7_75t_L g465 ( .A(n_417), .Y(n_465) );
INVx2_ASAP7_75t_SL g536 ( .A(n_417), .Y(n_536) );
INVx4_ASAP7_75t_L g563 ( .A(n_417), .Y(n_563) );
INVx4_ASAP7_75t_L g608 ( .A(n_417), .Y(n_608) );
INVx1_ASAP7_75t_L g656 ( .A(n_417), .Y(n_656) );
INVx8_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
HB1xp67_ASAP7_75t_L g420 ( .A(n_421), .Y(n_420) );
INVx1_ASAP7_75t_L g457 ( .A(n_421), .Y(n_457) );
HB1xp67_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
XNOR2x1_ASAP7_75t_L g422 ( .A(n_423), .B(n_455), .Y(n_422) );
NAND4xp75_ASAP7_75t_L g423 ( .A(n_424), .B(n_430), .C(n_436), .D(n_444), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_425), .B(n_429), .Y(n_424) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
INVx1_ASAP7_75t_L g569 ( .A(n_427), .Y(n_569) );
INVx2_ASAP7_75t_L g677 ( .A(n_427), .Y(n_677) );
AND2x2_ASAP7_75t_L g430 ( .A(n_431), .B(n_433), .Y(n_430) );
AND2x2_ASAP7_75t_L g436 ( .A(n_437), .B(n_440), .Y(n_436) );
INVx3_ASAP7_75t_SL g438 ( .A(n_439), .Y(n_438) );
INVx2_ASAP7_75t_L g476 ( .A(n_439), .Y(n_476) );
INVx2_ASAP7_75t_L g643 ( .A(n_439), .Y(n_643) );
INVx2_ASAP7_75t_L g672 ( .A(n_439), .Y(n_672) );
INVx2_ASAP7_75t_L g1062 ( .A(n_439), .Y(n_1062) );
INVx1_ASAP7_75t_L g597 ( .A(n_442), .Y(n_597) );
INVx3_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g487 ( .A(n_443), .Y(n_487) );
INVx2_ASAP7_75t_L g1063 ( .A(n_443), .Y(n_1063) );
AND2x2_ASAP7_75t_L g444 ( .A(n_445), .B(n_448), .Y(n_444) );
INVx3_ASAP7_75t_L g710 ( .A(n_446), .Y(n_710) );
INVx4_ASAP7_75t_L g595 ( .A(n_449), .Y(n_595) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_451), .B(n_452), .Y(n_450) );
NOR2xp33_ASAP7_75t_SL g589 ( .A(n_452), .B(n_590), .Y(n_589) );
INVx3_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
BUFx6f_ASAP7_75t_L g549 ( .A(n_454), .Y(n_549) );
BUFx6f_ASAP7_75t_L g722 ( .A(n_454), .Y(n_722) );
NOR2xp33_ASAP7_75t_L g774 ( .A(n_454), .B(n_775), .Y(n_774) );
NOR2xp33_ASAP7_75t_L g1039 ( .A(n_454), .B(n_1040), .Y(n_1039) );
INVx2_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
OA22x2_ASAP7_75t_L g459 ( .A1(n_460), .A2(n_493), .B1(n_494), .B2(n_552), .Y(n_459) );
HB1xp67_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g552 ( .A(n_461), .Y(n_552) );
XNOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_492), .Y(n_461) );
NAND2x1_ASAP7_75t_L g462 ( .A(n_463), .B(n_472), .Y(n_462) );
AND4x1_ASAP7_75t_L g463 ( .A(n_464), .B(n_466), .C(n_468), .D(n_469), .Y(n_463) );
OAI21xp5_ASAP7_75t_L g473 ( .A1(n_474), .A2(n_475), .B(n_477), .Y(n_473) );
INVx2_ASAP7_75t_L g475 ( .A(n_476), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
OAI21xp5_ASAP7_75t_SL g478 ( .A1(n_479), .A2(n_480), .B(n_481), .Y(n_478) );
INVx4_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI22xp5_ASAP7_75t_L g485 ( .A1(n_486), .A2(n_488), .B1(n_489), .B2(n_491), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_487), .Y(n_486) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
AOI22x1_ASAP7_75t_L g494 ( .A1(n_495), .A2(n_523), .B1(n_550), .B2(n_551), .Y(n_494) );
INVx2_ASAP7_75t_L g551 ( .A(n_495), .Y(n_551) );
INVx3_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
XNOR2x1_ASAP7_75t_L g496 ( .A(n_497), .B(n_498), .Y(n_496) );
OR2x2_ASAP7_75t_L g498 ( .A(n_499), .B(n_510), .Y(n_498) );
NAND4xp25_ASAP7_75t_L g499 ( .A(n_500), .B(n_503), .C(n_506), .D(n_508), .Y(n_499) );
INVx2_ASAP7_75t_L g690 ( .A(n_501), .Y(n_690) );
INVx2_ASAP7_75t_L g692 ( .A(n_504), .Y(n_692) );
INVx2_ASAP7_75t_L g687 ( .A(n_505), .Y(n_687) );
NAND4xp25_ASAP7_75t_L g510 ( .A(n_511), .B(n_514), .C(n_517), .D(n_520), .Y(n_510) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_519), .Y(n_1067) );
INVxp67_ASAP7_75t_SL g523 ( .A(n_524), .Y(n_523) );
BUFx2_ASAP7_75t_L g550 ( .A(n_524), .Y(n_550) );
XNOR2x1_ASAP7_75t_L g524 ( .A(n_525), .B(n_527), .Y(n_524) );
CKINVDCx5p33_ASAP7_75t_R g525 ( .A(n_526), .Y(n_525) );
NOR2x1_ASAP7_75t_L g527 ( .A(n_528), .B(n_541), .Y(n_527) );
NAND4xp25_ASAP7_75t_L g528 ( .A(n_529), .B(n_533), .C(n_537), .D(n_539), .Y(n_528) );
INVx2_ASAP7_75t_L g531 ( .A(n_532), .Y(n_531) );
INVx3_ASAP7_75t_L g567 ( .A(n_532), .Y(n_567) );
INVx2_ASAP7_75t_L g654 ( .A(n_532), .Y(n_654) );
INVx5_ASAP7_75t_L g743 ( .A(n_532), .Y(n_743) );
BUFx4f_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
BUFx6f_ASAP7_75t_L g661 ( .A(n_535), .Y(n_661) );
NAND4xp25_ASAP7_75t_L g541 ( .A(n_542), .B(n_543), .C(n_545), .D(n_546), .Y(n_541) );
INVx3_ASAP7_75t_L g716 ( .A(n_544), .Y(n_716) );
NOR2xp33_ASAP7_75t_L g547 ( .A(n_548), .B(n_549), .Y(n_547) );
NOR2xp33_ASAP7_75t_L g573 ( .A(n_549), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g624 ( .A(n_549), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g647 ( .A(n_549), .B(n_648), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g753 ( .A(n_549), .B(n_754), .Y(n_753) );
NOR2xp33_ASAP7_75t_L g791 ( .A(n_549), .B(n_792), .Y(n_791) );
NOR2xp67_ASAP7_75t_SL g1059 ( .A(n_549), .B(n_1060), .Y(n_1059) );
OAI22xp5_ASAP7_75t_L g554 ( .A1(n_555), .A2(n_634), .B1(n_801), .B2(n_802), .Y(n_554) );
INVx1_ASAP7_75t_L g802 ( .A(n_555), .Y(n_802) );
AOI22xp5_ASAP7_75t_L g555 ( .A1(n_556), .A2(n_557), .B1(n_578), .B2(n_579), .Y(n_555) );
INVx1_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
BUFx2_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
XNOR2x1_ASAP7_75t_L g558 ( .A(n_559), .B(n_560), .Y(n_558) );
NOR2x1_ASAP7_75t_L g560 ( .A(n_561), .B(n_571), .Y(n_560) );
NAND4xp25_ASAP7_75t_SL g561 ( .A(n_562), .B(n_564), .C(n_566), .D(n_568), .Y(n_561) );
NAND3xp33_ASAP7_75t_L g571 ( .A(n_572), .B(n_575), .C(n_576), .Y(n_571) );
INVx1_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
OAI22xp5_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .B1(n_610), .B2(n_632), .Y(n_579) );
INVx2_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
INVx2_ASAP7_75t_L g581 ( .A(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_586), .B(n_603), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_587), .B(n_593), .C(n_598), .Y(n_586) );
NAND2xp5_ASAP7_75t_SL g587 ( .A(n_588), .B(n_591), .Y(n_587) );
OAI22xp5_ASAP7_75t_L g593 ( .A1(n_594), .A2(n_595), .B1(n_596), .B2(n_597), .Y(n_593) );
OAI21xp33_ASAP7_75t_L g598 ( .A1(n_599), .A2(n_600), .B(n_601), .Y(n_598) );
AND4x1_ASAP7_75t_L g603 ( .A(n_604), .B(n_605), .C(n_606), .D(n_607), .Y(n_603) );
INVx1_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g633 ( .A(n_612), .Y(n_633) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
XOR2x2_ASAP7_75t_L g614 ( .A(n_615), .B(n_631), .Y(n_614) );
NOR2x1_ASAP7_75t_L g615 ( .A(n_616), .B(n_625), .Y(n_615) );
NAND4xp25_ASAP7_75t_L g616 ( .A(n_617), .B(n_619), .C(n_620), .D(n_622), .Y(n_616) );
INVx1_ASAP7_75t_L g708 ( .A(n_621), .Y(n_708) );
INVx2_ASAP7_75t_L g719 ( .A(n_623), .Y(n_719) );
NAND4xp25_ASAP7_75t_L g625 ( .A(n_626), .B(n_628), .C(n_629), .D(n_630), .Y(n_625) );
BUFx2_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
INVx1_ASAP7_75t_L g801 ( .A(n_634), .Y(n_801) );
OAI22xp5_ASAP7_75t_L g634 ( .A1(n_635), .A2(n_733), .B1(n_734), .B2(n_799), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
INVx2_ASAP7_75t_SL g800 ( .A(n_636), .Y(n_800) );
AO22x2_ASAP7_75t_L g636 ( .A1(n_637), .A2(n_700), .B1(n_730), .B2(n_731), .Y(n_636) );
INVx1_ASAP7_75t_L g730 ( .A(n_637), .Y(n_730) );
XNOR2xp5_ASAP7_75t_L g637 ( .A(n_638), .B(n_665), .Y(n_637) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_639), .A2(n_640), .B(n_662), .Y(n_638) );
AND2x2_ASAP7_75t_L g640 ( .A(n_641), .B(n_651), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g662 ( .A(n_641), .B(n_663), .C(n_664), .Y(n_662) );
AND4x1_ASAP7_75t_L g641 ( .A(n_642), .B(n_644), .C(n_649), .D(n_650), .Y(n_641) );
INVx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_652), .B(n_658), .Y(n_651) );
INVxp67_ASAP7_75t_SL g664 ( .A(n_652), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g652 ( .A(n_653), .B(n_655), .Y(n_652) );
NAND2xp5_ASAP7_75t_L g658 ( .A(n_659), .B(n_660), .Y(n_658) );
NAND2x1_ASAP7_75t_L g665 ( .A(n_666), .B(n_693), .Y(n_665) );
NOR3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_674), .C(n_679), .Y(n_666) );
OAI22xp33_ASAP7_75t_L g667 ( .A1(n_668), .A2(n_669), .B1(n_670), .B2(n_1077), .Y(n_667) );
INVx1_ASAP7_75t_L g698 ( .A(n_668), .Y(n_698) );
NOR2xp67_ASAP7_75t_L g674 ( .A(n_669), .B(n_675), .Y(n_674) );
OAI22xp5_ASAP7_75t_L g679 ( .A1(n_669), .A2(n_680), .B1(n_681), .B2(n_1078), .Y(n_679) );
INVx1_ASAP7_75t_L g695 ( .A(n_670), .Y(n_695) );
NAND3xp33_ASAP7_75t_L g693 ( .A(n_675), .B(n_694), .C(n_697), .Y(n_693) );
AND2x2_ASAP7_75t_L g675 ( .A(n_676), .B(n_678), .Y(n_675) );
INVx1_ASAP7_75t_L g699 ( .A(n_680), .Y(n_699) );
INVx1_ASAP7_75t_L g696 ( .A(n_681), .Y(n_696) );
NOR2x1_ASAP7_75t_L g681 ( .A(n_682), .B(n_688), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_683), .A2(n_684), .B1(n_686), .B2(n_687), .Y(n_682) );
INVx4_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B1(n_691), .B2(n_692), .Y(n_688) );
NOR2xp33_ASAP7_75t_L g694 ( .A(n_695), .B(n_696), .Y(n_694) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g732 ( .A(n_701), .Y(n_732) );
INVx1_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_705), .B(n_723), .Y(n_704) );
NOR3xp33_ASAP7_75t_SL g705 ( .A(n_706), .B(n_711), .C(n_717), .Y(n_705) );
OAI22xp5_ASAP7_75t_L g706 ( .A1(n_707), .A2(n_708), .B1(n_709), .B2(n_710), .Y(n_706) );
OAI22xp5_ASAP7_75t_L g711 ( .A1(n_712), .A2(n_713), .B1(n_715), .B2(n_716), .Y(n_711) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
OAI21xp33_ASAP7_75t_L g717 ( .A1(n_718), .A2(n_719), .B(n_720), .Y(n_717) );
INVx1_ASAP7_75t_L g721 ( .A(n_722), .Y(n_721) );
NOR2xp33_ASAP7_75t_L g723 ( .A(n_724), .B(n_727), .Y(n_723) );
NAND2xp5_ASAP7_75t_L g724 ( .A(n_725), .B(n_726), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
XNOR2xp5_ASAP7_75t_L g734 ( .A(n_735), .B(n_777), .Y(n_734) );
OA22x2_ASAP7_75t_L g735 ( .A1(n_736), .A2(n_760), .B1(n_761), .B2(n_776), .Y(n_735) );
INVx2_ASAP7_75t_L g776 ( .A(n_736), .Y(n_776) );
INVx2_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
AND2x2_ASAP7_75t_L g738 ( .A(n_739), .B(n_747), .Y(n_738) );
NOR3xp33_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .C(n_744), .Y(n_739) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
NOR3xp33_ASAP7_75t_L g758 ( .A(n_742), .B(n_751), .C(n_759), .Y(n_758) );
NOR2xp33_ASAP7_75t_L g757 ( .A(n_744), .B(n_748), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g744 ( .A(n_745), .B(n_746), .Y(n_744) );
NOR2xp33_ASAP7_75t_L g747 ( .A(n_748), .B(n_751), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g748 ( .A(n_749), .B(n_750), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_755), .Y(n_751) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
INVx2_ASAP7_75t_L g760 ( .A(n_761), .Y(n_760) );
BUFx3_ASAP7_75t_L g761 ( .A(n_762), .Y(n_761) );
AOI22xp5_ASAP7_75t_L g778 ( .A1(n_762), .A2(n_779), .B1(n_780), .B2(n_797), .Y(n_778) );
OR2x2_ASAP7_75t_L g763 ( .A(n_764), .B(n_769), .Y(n_763) );
NAND4xp25_ASAP7_75t_L g764 ( .A(n_765), .B(n_766), .C(n_767), .D(n_768), .Y(n_764) );
NAND4xp25_ASAP7_75t_L g769 ( .A(n_770), .B(n_771), .C(n_772), .D(n_773), .Y(n_769) );
INVxp67_ASAP7_75t_SL g777 ( .A(n_778), .Y(n_777) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
XNOR2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_796), .Y(n_780) );
NOR3xp33_ASAP7_75t_SL g781 ( .A(n_782), .B(n_785), .C(n_788), .Y(n_781) );
NAND2xp5_ASAP7_75t_L g782 ( .A(n_783), .B(n_784), .Y(n_782) );
NAND2xp5_ASAP7_75t_L g785 ( .A(n_786), .B(n_787), .Y(n_785) );
NAND4xp25_ASAP7_75t_L g788 ( .A(n_789), .B(n_790), .C(n_793), .D(n_794), .Y(n_788) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_SL g799 ( .A(n_800), .Y(n_799) );
OAI221xp5_ASAP7_75t_L g803 ( .A1(n_804), .A2(n_1026), .B1(n_1029), .B2(n_1046), .C(n_1051), .Y(n_803) );
NOR4xp25_ASAP7_75t_L g804 ( .A(n_805), .B(n_957), .C(n_1000), .D(n_1012), .Y(n_804) );
OAI221xp5_ASAP7_75t_L g805 ( .A1(n_806), .A2(n_900), .B1(n_905), .B2(n_922), .C(n_1079), .Y(n_805) );
O2A1O1Ixp33_ASAP7_75t_L g806 ( .A1(n_807), .A2(n_849), .B(n_855), .C(n_864), .Y(n_806) );
AOI211xp5_ASAP7_75t_SL g950 ( .A1(n_807), .A2(n_856), .B(n_951), .C(n_953), .Y(n_950) );
AND2x2_ASAP7_75t_L g807 ( .A(n_808), .B(n_830), .Y(n_807) );
INVx1_ASAP7_75t_L g808 ( .A(n_809), .Y(n_808) );
A2O1A1Ixp33_ASAP7_75t_L g893 ( .A1(n_809), .A2(n_894), .B(n_896), .C(n_898), .Y(n_893) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_809), .B(n_913), .Y(n_912) );
AOI21xp33_ASAP7_75t_L g925 ( .A1(n_809), .A2(n_889), .B(n_926), .Y(n_925) );
NOR2xp33_ASAP7_75t_L g997 ( .A(n_809), .B(n_998), .Y(n_997) );
NOR2xp33_ASAP7_75t_L g1018 ( .A(n_809), .B(n_884), .Y(n_1018) );
INVx2_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx3_ASAP7_75t_L g854 ( .A(n_810), .Y(n_854) );
NAND2xp5_ASAP7_75t_L g891 ( .A(n_810), .B(n_859), .Y(n_891) );
NAND2xp5_ASAP7_75t_L g931 ( .A(n_810), .B(n_831), .Y(n_931) );
NOR2xp33_ASAP7_75t_L g936 ( .A(n_810), .B(n_856), .Y(n_936) );
NOR2xp33_ASAP7_75t_L g947 ( .A(n_810), .B(n_884), .Y(n_947) );
NAND2xp5_ASAP7_75t_L g952 ( .A(n_810), .B(n_860), .Y(n_952) );
NAND2xp5_ASAP7_75t_L g955 ( .A(n_810), .B(n_956), .Y(n_955) );
NAND2xp5_ASAP7_75t_L g1009 ( .A(n_810), .B(n_855), .Y(n_1009) );
OR2x2_ASAP7_75t_L g810 ( .A(n_811), .B(n_822), .Y(n_810) );
OAI22xp5_ASAP7_75t_L g811 ( .A1(n_812), .A2(n_817), .B1(n_818), .B2(n_821), .Y(n_811) );
OAI22xp5_ASAP7_75t_L g902 ( .A1(n_812), .A2(n_818), .B1(n_903), .B2(n_904), .Y(n_902) );
INVx3_ASAP7_75t_L g812 ( .A(n_813), .Y(n_812) );
AND2x4_ASAP7_75t_L g813 ( .A(n_814), .B(n_816), .Y(n_813) );
AND2x4_ASAP7_75t_L g824 ( .A(n_814), .B(n_825), .Y(n_824) );
AND2x2_ASAP7_75t_L g843 ( .A(n_814), .B(n_816), .Y(n_843) );
AND2x2_ASAP7_75t_L g847 ( .A(n_814), .B(n_816), .Y(n_847) );
AND2x4_ASAP7_75t_L g819 ( .A(n_816), .B(n_820), .Y(n_819) );
AND2x2_ASAP7_75t_L g834 ( .A(n_816), .B(n_820), .Y(n_834) );
AND2x2_ASAP7_75t_L g862 ( .A(n_816), .B(n_820), .Y(n_862) );
INVx2_ASAP7_75t_L g818 ( .A(n_819), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g828 ( .A(n_820), .B(n_825), .Y(n_828) );
AND2x4_ASAP7_75t_L g836 ( .A(n_820), .B(n_825), .Y(n_836) );
AND2x4_ASAP7_75t_L g871 ( .A(n_820), .B(n_825), .Y(n_871) );
OAI22xp5_ASAP7_75t_L g822 ( .A1(n_823), .A2(n_827), .B1(n_828), .B2(n_829), .Y(n_822) );
INVx1_ASAP7_75t_L g901 ( .A(n_823), .Y(n_901) );
INVx3_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
CKINVDCx5p33_ASAP7_75t_R g1075 ( .A(n_825), .Y(n_1075) );
BUFx2_ASAP7_75t_L g1028 ( .A(n_828), .Y(n_1028) );
INVx1_ASAP7_75t_L g927 ( .A(n_830), .Y(n_927) );
AND2x2_ASAP7_75t_L g830 ( .A(n_831), .B(n_837), .Y(n_830) );
OR2x2_ASAP7_75t_L g877 ( .A(n_831), .B(n_878), .Y(n_877) );
NOR2xp33_ASAP7_75t_L g883 ( .A(n_831), .B(n_884), .Y(n_883) );
HB1xp67_ASAP7_75t_L g895 ( .A(n_831), .Y(n_895) );
NAND2xp5_ASAP7_75t_L g911 ( .A(n_831), .B(n_878), .Y(n_911) );
AND2x2_ASAP7_75t_L g913 ( .A(n_831), .B(n_887), .Y(n_913) );
NAND2xp5_ASAP7_75t_L g946 ( .A(n_831), .B(n_947), .Y(n_946) );
OR2x2_ASAP7_75t_L g948 ( .A(n_831), .B(n_838), .Y(n_948) );
NOR2xp33_ASAP7_75t_L g974 ( .A(n_831), .B(n_845), .Y(n_974) );
INVx3_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g853 ( .A(n_832), .B(n_854), .Y(n_853) );
INVx1_ASAP7_75t_L g918 ( .A(n_832), .Y(n_918) );
OR2x2_ASAP7_75t_L g998 ( .A(n_832), .B(n_845), .Y(n_998) );
AND2x2_ASAP7_75t_L g832 ( .A(n_833), .B(n_835), .Y(n_832) );
INVx1_ASAP7_75t_L g837 ( .A(n_838), .Y(n_837) );
NOR2xp33_ASAP7_75t_L g965 ( .A(n_838), .B(n_853), .Y(n_965) );
NOR2xp33_ASAP7_75t_L g1006 ( .A(n_838), .B(n_854), .Y(n_1006) );
OR2x2_ASAP7_75t_L g838 ( .A(n_839), .B(n_845), .Y(n_838) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_839), .Y(n_878) );
AND2x2_ASAP7_75t_L g887 ( .A(n_839), .B(n_845), .Y(n_887) );
OAI221xp5_ASAP7_75t_SL g988 ( .A1(n_839), .A2(n_989), .B1(n_991), .B2(n_993), .C(n_994), .Y(n_988) );
AND2x2_ASAP7_75t_L g839 ( .A(n_840), .B(n_844), .Y(n_839) );
INVx1_ASAP7_75t_L g851 ( .A(n_845), .Y(n_851) );
OR2x2_ASAP7_75t_L g884 ( .A(n_845), .B(n_878), .Y(n_884) );
AND2x2_ASAP7_75t_L g894 ( .A(n_845), .B(n_895), .Y(n_894) );
AND2x2_ASAP7_75t_L g897 ( .A(n_845), .B(n_878), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g954 ( .A(n_845), .B(n_917), .Y(n_954) );
AND2x2_ASAP7_75t_L g845 ( .A(n_846), .B(n_848), .Y(n_845) );
INVx1_ASAP7_75t_L g849 ( .A(n_850), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g850 ( .A(n_851), .B(n_852), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g938 ( .A(n_852), .B(n_939), .Y(n_938) );
AOI211xp5_ASAP7_75t_L g989 ( .A1(n_852), .A2(n_884), .B(n_916), .C(n_990), .Y(n_989) );
INVx1_ASAP7_75t_L g852 ( .A(n_853), .Y(n_852) );
INVx1_ASAP7_75t_SL g875 ( .A(n_854), .Y(n_875) );
AND2x2_ASAP7_75t_L g916 ( .A(n_854), .B(n_897), .Y(n_916) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_854), .B(n_860), .Y(n_921) );
AND2x2_ASAP7_75t_L g979 ( .A(n_854), .B(n_971), .Y(n_979) );
A2O1A1Ixp33_ASAP7_75t_SL g923 ( .A1(n_855), .A2(n_924), .B(n_925), .C(n_928), .Y(n_923) );
INVx1_ASAP7_75t_L g949 ( .A(n_855), .Y(n_949) );
NOR2xp33_ASAP7_75t_L g963 ( .A(n_855), .B(n_892), .Y(n_963) );
AND2x2_ASAP7_75t_L g855 ( .A(n_856), .B(n_859), .Y(n_855) );
CKINVDCx6p67_ASAP7_75t_R g873 ( .A(n_856), .Y(n_873) );
INVx1_ASAP7_75t_L g882 ( .A(n_856), .Y(n_882) );
OR2x2_ASAP7_75t_L g889 ( .A(n_856), .B(n_860), .Y(n_889) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_856), .A2(n_873), .B1(n_906), .B2(n_920), .Y(n_905) );
AND2x2_ASAP7_75t_L g956 ( .A(n_856), .B(n_860), .Y(n_956) );
OR2x2_ASAP7_75t_L g996 ( .A(n_856), .B(n_866), .Y(n_996) );
OR2x6_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
INVx1_ASAP7_75t_L g908 ( .A(n_859), .Y(n_908) );
CKINVDCx5p33_ASAP7_75t_R g859 ( .A(n_860), .Y(n_859) );
BUFx2_ASAP7_75t_L g899 ( .A(n_860), .Y(n_899) );
HB1xp67_ASAP7_75t_L g977 ( .A(n_860), .Y(n_977) );
AND2x4_ASAP7_75t_L g860 ( .A(n_861), .B(n_863), .Y(n_860) );
OAI211xp5_ASAP7_75t_L g864 ( .A1(n_865), .A2(n_874), .B(n_879), .C(n_893), .Y(n_864) );
NAND2xp5_ASAP7_75t_L g865 ( .A(n_866), .B(n_873), .Y(n_865) );
AND2x2_ASAP7_75t_L g880 ( .A(n_866), .B(n_881), .Y(n_880) );
INVx3_ASAP7_75t_L g892 ( .A(n_866), .Y(n_892) );
AND2x2_ASAP7_75t_L g898 ( .A(n_866), .B(n_899), .Y(n_898) );
INVx3_ASAP7_75t_L g866 ( .A(n_867), .Y(n_866) );
OR2x2_ASAP7_75t_L g888 ( .A(n_867), .B(n_889), .Y(n_888) );
OR2x2_ASAP7_75t_L g960 ( .A(n_867), .B(n_961), .Y(n_960) );
NOR2xp33_ASAP7_75t_L g969 ( .A(n_867), .B(n_900), .Y(n_969) );
AND2x2_ASAP7_75t_L g992 ( .A(n_867), .B(n_881), .Y(n_992) );
NAND2xp5_ASAP7_75t_L g867 ( .A(n_868), .B(n_872), .Y(n_867) );
INVx2_ASAP7_75t_L g869 ( .A(n_870), .Y(n_869) );
INVx2_ASAP7_75t_SL g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g934 ( .A(n_873), .Y(n_934) );
AND2x2_ASAP7_75t_L g985 ( .A(n_873), .B(n_899), .Y(n_985) );
OAI222xp33_ASAP7_75t_SL g1000 ( .A1(n_873), .A2(n_968), .B1(n_1001), .B2(n_1002), .C1(n_1004), .C2(n_1011), .Y(n_1000) );
A2O1A1Ixp33_ASAP7_75t_L g975 ( .A1(n_874), .A2(n_976), .B(n_977), .C(n_978), .Y(n_975) );
AOI21xp33_ASAP7_75t_SL g1010 ( .A1(n_874), .A2(n_889), .B(n_973), .Y(n_1010) );
NAND2xp5_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .Y(n_874) );
NAND2xp5_ASAP7_75t_L g909 ( .A(n_875), .B(n_910), .Y(n_909) );
NAND2xp5_ASAP7_75t_L g973 ( .A(n_875), .B(n_974), .Y(n_973) );
AND2x2_ASAP7_75t_L g983 ( .A(n_875), .B(n_897), .Y(n_983) );
NAND2xp5_ASAP7_75t_L g993 ( .A(n_875), .B(n_985), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g1022 ( .A(n_875), .B(n_1023), .Y(n_1022) );
INVx1_ASAP7_75t_L g876 ( .A(n_877), .Y(n_876) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_877), .B(n_927), .Y(n_926) );
NOR2xp33_ASAP7_75t_L g1023 ( .A(n_878), .B(n_917), .Y(n_1023) );
AOI211xp5_ASAP7_75t_L g879 ( .A1(n_880), .A2(n_883), .B(n_885), .C(n_890), .Y(n_879) );
AOI21xp5_ASAP7_75t_L g966 ( .A1(n_880), .A2(n_967), .B(n_968), .Y(n_966) );
INVx1_ASAP7_75t_L g1015 ( .A(n_880), .Y(n_1015) );
INVx2_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g976 ( .A(n_883), .Y(n_976) );
INVx1_ASAP7_75t_L g939 ( .A(n_884), .Y(n_939) );
NOR2xp33_ASAP7_75t_L g964 ( .A(n_884), .B(n_931), .Y(n_964) );
NOR2xp33_ASAP7_75t_L g885 ( .A(n_886), .B(n_888), .Y(n_885) );
NOR3xp33_ASAP7_75t_L g890 ( .A(n_886), .B(n_891), .C(n_892), .Y(n_890) );
NOR2xp33_ASAP7_75t_L g990 ( .A(n_886), .B(n_952), .Y(n_990) );
INVx1_ASAP7_75t_L g886 ( .A(n_887), .Y(n_886) );
INVx2_ASAP7_75t_L g971 ( .A(n_889), .Y(n_971) );
NAND2xp5_ASAP7_75t_L g940 ( .A(n_892), .B(n_900), .Y(n_940) );
INVx5_ASAP7_75t_L g942 ( .A(n_892), .Y(n_942) );
INVx3_ASAP7_75t_L g999 ( .A(n_892), .Y(n_999) );
OAI21xp33_ASAP7_75t_L g978 ( .A1(n_894), .A2(n_939), .B(n_979), .Y(n_978) );
AND2x2_ASAP7_75t_L g896 ( .A(n_895), .B(n_897), .Y(n_896) );
OAI21xp5_ASAP7_75t_L g1001 ( .A1(n_896), .A2(n_939), .B(n_979), .Y(n_1001) );
AND2x2_ASAP7_75t_L g929 ( .A(n_897), .B(n_930), .Y(n_929) );
AND2x2_ASAP7_75t_L g967 ( .A(n_897), .B(n_917), .Y(n_967) );
INVx1_ASAP7_75t_L g1008 ( .A(n_897), .Y(n_1008) );
AOI22xp5_ASAP7_75t_L g962 ( .A1(n_898), .A2(n_963), .B1(n_964), .B2(n_965), .Y(n_962) );
OAI21xp33_ASAP7_75t_L g994 ( .A1(n_899), .A2(n_995), .B(n_997), .Y(n_994) );
INVx2_ASAP7_75t_L g968 ( .A(n_900), .Y(n_968) );
HB1xp67_ASAP7_75t_SL g1003 ( .A(n_900), .Y(n_1003) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_900), .B(n_985), .Y(n_1020) );
OAI211xp5_ASAP7_75t_L g906 ( .A1(n_907), .A2(n_909), .B(n_912), .C(n_914), .Y(n_906) );
AOI211xp5_ASAP7_75t_L g935 ( .A1(n_907), .A2(n_926), .B(n_936), .C(n_937), .Y(n_935) );
INVx1_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g919 ( .A(n_908), .Y(n_919) );
INVx1_ASAP7_75t_L g910 ( .A(n_911), .Y(n_910) );
NOR2xp33_ASAP7_75t_L g920 ( .A(n_911), .B(n_921), .Y(n_920) );
O2A1O1Ixp33_ASAP7_75t_SL g932 ( .A1(n_912), .A2(n_933), .B(n_935), .C(n_940), .Y(n_932) );
INVx1_ASAP7_75t_L g924 ( .A(n_913), .Y(n_924) );
INVx1_ASAP7_75t_L g914 ( .A(n_915), .Y(n_914) );
O2A1O1Ixp33_ASAP7_75t_L g944 ( .A1(n_915), .A2(n_933), .B(n_937), .C(n_945), .Y(n_944) );
AND3x1_ASAP7_75t_L g915 ( .A(n_916), .B(n_917), .C(n_919), .Y(n_915) );
AND2x2_ASAP7_75t_L g987 ( .A(n_917), .B(n_983), .Y(n_987) );
NAND2xp5_ASAP7_75t_L g1017 ( .A(n_917), .B(n_1018), .Y(n_1017) );
INVx3_ASAP7_75t_L g917 ( .A(n_918), .Y(n_917) );
AOI22xp5_ASAP7_75t_L g922 ( .A1(n_923), .A2(n_932), .B1(n_941), .B2(n_943), .Y(n_922) );
NOR2xp33_ASAP7_75t_L g951 ( .A(n_927), .B(n_952), .Y(n_951) );
INVx1_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
CKINVDCx14_ASAP7_75t_R g933 ( .A(n_934), .Y(n_933) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
CKINVDCx14_ASAP7_75t_R g941 ( .A(n_942), .Y(n_941) );
NAND2xp5_ASAP7_75t_L g943 ( .A(n_944), .B(n_950), .Y(n_943) );
AOI21xp5_ASAP7_75t_SL g945 ( .A1(n_946), .A2(n_948), .B(n_949), .Y(n_945) );
OAI211xp5_ASAP7_75t_SL g1012 ( .A1(n_946), .A2(n_960), .B(n_1013), .C(n_1024), .Y(n_1012) );
NOR2xp33_ASAP7_75t_L g953 ( .A(n_954), .B(n_955), .Y(n_953) );
OAI211xp5_ASAP7_75t_L g959 ( .A1(n_954), .A2(n_960), .B(n_962), .C(n_966), .Y(n_959) );
INVx2_ASAP7_75t_L g961 ( .A(n_956), .Y(n_961) );
O2A1O1Ixp33_ASAP7_75t_SL g957 ( .A1(n_958), .A2(n_969), .B(n_970), .C(n_986), .Y(n_957) );
INVxp67_ASAP7_75t_L g958 ( .A(n_959), .Y(n_958) );
O2A1O1Ixp33_ASAP7_75t_L g986 ( .A1(n_959), .A2(n_987), .B(n_988), .C(n_999), .Y(n_986) );
INVx1_ASAP7_75t_L g1025 ( .A(n_960), .Y(n_1025) );
INVx1_ASAP7_75t_L g1005 ( .A(n_961), .Y(n_1005) );
INVx1_ASAP7_75t_L g981 ( .A(n_965), .Y(n_981) );
NAND2xp5_ASAP7_75t_L g1024 ( .A(n_967), .B(n_1025), .Y(n_1024) );
AOI211xp5_ASAP7_75t_L g970 ( .A1(n_971), .A2(n_972), .B(n_975), .C(n_980), .Y(n_970) );
INVx1_ASAP7_75t_L g972 ( .A(n_973), .Y(n_972) );
NAND2xp33_ASAP7_75t_SL g1014 ( .A(n_977), .B(n_1015), .Y(n_1014) );
AOI21xp33_ASAP7_75t_L g980 ( .A1(n_981), .A2(n_982), .B(n_984), .Y(n_980) );
INVx1_ASAP7_75t_L g982 ( .A(n_983), .Y(n_982) );
INVx1_ASAP7_75t_L g984 ( .A(n_985), .Y(n_984) );
INVx1_ASAP7_75t_L g1011 ( .A(n_987), .Y(n_1011) );
INVx1_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
INVx1_ASAP7_75t_L g995 ( .A(n_996), .Y(n_995) );
INVxp67_ASAP7_75t_L g1002 ( .A(n_1003), .Y(n_1002) );
AOI211xp5_ASAP7_75t_L g1004 ( .A1(n_1005), .A2(n_1006), .B(n_1007), .C(n_1010), .Y(n_1004) );
NOR2xp33_ASAP7_75t_L g1007 ( .A(n_1008), .B(n_1009), .Y(n_1007) );
AOI22xp33_ASAP7_75t_L g1013 ( .A1(n_1014), .A2(n_1016), .B1(n_1019), .B2(n_1021), .Y(n_1013) );
INVx1_ASAP7_75t_L g1016 ( .A(n_1017), .Y(n_1016) );
INVxp33_ASAP7_75t_L g1019 ( .A(n_1020), .Y(n_1019) );
INVxp33_ASAP7_75t_SL g1021 ( .A(n_1022), .Y(n_1021) );
CKINVDCx5p33_ASAP7_75t_R g1026 ( .A(n_1027), .Y(n_1026) );
INVx1_ASAP7_75t_L g1027 ( .A(n_1028), .Y(n_1027) );
INVx1_ASAP7_75t_L g1029 ( .A(n_1030), .Y(n_1029) );
HB1xp67_ASAP7_75t_SL g1030 ( .A(n_1031), .Y(n_1030) );
INVx2_ASAP7_75t_L g1031 ( .A(n_1032), .Y(n_1031) );
OR2x2_ASAP7_75t_L g1033 ( .A(n_1034), .B(n_1041), .Y(n_1033) );
NAND4xp25_ASAP7_75t_L g1034 ( .A(n_1035), .B(n_1036), .C(n_1037), .D(n_1038), .Y(n_1034) );
NAND4xp25_ASAP7_75t_L g1041 ( .A(n_1042), .B(n_1043), .C(n_1044), .D(n_1045), .Y(n_1041) );
INVx1_ASAP7_75t_L g1046 ( .A(n_1047), .Y(n_1046) );
HB1xp67_ASAP7_75t_L g1047 ( .A(n_1048), .Y(n_1047) );
INVx1_ASAP7_75t_L g1054 ( .A(n_1055), .Y(n_1054) );
HB1xp67_ASAP7_75t_L g1055 ( .A(n_1056), .Y(n_1055) );
NOR2x1_ASAP7_75t_L g1056 ( .A(n_1057), .B(n_1065), .Y(n_1056) );
NAND3xp33_ASAP7_75t_L g1057 ( .A(n_1058), .B(n_1061), .C(n_1064), .Y(n_1057) );
NAND4xp25_ASAP7_75t_L g1065 ( .A(n_1066), .B(n_1068), .C(n_1069), .D(n_1070), .Y(n_1065) );
BUFx2_ASAP7_75t_SL g1071 ( .A(n_1072), .Y(n_1071) );
BUFx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
endmodule