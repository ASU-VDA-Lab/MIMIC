module real_jpeg_26015_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_13;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_16;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_14;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_15;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_0),
.A2(n_52),
.B1(n_56),
.B2(n_57),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_0),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_0),
.A2(n_42),
.B1(n_43),
.B2(n_56),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_0),
.A2(n_22),
.B1(n_26),
.B2(n_56),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_0),
.A2(n_28),
.B1(n_30),
.B2(n_56),
.Y(n_164)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx8_ASAP7_75t_SL g60 ( 
.A(n_4),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g33 ( 
.A1(n_5),
.A2(n_22),
.B1(n_26),
.B2(n_34),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_5),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_5),
.A2(n_34),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_5),
.A2(n_34),
.B1(n_57),
.B2(n_58),
.Y(n_77)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_5),
.A2(n_28),
.B1(n_30),
.B2(n_34),
.Y(n_108)
);

O2A1O1Ixp33_ASAP7_75t_L g201 ( 
.A1(n_5),
.A2(n_61),
.B(n_202),
.C(n_203),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_5),
.B(n_59),
.Y(n_217)
);

O2A1O1Ixp33_ASAP7_75t_L g227 ( 
.A1(n_5),
.A2(n_38),
.B(n_43),
.C(n_228),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_5),
.B(n_25),
.C(n_28),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g249 ( 
.A(n_5),
.B(n_87),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_5),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_5),
.B(n_27),
.Y(n_275)
);

BUFx5_ASAP7_75t_L g38 ( 
.A(n_6),
.Y(n_38)
);

OAI22xp33_ASAP7_75t_SL g138 ( 
.A1(n_7),
.A2(n_55),
.B1(n_66),
.B2(n_139),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_7),
.Y(n_139)
);

OAI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_7),
.A2(n_42),
.B1(n_43),
.B2(n_139),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g232 ( 
.A1(n_7),
.A2(n_22),
.B1(n_26),
.B2(n_139),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_SL g257 ( 
.A1(n_7),
.A2(n_28),
.B1(n_30),
.B2(n_139),
.Y(n_257)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_8),
.A2(n_42),
.B1(n_43),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_8),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_8),
.A2(n_49),
.B1(n_55),
.B2(n_58),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_8),
.A2(n_22),
.B1(n_26),
.B2(n_49),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g130 ( 
.A1(n_8),
.A2(n_28),
.B1(n_30),
.B2(n_49),
.Y(n_130)
);

INVx13_ASAP7_75t_L g55 ( 
.A(n_9),
.Y(n_55)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g107 ( 
.A(n_11),
.Y(n_107)
);

INVx3_ASAP7_75t_L g206 ( 
.A(n_11),
.Y(n_206)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_11),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_80),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_78),
.Y(n_13)
);

NAND2xp5_ASAP7_75t_SL g14 ( 
.A(n_15),
.B(n_74),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_15),
.B(n_74),
.Y(n_79)
);

MAJIxp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_68),
.C(n_69),
.Y(n_15)
);

AOI22xp33_ASAP7_75t_SL g318 ( 
.A1(n_16),
.A2(n_17),
.B1(n_319),
.B2(n_320),
.Y(n_318)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

MAJIxp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_35),
.C(n_50),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g96 ( 
.A1(n_18),
.A2(n_97),
.B1(n_98),
.B2(n_101),
.Y(n_96)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_18),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_18),
.A2(n_35),
.B1(n_101),
.B2(n_147),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_18),
.A2(n_101),
.B1(n_186),
.B2(n_213),
.Y(n_212)
);

AOI21xp5_ASAP7_75t_SL g18 ( 
.A1(n_19),
.A2(n_31),
.B(n_32),
.Y(n_18)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_19),
.A2(n_111),
.B(n_112),
.Y(n_110)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_20),
.B(n_92),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_20),
.B(n_33),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_20),
.B(n_232),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_27),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_24),
.B1(n_25),
.B2(n_26),
.Y(n_21)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_22),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_22),
.A2(n_26),
.B1(n_38),
.B2(n_39),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_22),
.B(n_245),
.Y(n_244)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_24),
.A2(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_27)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

OAI21xp33_ASAP7_75t_L g228 ( 
.A1(n_26),
.A2(n_34),
.B(n_39),
.Y(n_228)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_27),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_27),
.B(n_92),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_27),
.B(n_232),
.Y(n_242)
);

INVx6_ASAP7_75t_SL g30 ( 
.A(n_28),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_28),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g268 ( 
.A(n_28),
.B(n_269),
.Y(n_268)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_31),
.B(n_32),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_31),
.A2(n_91),
.B(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

OAI21xp33_ASAP7_75t_L g202 ( 
.A1(n_34),
.A2(n_43),
.B(n_60),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_35),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_36),
.B(n_45),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g194 ( 
.A(n_36),
.B(n_195),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_47),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_40),
.B(n_46),
.Y(n_68)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_SL g100 ( 
.A(n_37),
.B(n_48),
.Y(n_100)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_38),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_38),
.A2(n_39),
.B1(n_42),
.B2(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_41),
.B(n_99),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_42),
.A2(n_43),
.B1(n_60),
.B2(n_61),
.Y(n_59)
);

INVx3_ASAP7_75t_SL g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g85 ( 
.A1(n_45),
.A2(n_86),
.B(n_87),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g186 ( 
.A(n_45),
.B(n_187),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_46),
.B(n_48),
.Y(n_45)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_46),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_46),
.B(n_196),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_50),
.B(n_146),
.Y(n_145)
);

AOI21xp5_ASAP7_75t_L g50 ( 
.A1(n_51),
.A2(n_59),
.B(n_62),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_51),
.Y(n_72)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_55),
.Y(n_58)
);

INVx11_ASAP7_75t_L g66 ( 
.A(n_55),
.Y(n_66)
);

INVx8_ASAP7_75t_L g204 ( 
.A(n_55),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_60),
.B1(n_61),
.B2(n_66),
.Y(n_65)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_59),
.B(n_67),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_59),
.B(n_77),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_59),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_59),
.B(n_138),
.Y(n_172)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_60),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_62),
.B(n_75),
.Y(n_74)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_63),
.B(n_172),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_67),
.Y(n_63)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_64),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_64),
.B(n_77),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_64),
.B(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_68),
.B(n_161),
.C(n_171),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_68),
.A2(n_171),
.B1(n_304),
.B2(n_305),
.Y(n_303)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_68),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_68),
.A2(n_69),
.B1(n_70),
.B2(n_304),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_70),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_71),
.A2(n_72),
.B(n_73),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_71),
.A2(n_115),
.B(n_116),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_73),
.B(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_73),
.B(n_137),
.Y(n_197)
);

INVxp33_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_76),
.B(n_137),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_77),
.Y(n_116)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_317),
.B(n_322),
.Y(n_80)
);

OAI211xp5_ASAP7_75t_L g81 ( 
.A1(n_82),
.A2(n_140),
.B(n_150),
.C(n_316),
.Y(n_81)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_117),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_83),
.B(n_117),
.Y(n_151)
);

BUFx24_ASAP7_75t_SL g323 ( 
.A(n_83),
.Y(n_323)
);

FAx1_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_93),
.CI(n_104),
.CON(n_83),
.SN(n_83)
);

OAI21xp5_ASAP7_75t_SL g122 ( 
.A1(n_84),
.A2(n_85),
.B(n_88),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_84),
.B(n_93),
.C(n_104),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_88),
.Y(n_84)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_86),
.A2(n_99),
.B(n_100),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_87),
.B(n_189),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_90),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_89),
.B(n_230),
.Y(n_229)
);

INVxp33_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_91),
.B(n_242),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_96),
.B1(n_102),
.B2(n_103),
.Y(n_93)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_94),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_L g144 ( 
.A1(n_94),
.A2(n_102),
.B1(n_145),
.B2(n_148),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_94),
.B(n_98),
.C(n_101),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_94),
.B(n_145),
.C(n_149),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_95),
.B(n_172),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_96),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_100),
.B(n_133),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_100),
.B(n_195),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_101),
.B(n_184),
.C(n_186),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_105),
.A2(n_109),
.B(n_113),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_110),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_105),
.A2(n_113),
.B1(n_114),
.B2(n_121),
.Y(n_120)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_105),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_105),
.A2(n_110),
.B1(n_121),
.B2(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_105),
.B(n_227),
.Y(n_226)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_105),
.A2(n_121),
.B1(n_227),
.B2(n_287),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_107),
.B(n_108),
.Y(n_105)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_106),
.B(n_130),
.Y(n_129)
);

OAI21xp5_ASAP7_75t_SL g163 ( 
.A1(n_106),
.A2(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g219 ( 
.A(n_106),
.B(n_108),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_106),
.B(n_256),
.Y(n_255)
);

INVx3_ASAP7_75t_SL g127 ( 
.A(n_107),
.Y(n_127)
);

INVx5_ASAP7_75t_L g168 ( 
.A(n_107),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g128 ( 
.A(n_108),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_110),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_112),
.B(n_170),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_112),
.B(n_231),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_122),
.C(n_123),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_118),
.A2(n_119),
.B1(n_122),
.B2(n_175),
.Y(n_174)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_122),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_174),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_132),
.C(n_135),
.Y(n_123)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_124),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_131),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_125),
.B(n_131),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_129),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_126),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_128),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_129),
.A2(n_164),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_129),
.B(n_262),
.Y(n_261)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_130),
.B(n_167),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_132),
.A2(n_135),
.B1(n_136),
.B2(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_132),
.Y(n_157)
);

CKINVDCx14_ASAP7_75t_R g133 ( 
.A(n_134),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_134),
.B(n_188),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

NAND3xp33_ASAP7_75t_SL g150 ( 
.A(n_141),
.B(n_151),
.C(n_152),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_143),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g316 ( 
.A(n_142),
.B(n_143),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g143 ( 
.A(n_144),
.B(n_149),
.Y(n_143)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_145),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_153),
.A2(n_176),
.B(n_315),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_173),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g315 ( 
.A(n_154),
.B(n_173),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.C(n_160),
.Y(n_154)
);

XOR2xp5_ASAP7_75t_L g313 ( 
.A(n_155),
.B(n_158),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_160),
.B(n_313),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_161),
.A2(n_162),
.B1(n_302),
.B2(n_303),
.Y(n_301)
);

CKINVDCx16_ASAP7_75t_R g161 ( 
.A(n_162),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_169),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g182 ( 
.A(n_163),
.B(n_169),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_166),
.B(n_219),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_166),
.B(n_255),
.Y(n_276)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_170),
.B(n_242),
.Y(n_241)
);

CKINVDCx14_ASAP7_75t_R g305 ( 
.A(n_171),
.Y(n_305)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_310),
.B(n_314),
.Y(n_176)
);

A2O1A1Ixp33_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_220),
.B(n_296),
.C(n_309),
.Y(n_177)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_208),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_179),
.B(n_208),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_181),
.B1(n_192),
.B2(n_207),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_190),
.B2(n_191),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g190 ( 
.A(n_182),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_182),
.B(n_191),
.C(n_207),
.Y(n_297)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_183),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_184),
.A2(n_185),
.B1(n_211),
.B2(n_212),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_186),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_188),
.Y(n_187)
);

INVxp67_ASAP7_75t_SL g196 ( 
.A(n_189),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_192),
.Y(n_207)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_200),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_194),
.A2(n_197),
.B1(n_198),
.B2(n_199),
.Y(n_193)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_194),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_194),
.B(n_199),
.C(n_200),
.Y(n_308)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_197),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_201),
.B(n_205),
.Y(n_214)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx3_ASAP7_75t_L g263 ( 
.A(n_206),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_214),
.C(n_215),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_209),
.A2(n_210),
.B1(n_234),
.B2(n_235),
.Y(n_233)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_215),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.C(n_218),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_216),
.B(n_225),
.Y(n_224)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_217),
.B(n_218),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_219),
.B(n_273),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_221),
.B(n_295),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g221 ( 
.A1(n_222),
.A2(n_236),
.B(n_294),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_233),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_223),
.B(n_233),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.C(n_229),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_224),
.B(n_292),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_226),
.B(n_229),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g287 ( 
.A(n_227),
.Y(n_287)
);

INVxp33_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_289),
.B(n_293),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_238),
.A2(n_280),
.B(n_288),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g238 ( 
.A1(n_239),
.A2(n_259),
.B(n_279),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_246),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_240),
.B(n_246),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_241),
.A2(n_243),
.B1(n_244),
.B2(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g243 ( 
.A(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_253),
.B2(n_258),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_250),
.B1(n_251),
.B2(n_252),
.Y(n_248)
);

CKINVDCx14_ASAP7_75t_R g251 ( 
.A(n_249),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_249),
.B(n_252),
.C(n_258),
.Y(n_281)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_253),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g256 ( 
.A(n_257),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_257),
.B(n_263),
.Y(n_262)
);

OAI21xp5_ASAP7_75t_SL g259 ( 
.A1(n_260),
.A2(n_266),
.B(n_278),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_264),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_261),
.B(n_264),
.Y(n_278)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_262),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_267),
.A2(n_274),
.B(n_277),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_272),
.Y(n_267)
);

INVx5_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_275),
.B(n_276),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_282),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_283),
.B(n_286),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_284),
.B(n_285),
.C(n_286),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_291),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g293 ( 
.A(n_290),
.B(n_291),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_298),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g309 ( 
.A(n_297),
.B(n_298),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_308),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g299 ( 
.A1(n_300),
.A2(n_301),
.B1(n_306),
.B2(n_307),
.Y(n_299)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_300),
.B(n_307),
.C(n_308),
.Y(n_311)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_312),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_311),
.B(n_312),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_321),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g322 ( 
.A(n_318),
.B(n_321),
.Y(n_322)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_319),
.Y(n_320)
);


endmodule