module fake_jpeg_22442_n_301 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_301);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_301;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_300;
wire n_211;
wire n_299;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_91;
wire n_93;
wire n_54;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_270;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_265;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

BUFx12f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_15),
.B(n_12),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx11_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_6),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

INVx8_ASAP7_75t_L g35 ( 
.A(n_22),
.Y(n_35)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_22),
.Y(n_36)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_37),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_21),
.B(n_7),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_23),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

BUFx24_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx2_ASAP7_75t_SL g59 ( 
.A(n_41),
.Y(n_59)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_42),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_19),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_44),
.B(n_46),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g46 ( 
.A(n_41),
.B(n_23),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_36),
.A2(n_25),
.B1(n_31),
.B2(n_23),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_47),
.A2(n_51),
.B1(n_36),
.B2(n_35),
.Y(n_67)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_43),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_49),
.B(n_62),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_36),
.A2(n_31),
.B1(n_23),
.B2(n_27),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_53),
.B(n_64),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_43),
.Y(n_56)
);

INVx8_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_58),
.Y(n_89)
);

OA22x2_ASAP7_75t_L g60 ( 
.A1(n_41),
.A2(n_18),
.B1(n_33),
.B2(n_23),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_60),
.A2(n_42),
.B1(n_35),
.B2(n_41),
.Y(n_75)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_L g63 ( 
.A1(n_36),
.A2(n_27),
.B1(n_17),
.B2(n_32),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g72 ( 
.A1(n_63),
.A2(n_29),
.B1(n_24),
.B2(n_34),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_34),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_38),
.B(n_17),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_24),
.Y(n_81)
);

AOI21xp33_ASAP7_75t_SL g66 ( 
.A1(n_41),
.A2(n_43),
.B(n_39),
.Y(n_66)
);

AOI22xp5_ASAP7_75t_SL g68 ( 
.A1(n_66),
.A2(n_36),
.B1(n_42),
.B2(n_35),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_67),
.A2(n_80),
.B1(n_59),
.B2(n_40),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_68),
.A2(n_82),
.B1(n_88),
.B2(n_67),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_59),
.A2(n_34),
.B1(n_19),
.B2(n_31),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g102 ( 
.A1(n_69),
.A2(n_71),
.B1(n_75),
.B2(n_79),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_66),
.A2(n_35),
.B1(n_42),
.B2(n_37),
.Y(n_71)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_72),
.A2(n_78),
.B1(n_40),
.B2(n_20),
.Y(n_109)
);

BUFx2_ASAP7_75t_L g74 ( 
.A(n_61),
.Y(n_74)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_74),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_44),
.B(n_35),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_77),
.B(n_85),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_57),
.A2(n_42),
.B1(n_37),
.B2(n_45),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_57),
.A2(n_42),
.B1(n_37),
.B2(n_43),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_18),
.B1(n_33),
.B2(n_29),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_81),
.B(n_83),
.Y(n_103)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_46),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_64),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_45),
.B(n_26),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_45),
.B(n_26),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_55),
.Y(n_108)
);

INVx5_ASAP7_75t_L g87 ( 
.A(n_48),
.Y(n_87)
);

INVx4_ASAP7_75t_L g120 ( 
.A(n_87),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_37),
.B1(n_41),
.B2(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_48),
.Y(n_91)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_91),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_28),
.Y(n_92)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_92),
.Y(n_114)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_55),
.Y(n_93)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_93),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_95),
.B(n_111),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_77),
.B(n_46),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_96),
.B(n_104),
.Y(n_126)
);

AOI21xp5_ASAP7_75t_L g127 ( 
.A1(n_97),
.A2(n_69),
.B(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_68),
.A2(n_50),
.B1(n_52),
.B2(n_62),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g125 ( 
.A1(n_98),
.A2(n_101),
.B1(n_106),
.B2(n_109),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_33),
.B1(n_60),
.B2(n_41),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g124 ( 
.A(n_99),
.Y(n_124)
);

OR2x4_ASAP7_75t_L g100 ( 
.A(n_68),
.B(n_41),
.Y(n_100)
);

XNOR2xp5_ASAP7_75t_SL g144 ( 
.A(n_100),
.B(n_113),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_71),
.A2(n_75),
.B1(n_73),
.B2(n_82),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_90),
.B(n_49),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_75),
.A2(n_52),
.B1(n_60),
.B2(n_40),
.Y(n_106)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_80),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_107),
.B(n_117),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_108),
.B(n_70),
.Y(n_141)
);

AND2x2_ASAP7_75t_SL g110 ( 
.A(n_83),
.B(n_60),
.Y(n_110)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_110),
.B(n_112),
.C(n_79),
.Y(n_132)
);

AND2x4_ASAP7_75t_L g111 ( 
.A(n_88),
.B(n_60),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_88),
.B(n_39),
.C(n_58),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_85),
.B(n_0),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_72),
.A2(n_40),
.B1(n_28),
.B2(n_32),
.Y(n_115)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_115),
.Y(n_135)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_76),
.Y(n_117)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_76),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_91),
.Y(n_130)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_108),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_121),
.B(n_122),
.Y(n_168)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_103),
.Y(n_122)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_120),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_123),
.B(n_129),
.Y(n_174)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_128),
.B(n_124),
.Y(n_166)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_120),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_SL g154 ( 
.A(n_130),
.B(n_142),
.Y(n_154)
);

O2A1O1Ixp33_ASAP7_75t_L g131 ( 
.A1(n_102),
.A2(n_78),
.B(n_86),
.C(n_89),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_131),
.A2(n_84),
.B1(n_55),
.B2(n_26),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_137),
.C(n_149),
.Y(n_150)
);

AOI22x1_ASAP7_75t_SL g134 ( 
.A1(n_100),
.A2(n_89),
.B1(n_79),
.B2(n_90),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_134),
.A2(n_94),
.B1(n_116),
.B2(n_118),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_92),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_141),
.Y(n_178)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_96),
.B(n_81),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_105),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_138),
.B(n_139),
.Y(n_162)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_140),
.B(n_147),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_103),
.B(n_30),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_56),
.Y(n_143)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_143),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g145 ( 
.A(n_117),
.B(n_20),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_114),
.B(n_110),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_113),
.B(n_56),
.Y(n_146)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_146),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_114),
.B(n_87),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_84),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_101),
.B(n_39),
.C(n_58),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_127),
.A2(n_111),
.B1(n_99),
.B2(n_102),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_151),
.A2(n_153),
.B1(n_156),
.B2(n_164),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_130),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_149),
.A2(n_111),
.B1(n_95),
.B2(n_98),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_133),
.A2(n_111),
.B1(n_110),
.B2(n_106),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_110),
.C(n_119),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_157),
.B(n_159),
.C(n_161),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_SL g187 ( 
.A(n_158),
.B(n_163),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_111),
.C(n_94),
.Y(n_159)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_160),
.B(n_169),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_137),
.B(n_39),
.Y(n_161)
);

FAx1_ASAP7_75t_SL g163 ( 
.A(n_126),
.B(n_39),
.CI(n_54),
.CON(n_163),
.SN(n_163)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_133),
.A2(n_93),
.B1(n_87),
.B2(n_116),
.Y(n_164)
);

AOI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_126),
.A2(n_118),
.B(n_30),
.Y(n_165)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_165),
.A2(n_166),
.B(n_179),
.Y(n_203)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_132),
.B(n_54),
.C(n_39),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_170),
.B(n_175),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_144),
.B(n_54),
.C(n_74),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_171),
.B(n_146),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_173),
.A2(n_129),
.B1(n_123),
.B2(n_122),
.Y(n_186)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_147),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_141),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_176),
.B(n_145),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_148),
.A2(n_84),
.B1(n_26),
.B2(n_22),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_131),
.B1(n_125),
.B2(n_142),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_128),
.A2(n_74),
.B(n_2),
.Y(n_179)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_180),
.B(n_196),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g181 ( 
.A1(n_160),
.A2(n_133),
.B1(n_131),
.B2(n_134),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_181),
.A2(n_186),
.B1(n_194),
.B2(n_197),
.Y(n_207)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_174),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_185),
.Y(n_215)
);

HB1xp67_ASAP7_75t_L g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_184),
.Y(n_228)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_168),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_162),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_189),
.B(n_190),
.Y(n_225)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_178),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_192),
.A2(n_205),
.B(n_163),
.Y(n_219)
);

OAI322xp33_ASAP7_75t_L g193 ( 
.A1(n_178),
.A2(n_136),
.A3(n_144),
.B1(n_143),
.B2(n_139),
.C1(n_134),
.C2(n_121),
.Y(n_193)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_193),
.B(n_9),
.Y(n_221)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_195),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_164),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_173),
.A2(n_133),
.B1(n_125),
.B2(n_135),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g198 ( 
.A(n_177),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_198),
.B(n_200),
.Y(n_212)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_155),
.A2(n_172),
.B1(n_151),
.B2(n_153),
.Y(n_199)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_199),
.Y(n_214)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_157),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_176),
.B(n_144),
.Y(n_204)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_204),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_152),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_202),
.B(n_150),
.Y(n_206)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_206),
.B(n_208),
.C(n_211),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_202),
.B(n_150),
.C(n_161),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_159),
.C(n_169),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_182),
.B(n_171),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_213),
.B(n_221),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_192),
.B(n_172),
.C(n_155),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_223),
.C(n_224),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_196),
.A2(n_166),
.B1(n_175),
.B2(n_156),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_218),
.Y(n_231)
);

AOI322xp5_ASAP7_75t_L g218 ( 
.A1(n_181),
.A2(n_158),
.A3(n_163),
.B1(n_154),
.B2(n_165),
.C1(n_179),
.C2(n_12),
.Y(n_218)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_219),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_198),
.A2(n_154),
.B1(n_10),
.B2(n_11),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_220),
.B(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_182),
.B(n_1),
.C(n_2),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_204),
.B(n_1),
.C(n_2),
.Y(n_224)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_187),
.B(n_9),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_199),
.B(n_10),
.Y(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_225),
.B(n_190),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

INVxp67_ASAP7_75t_SL g230 ( 
.A(n_210),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_203),
.B1(n_227),
.B2(n_226),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_236),
.Y(n_258)
);

NAND4xp25_ASAP7_75t_L g235 ( 
.A(n_217),
.B(n_205),
.C(n_201),
.D(n_191),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_235),
.A2(n_239),
.B1(n_240),
.B2(n_247),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_212),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_214),
.A2(n_197),
.B1(n_191),
.B2(n_180),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_222),
.A2(n_201),
.B(n_183),
.Y(n_240)
);

NOR3xp33_ASAP7_75t_L g242 ( 
.A(n_209),
.B(n_189),
.C(n_185),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_242),
.B(n_246),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_220),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_244),
.B(n_245),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_SL g245 ( 
.A(n_228),
.B(n_186),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_216),
.Y(n_246)
);

AO21x1_ASAP7_75t_L g247 ( 
.A1(n_207),
.A2(n_203),
.B(n_194),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_234),
.B(n_208),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_248),
.B(n_256),
.Y(n_265)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_249),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_234),
.B(n_206),
.C(n_211),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_251),
.B(n_254),
.C(n_255),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g253 ( 
.A(n_233),
.B(n_235),
.Y(n_253)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_253),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_246),
.B(n_223),
.C(n_213),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_237),
.B(n_240),
.C(n_243),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_237),
.B(n_224),
.C(n_188),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_243),
.B(n_1),
.C(n_2),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_257),
.B(n_261),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_239),
.B(n_10),
.Y(n_259)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_259),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g261 ( 
.A(n_238),
.B(n_11),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g264 ( 
.A(n_258),
.B(n_232),
.Y(n_264)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_264),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_250),
.A2(n_232),
.B1(n_229),
.B2(n_247),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g279 ( 
.A1(n_270),
.A2(n_271),
.B1(n_263),
.B2(n_274),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_260),
.A2(n_244),
.B1(n_247),
.B2(n_231),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g272 ( 
.A(n_262),
.B(n_241),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g280 ( 
.A(n_272),
.B(n_13),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g273 ( 
.A(n_252),
.B(n_238),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_273),
.B(n_14),
.Y(n_283)
);

A2O1A1Ixp33_ASAP7_75t_SL g274 ( 
.A1(n_253),
.A2(n_1),
.B(n_3),
.C(n_4),
.Y(n_274)
);

AOI21xp5_ASAP7_75t_L g276 ( 
.A1(n_274),
.A2(n_257),
.B(n_4),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_276),
.B(n_281),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_269),
.B(n_251),
.C(n_255),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_277),
.B(n_265),
.C(n_274),
.Y(n_288)
);

AOI221xp5_ASAP7_75t_L g278 ( 
.A1(n_267),
.A2(n_254),
.B1(n_261),
.B2(n_13),
.C(n_12),
.Y(n_278)
);

OAI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_278),
.A2(n_274),
.B(n_266),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g281 ( 
.A(n_271),
.B(n_13),
.Y(n_281)
);

AOI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_270),
.A2(n_14),
.B(n_16),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_284),
.B(n_16),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_283),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_L g284 ( 
.A1(n_269),
.A2(n_16),
.B(n_4),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_268),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_286),
.B(n_285),
.Y(n_294)
);

AOI321xp33_ASAP7_75t_L g296 ( 
.A1(n_287),
.A2(n_3),
.A3(n_4),
.B1(n_5),
.B2(n_6),
.C(n_260),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_288),
.B(n_277),
.C(n_278),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_291),
.B(n_292),
.Y(n_297)
);

INVxp33_ASAP7_75t_L g292 ( 
.A(n_275),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_293),
.B(n_294),
.Y(n_298)
);

AO21x1_ASAP7_75t_L g295 ( 
.A1(n_292),
.A2(n_289),
.B(n_290),
.Y(n_295)
);

NAND2x1_ASAP7_75t_L g299 ( 
.A(n_295),
.B(n_296),
.Y(n_299)
);

NOR3xp33_ASAP7_75t_L g300 ( 
.A(n_298),
.B(n_297),
.C(n_6),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_300),
.B(n_299),
.Y(n_301)
);


endmodule