module fake_netlist_5_586_n_1987 (n_137, n_168, n_164, n_91, n_82, n_122, n_142, n_176, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_165, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_173, n_25, n_53, n_160, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_55, n_99, n_2, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_171, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_1987);

input n_137;
input n_168;
input n_164;
input n_91;
input n_82;
input n_122;
input n_142;
input n_176;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_165;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_173;
input n_25;
input n_53;
input n_160;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_1987;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_1021;
wire n_1960;
wire n_551;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_447;
wire n_247;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_877;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_929;
wire n_1124;
wire n_1818;
wire n_902;
wire n_1576;
wire n_191;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_320;
wire n_1154;
wire n_1242;
wire n_1135;
wire n_406;
wire n_519;
wire n_1016;
wire n_1243;
wire n_546;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_1778;
wire n_227;
wire n_920;
wire n_1289;
wire n_1517;
wire n_335;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_297;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_1374;
wire n_1328;
wire n_223;
wire n_1948;
wire n_1984;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1097;
wire n_1036;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_1040;
wire n_1872;
wire n_1852;
wire n_578;
wire n_926;
wire n_344;
wire n_1218;
wire n_1931;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_845;
wire n_663;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_923;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_213;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_1471;
wire n_1986;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_1377;
wire n_190;
wire n_989;
wire n_1039;
wire n_228;
wire n_283;
wire n_1403;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_310;
wire n_593;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_1819;
wire n_476;
wire n_1527;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_832;
wire n_857;
wire n_207;
wire n_561;
wire n_1319;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_1532;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_1175;
wire n_817;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_759;
wire n_1892;
wire n_806;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_1571;
wire n_1189;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_776;
wire n_1798;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_526;
wire n_1916;
wire n_372;
wire n_293;
wire n_677;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_1933;
wire n_1656;
wire n_1158;
wire n_1509;
wire n_1874;
wire n_563;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_658;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_978;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_636;
wire n_660;
wire n_1640;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_742;
wire n_750;
wire n_995;
wire n_454;
wire n_1609;
wire n_374;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_218;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_743;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_1240;
wire n_1820;
wire n_829;
wire n_1612;
wire n_1416;
wire n_1724;
wire n_361;
wire n_1237;
wire n_700;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_1390;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_1941;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_1351;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_634;
wire n_199;
wire n_1958;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_302;
wire n_1343;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_212;
wire n_507;
wire n_1560;
wire n_1605;
wire n_330;
wire n_1228;
wire n_972;
wire n_692;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_286;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_918;
wire n_942;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_323;
wire n_195;
wire n_356;
wire n_894;
wire n_1636;
wire n_1730;
wire n_831;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_1940;
wire n_814;
wire n_192;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_1616;
wire n_1446;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_211;
wire n_1824;
wire n_1917;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_336;
wire n_681;
wire n_584;
wire n_1638;
wire n_1786;
wire n_430;
wire n_510;
wire n_216;
wire n_311;
wire n_830;
wire n_1296;
wire n_1413;
wire n_801;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_304;
wire n_1338;
wire n_577;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_1572;
wire n_1968;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_1661;
wire n_1212;
wire n_1541;
wire n_206;
wire n_217;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_1904;
wire n_774;
wire n_1628;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_527;
wire n_1168;
wire n_707;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_421;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_1803;
wire n_202;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_193;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_1117;
wire n_799;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_1782;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_676;
wire n_294;
wire n_318;
wire n_653;
wire n_642;
wire n_1602;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_664;
wire n_503;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_867;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_518;
wire n_505;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_826;
wire n_1813;
wire n_886;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_848;
wire n_1550;
wire n_1498;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_328;
wire n_1250;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_928;
wire n_608;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_402;
wire n_413;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_1502;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_203;
wire n_384;
wire n_1404;
wire n_1794;
wire n_1315;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_462;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_188;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_1321;
wire n_362;
wire n_1975;
wire n_273;
wire n_1937;
wire n_585;
wire n_1739;
wire n_270;
wire n_616;
wire n_1914;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_1325;
wire n_1595;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_403;
wire n_453;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_1621;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_651;
wire n_1340;
wire n_334;
wire n_811;
wire n_1558;
wire n_807;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_1254;
wire n_1026;
wire n_1969;
wire n_1234;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_1681;
wire n_1018;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;

INVx1_ASAP7_75t_L g188 ( 
.A(n_131),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_144),
.Y(n_189)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_154),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_150),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_14),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g194 ( 
.A(n_15),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_14),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_128),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_138),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_22),
.Y(n_198)
);

BUFx5_ASAP7_75t_L g199 ( 
.A(n_130),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_123),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_93),
.Y(n_201)
);

BUFx10_ASAP7_75t_L g202 ( 
.A(n_47),
.Y(n_202)
);

BUFx10_ASAP7_75t_L g203 ( 
.A(n_184),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_117),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_107),
.Y(n_205)
);

INVx1_ASAP7_75t_SL g206 ( 
.A(n_110),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g207 ( 
.A(n_139),
.Y(n_207)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_174),
.Y(n_208)
);

BUFx10_ASAP7_75t_L g209 ( 
.A(n_187),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_141),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_60),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_127),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_1),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_146),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_62),
.Y(n_215)
);

INVx2_ASAP7_75t_SL g216 ( 
.A(n_64),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_158),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_68),
.Y(n_218)
);

BUFx10_ASAP7_75t_L g219 ( 
.A(n_96),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_3),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_133),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_54),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_160),
.Y(n_223)
);

INVxp67_ASAP7_75t_SL g224 ( 
.A(n_162),
.Y(n_224)
);

BUFx10_ASAP7_75t_L g225 ( 
.A(n_39),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_84),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_61),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g228 ( 
.A(n_132),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_113),
.Y(n_229)
);

BUFx10_ASAP7_75t_L g230 ( 
.A(n_73),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_163),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_80),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_148),
.Y(n_233)
);

INVx1_ASAP7_75t_SL g234 ( 
.A(n_8),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_104),
.Y(n_235)
);

BUFx6f_ASAP7_75t_L g236 ( 
.A(n_134),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_99),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_143),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_19),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_124),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_78),
.Y(n_241)
);

BUFx10_ASAP7_75t_L g242 ( 
.A(n_81),
.Y(n_242)
);

BUFx10_ASAP7_75t_L g243 ( 
.A(n_151),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_92),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_36),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_85),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_75),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_71),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_5),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_166),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g251 ( 
.A(n_19),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_126),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_33),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_168),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_53),
.Y(n_255)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_77),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_100),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_87),
.Y(n_258)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_103),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_161),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_79),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_94),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_121),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_46),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_147),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_18),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_66),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_24),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_178),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_136),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_53),
.Y(n_271)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_89),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_67),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_28),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_41),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_9),
.Y(n_276)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_55),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_25),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_185),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_91),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_135),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_86),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_24),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_29),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_153),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_165),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_13),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_83),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_155),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_27),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_18),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_38),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_172),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_137),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_34),
.Y(n_295)
);

BUFx10_ASAP7_75t_L g296 ( 
.A(n_98),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_55),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g298 ( 
.A(n_102),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_38),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_44),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_9),
.Y(n_301)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_32),
.Y(n_302)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_170),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_118),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_145),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_159),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_176),
.Y(n_307)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_13),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_116),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_2),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_182),
.Y(n_311)
);

BUFx10_ASAP7_75t_L g312 ( 
.A(n_171),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_164),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_74),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_76),
.Y(n_315)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_186),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_122),
.Y(n_317)
);

CKINVDCx16_ASAP7_75t_R g318 ( 
.A(n_48),
.Y(n_318)
);

CKINVDCx5p33_ASAP7_75t_R g319 ( 
.A(n_95),
.Y(n_319)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_69),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_149),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_51),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_31),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_57),
.Y(n_324)
);

BUFx10_ASAP7_75t_L g325 ( 
.A(n_34),
.Y(n_325)
);

CKINVDCx5p33_ASAP7_75t_R g326 ( 
.A(n_46),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_26),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_7),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_21),
.Y(n_329)
);

CKINVDCx5p33_ASAP7_75t_R g330 ( 
.A(n_112),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_48),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_179),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_30),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_15),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_44),
.Y(n_335)
);

BUFx6f_ASAP7_75t_L g336 ( 
.A(n_59),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_49),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_57),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_120),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_7),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_35),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_30),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_20),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_114),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_45),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_27),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_72),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_115),
.Y(n_348)
);

CKINVDCx5p33_ASAP7_75t_R g349 ( 
.A(n_8),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_88),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_0),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_142),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_1),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g354 ( 
.A(n_65),
.Y(n_354)
);

BUFx3_ASAP7_75t_L g355 ( 
.A(n_54),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_157),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_58),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_25),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_42),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_56),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_47),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_21),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_106),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_175),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_183),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_26),
.Y(n_366)
);

BUFx6f_ASAP7_75t_L g367 ( 
.A(n_0),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_61),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g369 ( 
.A(n_12),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g370 ( 
.A(n_5),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_111),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_33),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_181),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_90),
.Y(n_374)
);

BUFx10_ASAP7_75t_L g375 ( 
.A(n_2),
.Y(n_375)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_45),
.Y(n_376)
);

INVxp33_ASAP7_75t_L g377 ( 
.A(n_193),
.Y(n_377)
);

BUFx6f_ASAP7_75t_L g378 ( 
.A(n_236),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_196),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_336),
.Y(n_380)
);

CKINVDCx20_ASAP7_75t_R g381 ( 
.A(n_228),
.Y(n_381)
);

CKINVDCx5p33_ASAP7_75t_R g382 ( 
.A(n_200),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_228),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_336),
.Y(n_384)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_252),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_221),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_252),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_267),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_229),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_336),
.Y(n_390)
);

HB1xp67_ASAP7_75t_L g391 ( 
.A(n_251),
.Y(n_391)
);

INVx2_ASAP7_75t_L g392 ( 
.A(n_199),
.Y(n_392)
);

INVx2_ASAP7_75t_SL g393 ( 
.A(n_355),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_336),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_358),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_202),
.Y(n_397)
);

HB1xp67_ASAP7_75t_L g398 ( 
.A(n_308),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_358),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_358),
.Y(n_400)
);

INVxp67_ASAP7_75t_SL g401 ( 
.A(n_207),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_367),
.Y(n_402)
);

CKINVDCx16_ASAP7_75t_R g403 ( 
.A(n_318),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_267),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_367),
.Y(n_405)
);

BUFx2_ASAP7_75t_L g406 ( 
.A(n_355),
.Y(n_406)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_270),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_367),
.Y(n_408)
);

INVxp67_ASAP7_75t_L g409 ( 
.A(n_202),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_231),
.Y(n_410)
);

INVxp67_ASAP7_75t_L g411 ( 
.A(n_202),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_367),
.Y(n_412)
);

INVxp67_ASAP7_75t_SL g413 ( 
.A(n_208),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_376),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_233),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_376),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_235),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_376),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_211),
.Y(n_420)
);

INVxp33_ASAP7_75t_L g421 ( 
.A(n_213),
.Y(n_421)
);

INVxp33_ASAP7_75t_SL g422 ( 
.A(n_341),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_237),
.Y(n_423)
);

CKINVDCx5p33_ASAP7_75t_R g424 ( 
.A(n_238),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_211),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_255),
.Y(n_426)
);

BUFx3_ASAP7_75t_L g427 ( 
.A(n_272),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_255),
.Y(n_428)
);

INVxp67_ASAP7_75t_SL g429 ( 
.A(n_272),
.Y(n_429)
);

INVxp67_ASAP7_75t_SL g430 ( 
.A(n_314),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_270),
.Y(n_431)
);

HB1xp67_ASAP7_75t_L g432 ( 
.A(n_341),
.Y(n_432)
);

INVxp67_ASAP7_75t_L g433 ( 
.A(n_225),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_241),
.Y(n_434)
);

CKINVDCx20_ASAP7_75t_R g435 ( 
.A(n_279),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_266),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_277),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_290),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_291),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_314),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_327),
.Y(n_441)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_279),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_244),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_328),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_199),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_345),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_353),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_362),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_368),
.Y(n_449)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_199),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_372),
.Y(n_451)
);

HB1xp67_ASAP7_75t_L g452 ( 
.A(n_342),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_246),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_310),
.Y(n_454)
);

CKINVDCx5p33_ASAP7_75t_R g455 ( 
.A(n_248),
.Y(n_455)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_298),
.Y(n_456)
);

CKINVDCx20_ASAP7_75t_R g457 ( 
.A(n_298),
.Y(n_457)
);

CKINVDCx14_ASAP7_75t_R g458 ( 
.A(n_225),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_310),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_217),
.Y(n_460)
);

BUFx3_ASAP7_75t_L g461 ( 
.A(n_203),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_217),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_232),
.Y(n_463)
);

CKINVDCx20_ASAP7_75t_R g464 ( 
.A(n_316),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_232),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g466 ( 
.A(n_316),
.Y(n_466)
);

CKINVDCx5p33_ASAP7_75t_R g467 ( 
.A(n_250),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_286),
.Y(n_468)
);

CKINVDCx16_ASAP7_75t_R g469 ( 
.A(n_354),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_286),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_188),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_380),
.Y(n_472)
);

BUFx6f_ASAP7_75t_L g473 ( 
.A(n_378),
.Y(n_473)
);

INVx2_ASAP7_75t_L g474 ( 
.A(n_378),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_378),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_378),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_SL g477 ( 
.A1(n_381),
.A2(n_302),
.B1(n_340),
.B2(n_222),
.Y(n_477)
);

AND2x6_ASAP7_75t_L g478 ( 
.A(n_378),
.B(n_236),
.Y(n_478)
);

INVx3_ASAP7_75t_L g479 ( 
.A(n_392),
.Y(n_479)
);

INVx2_ASAP7_75t_L g480 ( 
.A(n_392),
.Y(n_480)
);

AND2x2_ASAP7_75t_L g481 ( 
.A(n_429),
.B(n_216),
.Y(n_481)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_430),
.B(n_216),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_384),
.Y(n_484)
);

NAND2xp33_ASAP7_75t_L g485 ( 
.A(n_471),
.B(n_236),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_445),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_L g488 ( 
.A(n_401),
.B(n_259),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_390),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_440),
.B(n_204),
.Y(n_490)
);

AND2x2_ASAP7_75t_L g491 ( 
.A(n_427),
.B(n_189),
.Y(n_491)
);

NOR2xp33_ASAP7_75t_R g492 ( 
.A(n_458),
.B(n_254),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_390),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_394),
.Y(n_494)
);

INVx2_ASAP7_75t_L g495 ( 
.A(n_445),
.Y(n_495)
);

NOR2x1_ASAP7_75t_L g496 ( 
.A(n_460),
.B(n_190),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_397),
.A2(n_334),
.B1(n_302),
.B2(n_340),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_450),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_395),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_391),
.Y(n_500)
);

AND2x6_ASAP7_75t_L g501 ( 
.A(n_450),
.B(n_236),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_460),
.Y(n_502)
);

AND2x2_ASAP7_75t_L g503 ( 
.A(n_427),
.B(n_191),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_379),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_395),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_414),
.B(n_204),
.Y(n_506)
);

HB1xp67_ASAP7_75t_L g507 ( 
.A(n_398),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_396),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_403),
.B(n_203),
.Y(n_509)
);

OAI22xp5_ASAP7_75t_L g510 ( 
.A1(n_409),
.A2(n_334),
.B1(n_300),
.B2(n_222),
.Y(n_510)
);

INVx3_ASAP7_75t_L g511 ( 
.A(n_396),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_399),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_399),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_400),
.Y(n_514)
);

AND2x2_ASAP7_75t_L g515 ( 
.A(n_471),
.B(n_192),
.Y(n_515)
);

OAI22xp5_ASAP7_75t_SL g516 ( 
.A1(n_383),
.A2(n_300),
.B1(n_387),
.B2(n_385),
.Y(n_516)
);

CKINVDCx11_ASAP7_75t_R g517 ( 
.A(n_388),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_400),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_416),
.B(n_210),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_417),
.B(n_210),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_393),
.B(n_197),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_402),
.Y(n_522)
);

INVx3_ASAP7_75t_L g523 ( 
.A(n_402),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_405),
.Y(n_524)
);

INVx2_ASAP7_75t_L g525 ( 
.A(n_405),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_R g526 ( 
.A(n_382),
.B(n_260),
.Y(n_526)
);

INVx2_ASAP7_75t_SL g527 ( 
.A(n_393),
.Y(n_527)
);

CKINVDCx5p33_ASAP7_75t_R g528 ( 
.A(n_386),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_432),
.Y(n_529)
);

BUFx2_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_408),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_408),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_412),
.Y(n_533)
);

BUFx3_ASAP7_75t_L g534 ( 
.A(n_412),
.Y(n_534)
);

AND2x2_ASAP7_75t_L g535 ( 
.A(n_406),
.B(n_201),
.Y(n_535)
);

INVx1_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

INVx6_ASAP7_75t_L g537 ( 
.A(n_461),
.Y(n_537)
);

AND2x4_ASAP7_75t_L g538 ( 
.A(n_462),
.B(n_205),
.Y(n_538)
);

INVx2_ASAP7_75t_L g539 ( 
.A(n_419),
.Y(n_539)
);

AND2x4_ASAP7_75t_L g540 ( 
.A(n_462),
.B(n_212),
.Y(n_540)
);

OAI21x1_ASAP7_75t_L g541 ( 
.A1(n_463),
.A2(n_218),
.B(n_215),
.Y(n_541)
);

INVx2_ASAP7_75t_L g542 ( 
.A(n_463),
.Y(n_542)
);

BUFx8_ASAP7_75t_L g543 ( 
.A(n_461),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_389),
.Y(n_544)
);

NAND2xp5_ASAP7_75t_SL g545 ( 
.A(n_410),
.B(n_203),
.Y(n_545)
);

AND2x2_ASAP7_75t_L g546 ( 
.A(n_465),
.B(n_223),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_465),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_470),
.Y(n_548)
);

INVx1_ASAP7_75t_L g549 ( 
.A(n_470),
.Y(n_549)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_481),
.B(n_415),
.Y(n_550)
);

AOI22xp33_ASAP7_75t_L g551 ( 
.A1(n_481),
.A2(n_413),
.B1(n_422),
.B2(n_452),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_534),
.Y(n_552)
);

INVx2_ASAP7_75t_L g553 ( 
.A(n_480),
.Y(n_553)
);

INVx2_ASAP7_75t_L g554 ( 
.A(n_480),
.Y(n_554)
);

INVx2_ASAP7_75t_L g555 ( 
.A(n_480),
.Y(n_555)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_534),
.Y(n_556)
);

OAI22xp5_ASAP7_75t_L g557 ( 
.A1(n_488),
.A2(n_423),
.B1(n_424),
.B2(n_418),
.Y(n_557)
);

INVx2_ASAP7_75t_SL g558 ( 
.A(n_530),
.Y(n_558)
);

CKINVDCx20_ASAP7_75t_R g559 ( 
.A(n_517),
.Y(n_559)
);

INVx1_ASAP7_75t_L g560 ( 
.A(n_534),
.Y(n_560)
);

INVx2_ASAP7_75t_L g561 ( 
.A(n_480),
.Y(n_561)
);

CKINVDCx5p33_ASAP7_75t_R g562 ( 
.A(n_492),
.Y(n_562)
);

AOI22xp33_ASAP7_75t_L g563 ( 
.A1(n_481),
.A2(n_468),
.B1(n_451),
.B2(n_421),
.Y(n_563)
);

CKINVDCx5p33_ASAP7_75t_R g564 ( 
.A(n_492),
.Y(n_564)
);

NOR2x1p5_ASAP7_75t_L g565 ( 
.A(n_504),
.B(n_342),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_L g566 ( 
.A(n_483),
.B(n_434),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_R g567 ( 
.A(n_528),
.B(n_443),
.Y(n_567)
);

AOI22xp33_ASAP7_75t_L g568 ( 
.A1(n_483),
.A2(n_468),
.B1(n_377),
.B2(n_437),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_487),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_530),
.Y(n_570)
);

INVx1_ASAP7_75t_L g571 ( 
.A(n_487),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_487),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_487),
.Y(n_573)
);

AND2x4_ASAP7_75t_L g574 ( 
.A(n_546),
.B(n_224),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_495),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_526),
.B(n_453),
.Y(n_576)
);

INVx1_ASAP7_75t_L g577 ( 
.A(n_495),
.Y(n_577)
);

INVx2_ASAP7_75t_L g578 ( 
.A(n_495),
.Y(n_578)
);

NAND2xp33_ASAP7_75t_SL g579 ( 
.A(n_509),
.B(n_354),
.Y(n_579)
);

INVx2_ASAP7_75t_L g580 ( 
.A(n_495),
.Y(n_580)
);

BUFx6f_ASAP7_75t_L g581 ( 
.A(n_473),
.Y(n_581)
);

INVx1_ASAP7_75t_L g582 ( 
.A(n_479),
.Y(n_582)
);

INVx2_ASAP7_75t_SL g583 ( 
.A(n_530),
.Y(n_583)
);

INVx2_ASAP7_75t_L g584 ( 
.A(n_518),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_518),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_479),
.Y(n_586)
);

INVx2_ASAP7_75t_L g587 ( 
.A(n_518),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g588 ( 
.A1(n_488),
.A2(n_234),
.B1(n_369),
.B2(n_194),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_518),
.Y(n_589)
);

INVx2_ASAP7_75t_L g590 ( 
.A(n_524),
.Y(n_590)
);

INVx2_ASAP7_75t_L g591 ( 
.A(n_524),
.Y(n_591)
);

INVx2_ASAP7_75t_L g592 ( 
.A(n_524),
.Y(n_592)
);

INVx1_ASAP7_75t_L g593 ( 
.A(n_479),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_524),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_490),
.B(n_455),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_525),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_473),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_483),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_525),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_490),
.B(n_467),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_479),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_525),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_525),
.Y(n_603)
);

INVx2_ASAP7_75t_L g604 ( 
.A(n_532),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_479),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_532),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g607 ( 
.A(n_545),
.B(n_411),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_491),
.B(n_206),
.Y(n_608)
);

INVx2_ASAP7_75t_L g609 ( 
.A(n_532),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_515),
.B(n_546),
.C(n_521),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_498),
.Y(n_611)
);

AOI22xp5_ASAP7_75t_L g612 ( 
.A1(n_535),
.A2(n_343),
.B1(n_346),
.B2(n_349),
.Y(n_612)
);

NAND3xp33_ASAP7_75t_L g613 ( 
.A(n_515),
.B(n_437),
.C(n_436),
.Y(n_613)
);

AOI22xp33_ASAP7_75t_L g614 ( 
.A1(n_535),
.A2(n_436),
.B1(n_438),
.B2(n_439),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_SL g615 ( 
.A(n_544),
.B(n_442),
.Y(n_615)
);

AOI22xp5_ASAP7_75t_L g616 ( 
.A1(n_535),
.A2(n_343),
.B1(n_346),
.B2(n_349),
.Y(n_616)
);

OAI22xp33_ASAP7_75t_L g617 ( 
.A1(n_545),
.A2(n_301),
.B1(n_271),
.B2(n_268),
.Y(n_617)
);

AOI22xp5_ASAP7_75t_L g618 ( 
.A1(n_529),
.A2(n_351),
.B1(n_220),
.B2(n_326),
.Y(n_618)
);

AND2x2_ASAP7_75t_SL g619 ( 
.A(n_485),
.B(n_226),
.Y(n_619)
);

NOR2xp67_ASAP7_75t_L g620 ( 
.A(n_498),
.B(n_261),
.Y(n_620)
);

INVx2_ASAP7_75t_L g621 ( 
.A(n_532),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_498),
.Y(n_622)
);

AND2x4_ASAP7_75t_L g623 ( 
.A(n_546),
.B(n_240),
.Y(n_623)
);

INVx3_ASAP7_75t_L g624 ( 
.A(n_473),
.Y(n_624)
);

INVx1_ASAP7_75t_L g625 ( 
.A(n_498),
.Y(n_625)
);

INVx5_ASAP7_75t_L g626 ( 
.A(n_501),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_537),
.B(n_247),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_498),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_533),
.Y(n_629)
);

INVx5_ASAP7_75t_L g630 ( 
.A(n_501),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_533),
.Y(n_631)
);

BUFx3_ASAP7_75t_L g632 ( 
.A(n_537),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_526),
.B(n_469),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_472),
.Y(n_634)
);

BUFx6f_ASAP7_75t_L g635 ( 
.A(n_473),
.Y(n_635)
);

INVx2_ASAP7_75t_L g636 ( 
.A(n_533),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_SL g637 ( 
.A(n_543),
.B(n_509),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_473),
.Y(n_638)
);

BUFx3_ASAP7_75t_L g639 ( 
.A(n_537),
.Y(n_639)
);

NOR2xp33_ASAP7_75t_L g640 ( 
.A(n_537),
.B(n_433),
.Y(n_640)
);

CKINVDCx5p33_ASAP7_75t_R g641 ( 
.A(n_517),
.Y(n_641)
);

BUFx3_ASAP7_75t_L g642 ( 
.A(n_537),
.Y(n_642)
);

BUFx3_ASAP7_75t_L g643 ( 
.A(n_537),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_533),
.Y(n_644)
);

NAND2xp5_ASAP7_75t_L g645 ( 
.A(n_491),
.B(n_320),
.Y(n_645)
);

INVx2_ASAP7_75t_L g646 ( 
.A(n_539),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_472),
.Y(n_647)
);

INVx1_ASAP7_75t_L g648 ( 
.A(n_482),
.Y(n_648)
);

OR2x2_ASAP7_75t_L g649 ( 
.A(n_500),
.B(n_454),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_543),
.B(n_527),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_SL g651 ( 
.A(n_543),
.B(n_209),
.Y(n_651)
);

AND2x2_ASAP7_75t_L g652 ( 
.A(n_521),
.B(n_420),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_539),
.Y(n_653)
);

AND2x2_ASAP7_75t_L g654 ( 
.A(n_521),
.B(n_420),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_482),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_484),
.Y(n_656)
);

BUFx10_ASAP7_75t_L g657 ( 
.A(n_529),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_539),
.Y(n_658)
);

INVx3_ASAP7_75t_L g659 ( 
.A(n_473),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_539),
.Y(n_660)
);

BUFx3_ASAP7_75t_L g661 ( 
.A(n_538),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_491),
.B(n_262),
.Y(n_662)
);

BUFx6f_ASAP7_75t_L g663 ( 
.A(n_473),
.Y(n_663)
);

INVx2_ASAP7_75t_L g664 ( 
.A(n_542),
.Y(n_664)
);

INVx8_ASAP7_75t_L g665 ( 
.A(n_501),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_543),
.B(n_209),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_SL g667 ( 
.A(n_543),
.B(n_209),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_542),
.Y(n_668)
);

INVx6_ASAP7_75t_L g669 ( 
.A(n_538),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_484),
.Y(n_670)
);

INVx1_ASAP7_75t_L g671 ( 
.A(n_486),
.Y(n_671)
);

INVx3_ASAP7_75t_L g672 ( 
.A(n_473),
.Y(n_672)
);

BUFx8_ASAP7_75t_SL g673 ( 
.A(n_477),
.Y(n_673)
);

OR2x2_ASAP7_75t_L g674 ( 
.A(n_500),
.B(n_454),
.Y(n_674)
);

INVx2_ASAP7_75t_L g675 ( 
.A(n_542),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_486),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_474),
.Y(n_677)
);

OAI22xp33_ASAP7_75t_L g678 ( 
.A1(n_506),
.A2(n_292),
.B1(n_287),
.B2(n_284),
.Y(n_678)
);

BUFx6f_ASAP7_75t_L g679 ( 
.A(n_474),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_542),
.Y(n_680)
);

INVx1_ASAP7_75t_SL g681 ( 
.A(n_516),
.Y(n_681)
);

INVx2_ASAP7_75t_SL g682 ( 
.A(n_503),
.Y(n_682)
);

INVx3_ASAP7_75t_L g683 ( 
.A(n_474),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_508),
.Y(n_684)
);

BUFx6f_ASAP7_75t_L g685 ( 
.A(n_474),
.Y(n_685)
);

AND2x2_ASAP7_75t_L g686 ( 
.A(n_503),
.B(n_425),
.Y(n_686)
);

CKINVDCx5p33_ASAP7_75t_R g687 ( 
.A(n_516),
.Y(n_687)
);

OR2x2_ASAP7_75t_L g688 ( 
.A(n_507),
.B(n_459),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_489),
.Y(n_689)
);

AOI22xp5_ASAP7_75t_L g690 ( 
.A1(n_497),
.A2(n_351),
.B1(n_274),
.B2(n_331),
.Y(n_690)
);

NAND2xp5_ASAP7_75t_L g691 ( 
.A(n_503),
.B(n_527),
.Y(n_691)
);

INVx1_ASAP7_75t_L g692 ( 
.A(n_489),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_508),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_493),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_493),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_SL g696 ( 
.A(n_527),
.B(n_219),
.Y(n_696)
);

NAND2xp5_ASAP7_75t_L g697 ( 
.A(n_515),
.B(n_265),
.Y(n_697)
);

INVx3_ASAP7_75t_L g698 ( 
.A(n_475),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_506),
.B(n_219),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_475),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_508),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_552),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_L g703 ( 
.A(n_595),
.B(n_538),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_686),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_556),
.Y(n_705)
);

INVx2_ASAP7_75t_SL g706 ( 
.A(n_649),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_556),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_598),
.B(n_519),
.Y(n_708)
);

AOI22xp5_ASAP7_75t_L g709 ( 
.A1(n_607),
.A2(n_519),
.B1(n_520),
.B2(n_538),
.Y(n_709)
);

OAI221xp5_ASAP7_75t_L g710 ( 
.A1(n_588),
.A2(n_370),
.B1(n_520),
.B2(n_363),
.C(n_303),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_598),
.B(n_538),
.Y(n_711)
);

INVx1_ASAP7_75t_SL g712 ( 
.A(n_657),
.Y(n_712)
);

AND2x6_ASAP7_75t_L g713 ( 
.A(n_661),
.B(n_600),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_L g714 ( 
.A(n_574),
.B(n_540),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_558),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_574),
.B(n_540),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_550),
.B(n_507),
.Y(n_717)
);

A2O1A1Ixp33_ASAP7_75t_L g718 ( 
.A1(n_610),
.A2(n_541),
.B(n_540),
.C(n_496),
.Y(n_718)
);

OAI22xp5_ASAP7_75t_L g719 ( 
.A1(n_610),
.A2(n_304),
.B1(n_309),
.B2(n_256),
.Y(n_719)
);

NOR2xp33_ASAP7_75t_L g720 ( 
.A(n_566),
.B(n_214),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_574),
.B(n_540),
.Y(n_721)
);

AOI22xp33_ASAP7_75t_L g722 ( 
.A1(n_574),
.A2(n_540),
.B1(n_541),
.B2(n_258),
.Y(n_722)
);

AND2x4_ASAP7_75t_L g723 ( 
.A(n_682),
.B(n_438),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_558),
.B(n_497),
.Y(n_724)
);

NAND2xp5_ASAP7_75t_L g725 ( 
.A(n_682),
.B(n_496),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_560),
.Y(n_726)
);

NOR2xp33_ASAP7_75t_L g727 ( 
.A(n_557),
.B(n_214),
.Y(n_727)
);

AOI22xp5_ASAP7_75t_L g728 ( 
.A1(n_579),
.A2(n_435),
.B1(n_431),
.B2(n_456),
.Y(n_728)
);

BUFx3_ASAP7_75t_L g729 ( 
.A(n_686),
.Y(n_729)
);

INVx3_ASAP7_75t_R g730 ( 
.A(n_649),
.Y(n_730)
);

INVx2_ASAP7_75t_SL g731 ( 
.A(n_674),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_SL g732 ( 
.A(n_640),
.B(n_344),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_560),
.Y(n_733)
);

INVx1_ASAP7_75t_L g734 ( 
.A(n_634),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_691),
.B(n_508),
.Y(n_735)
);

INVx2_ASAP7_75t_L g736 ( 
.A(n_553),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_634),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_562),
.B(n_344),
.Y(n_738)
);

INVx2_ASAP7_75t_L g739 ( 
.A(n_553),
.Y(n_739)
);

AOI22xp5_ASAP7_75t_L g740 ( 
.A1(n_669),
.A2(n_404),
.B1(n_407),
.B2(n_457),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_608),
.B(n_347),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_697),
.B(n_623),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_623),
.B(n_511),
.Y(n_743)
);

INVx2_ASAP7_75t_L g744 ( 
.A(n_554),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_619),
.A2(n_541),
.B1(n_311),
.B2(n_313),
.Y(n_745)
);

INVx3_ASAP7_75t_L g746 ( 
.A(n_661),
.Y(n_746)
);

NOR2xp33_ASAP7_75t_L g747 ( 
.A(n_645),
.B(n_347),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_623),
.B(n_511),
.Y(n_748)
);

BUFx3_ASAP7_75t_L g749 ( 
.A(n_559),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_SL g750 ( 
.A(n_661),
.B(n_199),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_647),
.B(n_511),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_647),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_648),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_554),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_L g755 ( 
.A(n_648),
.B(n_511),
.Y(n_755)
);

INVx1_ASAP7_75t_L g756 ( 
.A(n_655),
.Y(n_756)
);

OAI22xp5_ASAP7_75t_L g757 ( 
.A1(n_669),
.A2(n_257),
.B1(n_315),
.B2(n_317),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_555),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_655),
.B(n_523),
.Y(n_759)
);

BUFx3_ASAP7_75t_L g760 ( 
.A(n_652),
.Y(n_760)
);

OAI221xp5_ASAP7_75t_L g761 ( 
.A1(n_588),
.A2(n_285),
.B1(n_263),
.B2(n_269),
.C(n_371),
.Y(n_761)
);

OAI22xp5_ASAP7_75t_SL g762 ( 
.A1(n_687),
.A2(n_464),
.B1(n_466),
.B2(n_510),
.Y(n_762)
);

INVx2_ASAP7_75t_SL g763 ( 
.A(n_674),
.Y(n_763)
);

NOR2xp33_ASAP7_75t_L g764 ( 
.A(n_570),
.B(n_348),
.Y(n_764)
);

BUFx6f_ASAP7_75t_L g765 ( 
.A(n_632),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_656),
.Y(n_766)
);

AOI22xp5_ASAP7_75t_L g767 ( 
.A1(n_669),
.A2(n_650),
.B1(n_637),
.B2(n_662),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_570),
.B(n_348),
.Y(n_768)
);

BUFx3_ASAP7_75t_L g769 ( 
.A(n_652),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_583),
.B(n_510),
.Y(n_770)
);

OAI22xp5_ASAP7_75t_L g771 ( 
.A1(n_669),
.A2(n_273),
.B1(n_332),
.B2(n_339),
.Y(n_771)
);

INVxp67_ASAP7_75t_L g772 ( 
.A(n_583),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_656),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_670),
.B(n_523),
.Y(n_774)
);

NOR2xp33_ASAP7_75t_L g775 ( 
.A(n_688),
.B(n_350),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_670),
.B(n_523),
.Y(n_776)
);

AOI22xp5_ASAP7_75t_L g777 ( 
.A1(n_699),
.A2(n_282),
.B1(n_280),
.B2(n_374),
.Y(n_777)
);

AOI22xp5_ASAP7_75t_L g778 ( 
.A1(n_565),
.A2(n_281),
.B1(n_289),
.B2(n_373),
.Y(n_778)
);

BUFx3_ASAP7_75t_L g779 ( 
.A(n_654),
.Y(n_779)
);

AOI22xp5_ASAP7_75t_L g780 ( 
.A1(n_565),
.A2(n_307),
.B1(n_364),
.B2(n_352),
.Y(n_780)
);

BUFx6f_ASAP7_75t_L g781 ( 
.A(n_632),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_688),
.B(n_195),
.Y(n_782)
);

INVx2_ASAP7_75t_L g783 ( 
.A(n_555),
.Y(n_783)
);

AOI221xp5_ASAP7_75t_L g784 ( 
.A1(n_617),
.A2(n_690),
.B1(n_612),
.B2(n_616),
.C(n_681),
.Y(n_784)
);

BUFx3_ASAP7_75t_L g785 ( 
.A(n_654),
.Y(n_785)
);

INVx2_ASAP7_75t_L g786 ( 
.A(n_561),
.Y(n_786)
);

NOR2xp33_ASAP7_75t_L g787 ( 
.A(n_678),
.B(n_198),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_619),
.B(n_199),
.Y(n_788)
);

NAND2xp5_ASAP7_75t_SL g789 ( 
.A(n_564),
.B(n_288),
.Y(n_789)
);

INVxp67_ASAP7_75t_L g790 ( 
.A(n_613),
.Y(n_790)
);

BUFx2_ASAP7_75t_L g791 ( 
.A(n_567),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_613),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_SL g793 ( 
.A(n_651),
.B(n_227),
.Y(n_793)
);

INVxp67_ASAP7_75t_L g794 ( 
.A(n_657),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_612),
.B(n_239),
.Y(n_795)
);

INVxp67_ASAP7_75t_L g796 ( 
.A(n_657),
.Y(n_796)
);

NAND2xp5_ASAP7_75t_L g797 ( 
.A(n_671),
.B(n_523),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_564),
.B(n_219),
.Y(n_798)
);

NAND2xp33_ASAP7_75t_L g799 ( 
.A(n_665),
.B(n_199),
.Y(n_799)
);

BUFx12f_ASAP7_75t_SL g800 ( 
.A(n_641),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_671),
.B(n_494),
.Y(n_801)
);

AO22x2_ASAP7_75t_L g802 ( 
.A1(n_666),
.A2(n_477),
.B1(n_356),
.B2(n_365),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_676),
.B(n_494),
.Y(n_803)
);

NAND3xp33_ASAP7_75t_L g804 ( 
.A(n_551),
.B(n_616),
.C(n_618),
.Y(n_804)
);

NAND2xp5_ASAP7_75t_SL g805 ( 
.A(n_568),
.B(n_293),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_689),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_561),
.Y(n_807)
);

NOR2xp67_ASAP7_75t_L g808 ( 
.A(n_576),
.B(n_547),
.Y(n_808)
);

INVx2_ASAP7_75t_SL g809 ( 
.A(n_657),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_SL g810 ( 
.A(n_563),
.B(n_294),
.Y(n_810)
);

NOR2xp67_ASAP7_75t_L g811 ( 
.A(n_667),
.B(n_547),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_692),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_569),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_614),
.B(n_459),
.Y(n_814)
);

OAI21xp33_ASAP7_75t_L g815 ( 
.A1(n_690),
.A2(n_439),
.B(n_441),
.Y(n_815)
);

AOI22xp33_ASAP7_75t_L g816 ( 
.A1(n_619),
.A2(n_321),
.B1(n_199),
.B2(n_549),
.Y(n_816)
);

BUFx6f_ASAP7_75t_SL g817 ( 
.A(n_673),
.Y(n_817)
);

NOR2xp33_ASAP7_75t_L g818 ( 
.A(n_692),
.B(n_694),
.Y(n_818)
);

INVx3_ASAP7_75t_L g819 ( 
.A(n_679),
.Y(n_819)
);

NAND2xp5_ASAP7_75t_L g820 ( 
.A(n_694),
.B(n_695),
.Y(n_820)
);

AOI22xp5_ASAP7_75t_L g821 ( 
.A1(n_620),
.A2(n_330),
.B1(n_319),
.B2(n_306),
.Y(n_821)
);

NOR2xp33_ASAP7_75t_R g822 ( 
.A(n_641),
.B(n_615),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_620),
.B(n_499),
.Y(n_823)
);

NAND2xp33_ASAP7_75t_L g824 ( 
.A(n_665),
.B(n_305),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_684),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_L g826 ( 
.A(n_582),
.B(n_505),
.Y(n_826)
);

NOR2xp33_ASAP7_75t_L g827 ( 
.A(n_696),
.B(n_245),
.Y(n_827)
);

INVx3_ASAP7_75t_L g828 ( 
.A(n_679),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_586),
.B(n_512),
.Y(n_829)
);

INVx1_ASAP7_75t_L g830 ( 
.A(n_684),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_586),
.B(n_512),
.Y(n_831)
);

NAND2xp5_ASAP7_75t_L g832 ( 
.A(n_593),
.B(n_513),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_693),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_593),
.B(n_513),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_601),
.B(n_514),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_SL g836 ( 
.A(n_626),
.B(n_502),
.Y(n_836)
);

NOR2xp67_ASAP7_75t_L g837 ( 
.A(n_633),
.B(n_548),
.Y(n_837)
);

INVxp67_ASAP7_75t_SL g838 ( 
.A(n_569),
.Y(n_838)
);

NAND2xp33_ASAP7_75t_L g839 ( 
.A(n_665),
.B(n_478),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_SL g840 ( 
.A(n_626),
.B(n_502),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_SL g841 ( 
.A(n_618),
.B(n_230),
.Y(n_841)
);

AND2x2_ASAP7_75t_L g842 ( 
.A(n_687),
.B(n_225),
.Y(n_842)
);

INVxp67_ASAP7_75t_L g843 ( 
.A(n_693),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_701),
.Y(n_844)
);

AND2x4_ASAP7_75t_L g845 ( 
.A(n_642),
.B(n_441),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_626),
.B(n_230),
.Y(n_846)
);

BUFx6f_ASAP7_75t_L g847 ( 
.A(n_642),
.Y(n_847)
);

INVx2_ASAP7_75t_L g848 ( 
.A(n_578),
.Y(n_848)
);

AND2x4_ASAP7_75t_L g849 ( 
.A(n_639),
.B(n_444),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_701),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_601),
.Y(n_851)
);

INVx4_ASAP7_75t_L g852 ( 
.A(n_665),
.Y(n_852)
);

INVx1_ASAP7_75t_L g853 ( 
.A(n_605),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_605),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_639),
.A2(n_476),
.B(n_475),
.Y(n_855)
);

INVx2_ASAP7_75t_L g856 ( 
.A(n_578),
.Y(n_856)
);

AOI22xp5_ASAP7_75t_L g857 ( 
.A1(n_627),
.A2(n_501),
.B1(n_548),
.B2(n_549),
.Y(n_857)
);

OAI22xp33_ASAP7_75t_L g858 ( 
.A1(n_627),
.A2(n_361),
.B1(n_360),
.B2(n_359),
.Y(n_858)
);

INVx1_ASAP7_75t_L g859 ( 
.A(n_611),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_626),
.B(n_502),
.Y(n_860)
);

NAND3xp33_ASAP7_75t_L g861 ( 
.A(n_627),
.B(n_335),
.C(n_249),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_L g862 ( 
.A(n_611),
.B(n_514),
.Y(n_862)
);

INVx2_ASAP7_75t_SL g863 ( 
.A(n_677),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_622),
.B(n_522),
.Y(n_864)
);

BUFx4f_ASAP7_75t_L g865 ( 
.A(n_791),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_818),
.B(n_622),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_703),
.A2(n_639),
.B1(n_643),
.B2(n_627),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_702),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_765),
.Y(n_869)
);

AND2x6_ASAP7_75t_L g870 ( 
.A(n_767),
.B(n_742),
.Y(n_870)
);

INVx2_ASAP7_75t_L g871 ( 
.A(n_705),
.Y(n_871)
);

AOI22xp33_ASAP7_75t_SL g872 ( 
.A1(n_804),
.A2(n_325),
.B1(n_375),
.B2(n_243),
.Y(n_872)
);

OR2x6_ASAP7_75t_L g873 ( 
.A(n_809),
.B(n_665),
.Y(n_873)
);

AND2x4_ASAP7_75t_L g874 ( 
.A(n_704),
.B(n_643),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_818),
.B(n_741),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_707),
.Y(n_876)
);

O2A1O1Ixp33_ASAP7_75t_L g877 ( 
.A1(n_790),
.A2(n_485),
.B(n_628),
.C(n_625),
.Y(n_877)
);

INVx2_ASAP7_75t_L g878 ( 
.A(n_825),
.Y(n_878)
);

INVx3_ASAP7_75t_L g879 ( 
.A(n_746),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_741),
.B(n_643),
.Y(n_880)
);

INVx3_ASAP7_75t_L g881 ( 
.A(n_746),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_726),
.Y(n_882)
);

AND2x2_ASAP7_75t_L g883 ( 
.A(n_760),
.B(n_769),
.Y(n_883)
);

INVxp67_ASAP7_75t_L g884 ( 
.A(n_706),
.Y(n_884)
);

INVx5_ASAP7_75t_L g885 ( 
.A(n_713),
.Y(n_885)
);

OR2x2_ASAP7_75t_L g886 ( 
.A(n_731),
.B(n_444),
.Y(n_886)
);

INVx3_ASAP7_75t_L g887 ( 
.A(n_765),
.Y(n_887)
);

OR2x6_ASAP7_75t_L g888 ( 
.A(n_715),
.B(n_627),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_733),
.Y(n_889)
);

NAND2xp5_ASAP7_75t_SL g890 ( 
.A(n_709),
.B(n_626),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_830),
.Y(n_891)
);

INVx2_ASAP7_75t_L g892 ( 
.A(n_833),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_747),
.B(n_597),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_714),
.B(n_630),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_L g895 ( 
.A(n_747),
.B(n_720),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_844),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_851),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_SL g898 ( 
.A(n_716),
.B(n_630),
.Y(n_898)
);

BUFx6f_ASAP7_75t_L g899 ( 
.A(n_765),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_779),
.Y(n_900)
);

CKINVDCx20_ASAP7_75t_R g901 ( 
.A(n_800),
.Y(n_901)
);

INVx2_ASAP7_75t_L g902 ( 
.A(n_850),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_720),
.B(n_597),
.Y(n_903)
);

AOI22xp5_ASAP7_75t_L g904 ( 
.A1(n_708),
.A2(n_624),
.B1(n_659),
.B2(n_597),
.Y(n_904)
);

AND2x2_ASAP7_75t_L g905 ( 
.A(n_785),
.B(n_325),
.Y(n_905)
);

NAND2xp5_ASAP7_75t_L g906 ( 
.A(n_734),
.B(n_624),
.Y(n_906)
);

INVx5_ASAP7_75t_L g907 ( 
.A(n_713),
.Y(n_907)
);

INVx3_ASAP7_75t_L g908 ( 
.A(n_781),
.Y(n_908)
);

AND2x2_ASAP7_75t_L g909 ( 
.A(n_715),
.B(n_325),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_737),
.B(n_624),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_853),
.Y(n_911)
);

INVx3_ASAP7_75t_L g912 ( 
.A(n_781),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_854),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_752),
.B(n_638),
.Y(n_914)
);

HB1xp67_ASAP7_75t_L g915 ( 
.A(n_772),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_753),
.Y(n_916)
);

NAND3xp33_ASAP7_75t_SL g917 ( 
.A(n_784),
.B(n_264),
.C(n_253),
.Y(n_917)
);

BUFx3_ASAP7_75t_L g918 ( 
.A(n_729),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_859),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_722),
.B(n_630),
.Y(n_920)
);

BUFx2_ASAP7_75t_L g921 ( 
.A(n_772),
.Y(n_921)
);

NOR2xp33_ASAP7_75t_L g922 ( 
.A(n_763),
.B(n_638),
.Y(n_922)
);

AOI22xp33_ASAP7_75t_SL g923 ( 
.A1(n_795),
.A2(n_375),
.B1(n_242),
.B2(n_243),
.Y(n_923)
);

INVx4_ASAP7_75t_L g924 ( 
.A(n_781),
.Y(n_924)
);

INVx2_ASAP7_75t_SL g925 ( 
.A(n_723),
.Y(n_925)
);

INVx2_ASAP7_75t_L g926 ( 
.A(n_736),
.Y(n_926)
);

AND2x4_ASAP7_75t_L g927 ( 
.A(n_723),
.B(n_446),
.Y(n_927)
);

INVx1_ASAP7_75t_L g928 ( 
.A(n_756),
.Y(n_928)
);

INVx2_ASAP7_75t_L g929 ( 
.A(n_739),
.Y(n_929)
);

NAND2xp5_ASAP7_75t_L g930 ( 
.A(n_766),
.B(n_773),
.Y(n_930)
);

AND3x1_ASAP7_75t_L g931 ( 
.A(n_795),
.B(n_447),
.C(n_446),
.Y(n_931)
);

OR2x6_ASAP7_75t_L g932 ( 
.A(n_762),
.B(n_447),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_806),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_745),
.A2(n_638),
.B1(n_659),
.B2(n_672),
.Y(n_934)
);

INVx1_ASAP7_75t_L g935 ( 
.A(n_812),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_790),
.B(n_792),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_843),
.Y(n_937)
);

NAND2x1p5_ASAP7_75t_L g938 ( 
.A(n_852),
.B(n_630),
.Y(n_938)
);

OR2x2_ASAP7_75t_L g939 ( 
.A(n_724),
.B(n_448),
.Y(n_939)
);

INVx3_ASAP7_75t_L g940 ( 
.A(n_781),
.Y(n_940)
);

AND2x4_ASAP7_75t_L g941 ( 
.A(n_837),
.B(n_448),
.Y(n_941)
);

AND2x4_ASAP7_75t_SL g942 ( 
.A(n_770),
.B(n_230),
.Y(n_942)
);

NAND2xp5_ASAP7_75t_L g943 ( 
.A(n_792),
.B(n_659),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_719),
.A2(n_788),
.B(n_710),
.C(n_761),
.Y(n_944)
);

NAND2xp5_ASAP7_75t_L g945 ( 
.A(n_725),
.B(n_672),
.Y(n_945)
);

NOR2x1_ASAP7_75t_R g946 ( 
.A(n_749),
.B(n_275),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_820),
.B(n_672),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_788),
.A2(n_577),
.B(n_575),
.C(n_573),
.Y(n_948)
);

BUFx3_ASAP7_75t_L g949 ( 
.A(n_845),
.Y(n_949)
);

AOI22xp33_ASAP7_75t_L g950 ( 
.A1(n_816),
.A2(n_745),
.B1(n_787),
.B2(n_727),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_843),
.Y(n_951)
);

BUFx5_ASAP7_75t_L g952 ( 
.A(n_713),
.Y(n_952)
);

OR2x2_ASAP7_75t_L g953 ( 
.A(n_842),
.B(n_449),
.Y(n_953)
);

AND3x1_ASAP7_75t_SL g954 ( 
.A(n_730),
.B(n_449),
.C(n_425),
.Y(n_954)
);

INVx2_ASAP7_75t_L g955 ( 
.A(n_744),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_711),
.B(n_571),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_775),
.B(n_572),
.Y(n_957)
);

NOR2xp33_ASAP7_75t_L g958 ( 
.A(n_717),
.B(n_775),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_L g959 ( 
.A(n_782),
.B(n_573),
.Y(n_959)
);

INVx2_ASAP7_75t_L g960 ( 
.A(n_754),
.Y(n_960)
);

NAND3xp33_ASAP7_75t_SL g961 ( 
.A(n_727),
.B(n_787),
.C(n_798),
.Y(n_961)
);

AOI22xp5_ASAP7_75t_L g962 ( 
.A1(n_721),
.A2(n_713),
.B1(n_750),
.B2(n_808),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_758),
.Y(n_963)
);

INVx1_ASAP7_75t_L g964 ( 
.A(n_849),
.Y(n_964)
);

NAND2xp5_ASAP7_75t_L g965 ( 
.A(n_735),
.B(n_577),
.Y(n_965)
);

INVx1_ASAP7_75t_L g966 ( 
.A(n_801),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_721),
.A2(n_635),
.B(n_581),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_803),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_783),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_847),
.Y(n_970)
);

AOI22xp5_ASAP7_75t_L g971 ( 
.A1(n_713),
.A2(n_677),
.B1(n_698),
.B2(n_683),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_822),
.Y(n_972)
);

HB1xp67_ASAP7_75t_L g973 ( 
.A(n_743),
.Y(n_973)
);

AND2x2_ASAP7_75t_L g974 ( 
.A(n_764),
.B(n_375),
.Y(n_974)
);

INVxp67_ASAP7_75t_L g975 ( 
.A(n_764),
.Y(n_975)
);

INVx2_ASAP7_75t_L g976 ( 
.A(n_786),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_SL g977 ( 
.A(n_722),
.B(n_852),
.Y(n_977)
);

NOR2xp33_ASAP7_75t_L g978 ( 
.A(n_768),
.B(n_276),
.Y(n_978)
);

BUFx2_ASAP7_75t_L g979 ( 
.A(n_740),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_838),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_838),
.B(n_580),
.Y(n_981)
);

AOI22xp5_ASAP7_75t_L g982 ( 
.A1(n_750),
.A2(n_677),
.B1(n_698),
.B2(n_683),
.Y(n_982)
);

INVx2_ASAP7_75t_L g983 ( 
.A(n_807),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_826),
.Y(n_984)
);

OAI21xp5_ASAP7_75t_L g985 ( 
.A1(n_718),
.A2(n_580),
.B(n_664),
.Y(n_985)
);

INVx2_ASAP7_75t_L g986 ( 
.A(n_813),
.Y(n_986)
);

NAND2xp5_ASAP7_75t_L g987 ( 
.A(n_816),
.B(n_683),
.Y(n_987)
);

AOI21xp5_ASAP7_75t_L g988 ( 
.A1(n_748),
.A2(n_635),
.B(n_581),
.Y(n_988)
);

AND2x2_ASAP7_75t_L g989 ( 
.A(n_712),
.B(n_426),
.Y(n_989)
);

OAI22xp5_ASAP7_75t_L g990 ( 
.A1(n_811),
.A2(n_698),
.B1(n_675),
.B2(n_664),
.Y(n_990)
);

AOI22xp33_ASAP7_75t_L g991 ( 
.A1(n_815),
.A2(n_668),
.B1(n_680),
.B2(n_675),
.Y(n_991)
);

INVx3_ASAP7_75t_L g992 ( 
.A(n_847),
.Y(n_992)
);

BUFx6f_ASAP7_75t_L g993 ( 
.A(n_847),
.Y(n_993)
);

BUFx3_ASAP7_75t_L g994 ( 
.A(n_847),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_SL g995 ( 
.A(n_858),
.B(n_630),
.Y(n_995)
);

INVx3_ASAP7_75t_L g996 ( 
.A(n_819),
.Y(n_996)
);

BUFx3_ASAP7_75t_L g997 ( 
.A(n_819),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_814),
.B(n_668),
.Y(n_998)
);

AND2x2_ASAP7_75t_SL g999 ( 
.A(n_799),
.B(n_827),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_858),
.B(n_630),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_732),
.B(n_680),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_848),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_863),
.B(n_679),
.Y(n_1003)
);

INVx3_ASAP7_75t_L g1004 ( 
.A(n_828),
.Y(n_1004)
);

INVx3_ASAP7_75t_L g1005 ( 
.A(n_828),
.Y(n_1005)
);

AND2x2_ASAP7_75t_SL g1006 ( 
.A(n_827),
.B(n_679),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_856),
.Y(n_1007)
);

NAND2xp5_ASAP7_75t_L g1008 ( 
.A(n_751),
.B(n_755),
.Y(n_1008)
);

AND2x4_ASAP7_75t_L g1009 ( 
.A(n_794),
.B(n_428),
.Y(n_1009)
);

NAND2xp5_ASAP7_75t_L g1010 ( 
.A(n_759),
.B(n_679),
.Y(n_1010)
);

NAND3xp33_ASAP7_75t_L g1011 ( 
.A(n_841),
.B(n_278),
.C(n_283),
.Y(n_1011)
);

BUFx6f_ASAP7_75t_L g1012 ( 
.A(n_774),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_794),
.B(n_428),
.Y(n_1013)
);

AND2x4_ASAP7_75t_L g1014 ( 
.A(n_796),
.B(n_685),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_829),
.Y(n_1015)
);

INVx4_ASAP7_75t_L g1016 ( 
.A(n_802),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_SL g1017 ( 
.A(n_823),
.B(n_685),
.Y(n_1017)
);

HB1xp67_ASAP7_75t_L g1018 ( 
.A(n_796),
.Y(n_1018)
);

NAND2xp5_ASAP7_75t_L g1019 ( 
.A(n_776),
.B(n_685),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_831),
.Y(n_1020)
);

INVx2_ASAP7_75t_L g1021 ( 
.A(n_832),
.Y(n_1021)
);

OR2x6_ASAP7_75t_L g1022 ( 
.A(n_802),
.B(n_581),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_797),
.B(n_834),
.Y(n_1023)
);

AOI22xp5_ASAP7_75t_L g1024 ( 
.A1(n_793),
.A2(n_700),
.B1(n_685),
.B2(n_602),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_835),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_862),
.B(n_685),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_864),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_857),
.Y(n_1028)
);

NOR3xp33_ASAP7_75t_SL g1029 ( 
.A(n_810),
.B(n_329),
.C(n_299),
.Y(n_1029)
);

NAND2xp5_ASAP7_75t_L g1030 ( 
.A(n_805),
.B(n_700),
.Y(n_1030)
);

OAI22xp33_ASAP7_75t_L g1031 ( 
.A1(n_728),
.A2(n_337),
.B1(n_295),
.B2(n_338),
.Y(n_1031)
);

BUFx3_ASAP7_75t_L g1032 ( 
.A(n_861),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_821),
.B(n_700),
.Y(n_1033)
);

AND2x2_ASAP7_75t_L g1034 ( 
.A(n_738),
.B(n_297),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_836),
.Y(n_1035)
);

NAND2x1p5_ASAP7_75t_L g1036 ( 
.A(n_836),
.B(n_581),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_802),
.Y(n_1037)
);

BUFx6f_ASAP7_75t_L g1038 ( 
.A(n_840),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_777),
.B(n_700),
.Y(n_1039)
);

INVx2_ASAP7_75t_L g1040 ( 
.A(n_840),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_757),
.Y(n_1041)
);

AOI22xp33_ASAP7_75t_SL g1042 ( 
.A1(n_822),
.A2(n_242),
.B1(n_243),
.B2(n_296),
.Y(n_1042)
);

INVx1_ASAP7_75t_L g1043 ( 
.A(n_771),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_778),
.B(n_700),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_891),
.Y(n_1045)
);

BUFx2_ASAP7_75t_L g1046 ( 
.A(n_918),
.Y(n_1046)
);

INVxp67_ASAP7_75t_L g1047 ( 
.A(n_915),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_895),
.A2(n_846),
.B(n_522),
.C(n_536),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_916),
.Y(n_1049)
);

INVx1_ASAP7_75t_L g1050 ( 
.A(n_916),
.Y(n_1050)
);

BUFx12f_ASAP7_75t_L g1051 ( 
.A(n_972),
.Y(n_1051)
);

AOI21xp33_ASAP7_75t_L g1052 ( 
.A1(n_978),
.A2(n_789),
.B(n_780),
.Y(n_1052)
);

INVx2_ASAP7_75t_SL g1053 ( 
.A(n_921),
.Y(n_1053)
);

NAND2xp5_ASAP7_75t_L g1054 ( 
.A(n_966),
.B(n_824),
.Y(n_1054)
);

AOI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_977),
.A2(n_839),
.B(n_581),
.Y(n_1055)
);

NOR2xp33_ASAP7_75t_R g1056 ( 
.A(n_901),
.B(n_817),
.Y(n_1056)
);

BUFx2_ASAP7_75t_L g1057 ( 
.A(n_918),
.Y(n_1057)
);

AO22x1_ASAP7_75t_L g1058 ( 
.A1(n_978),
.A2(n_357),
.B1(n_366),
.B2(n_333),
.Y(n_1058)
);

XOR2xp5_ASAP7_75t_L g1059 ( 
.A(n_961),
.B(n_817),
.Y(n_1059)
);

OA21x2_ASAP7_75t_L g1060 ( 
.A1(n_985),
.A2(n_855),
.B(n_594),
.Y(n_1060)
);

OAI22xp5_ASAP7_75t_L g1061 ( 
.A1(n_950),
.A2(n_860),
.B1(n_663),
.B2(n_635),
.Y(n_1061)
);

NOR2xp67_ASAP7_75t_L g1062 ( 
.A(n_961),
.B(n_63),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_871),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_968),
.B(n_531),
.Y(n_1064)
);

AOI21xp5_ASAP7_75t_L g1065 ( 
.A1(n_977),
.A2(n_635),
.B(n_663),
.Y(n_1065)
);

NAND3xp33_ASAP7_75t_L g1066 ( 
.A(n_923),
.B(n_324),
.C(n_322),
.Y(n_1066)
);

CKINVDCx11_ASAP7_75t_R g1067 ( 
.A(n_932),
.Y(n_1067)
);

O2A1O1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_917),
.A2(n_536),
.B(n_531),
.C(n_660),
.Y(n_1068)
);

OAI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_950),
.A2(n_860),
.B1(n_663),
.B2(n_635),
.Y(n_1069)
);

AOI22x1_ASAP7_75t_SL g1070 ( 
.A1(n_1016),
.A2(n_323),
.B1(n_312),
.B2(n_296),
.Y(n_1070)
);

NOR2xp33_ASAP7_75t_L g1071 ( 
.A(n_975),
.B(n_3),
.Y(n_1071)
);

AOI21xp5_ASAP7_75t_L g1072 ( 
.A1(n_920),
.A2(n_880),
.B(n_1023),
.Y(n_1072)
);

O2A1O1Ixp5_ASAP7_75t_L g1073 ( 
.A1(n_903),
.A2(n_599),
.B(n_584),
.C(n_660),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_920),
.A2(n_663),
.B(n_599),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_975),
.B(n_663),
.Y(n_1075)
);

OAI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_999),
.A2(n_596),
.B1(n_658),
.B2(n_653),
.Y(n_1076)
);

AOI21xp5_ASAP7_75t_L g1077 ( 
.A1(n_1026),
.A2(n_596),
.B(n_658),
.Y(n_1077)
);

OAI22xp5_ASAP7_75t_L g1078 ( 
.A1(n_999),
.A2(n_594),
.B1(n_653),
.B2(n_646),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_917),
.A2(n_592),
.B(n_646),
.C(n_644),
.Y(n_1079)
);

BUFx12f_ASAP7_75t_L g1080 ( 
.A(n_932),
.Y(n_1080)
);

INVx2_ASAP7_75t_L g1081 ( 
.A(n_892),
.Y(n_1081)
);

AOI21xp5_ASAP7_75t_L g1082 ( 
.A1(n_981),
.A2(n_592),
.B(n_644),
.Y(n_1082)
);

HB1xp67_ASAP7_75t_L g1083 ( 
.A(n_900),
.Y(n_1083)
);

INVx2_ASAP7_75t_L g1084 ( 
.A(n_892),
.Y(n_1084)
);

HB1xp67_ASAP7_75t_L g1085 ( 
.A(n_900),
.Y(n_1085)
);

INVx3_ASAP7_75t_L g1086 ( 
.A(n_869),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_SL g1087 ( 
.A(n_958),
.B(n_296),
.Y(n_1087)
);

BUFx12f_ASAP7_75t_L g1088 ( 
.A(n_932),
.Y(n_1088)
);

INVx8_ASAP7_75t_L g1089 ( 
.A(n_873),
.Y(n_1089)
);

AOI21xp33_ASAP7_75t_L g1090 ( 
.A1(n_944),
.A2(n_4),
.B(n_6),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_896),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_987),
.A2(n_591),
.B(n_636),
.Y(n_1092)
);

NAND2xp5_ASAP7_75t_SL g1093 ( 
.A(n_925),
.B(n_312),
.Y(n_1093)
);

NOR2xp33_ASAP7_75t_L g1094 ( 
.A(n_936),
.B(n_312),
.Y(n_1094)
);

INVx2_ASAP7_75t_SL g1095 ( 
.A(n_915),
.Y(n_1095)
);

AND2x2_ASAP7_75t_L g1096 ( 
.A(n_953),
.B(n_585),
.Y(n_1096)
);

NOR2xp33_ASAP7_75t_R g1097 ( 
.A(n_865),
.B(n_70),
.Y(n_1097)
);

INVx3_ASAP7_75t_L g1098 ( 
.A(n_869),
.Y(n_1098)
);

BUFx12f_ASAP7_75t_L g1099 ( 
.A(n_886),
.Y(n_1099)
);

AOI221x1_ASAP7_75t_L g1100 ( 
.A1(n_1016),
.A2(n_603),
.B1(n_636),
.B2(n_631),
.C(n_629),
.Y(n_1100)
);

A2O1A1Ixp33_ASAP7_75t_L g1101 ( 
.A1(n_984),
.A2(n_602),
.B(n_631),
.C(n_629),
.Y(n_1101)
);

BUFx2_ASAP7_75t_L g1102 ( 
.A(n_883),
.Y(n_1102)
);

NAND3xp33_ASAP7_75t_SL g1103 ( 
.A(n_923),
.B(n_591),
.C(n_609),
.Y(n_1103)
);

INVx2_ASAP7_75t_L g1104 ( 
.A(n_896),
.Y(n_1104)
);

AOI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_1008),
.A2(n_589),
.B(n_621),
.Y(n_1105)
);

HB1xp67_ASAP7_75t_L g1106 ( 
.A(n_884),
.Y(n_1106)
);

AND2x4_ASAP7_75t_L g1107 ( 
.A(n_949),
.B(n_97),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_1015),
.B(n_1020),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_867),
.A2(n_589),
.B(n_621),
.Y(n_1109)
);

OAI22xp5_ASAP7_75t_L g1110 ( 
.A1(n_1006),
.A2(n_590),
.B1(n_609),
.B2(n_606),
.Y(n_1110)
);

OAI21xp33_ASAP7_75t_L g1111 ( 
.A1(n_1042),
.A2(n_587),
.B(n_606),
.Y(n_1111)
);

NOR2xp33_ASAP7_75t_L g1112 ( 
.A(n_979),
.B(n_4),
.Y(n_1112)
);

INVx8_ASAP7_75t_L g1113 ( 
.A(n_873),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_931),
.B(n_604),
.Y(n_1114)
);

INVx3_ASAP7_75t_SL g1115 ( 
.A(n_1022),
.Y(n_1115)
);

NAND2xp33_ASAP7_75t_L g1116 ( 
.A(n_1038),
.B(n_478),
.Y(n_1116)
);

BUFx6f_ASAP7_75t_L g1117 ( 
.A(n_869),
.Y(n_1117)
);

AND2x2_ASAP7_75t_L g1118 ( 
.A(n_974),
.B(n_909),
.Y(n_1118)
);

BUFx2_ASAP7_75t_L g1119 ( 
.A(n_884),
.Y(n_1119)
);

INVx4_ASAP7_75t_L g1120 ( 
.A(n_869),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_938),
.A2(n_603),
.B(n_476),
.Y(n_1121)
);

NAND2xp5_ASAP7_75t_L g1122 ( 
.A(n_1025),
.B(n_502),
.Y(n_1122)
);

AO22x1_ASAP7_75t_L g1123 ( 
.A1(n_1037),
.A2(n_478),
.B1(n_501),
.B2(n_11),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_938),
.A2(n_476),
.B(n_475),
.Y(n_1124)
);

NOR2xp33_ASAP7_75t_L g1125 ( 
.A(n_939),
.B(n_6),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_876),
.Y(n_1126)
);

AOI21xp5_ASAP7_75t_L g1127 ( 
.A1(n_893),
.A2(n_476),
.B(n_502),
.Y(n_1127)
);

AOI22xp33_ASAP7_75t_L g1128 ( 
.A1(n_1028),
.A2(n_502),
.B1(n_501),
.B2(n_478),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_902),
.Y(n_1129)
);

BUFx12f_ASAP7_75t_L g1130 ( 
.A(n_927),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_973),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_1029),
.Y(n_1132)
);

BUFx4f_ASAP7_75t_SL g1133 ( 
.A(n_1032),
.Y(n_1133)
);

INVxp67_ASAP7_75t_L g1134 ( 
.A(n_905),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_L g1135 ( 
.A1(n_998),
.A2(n_478),
.B(n_501),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_902),
.Y(n_1136)
);

AOI21x1_ASAP7_75t_L g1137 ( 
.A1(n_1017),
.A2(n_501),
.B(n_478),
.Y(n_1137)
);

NOR2xp33_ASAP7_75t_L g1138 ( 
.A(n_1031),
.B(n_10),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1021),
.B(n_501),
.Y(n_1139)
);

NAND2xp5_ASAP7_75t_L g1140 ( 
.A(n_1021),
.B(n_10),
.Y(n_1140)
);

NOR2xp33_ASAP7_75t_L g1141 ( 
.A(n_1031),
.B(n_11),
.Y(n_1141)
);

OAI21xp33_ASAP7_75t_L g1142 ( 
.A1(n_1042),
.A2(n_12),
.B(n_16),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_965),
.A2(n_478),
.B(n_180),
.Y(n_1143)
);

O2A1O1Ixp33_ASAP7_75t_SL g1144 ( 
.A1(n_995),
.A2(n_177),
.B(n_173),
.C(n_169),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1027),
.B(n_16),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_928),
.Y(n_1146)
);

BUFx2_ASAP7_75t_L g1147 ( 
.A(n_1018),
.Y(n_1147)
);

NOR2xp33_ASAP7_75t_L g1148 ( 
.A(n_942),
.B(n_17),
.Y(n_1148)
);

BUFx2_ASAP7_75t_SL g1149 ( 
.A(n_927),
.Y(n_1149)
);

NAND2xp5_ASAP7_75t_L g1150 ( 
.A(n_1027),
.B(n_17),
.Y(n_1150)
);

BUFx6f_ASAP7_75t_L g1151 ( 
.A(n_899),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_933),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_935),
.Y(n_1153)
);

BUFx8_ASAP7_75t_L g1154 ( 
.A(n_1037),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_868),
.Y(n_1155)
);

AOI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_947),
.A2(n_478),
.B(n_167),
.Y(n_1156)
);

O2A1O1Ixp33_ASAP7_75t_L g1157 ( 
.A1(n_957),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_1157)
);

A2O1A1Ixp33_ASAP7_75t_L g1158 ( 
.A1(n_962),
.A2(n_23),
.B(n_28),
.C(n_29),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_980),
.B(n_31),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_949),
.B(n_152),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_937),
.B(n_951),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_973),
.Y(n_1162)
);

INVx3_ASAP7_75t_L g1163 ( 
.A(n_899),
.Y(n_1163)
);

BUFx6f_ASAP7_75t_L g1164 ( 
.A(n_899),
.Y(n_1164)
);

INVx1_ASAP7_75t_SL g1165 ( 
.A(n_1009),
.Y(n_1165)
);

NOR2xp33_ASAP7_75t_L g1166 ( 
.A(n_942),
.B(n_32),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_890),
.A2(n_478),
.B(n_140),
.Y(n_1167)
);

NAND2xp5_ASAP7_75t_L g1168 ( 
.A(n_930),
.B(n_35),
.Y(n_1168)
);

INVx3_ASAP7_75t_SL g1169 ( 
.A(n_1022),
.Y(n_1169)
);

O2A1O1Ixp5_ASAP7_75t_L g1170 ( 
.A1(n_1017),
.A2(n_129),
.B(n_125),
.C(n_119),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_SL g1171 ( 
.A(n_1006),
.B(n_109),
.Y(n_1171)
);

HB1xp67_ASAP7_75t_L g1172 ( 
.A(n_879),
.Y(n_1172)
);

INVx2_ASAP7_75t_SL g1173 ( 
.A(n_1009),
.Y(n_1173)
);

NAND3xp33_ASAP7_75t_SL g1174 ( 
.A(n_872),
.B(n_36),
.C(n_37),
.Y(n_1174)
);

HB1xp67_ASAP7_75t_L g1175 ( 
.A(n_879),
.Y(n_1175)
);

AOI21xp5_ASAP7_75t_L g1176 ( 
.A1(n_956),
.A2(n_108),
.B(n_105),
.Y(n_1176)
);

HB1xp67_ASAP7_75t_L g1177 ( 
.A(n_881),
.Y(n_1177)
);

NOR2xp33_ASAP7_75t_L g1178 ( 
.A(n_1018),
.B(n_1034),
.Y(n_1178)
);

OAI22xp5_ASAP7_75t_L g1179 ( 
.A1(n_959),
.A2(n_101),
.B1(n_82),
.B2(n_40),
.Y(n_1179)
);

AND2x4_ASAP7_75t_L g1180 ( 
.A(n_874),
.B(n_37),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_955),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1010),
.A2(n_60),
.B(n_40),
.Y(n_1182)
);

AOI21xp5_ASAP7_75t_L g1183 ( 
.A1(n_1019),
.A2(n_1033),
.B(n_1039),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_899),
.Y(n_1184)
);

AOI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_967),
.A2(n_59),
.B(n_41),
.Y(n_1185)
);

CKINVDCx6p67_ASAP7_75t_R g1186 ( 
.A(n_1032),
.Y(n_1186)
);

NOR2xp33_ASAP7_75t_L g1187 ( 
.A(n_1013),
.B(n_39),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_882),
.B(n_42),
.Y(n_1188)
);

AO21x1_ASAP7_75t_L g1189 ( 
.A1(n_1044),
.A2(n_43),
.B(n_49),
.Y(n_1189)
);

OAI21x1_ASAP7_75t_L g1190 ( 
.A1(n_988),
.A2(n_43),
.B(n_50),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_955),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_874),
.B(n_50),
.Y(n_1192)
);

NAND2x1_ASAP7_75t_L g1193 ( 
.A(n_924),
.B(n_51),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_1108),
.B(n_941),
.Y(n_1194)
);

CKINVDCx11_ASAP7_75t_R g1195 ( 
.A(n_1051),
.Y(n_1195)
);

INVx3_ASAP7_75t_L g1196 ( 
.A(n_1089),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_1138),
.A2(n_872),
.B1(n_870),
.B2(n_1013),
.Y(n_1197)
);

AOI221x1_ASAP7_75t_L g1198 ( 
.A1(n_1090),
.A2(n_1011),
.B1(n_1041),
.B2(n_1043),
.C(n_866),
.Y(n_1198)
);

A2O1A1Ixp33_ASAP7_75t_L g1199 ( 
.A1(n_1052),
.A2(n_1029),
.B(n_889),
.C(n_913),
.Y(n_1199)
);

NAND2x1_ASAP7_75t_L g1200 ( 
.A(n_1120),
.B(n_924),
.Y(n_1200)
);

NAND2x1p5_ASAP7_75t_L g1201 ( 
.A(n_1046),
.B(n_994),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1065),
.A2(n_1109),
.B(n_1055),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_1183),
.A2(n_945),
.B(n_1030),
.Y(n_1203)
);

NAND2xp5_ASAP7_75t_L g1204 ( 
.A(n_1118),
.B(n_1096),
.Y(n_1204)
);

OAI21xp5_ASAP7_75t_L g1205 ( 
.A1(n_1072),
.A2(n_870),
.B(n_948),
.Y(n_1205)
);

AOI211x1_ASAP7_75t_L g1206 ( 
.A1(n_1142),
.A2(n_911),
.B(n_897),
.C(n_943),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1054),
.A2(n_885),
.B(n_907),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_1146),
.Y(n_1208)
);

A2O1A1Ixp33_ASAP7_75t_L g1209 ( 
.A1(n_1094),
.A2(n_1141),
.B(n_1125),
.C(n_1066),
.Y(n_1209)
);

OAI21xp5_ASAP7_75t_L g1210 ( 
.A1(n_1073),
.A2(n_870),
.B(n_877),
.Y(n_1210)
);

AOI21x1_ASAP7_75t_L g1211 ( 
.A1(n_1100),
.A2(n_990),
.B(n_1001),
.Y(n_1211)
);

AO31x2_ASAP7_75t_L g1212 ( 
.A1(n_1189),
.A2(n_934),
.A3(n_922),
.B(n_906),
.Y(n_1212)
);

A2O1A1Ixp33_ASAP7_75t_L g1213 ( 
.A1(n_1125),
.A2(n_964),
.B(n_919),
.C(n_1000),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1131),
.B(n_870),
.Y(n_1214)
);

AOI21xp5_ASAP7_75t_L g1215 ( 
.A1(n_1105),
.A2(n_907),
.B(n_885),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1131),
.B(n_870),
.Y(n_1216)
);

NAND2xp5_ASAP7_75t_L g1217 ( 
.A(n_1162),
.B(n_1012),
.Y(n_1217)
);

AO31x2_ASAP7_75t_L g1218 ( 
.A1(n_1110),
.A2(n_910),
.A3(n_914),
.B(n_1003),
.Y(n_1218)
);

OAI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1115),
.A2(n_881),
.B1(n_888),
.B2(n_1022),
.Y(n_1219)
);

OR2x6_ASAP7_75t_SL g1220 ( 
.A(n_1132),
.B(n_878),
.Y(n_1220)
);

AND2x2_ASAP7_75t_L g1221 ( 
.A(n_1178),
.B(n_926),
.Y(n_1221)
);

NAND2xp5_ASAP7_75t_SL g1222 ( 
.A(n_1102),
.B(n_1014),
.Y(n_1222)
);

CKINVDCx8_ASAP7_75t_R g1223 ( 
.A(n_1149),
.Y(n_1223)
);

AOI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1061),
.A2(n_885),
.B(n_907),
.Y(n_1224)
);

HB1xp67_ASAP7_75t_L g1225 ( 
.A(n_1083),
.Y(n_1225)
);

AOI21xp5_ASAP7_75t_L g1226 ( 
.A1(n_1069),
.A2(n_898),
.B(n_894),
.Y(n_1226)
);

A2O1A1Ixp33_ASAP7_75t_L g1227 ( 
.A1(n_1103),
.A2(n_1024),
.B(n_976),
.C(n_929),
.Y(n_1227)
);

INVx1_ASAP7_75t_L g1228 ( 
.A(n_1152),
.Y(n_1228)
);

AOI221xp5_ASAP7_75t_L g1229 ( 
.A1(n_1112),
.A2(n_1012),
.B1(n_991),
.B2(n_986),
.C(n_983),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_1171),
.A2(n_894),
.B(n_1012),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1162),
.B(n_1012),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1082),
.A2(n_873),
.B(n_993),
.Y(n_1232)
);

OAI21x1_ASAP7_75t_L g1233 ( 
.A1(n_1127),
.A2(n_971),
.B(n_991),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_1117),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_1153),
.Y(n_1235)
);

NAND2xp33_ASAP7_75t_R g1236 ( 
.A(n_1097),
.B(n_888),
.Y(n_1236)
);

INVx2_ASAP7_75t_L g1237 ( 
.A(n_1045),
.Y(n_1237)
);

AND2x4_ASAP7_75t_L g1238 ( 
.A(n_1173),
.B(n_994),
.Y(n_1238)
);

NAND2xp5_ASAP7_75t_L g1239 ( 
.A(n_1161),
.B(n_1014),
.Y(n_1239)
);

AOI21xp5_ASAP7_75t_SL g1240 ( 
.A1(n_1107),
.A2(n_970),
.B(n_993),
.Y(n_1240)
);

AND2x2_ASAP7_75t_L g1241 ( 
.A(n_1165),
.B(n_888),
.Y(n_1241)
);

OAI21x1_ASAP7_75t_L g1242 ( 
.A1(n_1074),
.A2(n_1002),
.B(n_986),
.Y(n_1242)
);

INVxp67_ASAP7_75t_L g1243 ( 
.A(n_1106),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1077),
.A2(n_1007),
.B(n_983),
.Y(n_1244)
);

OAI22x1_ASAP7_75t_L g1245 ( 
.A1(n_1112),
.A2(n_954),
.B1(n_1036),
.B2(n_1035),
.Y(n_1245)
);

AO31x2_ASAP7_75t_L g1246 ( 
.A1(n_1076),
.A2(n_1035),
.A3(n_969),
.B(n_1007),
.Y(n_1246)
);

NOR2xp33_ASAP7_75t_L g1247 ( 
.A(n_1133),
.B(n_946),
.Y(n_1247)
);

HB1xp67_ASAP7_75t_L g1248 ( 
.A(n_1083),
.Y(n_1248)
);

AOI21xp5_ASAP7_75t_L g1249 ( 
.A1(n_1122),
.A2(n_970),
.B(n_993),
.Y(n_1249)
);

AOI221x1_ASAP7_75t_L g1250 ( 
.A1(n_1103),
.A2(n_940),
.B1(n_992),
.B2(n_912),
.C(n_887),
.Y(n_1250)
);

AND2x4_ASAP7_75t_L g1251 ( 
.A(n_1107),
.B(n_940),
.Y(n_1251)
);

INVx3_ASAP7_75t_L g1252 ( 
.A(n_1089),
.Y(n_1252)
);

NAND2xp5_ASAP7_75t_L g1253 ( 
.A(n_1064),
.B(n_1040),
.Y(n_1253)
);

INVx2_ASAP7_75t_SL g1254 ( 
.A(n_1057),
.Y(n_1254)
);

OAI21xp5_ASAP7_75t_L g1255 ( 
.A1(n_1079),
.A2(n_904),
.B(n_982),
.Y(n_1255)
);

INVx3_ASAP7_75t_L g1256 ( 
.A(n_1089),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1134),
.B(n_963),
.Y(n_1257)
);

NAND2xp33_ASAP7_75t_L g1258 ( 
.A(n_1113),
.B(n_952),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1071),
.B(n_963),
.Y(n_1259)
);

NOR2xp33_ASAP7_75t_L g1260 ( 
.A(n_1133),
.B(n_1038),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1058),
.B(n_1038),
.C(n_969),
.Y(n_1261)
);

INVx1_ASAP7_75t_L g1262 ( 
.A(n_1155),
.Y(n_1262)
);

AO21x1_ASAP7_75t_L g1263 ( 
.A1(n_1179),
.A2(n_1036),
.B(n_960),
.Y(n_1263)
);

BUFx8_ASAP7_75t_L g1264 ( 
.A(n_1130),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_L g1265 ( 
.A(n_1071),
.B(n_960),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1053),
.B(n_1038),
.Y(n_1266)
);

OAI22x1_ASAP7_75t_L g1267 ( 
.A1(n_1115),
.A2(n_954),
.B1(n_1002),
.B2(n_908),
.Y(n_1267)
);

INVx2_ASAP7_75t_SL g1268 ( 
.A(n_1119),
.Y(n_1268)
);

OR2x2_ASAP7_75t_L g1269 ( 
.A(n_1085),
.B(n_997),
.Y(n_1269)
);

INVx2_ASAP7_75t_SL g1270 ( 
.A(n_1106),
.Y(n_1270)
);

INVx3_ASAP7_75t_L g1271 ( 
.A(n_1113),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1092),
.A2(n_996),
.B(n_1004),
.Y(n_1272)
);

BUFx6f_ASAP7_75t_SL g1273 ( 
.A(n_1180),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_L g1274 ( 
.A(n_1168),
.B(n_1004),
.Y(n_1274)
);

OAI21x1_ASAP7_75t_L g1275 ( 
.A1(n_1137),
.A2(n_1005),
.B(n_952),
.Y(n_1275)
);

OAI21x1_ASAP7_75t_L g1276 ( 
.A1(n_1121),
.A2(n_1005),
.B(n_952),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1169),
.A2(n_952),
.B1(n_56),
.B2(n_58),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_1117),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1134),
.B(n_952),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1124),
.A2(n_52),
.B(n_1078),
.Y(n_1280)
);

AOI21xp5_ASAP7_75t_L g1281 ( 
.A1(n_1060),
.A2(n_52),
.B(n_1075),
.Y(n_1281)
);

NOR2xp67_ASAP7_75t_L g1282 ( 
.A(n_1120),
.B(n_1140),
.Y(n_1282)
);

OAI21x1_ASAP7_75t_L g1283 ( 
.A1(n_1079),
.A2(n_1190),
.B(n_1060),
.Y(n_1283)
);

AND2x2_ASAP7_75t_L g1284 ( 
.A(n_1180),
.B(n_1085),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1167),
.A2(n_1135),
.B(n_1170),
.Y(n_1285)
);

INVx4_ASAP7_75t_SL g1286 ( 
.A(n_1169),
.Y(n_1286)
);

AOI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1114),
.A2(n_1062),
.B(n_1150),
.Y(n_1287)
);

OAI21x1_ASAP7_75t_L g1288 ( 
.A1(n_1170),
.A2(n_1063),
.B(n_1126),
.Y(n_1288)
);

NAND2xp5_ASAP7_75t_L g1289 ( 
.A(n_1049),
.B(n_1050),
.Y(n_1289)
);

OAI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1101),
.A2(n_1068),
.B(n_1111),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1113),
.Y(n_1291)
);

AOI221xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1158),
.A2(n_1157),
.B1(n_1145),
.B2(n_1182),
.C(n_1188),
.Y(n_1292)
);

NAND3x1_ASAP7_75t_L g1293 ( 
.A(n_1148),
.B(n_1166),
.C(n_1187),
.Y(n_1293)
);

AOI21x1_ASAP7_75t_L g1294 ( 
.A1(n_1087),
.A2(n_1159),
.B(n_1156),
.Y(n_1294)
);

NOR2xp67_ASAP7_75t_L g1295 ( 
.A(n_1081),
.B(n_1136),
.Y(n_1295)
);

OAI21x1_ASAP7_75t_L g1296 ( 
.A1(n_1084),
.A2(n_1091),
.B(n_1129),
.Y(n_1296)
);

OAI21xp5_ASAP7_75t_L g1297 ( 
.A1(n_1068),
.A2(n_1048),
.B(n_1185),
.Y(n_1297)
);

OAI21xp5_ASAP7_75t_L g1298 ( 
.A1(n_1048),
.A2(n_1176),
.B(n_1139),
.Y(n_1298)
);

NAND2xp5_ASAP7_75t_L g1299 ( 
.A(n_1188),
.B(n_1095),
.Y(n_1299)
);

INVx3_ASAP7_75t_L g1300 ( 
.A(n_1117),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1104),
.B(n_1047),
.Y(n_1301)
);

BUFx6f_ASAP7_75t_L g1302 ( 
.A(n_1117),
.Y(n_1302)
);

CKINVDCx5p33_ASAP7_75t_R g1303 ( 
.A(n_1056),
.Y(n_1303)
);

OR2x2_ASAP7_75t_L g1304 ( 
.A(n_1147),
.B(n_1047),
.Y(n_1304)
);

OA21x2_ASAP7_75t_L g1305 ( 
.A1(n_1143),
.A2(n_1181),
.B(n_1191),
.Y(n_1305)
);

BUFx2_ASAP7_75t_R g1306 ( 
.A(n_1192),
.Y(n_1306)
);

NAND2xp33_ASAP7_75t_R g1307 ( 
.A(n_1070),
.B(n_1163),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1172),
.Y(n_1308)
);

NAND2xp5_ASAP7_75t_L g1309 ( 
.A(n_1172),
.B(n_1175),
.Y(n_1309)
);

BUFx6f_ASAP7_75t_L g1310 ( 
.A(n_1151),
.Y(n_1310)
);

AOI21xp33_ASAP7_75t_L g1311 ( 
.A1(n_1099),
.A2(n_1093),
.B(n_1157),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1177),
.Y(n_1312)
);

AOI21xp5_ASAP7_75t_L g1313 ( 
.A1(n_1144),
.A2(n_1116),
.B(n_1160),
.Y(n_1313)
);

AOI21x1_ASAP7_75t_L g1314 ( 
.A1(n_1193),
.A2(n_1123),
.B(n_1059),
.Y(n_1314)
);

A2O1A1Ixp33_ASAP7_75t_L g1315 ( 
.A1(n_1174),
.A2(n_1098),
.B(n_1163),
.C(n_1086),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1186),
.B(n_1086),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_1151),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_L g1318 ( 
.A(n_1098),
.B(n_1174),
.Y(n_1318)
);

BUFx6f_ASAP7_75t_L g1319 ( 
.A(n_1151),
.Y(n_1319)
);

AND2x2_ASAP7_75t_L g1320 ( 
.A(n_1067),
.B(n_1080),
.Y(n_1320)
);

INVx5_ASAP7_75t_L g1321 ( 
.A(n_1164),
.Y(n_1321)
);

A2O1A1Ixp33_ASAP7_75t_L g1322 ( 
.A1(n_1128),
.A2(n_1164),
.B(n_1184),
.C(n_1154),
.Y(n_1322)
);

INVx2_ASAP7_75t_SL g1323 ( 
.A(n_1154),
.Y(n_1323)
);

AOI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1164),
.A2(n_1184),
.B(n_1128),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1184),
.Y(n_1325)
);

NAND2xp5_ASAP7_75t_L g1326 ( 
.A(n_1184),
.B(n_1088),
.Y(n_1326)
);

NAND2xp5_ASAP7_75t_L g1327 ( 
.A(n_1108),
.B(n_875),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1108),
.B(n_875),
.Y(n_1328)
);

OAI21x1_ASAP7_75t_L g1329 ( 
.A1(n_1065),
.A2(n_1109),
.B(n_1055),
.Y(n_1329)
);

AOI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1183),
.A2(n_977),
.B(n_1072),
.Y(n_1330)
);

AND2x2_ASAP7_75t_L g1331 ( 
.A(n_1118),
.B(n_989),
.Y(n_1331)
);

OAI21xp5_ASAP7_75t_SL g1332 ( 
.A1(n_1138),
.A2(n_804),
.B(n_784),
.Y(n_1332)
);

NAND2x1p5_ASAP7_75t_L g1333 ( 
.A(n_1046),
.B(n_1057),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1099),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1108),
.B(n_875),
.Y(n_1335)
);

AOI21xp5_ASAP7_75t_L g1336 ( 
.A1(n_1183),
.A2(n_977),
.B(n_1072),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_1146),
.Y(n_1337)
);

OAI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1072),
.A2(n_895),
.B(n_1183),
.Y(n_1338)
);

BUFx6f_ASAP7_75t_L g1339 ( 
.A(n_1117),
.Y(n_1339)
);

NAND2xp5_ASAP7_75t_SL g1340 ( 
.A(n_1178),
.B(n_865),
.Y(n_1340)
);

AO31x2_ASAP7_75t_L g1341 ( 
.A1(n_1100),
.A2(n_1183),
.A3(n_1189),
.B(n_1072),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1072),
.A2(n_895),
.B(n_1183),
.Y(n_1342)
);

INVx1_ASAP7_75t_L g1343 ( 
.A(n_1146),
.Y(n_1343)
);

OAI21xp5_ASAP7_75t_L g1344 ( 
.A1(n_1072),
.A2(n_895),
.B(n_1183),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1146),
.Y(n_1345)
);

AOI21xp5_ASAP7_75t_L g1346 ( 
.A1(n_1183),
.A2(n_977),
.B(n_1072),
.Y(n_1346)
);

NAND2x1p5_ASAP7_75t_L g1347 ( 
.A(n_1046),
.B(n_1057),
.Y(n_1347)
);

INVx1_ASAP7_75t_L g1348 ( 
.A(n_1146),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1296),
.Y(n_1349)
);

INVx3_ASAP7_75t_L g1350 ( 
.A(n_1321),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1237),
.Y(n_1351)
);

AO21x2_ASAP7_75t_L g1352 ( 
.A1(n_1297),
.A2(n_1205),
.B(n_1210),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1215),
.A2(n_1224),
.B(n_1287),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1327),
.B(n_1328),
.Y(n_1354)
);

OR2x2_ASAP7_75t_L g1355 ( 
.A(n_1204),
.B(n_1304),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1331),
.B(n_1221),
.Y(n_1356)
);

OAI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1209),
.A2(n_1332),
.B(n_1199),
.Y(n_1357)
);

OA21x2_ASAP7_75t_L g1358 ( 
.A1(n_1297),
.A2(n_1250),
.B(n_1210),
.Y(n_1358)
);

BUFx3_ASAP7_75t_L g1359 ( 
.A(n_1333),
.Y(n_1359)
);

OA21x2_ASAP7_75t_L g1360 ( 
.A1(n_1283),
.A2(n_1342),
.B(n_1338),
.Y(n_1360)
);

INVx3_ASAP7_75t_L g1361 ( 
.A(n_1321),
.Y(n_1361)
);

INVx4_ASAP7_75t_L g1362 ( 
.A(n_1321),
.Y(n_1362)
);

OA21x2_ASAP7_75t_L g1363 ( 
.A1(n_1338),
.A2(n_1344),
.B(n_1342),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1208),
.Y(n_1364)
);

INVx4_ASAP7_75t_L g1365 ( 
.A(n_1286),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1336),
.A2(n_1346),
.B(n_1232),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1197),
.A2(n_1335),
.B1(n_1311),
.B2(n_1332),
.Y(n_1367)
);

OA21x2_ASAP7_75t_L g1368 ( 
.A1(n_1344),
.A2(n_1205),
.B(n_1290),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1228),
.Y(n_1369)
);

INVx2_ASAP7_75t_L g1370 ( 
.A(n_1235),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1262),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1337),
.Y(n_1372)
);

BUFx2_ASAP7_75t_L g1373 ( 
.A(n_1268),
.Y(n_1373)
);

AO21x2_ASAP7_75t_L g1374 ( 
.A1(n_1290),
.A2(n_1281),
.B(n_1263),
.Y(n_1374)
);

NOR2xp67_ASAP7_75t_L g1375 ( 
.A(n_1243),
.B(n_1270),
.Y(n_1375)
);

INVxp67_ASAP7_75t_SL g1376 ( 
.A(n_1225),
.Y(n_1376)
);

A2O1A1Ixp33_ASAP7_75t_L g1377 ( 
.A1(n_1197),
.A2(n_1292),
.B(n_1213),
.C(n_1194),
.Y(n_1377)
);

AO21x2_ASAP7_75t_L g1378 ( 
.A1(n_1298),
.A2(n_1255),
.B(n_1203),
.Y(n_1378)
);

NOR2xp33_ASAP7_75t_L g1379 ( 
.A(n_1299),
.B(n_1239),
.Y(n_1379)
);

OAI21x1_ASAP7_75t_SL g1380 ( 
.A1(n_1259),
.A2(n_1265),
.B(n_1314),
.Y(n_1380)
);

INVx4_ASAP7_75t_L g1381 ( 
.A(n_1286),
.Y(n_1381)
);

OAI21x1_ASAP7_75t_L g1382 ( 
.A1(n_1285),
.A2(n_1276),
.B(n_1244),
.Y(n_1382)
);

AO31x2_ASAP7_75t_L g1383 ( 
.A1(n_1198),
.A2(n_1245),
.A3(n_1226),
.B(n_1227),
.Y(n_1383)
);

NAND2xp33_ASAP7_75t_R g1384 ( 
.A(n_1260),
.B(n_1214),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1242),
.A2(n_1233),
.B(n_1288),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1275),
.A2(n_1280),
.B(n_1272),
.Y(n_1386)
);

CKINVDCx11_ASAP7_75t_R g1387 ( 
.A(n_1195),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1261),
.A2(n_1230),
.B(n_1298),
.Y(n_1388)
);

AOI22xp33_ASAP7_75t_L g1389 ( 
.A1(n_1277),
.A2(n_1340),
.B1(n_1253),
.B2(n_1318),
.Y(n_1389)
);

NAND2x1p5_ASAP7_75t_L g1390 ( 
.A(n_1196),
.B(n_1252),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1343),
.Y(n_1391)
);

AOI22xp33_ASAP7_75t_SL g1392 ( 
.A1(n_1273),
.A2(n_1241),
.B1(n_1334),
.B2(n_1261),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1345),
.Y(n_1393)
);

AO21x2_ASAP7_75t_L g1394 ( 
.A1(n_1255),
.A2(n_1294),
.B(n_1207),
.Y(n_1394)
);

INVx2_ASAP7_75t_L g1395 ( 
.A(n_1348),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1211),
.A2(n_1249),
.B(n_1324),
.Y(n_1396)
);

INVx1_ASAP7_75t_L g1397 ( 
.A(n_1301),
.Y(n_1397)
);

CKINVDCx6p67_ASAP7_75t_R g1398 ( 
.A(n_1273),
.Y(n_1398)
);

A2O1A1Ixp33_ASAP7_75t_L g1399 ( 
.A1(n_1229),
.A2(n_1258),
.B(n_1313),
.C(n_1322),
.Y(n_1399)
);

OAI21x1_ASAP7_75t_L g1400 ( 
.A1(n_1305),
.A2(n_1216),
.B(n_1279),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1305),
.A2(n_1274),
.B(n_1219),
.Y(n_1401)
);

NOR2xp33_ASAP7_75t_SL g1402 ( 
.A(n_1223),
.B(n_1303),
.Y(n_1402)
);

NAND2x1p5_ASAP7_75t_L g1403 ( 
.A(n_1252),
.B(n_1271),
.Y(n_1403)
);

OAI22xp5_ASAP7_75t_L g1404 ( 
.A1(n_1293),
.A2(n_1220),
.B1(n_1240),
.B2(n_1306),
.Y(n_1404)
);

INVx1_ASAP7_75t_L g1405 ( 
.A(n_1289),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1248),
.Y(n_1406)
);

A2O1A1Ixp33_ASAP7_75t_L g1407 ( 
.A1(n_1257),
.A2(n_1282),
.B(n_1315),
.C(n_1251),
.Y(n_1407)
);

OAI222xp33_ASAP7_75t_L g1408 ( 
.A1(n_1222),
.A2(n_1217),
.B1(n_1231),
.B2(n_1284),
.C1(n_1269),
.C2(n_1266),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1282),
.A2(n_1291),
.B(n_1271),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1256),
.A2(n_1291),
.B(n_1200),
.Y(n_1410)
);

OAI21x1_ASAP7_75t_L g1411 ( 
.A1(n_1256),
.A2(n_1300),
.B(n_1317),
.Y(n_1411)
);

NAND2xp5_ASAP7_75t_L g1412 ( 
.A(n_1309),
.B(n_1254),
.Y(n_1412)
);

AOI21xp5_ASAP7_75t_L g1413 ( 
.A1(n_1295),
.A2(n_1267),
.B(n_1341),
.Y(n_1413)
);

BUFx3_ASAP7_75t_L g1414 ( 
.A(n_1347),
.Y(n_1414)
);

BUFx2_ASAP7_75t_L g1415 ( 
.A(n_1201),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1325),
.A2(n_1312),
.B(n_1308),
.Y(n_1416)
);

NAND2x1_ASAP7_75t_L g1417 ( 
.A(n_1234),
.B(n_1302),
.Y(n_1417)
);

INVx8_ASAP7_75t_L g1418 ( 
.A(n_1234),
.Y(n_1418)
);

INVx1_ASAP7_75t_L g1419 ( 
.A(n_1206),
.Y(n_1419)
);

OR2x6_ASAP7_75t_L g1420 ( 
.A(n_1206),
.B(n_1323),
.Y(n_1420)
);

INVx5_ASAP7_75t_L g1421 ( 
.A(n_1234),
.Y(n_1421)
);

OAI21xp5_ASAP7_75t_L g1422 ( 
.A1(n_1316),
.A2(n_1238),
.B(n_1326),
.Y(n_1422)
);

OAI21xp5_ASAP7_75t_L g1423 ( 
.A1(n_1238),
.A2(n_1247),
.B(n_1236),
.Y(n_1423)
);

BUFx3_ASAP7_75t_L g1424 ( 
.A(n_1264),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1278),
.Y(n_1425)
);

AND2x4_ASAP7_75t_L g1426 ( 
.A(n_1278),
.B(n_1339),
.Y(n_1426)
);

INVx3_ASAP7_75t_L g1427 ( 
.A(n_1278),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1302),
.Y(n_1428)
);

OAI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1320),
.A2(n_1339),
.B1(n_1319),
.B2(n_1310),
.Y(n_1429)
);

INVxp67_ASAP7_75t_L g1430 ( 
.A(n_1307),
.Y(n_1430)
);

AO21x1_ASAP7_75t_L g1431 ( 
.A1(n_1212),
.A2(n_1341),
.B(n_1246),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1302),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1310),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1341),
.A2(n_1246),
.B(n_1218),
.Y(n_1434)
);

OAI21xp5_ASAP7_75t_L g1435 ( 
.A1(n_1212),
.A2(n_1218),
.B(n_1246),
.Y(n_1435)
);

OAI221xp5_ASAP7_75t_L g1436 ( 
.A1(n_1310),
.A2(n_1319),
.B1(n_1339),
.B2(n_1264),
.C(n_1212),
.Y(n_1436)
);

OAI21x1_ASAP7_75t_L g1437 ( 
.A1(n_1218),
.A2(n_1283),
.B(n_1202),
.Y(n_1437)
);

INVx4_ASAP7_75t_L g1438 ( 
.A(n_1319),
.Y(n_1438)
);

AO31x2_ASAP7_75t_L g1439 ( 
.A1(n_1250),
.A2(n_1263),
.A3(n_1336),
.B(n_1330),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1225),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1208),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1443)
);

OA21x2_ASAP7_75t_L g1444 ( 
.A1(n_1297),
.A2(n_1250),
.B(n_1210),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1321),
.B(n_1196),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1208),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1296),
.Y(n_1447)
);

HB1xp67_ASAP7_75t_L g1448 ( 
.A(n_1225),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1296),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1208),
.Y(n_1450)
);

BUFx6f_ASAP7_75t_L g1451 ( 
.A(n_1321),
.Y(n_1451)
);

BUFx12f_ASAP7_75t_L g1452 ( 
.A(n_1195),
.Y(n_1452)
);

OAI21xp5_ASAP7_75t_L g1453 ( 
.A1(n_1209),
.A2(n_895),
.B(n_978),
.Y(n_1453)
);

INVx3_ASAP7_75t_L g1454 ( 
.A(n_1321),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1208),
.Y(n_1455)
);

OAI21x1_ASAP7_75t_L g1456 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1331),
.B(n_1221),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1208),
.Y(n_1458)
);

OAI21x1_ASAP7_75t_L g1459 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1459)
);

AO21x1_ASAP7_75t_L g1460 ( 
.A1(n_1332),
.A2(n_895),
.B(n_1090),
.Y(n_1460)
);

OAI21x1_ASAP7_75t_L g1461 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1461)
);

OAI22xp33_ASAP7_75t_SL g1462 ( 
.A1(n_1197),
.A2(n_1138),
.B1(n_1141),
.B2(n_895),
.Y(n_1462)
);

NOR2xp33_ASAP7_75t_L g1463 ( 
.A(n_1332),
.B(n_961),
.Y(n_1463)
);

BUFx3_ASAP7_75t_L g1464 ( 
.A(n_1333),
.Y(n_1464)
);

HB1xp67_ASAP7_75t_L g1465 ( 
.A(n_1225),
.Y(n_1465)
);

BUFx3_ASAP7_75t_L g1466 ( 
.A(n_1333),
.Y(n_1466)
);

INVx2_ASAP7_75t_L g1467 ( 
.A(n_1296),
.Y(n_1467)
);

INVx2_ASAP7_75t_L g1468 ( 
.A(n_1296),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1469)
);

HB1xp67_ASAP7_75t_L g1470 ( 
.A(n_1225),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1208),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1208),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1473)
);

O2A1O1Ixp33_ASAP7_75t_SL g1474 ( 
.A1(n_1209),
.A2(n_1158),
.B(n_961),
.C(n_1052),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1475)
);

O2A1O1Ixp33_ASAP7_75t_SL g1476 ( 
.A1(n_1209),
.A2(n_1158),
.B(n_961),
.C(n_1052),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1296),
.Y(n_1477)
);

OAI21x1_ASAP7_75t_L g1478 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1478)
);

NAND2x1p5_ASAP7_75t_L g1479 ( 
.A(n_1321),
.B(n_1196),
.Y(n_1479)
);

OAI21x1_ASAP7_75t_L g1480 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1480)
);

AND2x4_ASAP7_75t_L g1481 ( 
.A(n_1251),
.B(n_1196),
.Y(n_1481)
);

CKINVDCx20_ASAP7_75t_R g1482 ( 
.A(n_1195),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1296),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1208),
.Y(n_1484)
);

AO21x2_ASAP7_75t_L g1485 ( 
.A1(n_1297),
.A2(n_1205),
.B(n_1210),
.Y(n_1485)
);

INVx1_ASAP7_75t_L g1486 ( 
.A(n_1208),
.Y(n_1486)
);

AOI22xp5_ASAP7_75t_L g1487 ( 
.A1(n_1332),
.A2(n_961),
.B1(n_607),
.B2(n_978),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1208),
.Y(n_1488)
);

AO31x2_ASAP7_75t_L g1489 ( 
.A1(n_1250),
.A2(n_1263),
.A3(n_1336),
.B(n_1330),
.Y(n_1489)
);

OAI22xp5_ASAP7_75t_L g1490 ( 
.A1(n_1209),
.A2(n_950),
.B1(n_895),
.B2(n_1327),
.Y(n_1490)
);

OAI22xp33_ASAP7_75t_L g1491 ( 
.A1(n_1332),
.A2(n_798),
.B1(n_895),
.B2(n_961),
.Y(n_1491)
);

OAI21x1_ASAP7_75t_L g1492 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1492)
);

OAI22xp5_ASAP7_75t_L g1493 ( 
.A1(n_1209),
.A2(n_950),
.B1(n_895),
.B2(n_1327),
.Y(n_1493)
);

INVx1_ASAP7_75t_L g1494 ( 
.A(n_1208),
.Y(n_1494)
);

INVx1_ASAP7_75t_SL g1495 ( 
.A(n_1304),
.Y(n_1495)
);

AOI21xp5_ASAP7_75t_SL g1496 ( 
.A1(n_1209),
.A2(n_977),
.B(n_895),
.Y(n_1496)
);

OAI21x1_ASAP7_75t_L g1497 ( 
.A1(n_1283),
.A2(n_1329),
.B(n_1202),
.Y(n_1497)
);

AOI21x1_ASAP7_75t_L g1498 ( 
.A1(n_1215),
.A2(n_1224),
.B(n_1287),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1208),
.Y(n_1499)
);

BUFx2_ASAP7_75t_L g1500 ( 
.A(n_1268),
.Y(n_1500)
);

O2A1O1Ixp33_ASAP7_75t_L g1501 ( 
.A1(n_1209),
.A2(n_961),
.B(n_1332),
.C(n_895),
.Y(n_1501)
);

INVx3_ASAP7_75t_L g1502 ( 
.A(n_1411),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1416),
.Y(n_1503)
);

O2A1O1Ixp33_ASAP7_75t_L g1504 ( 
.A1(n_1453),
.A2(n_1462),
.B(n_1491),
.C(n_1474),
.Y(n_1504)
);

NAND2xp5_ASAP7_75t_L g1505 ( 
.A(n_1379),
.B(n_1354),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1463),
.B(n_1357),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1463),
.B(n_1419),
.Y(n_1507)
);

BUFx3_ASAP7_75t_L g1508 ( 
.A(n_1373),
.Y(n_1508)
);

HB1xp67_ASAP7_75t_L g1509 ( 
.A(n_1406),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1352),
.B(n_1485),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1441),
.Y(n_1511)
);

HB1xp67_ASAP7_75t_L g1512 ( 
.A(n_1448),
.Y(n_1512)
);

O2A1O1Ixp33_ASAP7_75t_L g1513 ( 
.A1(n_1474),
.A2(n_1476),
.B(n_1501),
.C(n_1493),
.Y(n_1513)
);

A2O1A1Ixp33_ASAP7_75t_L g1514 ( 
.A1(n_1487),
.A2(n_1490),
.B(n_1377),
.C(n_1399),
.Y(n_1514)
);

INVx1_ASAP7_75t_SL g1515 ( 
.A(n_1356),
.Y(n_1515)
);

OAI22xp5_ASAP7_75t_L g1516 ( 
.A1(n_1367),
.A2(n_1404),
.B1(n_1389),
.B2(n_1392),
.Y(n_1516)
);

AND2x2_ASAP7_75t_L g1517 ( 
.A(n_1352),
.B(n_1485),
.Y(n_1517)
);

OR2x2_ASAP7_75t_L g1518 ( 
.A(n_1355),
.B(n_1495),
.Y(n_1518)
);

NOR2xp67_ASAP7_75t_L g1519 ( 
.A(n_1365),
.B(n_1381),
.Y(n_1519)
);

OA21x2_ASAP7_75t_L g1520 ( 
.A1(n_1435),
.A2(n_1434),
.B(n_1437),
.Y(n_1520)
);

OR2x2_ASAP7_75t_L g1521 ( 
.A(n_1457),
.B(n_1465),
.Y(n_1521)
);

OA21x2_ASAP7_75t_L g1522 ( 
.A1(n_1434),
.A2(n_1437),
.B(n_1388),
.Y(n_1522)
);

OA22x2_ASAP7_75t_L g1523 ( 
.A1(n_1422),
.A2(n_1380),
.B1(n_1420),
.B2(n_1496),
.Y(n_1523)
);

OA21x2_ASAP7_75t_L g1524 ( 
.A1(n_1385),
.A2(n_1366),
.B(n_1396),
.Y(n_1524)
);

NAND2xp5_ASAP7_75t_L g1525 ( 
.A(n_1379),
.B(n_1397),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1470),
.B(n_1376),
.Y(n_1526)
);

CKINVDCx20_ASAP7_75t_R g1527 ( 
.A(n_1482),
.Y(n_1527)
);

OA21x2_ASAP7_75t_L g1528 ( 
.A1(n_1385),
.A2(n_1366),
.B(n_1396),
.Y(n_1528)
);

HB1xp67_ASAP7_75t_L g1529 ( 
.A(n_1412),
.Y(n_1529)
);

BUFx3_ASAP7_75t_L g1530 ( 
.A(n_1500),
.Y(n_1530)
);

NAND2xp5_ASAP7_75t_L g1531 ( 
.A(n_1405),
.B(n_1367),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_1387),
.Y(n_1532)
);

CKINVDCx5p33_ASAP7_75t_R g1533 ( 
.A(n_1387),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1389),
.A2(n_1375),
.B1(n_1399),
.B2(n_1407),
.Y(n_1534)
);

NAND2xp5_ASAP7_75t_L g1535 ( 
.A(n_1351),
.B(n_1395),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1407),
.A2(n_1430),
.B1(n_1377),
.B2(n_1398),
.Y(n_1536)
);

OR2x2_ASAP7_75t_L g1537 ( 
.A(n_1364),
.B(n_1369),
.Y(n_1537)
);

AND2x2_ASAP7_75t_L g1538 ( 
.A(n_1368),
.B(n_1358),
.Y(n_1538)
);

O2A1O1Ixp5_ASAP7_75t_L g1539 ( 
.A1(n_1460),
.A2(n_1413),
.B(n_1431),
.C(n_1408),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1402),
.Y(n_1540)
);

AND2x2_ASAP7_75t_L g1541 ( 
.A(n_1368),
.B(n_1358),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1368),
.B(n_1358),
.Y(n_1542)
);

OAI22xp5_ASAP7_75t_L g1543 ( 
.A1(n_1398),
.A2(n_1423),
.B1(n_1420),
.B2(n_1464),
.Y(n_1543)
);

CKINVDCx5p33_ASAP7_75t_R g1544 ( 
.A(n_1452),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1444),
.B(n_1363),
.Y(n_1545)
);

AOI21xp5_ASAP7_75t_L g1546 ( 
.A1(n_1378),
.A2(n_1363),
.B(n_1476),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1444),
.B(n_1363),
.Y(n_1547)
);

NAND2xp5_ASAP7_75t_L g1548 ( 
.A(n_1351),
.B(n_1371),
.Y(n_1548)
);

NAND2xp5_ASAP7_75t_L g1549 ( 
.A(n_1372),
.B(n_1391),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1442),
.Y(n_1550)
);

OAI22xp5_ASAP7_75t_L g1551 ( 
.A1(n_1420),
.A2(n_1464),
.B1(n_1466),
.B2(n_1414),
.Y(n_1551)
);

OAI22xp5_ASAP7_75t_L g1552 ( 
.A1(n_1359),
.A2(n_1414),
.B1(n_1466),
.B2(n_1436),
.Y(n_1552)
);

OAI22xp5_ASAP7_75t_L g1553 ( 
.A1(n_1359),
.A2(n_1381),
.B1(n_1365),
.B2(n_1415),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1383),
.B(n_1446),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1450),
.Y(n_1555)
);

INVxp67_ASAP7_75t_L g1556 ( 
.A(n_1455),
.Y(n_1556)
);

HB1xp67_ASAP7_75t_L g1557 ( 
.A(n_1458),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1383),
.B(n_1471),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1383),
.B(n_1472),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1484),
.B(n_1486),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1488),
.B(n_1494),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1383),
.B(n_1499),
.Y(n_1562)
);

INVxp67_ASAP7_75t_L g1563 ( 
.A(n_1425),
.Y(n_1563)
);

BUFx2_ASAP7_75t_L g1564 ( 
.A(n_1426),
.Y(n_1564)
);

NOR2xp67_ASAP7_75t_L g1565 ( 
.A(n_1365),
.B(n_1381),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1374),
.B(n_1378),
.Y(n_1566)
);

O2A1O1Ixp5_ASAP7_75t_L g1567 ( 
.A1(n_1498),
.A2(n_1353),
.B(n_1429),
.C(n_1362),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1384),
.Y(n_1568)
);

NAND2x1p5_ASAP7_75t_L g1569 ( 
.A(n_1362),
.B(n_1409),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1374),
.B(n_1400),
.Y(n_1570)
);

OA21x2_ASAP7_75t_L g1571 ( 
.A1(n_1382),
.A2(n_1497),
.B(n_1492),
.Y(n_1571)
);

AOI211xp5_ASAP7_75t_SL g1572 ( 
.A1(n_1350),
.A2(n_1454),
.B(n_1361),
.C(n_1428),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1481),
.B(n_1432),
.Y(n_1573)
);

AND2x4_ASAP7_75t_L g1574 ( 
.A(n_1411),
.B(n_1409),
.Y(n_1574)
);

AND2x2_ASAP7_75t_L g1575 ( 
.A(n_1401),
.B(n_1360),
.Y(n_1575)
);

AND2x2_ASAP7_75t_L g1576 ( 
.A(n_1401),
.B(n_1360),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1433),
.B(n_1427),
.Y(n_1577)
);

BUFx4f_ASAP7_75t_SL g1578 ( 
.A(n_1452),
.Y(n_1578)
);

OA21x2_ASAP7_75t_L g1579 ( 
.A1(n_1440),
.A2(n_1497),
.B(n_1492),
.Y(n_1579)
);

CKINVDCx11_ASAP7_75t_R g1580 ( 
.A(n_1482),
.Y(n_1580)
);

O2A1O1Ixp33_ASAP7_75t_L g1581 ( 
.A1(n_1424),
.A2(n_1403),
.B(n_1390),
.C(n_1445),
.Y(n_1581)
);

BUFx3_ASAP7_75t_L g1582 ( 
.A(n_1418),
.Y(n_1582)
);

INVx3_ASAP7_75t_SL g1583 ( 
.A(n_1418),
.Y(n_1583)
);

O2A1O1Ixp5_ASAP7_75t_L g1584 ( 
.A1(n_1362),
.A2(n_1349),
.B(n_1483),
.C(n_1477),
.Y(n_1584)
);

NAND2xp5_ASAP7_75t_L g1585 ( 
.A(n_1427),
.B(n_1350),
.Y(n_1585)
);

OAI22xp5_ASAP7_75t_L g1586 ( 
.A1(n_1445),
.A2(n_1479),
.B1(n_1361),
.B2(n_1350),
.Y(n_1586)
);

AOI221xp5_ASAP7_75t_L g1587 ( 
.A1(n_1394),
.A2(n_1447),
.B1(n_1468),
.B2(n_1467),
.C(n_1449),
.Y(n_1587)
);

AOI22xp5_ASAP7_75t_L g1588 ( 
.A1(n_1451),
.A2(n_1438),
.B1(n_1410),
.B2(n_1418),
.Y(n_1588)
);

OAI211xp5_ASAP7_75t_L g1589 ( 
.A1(n_1417),
.A2(n_1438),
.B(n_1468),
.C(n_1467),
.Y(n_1589)
);

OA21x2_ASAP7_75t_L g1590 ( 
.A1(n_1440),
.A2(n_1459),
.B(n_1480),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1438),
.B(n_1451),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1451),
.B(n_1421),
.Y(n_1592)
);

AND2x2_ASAP7_75t_L g1593 ( 
.A(n_1439),
.B(n_1489),
.Y(n_1593)
);

INVx2_ASAP7_75t_L g1594 ( 
.A(n_1439),
.Y(n_1594)
);

AND2x2_ASAP7_75t_L g1595 ( 
.A(n_1386),
.B(n_1469),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1421),
.Y(n_1596)
);

AOI21xp5_ASAP7_75t_SL g1597 ( 
.A1(n_1421),
.A2(n_1443),
.B(n_1456),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1443),
.B(n_1469),
.Y(n_1598)
);

OA22x2_ASAP7_75t_L g1599 ( 
.A1(n_1461),
.A2(n_1473),
.B1(n_1475),
.B2(n_1478),
.Y(n_1599)
);

OA21x2_ASAP7_75t_L g1600 ( 
.A1(n_1480),
.A2(n_1478),
.B(n_1421),
.Y(n_1600)
);

NAND2xp5_ASAP7_75t_L g1601 ( 
.A(n_1379),
.B(n_1354),
.Y(n_1601)
);

INVx1_ASAP7_75t_L g1602 ( 
.A(n_1416),
.Y(n_1602)
);

AND2x4_ASAP7_75t_L g1603 ( 
.A(n_1370),
.B(n_1393),
.Y(n_1603)
);

INVx2_ASAP7_75t_SL g1604 ( 
.A(n_1359),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1451),
.Y(n_1605)
);

NOR2xp67_ASAP7_75t_L g1606 ( 
.A(n_1365),
.B(n_1051),
.Y(n_1606)
);

HB1xp67_ASAP7_75t_L g1607 ( 
.A(n_1406),
.Y(n_1607)
);

OA21x2_ASAP7_75t_L g1608 ( 
.A1(n_1435),
.A2(n_1434),
.B(n_1437),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1463),
.B(n_1357),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1463),
.B(n_1357),
.Y(n_1610)
);

OAI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1487),
.A2(n_950),
.B1(n_923),
.B2(n_1209),
.Y(n_1611)
);

AND2x2_ASAP7_75t_L g1612 ( 
.A(n_1510),
.B(n_1517),
.Y(n_1612)
);

OR2x6_ASAP7_75t_L g1613 ( 
.A(n_1546),
.B(n_1597),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1554),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1554),
.Y(n_1615)
);

INVx1_ASAP7_75t_L g1616 ( 
.A(n_1558),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1510),
.B(n_1517),
.Y(n_1617)
);

CKINVDCx5p33_ASAP7_75t_R g1618 ( 
.A(n_1580),
.Y(n_1618)
);

INVx1_ASAP7_75t_L g1619 ( 
.A(n_1558),
.Y(n_1619)
);

NOR2xp67_ASAP7_75t_SL g1620 ( 
.A(n_1568),
.B(n_1544),
.Y(n_1620)
);

INVx1_ASAP7_75t_L g1621 ( 
.A(n_1559),
.Y(n_1621)
);

OR2x2_ASAP7_75t_L g1622 ( 
.A(n_1562),
.B(n_1503),
.Y(n_1622)
);

AND2x2_ASAP7_75t_L g1623 ( 
.A(n_1507),
.B(n_1506),
.Y(n_1623)
);

AND2x4_ASAP7_75t_L g1624 ( 
.A(n_1574),
.B(n_1502),
.Y(n_1624)
);

INVx1_ASAP7_75t_L g1625 ( 
.A(n_1602),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1539),
.A2(n_1584),
.B(n_1587),
.Y(n_1626)
);

HB1xp67_ASAP7_75t_L g1627 ( 
.A(n_1509),
.Y(n_1627)
);

AOI222xp33_ASAP7_75t_L g1628 ( 
.A1(n_1611),
.A2(n_1609),
.B1(n_1506),
.B2(n_1610),
.C1(n_1514),
.C2(n_1516),
.Y(n_1628)
);

AND2x2_ASAP7_75t_L g1629 ( 
.A(n_1507),
.B(n_1609),
.Y(n_1629)
);

NAND2xp5_ASAP7_75t_L g1630 ( 
.A(n_1610),
.B(n_1525),
.Y(n_1630)
);

NAND2xp5_ASAP7_75t_L g1631 ( 
.A(n_1529),
.B(n_1505),
.Y(n_1631)
);

OR2x2_ASAP7_75t_L g1632 ( 
.A(n_1545),
.B(n_1547),
.Y(n_1632)
);

OAI221xp5_ASAP7_75t_SL g1633 ( 
.A1(n_1514),
.A2(n_1504),
.B1(n_1513),
.B2(n_1531),
.C(n_1601),
.Y(n_1633)
);

OR2x6_ASAP7_75t_L g1634 ( 
.A(n_1523),
.B(n_1574),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1580),
.Y(n_1635)
);

HB1xp67_ASAP7_75t_L g1636 ( 
.A(n_1511),
.Y(n_1636)
);

BUFx2_ASAP7_75t_L g1637 ( 
.A(n_1574),
.Y(n_1637)
);

OR2x2_ASAP7_75t_L g1638 ( 
.A(n_1547),
.B(n_1538),
.Y(n_1638)
);

AOI21x1_ASAP7_75t_L g1639 ( 
.A1(n_1589),
.A2(n_1536),
.B(n_1534),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1541),
.B(n_1542),
.Y(n_1640)
);

OAI21xp33_ASAP7_75t_SL g1641 ( 
.A1(n_1523),
.A2(n_1588),
.B(n_1550),
.Y(n_1641)
);

OA21x2_ASAP7_75t_L g1642 ( 
.A1(n_1575),
.A2(n_1576),
.B(n_1594),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1557),
.Y(n_1643)
);

OR2x6_ASAP7_75t_L g1644 ( 
.A(n_1569),
.B(n_1581),
.Y(n_1644)
);

BUFx6f_ASAP7_75t_L g1645 ( 
.A(n_1569),
.Y(n_1645)
);

INVxp67_ASAP7_75t_L g1646 ( 
.A(n_1512),
.Y(n_1646)
);

AO21x2_ASAP7_75t_L g1647 ( 
.A1(n_1575),
.A2(n_1576),
.B(n_1566),
.Y(n_1647)
);

HB1xp67_ASAP7_75t_L g1648 ( 
.A(n_1607),
.Y(n_1648)
);

AO21x2_ASAP7_75t_L g1649 ( 
.A1(n_1566),
.A2(n_1570),
.B(n_1595),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1551),
.B(n_1570),
.Y(n_1650)
);

AO21x2_ASAP7_75t_L g1651 ( 
.A1(n_1595),
.A2(n_1598),
.B(n_1593),
.Y(n_1651)
);

OR2x2_ASAP7_75t_L g1652 ( 
.A(n_1593),
.B(n_1526),
.Y(n_1652)
);

OR2x2_ASAP7_75t_L g1653 ( 
.A(n_1518),
.B(n_1521),
.Y(n_1653)
);

OAI21x1_ASAP7_75t_L g1654 ( 
.A1(n_1599),
.A2(n_1567),
.B(n_1579),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1564),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1555),
.Y(n_1656)
);

AO21x2_ASAP7_75t_L g1657 ( 
.A1(n_1598),
.A2(n_1543),
.B(n_1560),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1603),
.B(n_1556),
.Y(n_1658)
);

AO21x2_ASAP7_75t_L g1659 ( 
.A1(n_1549),
.A2(n_1561),
.B(n_1548),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1552),
.B(n_1586),
.Y(n_1660)
);

OA21x2_ASAP7_75t_L g1661 ( 
.A1(n_1535),
.A2(n_1585),
.B(n_1537),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1600),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1515),
.B(n_1522),
.Y(n_1663)
);

OA21x2_ASAP7_75t_L g1664 ( 
.A1(n_1563),
.A2(n_1608),
.B(n_1520),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1571),
.Y(n_1665)
);

INVx1_ASAP7_75t_L g1666 ( 
.A(n_1625),
.Y(n_1666)
);

HB1xp67_ASAP7_75t_L g1667 ( 
.A(n_1661),
.Y(n_1667)
);

INVx2_ASAP7_75t_L g1668 ( 
.A(n_1665),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1625),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1661),
.B(n_1522),
.Y(n_1670)
);

BUFx2_ASAP7_75t_L g1671 ( 
.A(n_1642),
.Y(n_1671)
);

AOI221xp5_ASAP7_75t_L g1672 ( 
.A1(n_1633),
.A2(n_1553),
.B1(n_1508),
.B2(n_1530),
.C(n_1540),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1640),
.B(n_1608),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1656),
.Y(n_1674)
);

AND2x2_ASAP7_75t_L g1675 ( 
.A(n_1640),
.B(n_1608),
.Y(n_1675)
);

OR2x2_ASAP7_75t_L g1676 ( 
.A(n_1647),
.B(n_1632),
.Y(n_1676)
);

NAND2xp5_ASAP7_75t_L g1677 ( 
.A(n_1661),
.B(n_1520),
.Y(n_1677)
);

INVx1_ASAP7_75t_SL g1678 ( 
.A(n_1643),
.Y(n_1678)
);

CKINVDCx5p33_ASAP7_75t_R g1679 ( 
.A(n_1618),
.Y(n_1679)
);

AND2x4_ASAP7_75t_SL g1680 ( 
.A(n_1644),
.B(n_1605),
.Y(n_1680)
);

INVx3_ASAP7_75t_L g1681 ( 
.A(n_1624),
.Y(n_1681)
);

AOI22xp33_ASAP7_75t_SL g1682 ( 
.A1(n_1628),
.A2(n_1578),
.B1(n_1527),
.B2(n_1532),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1656),
.Y(n_1683)
);

HB1xp67_ASAP7_75t_L g1684 ( 
.A(n_1661),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1654),
.A2(n_1573),
.B(n_1596),
.Y(n_1685)
);

AND2x2_ASAP7_75t_L g1686 ( 
.A(n_1647),
.B(n_1528),
.Y(n_1686)
);

AND2x2_ASAP7_75t_SL g1687 ( 
.A(n_1626),
.B(n_1664),
.Y(n_1687)
);

AND2x2_ASAP7_75t_L g1688 ( 
.A(n_1647),
.B(n_1528),
.Y(n_1688)
);

NAND2xp5_ASAP7_75t_L g1689 ( 
.A(n_1659),
.B(n_1524),
.Y(n_1689)
);

OR2x2_ASAP7_75t_L g1690 ( 
.A(n_1647),
.B(n_1524),
.Y(n_1690)
);

OR2x2_ASAP7_75t_L g1691 ( 
.A(n_1632),
.B(n_1524),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1628),
.B(n_1604),
.Y(n_1692)
);

OR2x2_ASAP7_75t_L g1693 ( 
.A(n_1638),
.B(n_1571),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1651),
.B(n_1612),
.Y(n_1694)
);

OAI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1639),
.A2(n_1527),
.B1(n_1508),
.B2(n_1530),
.Y(n_1695)
);

AND2x2_ASAP7_75t_L g1696 ( 
.A(n_1651),
.B(n_1571),
.Y(n_1696)
);

BUFx2_ASAP7_75t_L g1697 ( 
.A(n_1642),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1659),
.B(n_1572),
.Y(n_1698)
);

AOI21xp5_ASAP7_75t_L g1699 ( 
.A1(n_1613),
.A2(n_1579),
.B(n_1590),
.Y(n_1699)
);

AND2x2_ASAP7_75t_L g1700 ( 
.A(n_1651),
.B(n_1579),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1612),
.B(n_1590),
.Y(n_1701)
);

AND2x2_ASAP7_75t_L g1702 ( 
.A(n_1617),
.B(n_1577),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1649),
.B(n_1604),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1674),
.Y(n_1704)
);

BUFx2_ASAP7_75t_L g1705 ( 
.A(n_1681),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1674),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1681),
.B(n_1624),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1683),
.Y(n_1708)
);

AOI211xp5_ASAP7_75t_L g1709 ( 
.A1(n_1695),
.A2(n_1641),
.B(n_1620),
.C(n_1630),
.Y(n_1709)
);

AND2x4_ASAP7_75t_L g1710 ( 
.A(n_1681),
.B(n_1624),
.Y(n_1710)
);

OA222x2_ASAP7_75t_L g1711 ( 
.A1(n_1698),
.A2(n_1644),
.B1(n_1613),
.B2(n_1634),
.C1(n_1650),
.C2(n_1655),
.Y(n_1711)
);

BUFx2_ASAP7_75t_L g1712 ( 
.A(n_1703),
.Y(n_1712)
);

OAI33xp33_ASAP7_75t_L g1713 ( 
.A1(n_1698),
.A2(n_1630),
.A3(n_1646),
.B1(n_1631),
.B2(n_1652),
.B3(n_1658),
.Y(n_1713)
);

INVx2_ASAP7_75t_L g1714 ( 
.A(n_1671),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1676),
.B(n_1638),
.Y(n_1715)
);

OAI221xp5_ASAP7_75t_L g1716 ( 
.A1(n_1682),
.A2(n_1641),
.B1(n_1660),
.B2(n_1620),
.C(n_1639),
.Y(n_1716)
);

INVx3_ASAP7_75t_L g1717 ( 
.A(n_1681),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1683),
.Y(n_1718)
);

NAND3xp33_ASAP7_75t_L g1719 ( 
.A(n_1682),
.B(n_1660),
.C(n_1644),
.Y(n_1719)
);

AOI22xp5_ASAP7_75t_L g1720 ( 
.A1(n_1695),
.A2(n_1644),
.B1(n_1635),
.B2(n_1634),
.Y(n_1720)
);

OAI211xp5_ASAP7_75t_L g1721 ( 
.A1(n_1692),
.A2(n_1658),
.B(n_1627),
.C(n_1636),
.Y(n_1721)
);

OA21x2_ASAP7_75t_L g1722 ( 
.A1(n_1699),
.A2(n_1654),
.B(n_1662),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1671),
.B(n_1644),
.Y(n_1723)
);

AOI22xp5_ASAP7_75t_L g1724 ( 
.A1(n_1692),
.A2(n_1634),
.B1(n_1629),
.B2(n_1623),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1671),
.Y(n_1725)
);

INVx2_ASAP7_75t_L g1726 ( 
.A(n_1697),
.Y(n_1726)
);

BUFx3_ASAP7_75t_L g1727 ( 
.A(n_1679),
.Y(n_1727)
);

OAI221xp5_ASAP7_75t_L g1728 ( 
.A1(n_1672),
.A2(n_1653),
.B1(n_1634),
.B2(n_1648),
.C(n_1606),
.Y(n_1728)
);

AOI221xp5_ASAP7_75t_L g1729 ( 
.A1(n_1672),
.A2(n_1623),
.B1(n_1629),
.B2(n_1643),
.C(n_1614),
.Y(n_1729)
);

AO21x1_ASAP7_75t_SL g1730 ( 
.A1(n_1676),
.A2(n_1616),
.B(n_1621),
.Y(n_1730)
);

OAI22xp5_ASAP7_75t_L g1731 ( 
.A1(n_1680),
.A2(n_1634),
.B1(n_1653),
.B2(n_1650),
.Y(n_1731)
);

AOI22xp33_ASAP7_75t_L g1732 ( 
.A1(n_1687),
.A2(n_1626),
.B1(n_1657),
.B2(n_1650),
.Y(n_1732)
);

BUFx3_ASAP7_75t_L g1733 ( 
.A(n_1679),
.Y(n_1733)
);

NOR4xp25_ASAP7_75t_SL g1734 ( 
.A(n_1697),
.B(n_1533),
.C(n_1532),
.D(n_1544),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1666),
.Y(n_1735)
);

AOI221xp5_ASAP7_75t_L g1736 ( 
.A1(n_1694),
.A2(n_1678),
.B1(n_1703),
.B2(n_1667),
.C(n_1684),
.Y(n_1736)
);

OAI221xp5_ASAP7_75t_L g1737 ( 
.A1(n_1678),
.A2(n_1650),
.B1(n_1533),
.B2(n_1613),
.C(n_1519),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1666),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1694),
.B(n_1637),
.Y(n_1739)
);

HB1xp67_ASAP7_75t_L g1740 ( 
.A(n_1703),
.Y(n_1740)
);

AOI22xp33_ASAP7_75t_SL g1741 ( 
.A1(n_1680),
.A2(n_1650),
.B1(n_1657),
.B2(n_1626),
.Y(n_1741)
);

AND2x2_ASAP7_75t_L g1742 ( 
.A(n_1694),
.B(n_1681),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1702),
.B(n_1657),
.Y(n_1743)
);

INVx1_ASAP7_75t_SL g1744 ( 
.A(n_1702),
.Y(n_1744)
);

HB1xp67_ASAP7_75t_L g1745 ( 
.A(n_1685),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1697),
.Y(n_1746)
);

INVxp67_ASAP7_75t_L g1747 ( 
.A(n_1702),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1673),
.B(n_1659),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1668),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1667),
.A2(n_1616),
.B1(n_1621),
.B2(n_1615),
.C(n_1619),
.Y(n_1750)
);

HB1xp67_ASAP7_75t_L g1751 ( 
.A(n_1685),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1673),
.B(n_1637),
.Y(n_1752)
);

NAND3xp33_ASAP7_75t_L g1753 ( 
.A(n_1687),
.B(n_1645),
.C(n_1663),
.Y(n_1753)
);

OAI221xp5_ASAP7_75t_L g1754 ( 
.A1(n_1676),
.A2(n_1613),
.B1(n_1565),
.B2(n_1652),
.C(n_1684),
.Y(n_1754)
);

AOI211xp5_ASAP7_75t_SL g1755 ( 
.A1(n_1699),
.A2(n_1663),
.B(n_1592),
.C(n_1622),
.Y(n_1755)
);

OR2x6_ASAP7_75t_L g1756 ( 
.A(n_1691),
.B(n_1613),
.Y(n_1756)
);

INVx3_ASAP7_75t_L g1757 ( 
.A(n_1707),
.Y(n_1757)
);

NOR2xp33_ASAP7_75t_SL g1758 ( 
.A(n_1716),
.B(n_1680),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1704),
.Y(n_1759)
);

INVx2_ASAP7_75t_L g1760 ( 
.A(n_1714),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1706),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1723),
.Y(n_1762)
);

BUFx12f_ASAP7_75t_L g1763 ( 
.A(n_1727),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1742),
.B(n_1673),
.Y(n_1764)
);

OA21x2_ASAP7_75t_L g1765 ( 
.A1(n_1732),
.A2(n_1670),
.B(n_1677),
.Y(n_1765)
);

NAND2xp5_ASAP7_75t_SL g1766 ( 
.A(n_1709),
.B(n_1645),
.Y(n_1766)
);

INVx2_ASAP7_75t_L g1767 ( 
.A(n_1714),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1708),
.Y(n_1768)
);

HB1xp67_ASAP7_75t_L g1769 ( 
.A(n_1745),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1715),
.B(n_1748),
.Y(n_1770)
);

HB1xp67_ASAP7_75t_L g1771 ( 
.A(n_1751),
.Y(n_1771)
);

INVx1_ASAP7_75t_SL g1772 ( 
.A(n_1705),
.Y(n_1772)
);

INVx4_ASAP7_75t_L g1773 ( 
.A(n_1727),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_SL g1774 ( 
.A(n_1721),
.B(n_1696),
.C(n_1700),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1742),
.B(n_1675),
.Y(n_1775)
);

OR2x2_ASAP7_75t_L g1776 ( 
.A(n_1715),
.B(n_1691),
.Y(n_1776)
);

AND2x2_ASAP7_75t_L g1777 ( 
.A(n_1712),
.B(n_1675),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1740),
.B(n_1730),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1705),
.B(n_1675),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1725),
.Y(n_1780)
);

INVx2_ASAP7_75t_L g1781 ( 
.A(n_1725),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1718),
.Y(n_1782)
);

OR2x2_ASAP7_75t_L g1783 ( 
.A(n_1743),
.B(n_1691),
.Y(n_1783)
);

CKINVDCx5p33_ASAP7_75t_R g1784 ( 
.A(n_1733),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1735),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1719),
.B(n_1645),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1723),
.B(n_1645),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1738),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1749),
.Y(n_1789)
);

OAI21x1_ASAP7_75t_L g1790 ( 
.A1(n_1726),
.A2(n_1670),
.B(n_1677),
.Y(n_1790)
);

INVx2_ASAP7_75t_SL g1791 ( 
.A(n_1717),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1732),
.A2(n_1687),
.B(n_1626),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1747),
.Y(n_1794)
);

OA21x2_ASAP7_75t_L g1795 ( 
.A1(n_1726),
.A2(n_1689),
.B(n_1688),
.Y(n_1795)
);

INVx2_ASAP7_75t_SL g1796 ( 
.A(n_1717),
.Y(n_1796)
);

INVx1_ASAP7_75t_L g1797 ( 
.A(n_1746),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1746),
.Y(n_1798)
);

OR2x2_ASAP7_75t_L g1799 ( 
.A(n_1743),
.B(n_1693),
.Y(n_1799)
);

NAND2xp5_ASAP7_75t_SL g1800 ( 
.A(n_1758),
.B(n_1720),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1790),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1794),
.B(n_1736),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1782),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1762),
.B(n_1711),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1782),
.Y(n_1805)
);

NAND3x1_ASAP7_75t_L g1806 ( 
.A(n_1793),
.B(n_1717),
.C(n_1729),
.Y(n_1806)
);

AND2x4_ASAP7_75t_L g1807 ( 
.A(n_1778),
.B(n_1723),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1766),
.A2(n_1758),
.B1(n_1774),
.B2(n_1786),
.Y(n_1808)
);

NOR3xp33_ASAP7_75t_L g1809 ( 
.A(n_1774),
.B(n_1737),
.C(n_1728),
.Y(n_1809)
);

BUFx2_ASAP7_75t_L g1810 ( 
.A(n_1763),
.Y(n_1810)
);

OAI21xp33_ASAP7_75t_L g1811 ( 
.A1(n_1793),
.A2(n_1741),
.B(n_1724),
.Y(n_1811)
);

OR2x2_ASAP7_75t_L g1812 ( 
.A(n_1783),
.B(n_1693),
.Y(n_1812)
);

AND2x2_ASAP7_75t_L g1813 ( 
.A(n_1762),
.B(n_1707),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1794),
.B(n_1755),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1773),
.B(n_1744),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1773),
.B(n_1739),
.Y(n_1816)
);

AOI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1787),
.A2(n_1713),
.B(n_1753),
.Y(n_1817)
);

AND2x2_ASAP7_75t_L g1818 ( 
.A(n_1757),
.B(n_1707),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1759),
.Y(n_1819)
);

AND2x2_ASAP7_75t_L g1820 ( 
.A(n_1757),
.B(n_1778),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1821)
);

AOI21xp33_ASAP7_75t_SL g1822 ( 
.A1(n_1784),
.A2(n_1754),
.B(n_1731),
.Y(n_1822)
);

CKINVDCx20_ASAP7_75t_R g1823 ( 
.A(n_1763),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1757),
.B(n_1710),
.Y(n_1824)
);

NOR2xp33_ASAP7_75t_L g1825 ( 
.A(n_1763),
.B(n_1733),
.Y(n_1825)
);

AND2x2_ASAP7_75t_L g1826 ( 
.A(n_1778),
.B(n_1710),
.Y(n_1826)
);

NOR3xp33_ASAP7_75t_L g1827 ( 
.A(n_1773),
.B(n_1591),
.C(n_1750),
.Y(n_1827)
);

INVx1_ASAP7_75t_L g1828 ( 
.A(n_1759),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1773),
.B(n_1739),
.Y(n_1829)
);

OR2x2_ASAP7_75t_L g1830 ( 
.A(n_1783),
.B(n_1693),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1799),
.B(n_1752),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1777),
.B(n_1723),
.Y(n_1832)
);

AOI211xp5_ASAP7_75t_L g1833 ( 
.A1(n_1799),
.A2(n_1696),
.B(n_1700),
.C(n_1686),
.Y(n_1833)
);

NAND3xp33_ASAP7_75t_SL g1834 ( 
.A(n_1772),
.B(n_1734),
.C(n_1690),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1777),
.B(n_1752),
.Y(n_1835)
);

OAI31xp33_ASAP7_75t_L g1836 ( 
.A1(n_1772),
.A2(n_1680),
.A3(n_1700),
.B(n_1696),
.Y(n_1836)
);

HB1xp67_ASAP7_75t_L g1837 ( 
.A(n_1761),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1765),
.B(n_1657),
.Y(n_1838)
);

NAND2xp5_ASAP7_75t_L g1839 ( 
.A(n_1765),
.B(n_1701),
.Y(n_1839)
);

OAI22xp5_ASAP7_75t_SL g1840 ( 
.A1(n_1765),
.A2(n_1787),
.B1(n_1687),
.B2(n_1756),
.Y(n_1840)
);

INVx1_ASAP7_75t_L g1841 ( 
.A(n_1761),
.Y(n_1841)
);

OR2x2_ASAP7_75t_L g1842 ( 
.A(n_1770),
.B(n_1776),
.Y(n_1842)
);

NAND3xp33_ASAP7_75t_L g1843 ( 
.A(n_1765),
.B(n_1756),
.C(n_1685),
.Y(n_1843)
);

AND2x4_ASAP7_75t_L g1844 ( 
.A(n_1807),
.B(n_1787),
.Y(n_1844)
);

NAND2x1_ASAP7_75t_L g1845 ( 
.A(n_1807),
.B(n_1791),
.Y(n_1845)
);

INVx2_ASAP7_75t_L g1846 ( 
.A(n_1820),
.Y(n_1846)
);

NOR2xp33_ASAP7_75t_L g1847 ( 
.A(n_1823),
.B(n_1768),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1827),
.B(n_1768),
.Y(n_1848)
);

INVx2_ASAP7_75t_L g1849 ( 
.A(n_1820),
.Y(n_1849)
);

INVx1_ASAP7_75t_L g1850 ( 
.A(n_1837),
.Y(n_1850)
);

INVx1_ASAP7_75t_L g1851 ( 
.A(n_1828),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1828),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1841),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1813),
.B(n_1764),
.Y(n_1854)
);

INVx1_ASAP7_75t_SL g1855 ( 
.A(n_1823),
.Y(n_1855)
);

OR2x2_ASAP7_75t_L g1856 ( 
.A(n_1802),
.B(n_1770),
.Y(n_1856)
);

NOR2x1p5_ASAP7_75t_L g1857 ( 
.A(n_1814),
.B(n_1776),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1841),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1831),
.B(n_1765),
.Y(n_1859)
);

OAI21xp33_ASAP7_75t_SL g1860 ( 
.A1(n_1808),
.A2(n_1800),
.B(n_1804),
.Y(n_1860)
);

NAND2xp5_ASAP7_75t_L g1861 ( 
.A(n_1809),
.B(n_1785),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1810),
.B(n_1785),
.Y(n_1862)
);

AND2x4_ASAP7_75t_L g1863 ( 
.A(n_1807),
.B(n_1787),
.Y(n_1863)
);

NAND2xp5_ASAP7_75t_L g1864 ( 
.A(n_1810),
.B(n_1788),
.Y(n_1864)
);

OR2x2_ASAP7_75t_L g1865 ( 
.A(n_1816),
.B(n_1788),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1819),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1817),
.B(n_1764),
.Y(n_1867)
);

NOR2xp33_ASAP7_75t_L g1868 ( 
.A(n_1825),
.B(n_1822),
.Y(n_1868)
);

AND2x4_ASAP7_75t_L g1869 ( 
.A(n_1826),
.B(n_1787),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1805),
.Y(n_1870)
);

OR2x2_ASAP7_75t_L g1871 ( 
.A(n_1829),
.B(n_1797),
.Y(n_1871)
);

NAND2xp5_ASAP7_75t_L g1872 ( 
.A(n_1811),
.B(n_1804),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1805),
.Y(n_1873)
);

OR2x2_ASAP7_75t_L g1874 ( 
.A(n_1842),
.B(n_1797),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1803),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1815),
.B(n_1764),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1813),
.B(n_1775),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1835),
.B(n_1775),
.Y(n_1878)
);

AND2x2_ASAP7_75t_L g1879 ( 
.A(n_1826),
.B(n_1775),
.Y(n_1879)
);

AND2x2_ASAP7_75t_L g1880 ( 
.A(n_1818),
.B(n_1779),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1851),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_SL g1882 ( 
.A(n_1860),
.B(n_1836),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_L g1883 ( 
.A(n_1850),
.B(n_1835),
.Y(n_1883)
);

OAI21x1_ASAP7_75t_L g1884 ( 
.A1(n_1845),
.A2(n_1806),
.B(n_1838),
.Y(n_1884)
);

INVx2_ASAP7_75t_L g1885 ( 
.A(n_1846),
.Y(n_1885)
);

NAND2xp5_ASAP7_75t_L g1886 ( 
.A(n_1861),
.B(n_1806),
.Y(n_1886)
);

AOI22xp33_ASAP7_75t_L g1887 ( 
.A1(n_1868),
.A2(n_1840),
.B1(n_1834),
.B2(n_1843),
.Y(n_1887)
);

OA21x2_ASAP7_75t_L g1888 ( 
.A1(n_1872),
.A2(n_1801),
.B(n_1839),
.Y(n_1888)
);

HB1xp67_ASAP7_75t_L g1889 ( 
.A(n_1846),
.Y(n_1889)
);

INVx2_ASAP7_75t_L g1890 ( 
.A(n_1849),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1849),
.Y(n_1891)
);

NOR2xp67_ASAP7_75t_L g1892 ( 
.A(n_1844),
.B(n_1832),
.Y(n_1892)
);

NAND2xp5_ASAP7_75t_L g1893 ( 
.A(n_1875),
.B(n_1833),
.Y(n_1893)
);

AND2x2_ASAP7_75t_L g1894 ( 
.A(n_1879),
.B(n_1818),
.Y(n_1894)
);

AO21x2_ASAP7_75t_L g1895 ( 
.A1(n_1867),
.A2(n_1801),
.B(n_1769),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1870),
.B(n_1798),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1880),
.Y(n_1897)
);

AND2x4_ASAP7_75t_L g1898 ( 
.A(n_1844),
.B(n_1832),
.Y(n_1898)
);

NOR2x1_ASAP7_75t_L g1899 ( 
.A(n_1855),
.B(n_1868),
.Y(n_1899)
);

INVxp67_ASAP7_75t_L g1900 ( 
.A(n_1847),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1852),
.Y(n_1901)
);

INVxp67_ASAP7_75t_SL g1902 ( 
.A(n_1847),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1853),
.Y(n_1903)
);

AND2x4_ASAP7_75t_L g1904 ( 
.A(n_1844),
.B(n_1821),
.Y(n_1904)
);

AOI22xp33_ASAP7_75t_SL g1905 ( 
.A1(n_1848),
.A2(n_1771),
.B1(n_1769),
.B2(n_1795),
.Y(n_1905)
);

HB1xp67_ASAP7_75t_L g1906 ( 
.A(n_1857),
.Y(n_1906)
);

NAND2xp5_ASAP7_75t_L g1907 ( 
.A(n_1902),
.B(n_1862),
.Y(n_1907)
);

AOI22xp5_ASAP7_75t_L g1908 ( 
.A1(n_1899),
.A2(n_1864),
.B1(n_1856),
.B2(n_1873),
.Y(n_1908)
);

AOI322xp5_ASAP7_75t_L g1909 ( 
.A1(n_1899),
.A2(n_1877),
.A3(n_1854),
.B1(n_1878),
.B2(n_1879),
.C1(n_1880),
.C2(n_1876),
.Y(n_1909)
);

OR2x2_ASAP7_75t_L g1910 ( 
.A(n_1902),
.B(n_1865),
.Y(n_1910)
);

OR2x2_ASAP7_75t_L g1911 ( 
.A(n_1900),
.B(n_1871),
.Y(n_1911)
);

CKINVDCx16_ASAP7_75t_R g1912 ( 
.A(n_1906),
.Y(n_1912)
);

AOI22xp33_ASAP7_75t_L g1913 ( 
.A1(n_1882),
.A2(n_1863),
.B1(n_1869),
.B2(n_1859),
.Y(n_1913)
);

AOI221xp5_ASAP7_75t_L g1914 ( 
.A1(n_1886),
.A2(n_1866),
.B1(n_1863),
.B2(n_1858),
.C(n_1869),
.Y(n_1914)
);

INVx1_ASAP7_75t_L g1915 ( 
.A(n_1891),
.Y(n_1915)
);

AOI221xp5_ASAP7_75t_L g1916 ( 
.A1(n_1886),
.A2(n_1863),
.B1(n_1869),
.B2(n_1874),
.C(n_1771),
.Y(n_1916)
);

INVx2_ASAP7_75t_L g1917 ( 
.A(n_1904),
.Y(n_1917)
);

NAND4xp25_ASAP7_75t_L g1918 ( 
.A(n_1887),
.B(n_1842),
.C(n_1821),
.D(n_1824),
.Y(n_1918)
);

OAI32xp33_ASAP7_75t_L g1919 ( 
.A1(n_1893),
.A2(n_1830),
.A3(n_1812),
.B1(n_1824),
.B2(n_1690),
.Y(n_1919)
);

AOI21xp5_ASAP7_75t_L g1920 ( 
.A1(n_1900),
.A2(n_1787),
.B(n_1791),
.Y(n_1920)
);

INVx2_ASAP7_75t_L g1921 ( 
.A(n_1904),
.Y(n_1921)
);

INVx2_ASAP7_75t_SL g1922 ( 
.A(n_1904),
.Y(n_1922)
);

OAI21xp33_ASAP7_75t_SL g1923 ( 
.A1(n_1884),
.A2(n_1796),
.B(n_1791),
.Y(n_1923)
);

INVx1_ASAP7_75t_L g1924 ( 
.A(n_1891),
.Y(n_1924)
);

OAI221xp5_ASAP7_75t_L g1925 ( 
.A1(n_1905),
.A2(n_1830),
.B1(n_1812),
.B2(n_1756),
.C(n_1796),
.Y(n_1925)
);

INVx2_ASAP7_75t_SL g1926 ( 
.A(n_1904),
.Y(n_1926)
);

OR2x2_ASAP7_75t_L g1927 ( 
.A(n_1883),
.B(n_1760),
.Y(n_1927)
);

OR2x2_ASAP7_75t_L g1928 ( 
.A(n_1912),
.B(n_1883),
.Y(n_1928)
);

NAND2xp5_ASAP7_75t_SL g1929 ( 
.A(n_1908),
.B(n_1892),
.Y(n_1929)
);

NAND2xp33_ASAP7_75t_L g1930 ( 
.A(n_1910),
.B(n_1897),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1907),
.B(n_1897),
.Y(n_1931)
);

NOR2xp33_ASAP7_75t_L g1932 ( 
.A(n_1911),
.B(n_1898),
.Y(n_1932)
);

INVx1_ASAP7_75t_L g1933 ( 
.A(n_1915),
.Y(n_1933)
);

NAND2x1p5_ASAP7_75t_L g1934 ( 
.A(n_1922),
.B(n_1892),
.Y(n_1934)
);

NAND2xp5_ASAP7_75t_L g1935 ( 
.A(n_1924),
.B(n_1889),
.Y(n_1935)
);

AND2x2_ASAP7_75t_L g1936 ( 
.A(n_1926),
.B(n_1898),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1917),
.Y(n_1937)
);

NOR2xp33_ASAP7_75t_L g1938 ( 
.A(n_1918),
.B(n_1898),
.Y(n_1938)
);

AND2x2_ASAP7_75t_L g1939 ( 
.A(n_1921),
.B(n_1898),
.Y(n_1939)
);

NAND4xp25_ASAP7_75t_L g1940 ( 
.A(n_1938),
.B(n_1913),
.C(n_1914),
.D(n_1916),
.Y(n_1940)
);

OAI22xp33_ASAP7_75t_L g1941 ( 
.A1(n_1929),
.A2(n_1908),
.B1(n_1893),
.B2(n_1925),
.Y(n_1941)
);

NAND4xp25_ASAP7_75t_SL g1942 ( 
.A(n_1928),
.B(n_1909),
.C(n_1905),
.D(n_1923),
.Y(n_1942)
);

OAI22xp33_ASAP7_75t_L g1943 ( 
.A1(n_1934),
.A2(n_1897),
.B1(n_1888),
.B2(n_1920),
.Y(n_1943)
);

AOI22xp5_ASAP7_75t_L g1944 ( 
.A1(n_1932),
.A2(n_1884),
.B1(n_1888),
.B2(n_1923),
.Y(n_1944)
);

NOR3xp33_ASAP7_75t_L g1945 ( 
.A(n_1930),
.B(n_1884),
.C(n_1903),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1933),
.A2(n_1919),
.B1(n_1881),
.B2(n_1903),
.C(n_1901),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1936),
.B(n_1894),
.Y(n_1947)
);

AOI211xp5_ASAP7_75t_L g1948 ( 
.A1(n_1939),
.A2(n_1901),
.B(n_1881),
.C(n_1890),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_SL g1949 ( 
.A(n_1931),
.B(n_1927),
.Y(n_1949)
);

AOI211xp5_ASAP7_75t_L g1950 ( 
.A1(n_1937),
.A2(n_1890),
.B(n_1885),
.C(n_1894),
.Y(n_1950)
);

O2A1O1Ixp33_ASAP7_75t_L g1951 ( 
.A1(n_1945),
.A2(n_1935),
.B(n_1895),
.C(n_1888),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1947),
.Y(n_1952)
);

OAI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1944),
.A2(n_1941),
.B1(n_1935),
.B2(n_1946),
.Y(n_1953)
);

OAI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1942),
.A2(n_1940),
.B(n_1949),
.Y(n_1954)
);

A2O1A1Ixp33_ASAP7_75t_L g1955 ( 
.A1(n_1950),
.A2(n_1890),
.B(n_1885),
.C(n_1896),
.Y(n_1955)
);

AOI22xp5_ASAP7_75t_L g1956 ( 
.A1(n_1943),
.A2(n_1888),
.B1(n_1885),
.B2(n_1895),
.Y(n_1956)
);

AOI21xp33_ASAP7_75t_R g1957 ( 
.A1(n_1948),
.A2(n_1896),
.B(n_1888),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1952),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1954),
.B(n_1895),
.Y(n_1959)
);

XOR2x2_ASAP7_75t_L g1960 ( 
.A(n_1953),
.B(n_1895),
.Y(n_1960)
);

AND2x2_ASAP7_75t_L g1961 ( 
.A(n_1955),
.B(n_1779),
.Y(n_1961)
);

AND2x2_ASAP7_75t_L g1962 ( 
.A(n_1956),
.B(n_1779),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1951),
.Y(n_1963)
);

OAI221xp5_ASAP7_75t_L g1964 ( 
.A1(n_1957),
.A2(n_1796),
.B1(n_1760),
.B2(n_1767),
.C(n_1781),
.Y(n_1964)
);

OAI221xp5_ASAP7_75t_L g1965 ( 
.A1(n_1959),
.A2(n_1767),
.B1(n_1760),
.B2(n_1780),
.C(n_1781),
.Y(n_1965)
);

AND2x2_ASAP7_75t_L g1966 ( 
.A(n_1961),
.B(n_1777),
.Y(n_1966)
);

NAND2xp33_ASAP7_75t_SL g1967 ( 
.A(n_1959),
.B(n_1583),
.Y(n_1967)
);

NAND3xp33_ASAP7_75t_L g1968 ( 
.A(n_1963),
.B(n_1798),
.C(n_1780),
.Y(n_1968)
);

INVx3_ASAP7_75t_SL g1969 ( 
.A(n_1958),
.Y(n_1969)
);

OAI21xp33_ASAP7_75t_L g1970 ( 
.A1(n_1962),
.A2(n_1780),
.B(n_1781),
.Y(n_1970)
);

AOI21xp33_ASAP7_75t_SL g1971 ( 
.A1(n_1969),
.A2(n_1960),
.B(n_1964),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1966),
.Y(n_1972)
);

NAND4xp75_ASAP7_75t_L g1973 ( 
.A(n_1967),
.B(n_1795),
.C(n_1767),
.D(n_1722),
.Y(n_1973)
);

AND3x4_ASAP7_75t_L g1974 ( 
.A(n_1971),
.B(n_1968),
.C(n_1970),
.Y(n_1974)
);

AOI22xp33_ASAP7_75t_L g1975 ( 
.A1(n_1974),
.A2(n_1972),
.B1(n_1965),
.B2(n_1973),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1975),
.A2(n_1792),
.B1(n_1789),
.B2(n_1795),
.Y(n_1976)
);

INVx4_ASAP7_75t_L g1977 ( 
.A(n_1975),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1977),
.Y(n_1978)
);

INVx2_ASAP7_75t_L g1979 ( 
.A(n_1976),
.Y(n_1979)
);

OAI22xp5_ASAP7_75t_L g1980 ( 
.A1(n_1978),
.A2(n_1792),
.B1(n_1789),
.B2(n_1795),
.Y(n_1980)
);

AOI22xp5_ASAP7_75t_L g1981 ( 
.A1(n_1979),
.A2(n_1795),
.B1(n_1583),
.B2(n_1790),
.Y(n_1981)
);

BUFx2_ASAP7_75t_L g1982 ( 
.A(n_1981),
.Y(n_1982)
);

AOI21xp5_ASAP7_75t_L g1983 ( 
.A1(n_1982),
.A2(n_1980),
.B(n_1790),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_L g1984 ( 
.A(n_1983),
.B(n_1582),
.Y(n_1984)
);

NAND3xp33_ASAP7_75t_L g1985 ( 
.A(n_1984),
.B(n_1605),
.C(n_1582),
.Y(n_1985)
);

AOI221xp5_ASAP7_75t_L g1986 ( 
.A1(n_1985),
.A2(n_1605),
.B1(n_1645),
.B2(n_1669),
.C(n_1689),
.Y(n_1986)
);

AOI211xp5_ASAP7_75t_L g1987 ( 
.A1(n_1986),
.A2(n_1605),
.B(n_1645),
.C(n_1690),
.Y(n_1987)
);


endmodule