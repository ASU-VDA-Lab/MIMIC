module real_aes_411_n_335 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_14, n_194, n_137, n_225, n_16, n_39, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_335);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_335;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_887;
wire n_436;
wire n_684;
wire n_390;
wire n_821;
wire n_830;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_635;
wire n_357;
wire n_792;
wire n_673;
wire n_386;
wire n_503;
wire n_518;
wire n_905;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_900;
wire n_718;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_364;
wire n_421;
wire n_555;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_353;
wire n_431;
wire n_865;
wire n_666;
wire n_884;
wire n_537;
wire n_551;
wire n_560;
wire n_660;
wire n_814;
wire n_886;
wire n_856;
wire n_594;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_786;
wire n_388;
wire n_512;
wire n_395;
wire n_795;
wire n_626;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_462;
wire n_615;
wire n_550;
wire n_670;
wire n_818;
wire n_716;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_774;
wire n_813;
wire n_791;
wire n_559;
wire n_466;
wire n_636;
wire n_872;
wire n_906;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_801;
wire n_383;
wire n_529;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_659;
wire n_547;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_885;
wire n_381;
wire n_493;
wire n_664;
wire n_367;
wire n_819;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_609;
wire n_425;
wire n_879;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_783;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_617;
wire n_402;
wire n_552;
wire n_602;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_642;
wire n_613;
wire n_869;
wire n_387;
wire n_702;
wire n_912;
wire n_464;
wire n_351;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_358;
wire n_385;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_851;
wire n_470;
wire n_915;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_927;
wire n_723;
wire n_662;
wire n_382;
wire n_845;
wire n_850;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_907;
wire n_847;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_365;
wire n_526;
wire n_637;
wire n_899;
wire n_928;
wire n_692;
wire n_544;
wire n_789;
wire n_389;
wire n_738;
wire n_701;
wire n_344;
wire n_827;
wire n_809;
wire n_922;
wire n_482;
wire n_520;
wire n_633;
wire n_926;
wire n_679;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_741;
wire n_753;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_456;
wire n_359;
wire n_717;
wire n_712;
wire n_433;
wire n_516;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_583;
wire n_347;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_614;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_473;
wire n_465;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_640;
wire n_340;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_652;
wire n_703;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_0), .A2(n_203), .B1(n_610), .B2(n_673), .Y(n_672) );
AOI22xp5_ASAP7_75t_L g838 ( .A1(n_1), .A2(n_271), .B1(n_477), .B2(n_481), .Y(n_838) );
AOI22xp33_ASAP7_75t_L g634 ( .A1(n_2), .A2(n_53), .B1(n_418), .B2(n_635), .Y(n_634) );
AOI22xp5_ASAP7_75t_L g486 ( .A1(n_3), .A2(n_103), .B1(n_487), .B2(n_490), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g921 ( .A1(n_4), .A2(n_113), .B1(n_828), .B2(n_922), .Y(n_921) );
CKINVDCx20_ASAP7_75t_R g547 ( .A(n_5), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g790 ( .A(n_6), .Y(n_790) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_7), .A2(n_222), .B1(n_532), .B2(n_533), .Y(n_531) );
CKINVDCx20_ASAP7_75t_R g701 ( .A(n_8), .Y(n_701) );
CKINVDCx20_ASAP7_75t_R g837 ( .A(n_9), .Y(n_837) );
AOI22xp33_ASAP7_75t_SL g916 ( .A1(n_10), .A2(n_302), .B1(n_514), .B2(n_917), .Y(n_916) );
AOI22xp33_ASAP7_75t_L g748 ( .A1(n_11), .A2(n_44), .B1(n_446), .B2(n_577), .Y(n_748) );
AOI22xp33_ASAP7_75t_L g665 ( .A1(n_12), .A2(n_182), .B1(n_609), .B2(n_666), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g740 ( .A1(n_13), .A2(n_215), .B1(n_481), .B2(n_510), .Y(n_740) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_14), .A2(n_226), .B1(n_380), .B2(n_635), .Y(n_876) );
AOI22xp33_ASAP7_75t_L g682 ( .A1(n_15), .A2(n_122), .B1(n_418), .B2(n_635), .Y(n_682) );
AOI22xp5_ASAP7_75t_L g632 ( .A1(n_16), .A2(n_165), .B1(n_457), .B2(n_532), .Y(n_632) );
AOI22xp33_ASAP7_75t_L g539 ( .A1(n_17), .A2(n_292), .B1(n_371), .B2(n_375), .Y(n_539) );
AOI22xp33_ASAP7_75t_L g886 ( .A1(n_18), .A2(n_169), .B1(n_453), .B2(n_747), .Y(n_886) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_19), .A2(n_225), .B1(n_371), .B2(n_375), .Y(n_722) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_20), .B(n_472), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g661 ( .A1(n_21), .A2(n_259), .B1(n_662), .B2(n_663), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g741 ( .A1(n_22), .A2(n_195), .B1(n_516), .B2(n_517), .Y(n_741) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_23), .A2(n_125), .B1(n_516), .B2(n_517), .Y(n_515) );
INVx1_ASAP7_75t_SL g360 ( .A(n_24), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g903 ( .A(n_24), .B(n_36), .Y(n_903) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_25), .A2(n_104), .B1(n_386), .B2(n_420), .Y(n_419) );
AOI222xp33_ASAP7_75t_L g639 ( .A1(n_26), .A2(n_274), .B1(n_305), .B2(n_541), .C1(n_640), .C2(n_642), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_27), .B(n_519), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g545 ( .A(n_28), .Y(n_545) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_29), .A2(n_301), .B1(n_572), .B2(n_574), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g801 ( .A1(n_30), .A2(n_32), .B1(n_456), .B2(n_609), .Y(n_801) );
AOI22xp33_ASAP7_75t_L g848 ( .A1(n_31), .A2(n_209), .B1(n_530), .B2(n_849), .Y(n_848) );
AOI22xp5_ASAP7_75t_L g915 ( .A1(n_33), .A2(n_96), .B1(n_820), .B2(n_821), .Y(n_915) );
AOI22xp33_ASAP7_75t_L g749 ( .A1(n_34), .A2(n_88), .B1(n_530), .B2(n_567), .Y(n_749) );
AOI22xp33_ASAP7_75t_L g924 ( .A1(n_35), .A2(n_90), .B1(n_631), .B2(n_825), .Y(n_924) );
AO22x2_ASAP7_75t_L g362 ( .A1(n_36), .A2(n_311), .B1(n_359), .B2(n_363), .Y(n_362) );
AOI22xp33_ASAP7_75t_L g394 ( .A1(n_37), .A2(n_258), .B1(n_395), .B2(n_396), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g528 ( .A1(n_38), .A2(n_97), .B1(n_529), .B2(n_530), .Y(n_528) );
AOI22xp33_ASAP7_75t_L g710 ( .A1(n_39), .A2(n_82), .B1(n_395), .B2(n_396), .Y(n_710) );
AOI22xp33_ASAP7_75t_L g626 ( .A1(n_40), .A2(n_242), .B1(n_461), .B2(n_527), .Y(n_626) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_41), .A2(n_245), .B1(n_509), .B2(n_510), .Y(n_508) );
INVx1_ASAP7_75t_L g361 ( .A(n_42), .Y(n_361) );
AO222x2_ASAP7_75t_SL g415 ( .A1(n_43), .A2(n_183), .B1(n_252), .B2(n_355), .C1(n_371), .C2(n_375), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g913 ( .A1(n_45), .A2(n_303), .B1(n_584), .B2(n_810), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g731 ( .A1(n_46), .A2(n_220), .B1(n_407), .B2(n_408), .Y(n_731) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_47), .A2(n_86), .B1(n_609), .B2(n_610), .Y(n_608) );
AOI22xp33_ASAP7_75t_SL g763 ( .A1(n_48), .A2(n_284), .B1(n_395), .B2(n_396), .Y(n_763) );
AOI22xp33_ASAP7_75t_L g817 ( .A1(n_49), .A2(n_106), .B1(n_513), .B2(n_818), .Y(n_817) );
AO222x2_ASAP7_75t_SL g354 ( .A1(n_50), .A2(n_109), .B1(n_147), .B2(n_355), .C1(n_371), .C2(n_375), .Y(n_354) );
AOI22xp33_ASAP7_75t_L g864 ( .A1(n_51), .A2(n_261), .B1(n_488), .B2(n_589), .Y(n_864) );
AO22x2_ASAP7_75t_L g369 ( .A1(n_52), .A2(n_174), .B1(n_359), .B2(n_370), .Y(n_369) );
XNOR2x1_ASAP7_75t_L g430 ( .A(n_54), .B(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_55), .A2(n_61), .B1(n_404), .B2(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_56), .B(n_586), .Y(n_585) );
AOI22xp33_ASAP7_75t_L g868 ( .A1(n_57), .A2(n_285), .B1(n_615), .B2(n_666), .Y(n_868) );
INVx1_ASAP7_75t_L g592 ( .A(n_58), .Y(n_592) );
AOI22xp33_ASAP7_75t_L g493 ( .A1(n_59), .A2(n_309), .B1(n_494), .B2(n_497), .Y(n_493) );
AOI221x1_ASAP7_75t_L g452 ( .A1(n_60), .A2(n_69), .B1(n_453), .B2(n_456), .C(n_458), .Y(n_452) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_62), .A2(n_140), .B1(n_407), .B2(n_408), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g760 ( .A1(n_63), .A2(n_244), .B1(n_380), .B2(n_635), .Y(n_760) );
AOI22xp5_ASAP7_75t_L g660 ( .A1(n_64), .A2(n_294), .B1(n_488), .B2(n_589), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g813 ( .A1(n_65), .A2(n_114), .B1(n_526), .B2(n_814), .Y(n_813) );
AOI22xp33_ASAP7_75t_L g844 ( .A1(n_66), .A2(n_142), .B1(n_526), .B2(n_527), .Y(n_844) );
AOI22xp33_ASAP7_75t_L g426 ( .A1(n_67), .A2(n_289), .B1(n_401), .B2(n_404), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g712 ( .A1(n_68), .A2(n_231), .B1(n_532), .B2(n_667), .Y(n_712) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_70), .B(n_541), .Y(n_540) );
CKINVDCx20_ASAP7_75t_R g808 ( .A(n_71), .Y(n_808) );
AOI22xp33_ASAP7_75t_L g671 ( .A1(n_72), .A2(n_221), .B1(n_440), .B2(n_619), .Y(n_671) );
AOI22xp33_ASAP7_75t_L g767 ( .A1(n_73), .A2(n_240), .B1(n_404), .B2(n_620), .Y(n_767) );
INVx1_ASAP7_75t_L g464 ( .A(n_74), .Y(n_464) );
AOI22xp33_ASAP7_75t_L g406 ( .A1(n_75), .A2(n_333), .B1(n_407), .B2(n_408), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g579 ( .A1(n_76), .A2(n_219), .B1(n_487), .B2(n_580), .Y(n_579) );
AOI22xp5_ASAP7_75t_L g850 ( .A1(n_77), .A2(n_102), .B1(n_457), .B2(n_631), .Y(n_850) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_78), .A2(n_228), .B1(n_401), .B2(n_532), .Y(n_687) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_79), .A2(n_290), .B1(n_522), .B2(n_747), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g841 ( .A1(n_80), .A2(n_178), .B1(n_513), .B2(n_514), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_81), .B(n_586), .Y(n_655) );
AOI22xp5_ASAP7_75t_L g553 ( .A1(n_83), .A2(n_123), .B1(n_451), .B2(n_532), .Y(n_553) );
INVx1_ASAP7_75t_L g479 ( .A(n_84), .Y(n_479) );
INVx1_ASAP7_75t_L g438 ( .A(n_85), .Y(n_438) );
AOI22xp33_ASAP7_75t_SL g724 ( .A1(n_87), .A2(n_276), .B1(n_386), .B2(n_389), .Y(n_724) );
AO22x2_ASAP7_75t_L g803 ( .A1(n_89), .A2(n_804), .B1(n_829), .B2(n_830), .Y(n_803) );
INVx1_ASAP7_75t_L g830 ( .A(n_89), .Y(n_830) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_91), .A2(n_212), .B1(n_399), .B2(n_405), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_92), .A2(n_293), .B1(n_383), .B2(n_418), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g809 ( .A1(n_93), .A2(n_313), .B1(n_584), .B2(n_810), .Y(n_809) );
AOI22xp33_ASAP7_75t_L g845 ( .A1(n_94), .A2(n_263), .B1(n_524), .B2(n_846), .Y(n_845) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_95), .A2(n_295), .B1(n_401), .B2(n_404), .Y(n_554) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_98), .A2(n_126), .B1(n_488), .B2(n_820), .Y(n_875) );
OAI22x1_ASAP7_75t_L g597 ( .A1(n_99), .A2(n_598), .B1(n_599), .B2(n_621), .Y(n_597) );
INVx1_ASAP7_75t_L g598 ( .A(n_99), .Y(n_598) );
CKINVDCx20_ASAP7_75t_R g792 ( .A(n_100), .Y(n_792) );
AOI22xp33_ASAP7_75t_L g869 ( .A1(n_101), .A2(n_223), .B1(n_440), .B2(n_619), .Y(n_869) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_105), .A2(n_287), .B1(n_669), .B2(n_670), .Y(n_668) );
AO22x2_ASAP7_75t_L g366 ( .A1(n_107), .A2(n_248), .B1(n_359), .B2(n_367), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g379 ( .A1(n_108), .A2(n_200), .B1(n_380), .B2(n_383), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g614 ( .A1(n_110), .A2(n_181), .B1(n_615), .B2(n_617), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g575 ( .A1(n_111), .A2(n_189), .B1(n_529), .B2(n_576), .Y(n_575) );
AOI22xp33_ASAP7_75t_L g743 ( .A1(n_112), .A2(n_329), .B1(n_744), .B2(n_745), .Y(n_743) );
AOI22xp5_ASAP7_75t_L g398 ( .A1(n_115), .A2(n_306), .B1(n_399), .B2(n_401), .Y(n_398) );
AOI22xp33_ASAP7_75t_L g681 ( .A1(n_116), .A2(n_158), .B1(n_371), .B2(n_375), .Y(n_681) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_117), .A2(n_234), .B1(n_572), .B2(n_814), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_118), .A2(n_132), .B1(n_495), .B2(n_603), .Y(n_602) );
AOI22xp33_ASAP7_75t_L g512 ( .A1(n_119), .A2(n_139), .B1(n_513), .B2(n_514), .Y(n_512) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_120), .A2(n_151), .B1(n_386), .B2(n_389), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g800 ( .A1(n_121), .A2(n_130), .B1(n_619), .B2(n_666), .Y(n_800) );
AOI22xp33_ASAP7_75t_L g680 ( .A1(n_124), .A2(n_188), .B1(n_386), .B2(n_420), .Y(n_680) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_127), .A2(n_278), .B1(n_371), .B2(n_642), .Y(n_757) );
AOI22xp33_ASAP7_75t_L g711 ( .A1(n_128), .A2(n_262), .B1(n_408), .B2(n_557), .Y(n_711) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_129), .A2(n_319), .B1(n_820), .B2(n_821), .Y(n_819) );
XOR2x2_ASAP7_75t_L g833 ( .A(n_131), .B(n_834), .Y(n_833) );
AOI22xp33_ASAP7_75t_L g766 ( .A1(n_133), .A2(n_279), .B1(n_407), .B2(n_408), .Y(n_766) );
CKINVDCx20_ASAP7_75t_R g543 ( .A(n_134), .Y(n_543) );
CKINVDCx20_ASAP7_75t_R g428 ( .A(n_135), .Y(n_428) );
AO22x1_ASAP7_75t_L g785 ( .A1(n_136), .A2(n_197), .B1(n_477), .B2(n_786), .Y(n_785) );
AOI22xp33_ASAP7_75t_L g858 ( .A1(n_137), .A2(n_155), .B1(n_662), .B2(n_663), .Y(n_858) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_138), .B(n_587), .Y(n_683) );
AOI22xp33_ASAP7_75t_SL g728 ( .A1(n_141), .A2(n_201), .B1(n_395), .B2(n_396), .Y(n_728) );
AOI22xp33_ASAP7_75t_L g732 ( .A1(n_143), .A2(n_160), .B1(n_399), .B2(n_405), .Y(n_732) );
AOI22xp33_ASAP7_75t_SL g759 ( .A1(n_144), .A2(n_312), .B1(n_386), .B2(n_389), .Y(n_759) );
OA22x2_ASAP7_75t_L g872 ( .A1(n_145), .A2(n_873), .B1(n_887), .B2(n_888), .Y(n_872) );
INVx1_ASAP7_75t_L g887 ( .A(n_145), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g823 ( .A1(n_146), .A2(n_255), .B1(n_824), .B2(n_825), .Y(n_823) );
INVx1_ASAP7_75t_L g437 ( .A(n_148), .Y(n_437) );
AOI22xp33_ASAP7_75t_L g565 ( .A1(n_149), .A2(n_227), .B1(n_435), .B2(n_524), .Y(n_565) );
AOI22xp33_ASAP7_75t_L g605 ( .A1(n_150), .A2(n_318), .B1(n_488), .B2(n_606), .Y(n_605) );
CKINVDCx20_ASAP7_75t_R g721 ( .A(n_152), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g630 ( .A1(n_153), .A2(n_213), .B1(n_569), .B2(n_631), .Y(n_630) );
AOI22xp33_ASAP7_75t_L g827 ( .A1(n_154), .A2(n_191), .B1(n_435), .B2(n_828), .Y(n_827) );
AOI22xp5_ASAP7_75t_L g627 ( .A1(n_156), .A2(n_249), .B1(n_522), .B2(n_628), .Y(n_627) );
XNOR2x1_ASAP7_75t_L g652 ( .A(n_157), .B(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g729 ( .A1(n_159), .A2(n_307), .B1(n_401), .B2(n_404), .Y(n_729) );
AOI22xp33_ASAP7_75t_L g558 ( .A1(n_161), .A2(n_193), .B1(n_395), .B2(n_396), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g549 ( .A(n_162), .Y(n_549) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_163), .A2(n_207), .B1(n_663), .B2(n_739), .Y(n_738) );
AOI22xp33_ASAP7_75t_L g521 ( .A1(n_164), .A2(n_216), .B1(n_522), .B2(n_524), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g618 ( .A1(n_166), .A2(n_218), .B1(n_619), .B2(n_620), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g756 ( .A(n_167), .B(n_587), .Y(n_756) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_168), .A2(n_206), .B1(n_609), .B2(n_610), .Y(n_866) );
AOI22xp33_ASAP7_75t_L g880 ( .A1(n_170), .A2(n_288), .B1(n_569), .B2(n_881), .Y(n_880) );
AOI22xp33_ASAP7_75t_L g877 ( .A1(n_171), .A2(n_254), .B1(n_659), .B2(n_810), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_172), .A2(n_324), .B1(n_395), .B2(n_396), .Y(n_423) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_173), .A2(n_235), .B1(n_404), .B2(n_667), .Y(n_688) );
INVx1_ASAP7_75t_L g902 ( .A(n_174), .Y(n_902) );
AOI22xp33_ASAP7_75t_L g725 ( .A1(n_175), .A2(n_232), .B1(n_380), .B2(n_383), .Y(n_725) );
INVx1_ASAP7_75t_L g447 ( .A(n_176), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g798 ( .A1(n_177), .A2(n_229), .B1(n_628), .B2(n_673), .Y(n_798) );
AOI22xp33_ASAP7_75t_L g556 ( .A1(n_179), .A2(n_316), .B1(n_408), .B2(n_557), .Y(n_556) );
CKINVDCx20_ASAP7_75t_R g690 ( .A(n_180), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g797 ( .A1(n_184), .A2(n_326), .B1(n_574), .B2(n_612), .Y(n_797) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_185), .A2(n_269), .B1(n_396), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_SL g920 ( .A1(n_186), .A2(n_321), .B1(n_573), .B2(n_670), .Y(n_920) );
AOI22xp33_ASAP7_75t_L g689 ( .A1(n_187), .A2(n_217), .B1(n_407), .B2(n_408), .Y(n_689) );
AOI22xp33_ASAP7_75t_L g925 ( .A1(n_190), .A2(n_330), .B1(n_530), .B2(n_846), .Y(n_925) );
AOI22xp33_ASAP7_75t_L g705 ( .A1(n_192), .A2(n_328), .B1(n_371), .B2(n_375), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g656 ( .A1(n_194), .A2(n_210), .B1(n_477), .B2(n_657), .Y(n_656) );
AOI22xp33_ASAP7_75t_L g525 ( .A1(n_196), .A2(n_334), .B1(n_526), .B2(n_527), .Y(n_525) );
INVx2_ASAP7_75t_L g342 ( .A(n_198), .Y(n_342) );
XOR2x2_ASAP7_75t_L g855 ( .A(n_199), .B(n_856), .Y(n_855) );
CKINVDCx20_ASAP7_75t_R g768 ( .A(n_202), .Y(n_768) );
AOI22xp5_ASAP7_75t_L g709 ( .A1(n_204), .A2(n_224), .B1(n_401), .B2(n_404), .Y(n_709) );
AOI22xp33_ASAP7_75t_SL g840 ( .A1(n_205), .A2(n_300), .B1(n_516), .B2(n_517), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g424 ( .A1(n_208), .A2(n_270), .B1(n_407), .B2(n_408), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g706 ( .A1(n_211), .A2(n_291), .B1(n_380), .B2(n_383), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g905 ( .A1(n_214), .A2(n_906), .B1(n_907), .B2(n_926), .Y(n_905) );
CKINVDCx20_ASAP7_75t_R g926 ( .A(n_214), .Y(n_926) );
NAND2xp5_ASAP7_75t_L g736 ( .A(n_230), .B(n_737), .Y(n_736) );
INVx1_ASAP7_75t_L g444 ( .A(n_233), .Y(n_444) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_236), .A2(n_283), .B1(n_861), .B2(n_862), .Y(n_860) );
OA22x2_ASAP7_75t_L g622 ( .A1(n_237), .A2(n_623), .B1(n_624), .B2(n_643), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_237), .Y(n_623) );
AO21x2_ASAP7_75t_L g646 ( .A1(n_237), .A2(n_624), .B(n_647), .Y(n_646) );
INVx1_ASAP7_75t_L g750 ( .A(n_238), .Y(n_750) );
XNOR2xp5_ASAP7_75t_L g716 ( .A(n_239), .B(n_717), .Y(n_716) );
AOI22x1_ASAP7_75t_L g351 ( .A1(n_241), .A2(n_352), .B1(n_409), .B2(n_410), .Y(n_351) );
INVx1_ASAP7_75t_L g410 ( .A(n_241), .Y(n_410) );
XNOR2x1_ASAP7_75t_L g505 ( .A(n_243), .B(n_506), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g588 ( .A1(n_246), .A2(n_251), .B1(n_495), .B2(n_589), .Y(n_588) );
AOI22xp33_ASAP7_75t_L g566 ( .A1(n_247), .A2(n_299), .B1(n_567), .B2(n_568), .Y(n_566) );
NOR2xp33_ASAP7_75t_L g900 ( .A(n_248), .B(n_901), .Y(n_900) );
AOI211xp5_ASAP7_75t_L g335 ( .A1(n_250), .A2(n_336), .B(n_345), .C(n_904), .Y(n_335) );
AOI22xp5_ASAP7_75t_L g764 ( .A1(n_253), .A2(n_275), .B1(n_401), .B2(n_532), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g878 ( .A(n_256), .B(n_473), .Y(n_878) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_257), .A2(n_322), .B1(n_386), .B2(n_420), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g812 ( .A1(n_260), .A2(n_298), .B1(n_450), .B2(n_631), .Y(n_812) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_264), .A2(n_327), .B1(n_574), .B2(n_612), .Y(n_611) );
OA22x2_ASAP7_75t_L g534 ( .A1(n_265), .A2(n_535), .B1(n_536), .B2(n_559), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g535 ( .A(n_265), .Y(n_535) );
AND2x2_ASAP7_75t_L g782 ( .A(n_266), .B(n_783), .Y(n_782) );
AOI22xp33_ASAP7_75t_L g883 ( .A1(n_267), .A2(n_282), .B1(n_670), .B2(n_884), .Y(n_883) );
INVx3_ASAP7_75t_L g359 ( .A(n_268), .Y(n_359) );
INVx1_ASAP7_75t_L g465 ( .A(n_272), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_273), .A2(n_304), .B1(n_582), .B2(n_583), .Y(n_581) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_277), .A2(n_286), .B1(n_477), .B2(n_509), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g636 ( .A1(n_280), .A2(n_323), .B1(n_517), .B2(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g777 ( .A(n_281), .Y(n_777) );
INVx1_ASAP7_75t_L g484 ( .A(n_296), .Y(n_484) );
CKINVDCx20_ASAP7_75t_R g912 ( .A(n_297), .Y(n_912) );
CKINVDCx20_ASAP7_75t_R g788 ( .A(n_308), .Y(n_788) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_310), .B(n_519), .Y(n_518) );
NAND2xp5_ASAP7_75t_L g859 ( .A(n_314), .B(n_586), .Y(n_859) );
NAND2xp5_ASAP7_75t_SL g343 ( .A(n_315), .B(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g898 ( .A(n_315), .Y(n_898) );
INVx1_ASAP7_75t_L g339 ( .A(n_317), .Y(n_339) );
AND2x2_ASAP7_75t_R g928 ( .A(n_317), .B(n_898), .Y(n_928) );
INVxp67_ASAP7_75t_L g344 ( .A(n_320), .Y(n_344) );
CKINVDCx20_ASAP7_75t_R g794 ( .A(n_325), .Y(n_794) );
INVx1_ASAP7_75t_L g470 ( .A(n_331), .Y(n_470) );
XOR2x2_ASAP7_75t_L g932 ( .A(n_332), .B(n_908), .Y(n_932) );
CKINVDCx20_ASAP7_75t_R g937 ( .A(n_332), .Y(n_937) );
BUFx2_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
NOR2x1_ASAP7_75t_R g337 ( .A(n_338), .B(n_340), .Y(n_337) );
OR2x2_ASAP7_75t_L g936 ( .A(n_338), .B(n_341), .Y(n_936) );
INVx1_ASAP7_75t_L g338 ( .A(n_339), .Y(n_338) );
NOR2xp33_ASAP7_75t_L g897 ( .A(n_339), .B(n_898), .Y(n_897) );
INVx1_ASAP7_75t_L g340 ( .A(n_341), .Y(n_340) );
NOR2xp33_ASAP7_75t_L g341 ( .A(n_342), .B(n_343), .Y(n_341) );
AOI221xp5_ASAP7_75t_L g345 ( .A1(n_346), .A2(n_696), .B1(n_893), .B2(n_894), .C(n_895), .Y(n_345) );
INVx1_ASAP7_75t_L g893 ( .A(n_346), .Y(n_893) );
AOI22xp5_ASAP7_75t_L g346 ( .A1(n_347), .A2(n_595), .B1(n_694), .B2(n_695), .Y(n_346) );
INVxp67_ASAP7_75t_SL g695 ( .A(n_347), .Y(n_695) );
AOI22xp5_ASAP7_75t_L g347 ( .A1(n_348), .A2(n_501), .B1(n_593), .B2(n_594), .Y(n_347) );
INVx2_ASAP7_75t_L g593 ( .A(n_348), .Y(n_593) );
OA22x2_ASAP7_75t_L g348 ( .A1(n_349), .A2(n_350), .B1(n_430), .B2(n_500), .Y(n_348) );
INVx2_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
AO22x2_ASAP7_75t_L g350 ( .A1(n_351), .A2(n_411), .B1(n_412), .B2(n_429), .Y(n_350) );
INVx1_ASAP7_75t_L g429 ( .A(n_351), .Y(n_429) );
INVx1_ASAP7_75t_L g409 ( .A(n_352), .Y(n_409) );
NAND2x1_ASAP7_75t_SL g352 ( .A(n_353), .B(n_392), .Y(n_352) );
NOR2xp67_ASAP7_75t_L g353 ( .A(n_354), .B(n_378), .Y(n_353) );
BUFx2_ASAP7_75t_L g541 ( .A(n_355), .Y(n_541) );
INVx2_ASAP7_75t_SL g720 ( .A(n_355), .Y(n_720) );
AND2x4_ASAP7_75t_L g355 ( .A(n_356), .B(n_364), .Y(n_355) );
AND2x2_ASAP7_75t_L g383 ( .A(n_356), .B(n_384), .Y(n_383) );
AND2x2_ASAP7_75t_L g389 ( .A(n_356), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g420 ( .A(n_356), .B(n_390), .Y(n_420) );
AND2x2_ASAP7_75t_L g475 ( .A(n_356), .B(n_364), .Y(n_475) );
AND2x4_ASAP7_75t_L g492 ( .A(n_356), .B(n_390), .Y(n_492) );
AND2x4_ASAP7_75t_L g499 ( .A(n_356), .B(n_384), .Y(n_499) );
AND2x2_ASAP7_75t_L g635 ( .A(n_356), .B(n_384), .Y(n_635) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_362), .Y(n_356) );
AND2x2_ASAP7_75t_L g373 ( .A(n_357), .B(n_374), .Y(n_373) );
HB1xp67_ASAP7_75t_L g376 ( .A(n_357), .Y(n_376) );
INVx2_ASAP7_75t_L g382 ( .A(n_357), .Y(n_382) );
OAI22x1_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g363 ( .A(n_359), .Y(n_363) );
INVx2_ASAP7_75t_L g367 ( .A(n_359), .Y(n_367) );
INVx1_ASAP7_75t_L g370 ( .A(n_359), .Y(n_370) );
INVx2_ASAP7_75t_L g374 ( .A(n_362), .Y(n_374) );
AND2x2_ASAP7_75t_L g381 ( .A(n_362), .B(n_382), .Y(n_381) );
BUFx2_ASAP7_75t_L g397 ( .A(n_362), .Y(n_397) );
AND2x2_ASAP7_75t_L g399 ( .A(n_364), .B(n_400), .Y(n_399) );
AND2x6_ASAP7_75t_L g404 ( .A(n_364), .B(n_381), .Y(n_404) );
AND2x2_ASAP7_75t_L g407 ( .A(n_364), .B(n_373), .Y(n_407) );
AND2x2_ASAP7_75t_L g436 ( .A(n_364), .B(n_381), .Y(n_436) );
AND2x4_ASAP7_75t_L g446 ( .A(n_364), .B(n_373), .Y(n_446) );
AND2x4_ASAP7_75t_L g455 ( .A(n_364), .B(n_400), .Y(n_455) );
AND2x2_ASAP7_75t_L g557 ( .A(n_364), .B(n_373), .Y(n_557) );
AND2x4_ASAP7_75t_L g364 ( .A(n_365), .B(n_368), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AND2x4_ASAP7_75t_L g372 ( .A(n_366), .B(n_368), .Y(n_372) );
AND2x2_ASAP7_75t_L g377 ( .A(n_366), .B(n_369), .Y(n_377) );
INVx1_ASAP7_75t_L g388 ( .A(n_366), .Y(n_388) );
INVxp67_ASAP7_75t_L g384 ( .A(n_368), .Y(n_384) );
INVx2_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AND2x2_ASAP7_75t_L g387 ( .A(n_369), .B(n_388), .Y(n_387) );
INVx1_ASAP7_75t_SL g641 ( .A(n_371), .Y(n_641) );
AND2x4_ASAP7_75t_L g371 ( .A(n_372), .B(n_373), .Y(n_371) );
AND2x2_ASAP7_75t_L g380 ( .A(n_372), .B(n_381), .Y(n_380) );
AND2x2_ASAP7_75t_L g405 ( .A(n_372), .B(n_400), .Y(n_405) );
AND2x2_ASAP7_75t_L g418 ( .A(n_372), .B(n_381), .Y(n_418) );
AND2x4_ASAP7_75t_L g451 ( .A(n_372), .B(n_400), .Y(n_451) );
AND2x2_ASAP7_75t_L g483 ( .A(n_372), .B(n_373), .Y(n_483) );
AND2x4_ASAP7_75t_L g496 ( .A(n_372), .B(n_381), .Y(n_496) );
AND2x4_ASAP7_75t_L g386 ( .A(n_373), .B(n_387), .Y(n_386) );
AND2x2_ASAP7_75t_L g489 ( .A(n_373), .B(n_387), .Y(n_489) );
AND2x4_ASAP7_75t_L g400 ( .A(n_374), .B(n_382), .Y(n_400) );
AND2x2_ASAP7_75t_SL g375 ( .A(n_376), .B(n_377), .Y(n_375) );
AND2x2_ASAP7_75t_L g478 ( .A(n_376), .B(n_377), .Y(n_478) );
AND2x2_ASAP7_75t_SL g642 ( .A(n_376), .B(n_377), .Y(n_642) );
AND2x4_ASAP7_75t_L g396 ( .A(n_377), .B(n_397), .Y(n_396) );
AND2x4_ASAP7_75t_L g408 ( .A(n_377), .B(n_400), .Y(n_408) );
AND2x4_ASAP7_75t_L g457 ( .A(n_377), .B(n_400), .Y(n_457) );
AND2x4_ASAP7_75t_L g467 ( .A(n_377), .B(n_397), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_379), .B(n_385), .Y(n_378) );
AND2x2_ASAP7_75t_SL g395 ( .A(n_381), .B(n_387), .Y(n_395) );
AND2x2_ASAP7_75t_L g463 ( .A(n_381), .B(n_387), .Y(n_463) );
AND2x2_ASAP7_75t_L g686 ( .A(n_381), .B(n_387), .Y(n_686) );
INVxp67_ASAP7_75t_L g550 ( .A(n_383), .Y(n_550) );
AND2x6_ASAP7_75t_L g401 ( .A(n_387), .B(n_400), .Y(n_401) );
AND2x4_ASAP7_75t_L g442 ( .A(n_387), .B(n_400), .Y(n_442) );
HB1xp67_ASAP7_75t_L g391 ( .A(n_388), .Y(n_391) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_393), .B(n_402), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_394), .B(n_398), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
INVx1_ASAP7_75t_L g882 ( .A(n_404), .Y(n_882) );
AO22x2_ASAP7_75t_L g832 ( .A1(n_411), .A2(n_412), .B1(n_833), .B2(n_851), .Y(n_832) );
INVx2_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
XOR2x2_ASAP7_75t_L g412 ( .A(n_413), .B(n_428), .Y(n_412) );
NAND2x1_ASAP7_75t_L g413 ( .A(n_414), .B(n_421), .Y(n_413) );
NOR2x1_ASAP7_75t_L g414 ( .A(n_415), .B(n_416), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g416 ( .A(n_417), .B(n_419), .Y(n_416) );
INVxp67_ASAP7_75t_L g548 ( .A(n_418), .Y(n_548) );
NOR2x1_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_423), .B(n_424), .Y(n_422) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_426), .B(n_427), .Y(n_425) );
INVx2_ASAP7_75t_L g500 ( .A(n_430), .Y(n_500) );
NAND3xp33_ASAP7_75t_L g431 ( .A(n_432), .B(n_452), .C(n_468), .Y(n_431) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_433), .B(n_443), .Y(n_432) );
OAI22xp33_ASAP7_75t_L g433 ( .A1(n_434), .A2(n_437), .B1(n_438), .B2(n_439), .Y(n_433) );
INVx2_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
BUFx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVx3_ASAP7_75t_L g523 ( .A(n_436), .Y(n_523) );
BUFx2_ASAP7_75t_L g849 ( .A(n_436), .Y(n_849) );
INVx1_ASAP7_75t_L g439 ( .A(n_440), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g524 ( .A(n_441), .Y(n_524) );
INVx1_ASAP7_75t_SL g617 ( .A(n_441), .Y(n_617) );
INVx2_ASAP7_75t_L g628 ( .A(n_441), .Y(n_628) );
INVx2_ASAP7_75t_SL g747 ( .A(n_441), .Y(n_747) );
INVx2_ASAP7_75t_L g828 ( .A(n_441), .Y(n_828) );
INVx8_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g443 ( .A1(n_444), .A2(n_445), .B1(n_447), .B2(n_448), .Y(n_443) );
INVx3_ASAP7_75t_L g529 ( .A(n_445), .Y(n_529) );
INVx2_ASAP7_75t_L g609 ( .A(n_445), .Y(n_609) );
INVx6_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
BUFx3_ASAP7_75t_L g631 ( .A(n_446), .Y(n_631) );
INVx1_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
BUFx2_ASAP7_75t_L g449 ( .A(n_450), .Y(n_449) );
BUFx3_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
BUFx6f_ASAP7_75t_L g530 ( .A(n_451), .Y(n_530) );
INVx2_ASAP7_75t_L g570 ( .A(n_451), .Y(n_570) );
BUFx6f_ASAP7_75t_L g667 ( .A(n_451), .Y(n_667) );
INVx3_ASAP7_75t_SL g453 ( .A(n_454), .Y(n_453) );
INVx3_ASAP7_75t_L g532 ( .A(n_454), .Y(n_532) );
INVx2_ASAP7_75t_L g567 ( .A(n_454), .Y(n_567) );
INVx4_ASAP7_75t_L g616 ( .A(n_454), .Y(n_616) );
INVx2_ASAP7_75t_SL g824 ( .A(n_454), .Y(n_824) );
INVx2_ASAP7_75t_SL g846 ( .A(n_454), .Y(n_846) );
INVx8_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
BUFx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
BUFx3_ASAP7_75t_L g533 ( .A(n_457), .Y(n_533) );
BUFx3_ASAP7_75t_L g577 ( .A(n_457), .Y(n_577) );
BUFx2_ASAP7_75t_SL g610 ( .A(n_457), .Y(n_610) );
INVx2_ASAP7_75t_L g826 ( .A(n_457), .Y(n_826) );
OAI22xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_464), .B1(n_465), .B2(n_466), .Y(n_458) );
HB1xp67_ASAP7_75t_L g459 ( .A(n_460), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g613 ( .A(n_461), .Y(n_613) );
BUFx6f_ASAP7_75t_L g669 ( .A(n_461), .Y(n_669) );
INVx2_ASAP7_75t_L g461 ( .A(n_462), .Y(n_461) );
INVx1_ASAP7_75t_L g573 ( .A(n_462), .Y(n_573) );
INVx1_ASAP7_75t_L g884 ( .A(n_462), .Y(n_884) );
INVx2_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
BUFx6f_ASAP7_75t_L g526 ( .A(n_463), .Y(n_526) );
BUFx3_ASAP7_75t_L g744 ( .A(n_463), .Y(n_744) );
INVx2_ASAP7_75t_L g527 ( .A(n_466), .Y(n_527) );
INVx2_ASAP7_75t_L g574 ( .A(n_466), .Y(n_574) );
INVx5_ASAP7_75t_SL g466 ( .A(n_467), .Y(n_466) );
BUFx2_ASAP7_75t_L g670 ( .A(n_467), .Y(n_670) );
BUFx3_ASAP7_75t_L g745 ( .A(n_467), .Y(n_745) );
BUFx2_ASAP7_75t_L g814 ( .A(n_467), .Y(n_814) );
NOR2xp33_ASAP7_75t_L g468 ( .A(n_469), .B(n_485), .Y(n_468) );
OAI222xp33_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B1(n_476), .B2(n_479), .C1(n_480), .C2(n_484), .Y(n_469) );
INVx3_ASAP7_75t_L g471 ( .A(n_472), .Y(n_471) );
BUFx6f_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
INVx2_ASAP7_75t_L g807 ( .A(n_473), .Y(n_807) );
INVx3_ASAP7_75t_SL g473 ( .A(n_474), .Y(n_473) );
INVx4_ASAP7_75t_SL g519 ( .A(n_474), .Y(n_519) );
INVx4_ASAP7_75t_SL g587 ( .A(n_474), .Y(n_587) );
INVx3_ASAP7_75t_L g737 ( .A(n_474), .Y(n_737) );
BUFx2_ASAP7_75t_L g784 ( .A(n_474), .Y(n_784) );
INVx6_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx2_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
BUFx12f_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx3_ASAP7_75t_L g511 ( .A(n_478), .Y(n_511) );
INVx1_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
INVx2_ASAP7_75t_L g509 ( .A(n_482), .Y(n_509) );
INVx1_ASAP7_75t_L g786 ( .A(n_482), .Y(n_786) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
BUFx3_ASAP7_75t_L g584 ( .A(n_483), .Y(n_584) );
BUFx3_ASAP7_75t_L g659 ( .A(n_483), .Y(n_659) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_486), .B(n_493), .Y(n_485) );
BUFx6f_ASAP7_75t_SL g487 ( .A(n_488), .Y(n_487) );
INVx1_ASAP7_75t_L g544 ( .A(n_488), .Y(n_544) );
BUFx6f_ASAP7_75t_L g488 ( .A(n_489), .Y(n_488) );
BUFx6f_ASAP7_75t_L g516 ( .A(n_489), .Y(n_516) );
INVx3_ASAP7_75t_L g638 ( .A(n_489), .Y(n_638) );
INVx2_ASAP7_75t_SL g490 ( .A(n_491), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g542 ( .A1(n_491), .A2(n_543), .B1(n_544), .B2(n_545), .Y(n_542) );
INVx1_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
BUFx3_ASAP7_75t_L g517 ( .A(n_492), .Y(n_517) );
INVx2_ASAP7_75t_L g591 ( .A(n_492), .Y(n_591) );
BUFx4f_ASAP7_75t_L g606 ( .A(n_492), .Y(n_606) );
BUFx6f_ASAP7_75t_SL g820 ( .A(n_492), .Y(n_820) );
BUFx2_ASAP7_75t_L g494 ( .A(n_495), .Y(n_494) );
BUFx2_ASAP7_75t_L g662 ( .A(n_495), .Y(n_662) );
INVx1_ASAP7_75t_L g793 ( .A(n_495), .Y(n_793) );
BUFx6f_ASAP7_75t_L g495 ( .A(n_496), .Y(n_495) );
BUFx3_ASAP7_75t_L g513 ( .A(n_496), .Y(n_513) );
BUFx2_ASAP7_75t_L g739 ( .A(n_496), .Y(n_739) );
BUFx2_ASAP7_75t_L g917 ( .A(n_496), .Y(n_917) );
INVx2_ASAP7_75t_L g497 ( .A(n_498), .Y(n_497) );
INVx2_ASAP7_75t_L g514 ( .A(n_498), .Y(n_514) );
INVx2_ASAP7_75t_SL g580 ( .A(n_498), .Y(n_580) );
INVx2_ASAP7_75t_L g603 ( .A(n_498), .Y(n_603) );
INVx2_ASAP7_75t_L g663 ( .A(n_498), .Y(n_663) );
OAI22xp5_ASAP7_75t_L g791 ( .A1(n_498), .A2(n_792), .B1(n_793), .B2(n_794), .Y(n_791) );
INVx2_ASAP7_75t_SL g818 ( .A(n_498), .Y(n_818) );
INVx6_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
INVx1_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
OA22x2_ASAP7_75t_L g501 ( .A1(n_502), .A2(n_503), .B1(n_561), .B2(n_562), .Y(n_501) );
INVx2_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
AO22x2_ASAP7_75t_L g503 ( .A1(n_504), .A2(n_505), .B1(n_534), .B2(n_560), .Y(n_503) );
INVx1_ASAP7_75t_SL g504 ( .A(n_505), .Y(n_504) );
OR2x2_ASAP7_75t_L g506 ( .A(n_507), .B(n_520), .Y(n_506) );
NAND4xp25_ASAP7_75t_L g507 ( .A(n_508), .B(n_512), .C(n_515), .D(n_518), .Y(n_507) );
BUFx2_ASAP7_75t_L g582 ( .A(n_510), .Y(n_582) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx2_ASAP7_75t_L g810 ( .A(n_511), .Y(n_810) );
INVx3_ASAP7_75t_L g863 ( .A(n_511), .Y(n_863) );
INVx1_ASAP7_75t_SL g911 ( .A(n_519), .Y(n_911) );
NAND4xp25_ASAP7_75t_L g520 ( .A(n_521), .B(n_525), .C(n_528), .D(n_531), .Y(n_520) );
INVx3_ASAP7_75t_L g522 ( .A(n_523), .Y(n_522) );
INVx2_ASAP7_75t_SL g619 ( .A(n_523), .Y(n_619) );
INVx2_ASAP7_75t_L g922 ( .A(n_523), .Y(n_922) );
INVx2_ASAP7_75t_L g560 ( .A(n_534), .Y(n_560) );
INVx1_ASAP7_75t_L g559 ( .A(n_536), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_537), .B(n_551), .Y(n_536) );
NOR3xp33_ASAP7_75t_L g537 ( .A(n_538), .B(n_542), .C(n_546), .Y(n_537) );
NAND2xp5_ASAP7_75t_SL g538 ( .A(n_539), .B(n_540), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g546 ( .A1(n_547), .A2(n_548), .B1(n_549), .B2(n_550), .Y(n_546) );
NOR2xp33_ASAP7_75t_L g551 ( .A(n_552), .B(n_555), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_553), .B(n_554), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_556), .B(n_558), .Y(n_555) );
INVx2_ASAP7_75t_L g561 ( .A(n_562), .Y(n_561) );
XNOR2x1_ASAP7_75t_L g562 ( .A(n_563), .B(n_592), .Y(n_562) );
NOR2xp67_ASAP7_75t_L g563 ( .A(n_564), .B(n_578), .Y(n_563) );
NAND4xp25_ASAP7_75t_L g564 ( .A(n_565), .B(n_566), .C(n_571), .D(n_575), .Y(n_564) );
HB1xp67_ASAP7_75t_L g568 ( .A(n_569), .Y(n_568) );
INVx2_ASAP7_75t_L g569 ( .A(n_570), .Y(n_569) );
INVx1_ASAP7_75t_L g620 ( .A(n_570), .Y(n_620) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
NAND4xp25_ASAP7_75t_L g578 ( .A(n_579), .B(n_581), .C(n_585), .D(n_588), .Y(n_578) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
BUFx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
INVx3_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_590), .A2(n_788), .B1(n_789), .B2(n_790), .Y(n_787) );
BUFx2_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx2_ASAP7_75t_SL g694 ( .A(n_595), .Y(n_694) );
AO22x2_ASAP7_75t_L g595 ( .A1(n_596), .A2(n_649), .B1(n_692), .B2(n_693), .Y(n_595) );
INVx2_ASAP7_75t_SL g692 ( .A(n_596), .Y(n_692) );
OA22x2_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_622), .B1(n_644), .B2(n_645), .Y(n_596) );
INVx1_ASAP7_75t_SL g644 ( .A(n_597), .Y(n_644) );
INVx2_ASAP7_75t_SL g621 ( .A(n_599), .Y(n_621) );
OR2x2_ASAP7_75t_L g599 ( .A(n_600), .B(n_607), .Y(n_599) );
NAND4xp25_ASAP7_75t_SL g600 ( .A(n_601), .B(n_602), .C(n_604), .D(n_605), .Y(n_600) );
NAND4xp25_ASAP7_75t_L g607 ( .A(n_608), .B(n_611), .C(n_614), .D(n_618), .Y(n_607) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
BUFx6f_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g674 ( .A(n_616), .Y(n_674) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_622), .A2(n_645), .B1(n_652), .B2(n_675), .Y(n_651) );
CKINVDCx20_ASAP7_75t_R g648 ( .A(n_623), .Y(n_648) );
INVx1_ASAP7_75t_L g643 ( .A(n_624), .Y(n_643) );
NOR2x1_ASAP7_75t_SL g647 ( .A(n_624), .B(n_648), .Y(n_647) );
NAND4xp75_ASAP7_75t_L g624 ( .A(n_625), .B(n_629), .C(n_633), .D(n_639), .Y(n_624) );
AND2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_627), .Y(n_625) );
AND2x2_ASAP7_75t_L g629 ( .A(n_630), .B(n_632), .Y(n_629) );
AND2x2_ASAP7_75t_L g633 ( .A(n_634), .B(n_636), .Y(n_633) );
INVx2_ASAP7_75t_SL g789 ( .A(n_637), .Y(n_789) );
INVx4_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVx2_ASAP7_75t_L g821 ( .A(n_638), .Y(n_821) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
INVx3_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx4_ASAP7_75t_L g693 ( .A(n_649), .Y(n_693) );
OA22x2_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .B1(n_676), .B2(n_691), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
INVx1_ASAP7_75t_SL g675 ( .A(n_652), .Y(n_675) );
OR2x2_ASAP7_75t_L g653 ( .A(n_654), .B(n_664), .Y(n_653) );
NAND4xp25_ASAP7_75t_L g654 ( .A(n_655), .B(n_656), .C(n_660), .D(n_661), .Y(n_654) );
INVx2_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
BUFx6f_ASAP7_75t_SL g861 ( .A(n_659), .Y(n_861) );
NAND4xp25_ASAP7_75t_L g664 ( .A(n_665), .B(n_668), .C(n_671), .D(n_672), .Y(n_664) );
BUFx6f_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g673 ( .A(n_674), .Y(n_673) );
INVx1_ASAP7_75t_L g691 ( .A(n_676), .Y(n_691) );
INVx2_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
XNOR2x2_ASAP7_75t_L g677 ( .A(n_678), .B(n_690), .Y(n_677) );
NOR2x1_ASAP7_75t_L g678 ( .A(n_679), .B(n_684), .Y(n_678) );
NAND4xp25_ASAP7_75t_L g679 ( .A(n_680), .B(n_681), .C(n_682), .D(n_683), .Y(n_679) );
NAND4xp25_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .C(n_688), .D(n_689), .Y(n_684) );
INVx1_ASAP7_75t_L g894 ( .A(n_696), .Y(n_894) );
AOI22xp5_ASAP7_75t_SL g696 ( .A1(n_697), .A2(n_698), .B1(n_771), .B2(n_892), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
AOI22xp33_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_713), .B1(n_714), .B2(n_770), .Y(n_698) );
INVx2_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_700), .Y(n_770) );
XNOR2x1_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .Y(n_700) );
NOR2x1_ASAP7_75t_L g702 ( .A(n_703), .B(n_708), .Y(n_702) );
NAND4xp25_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .C(n_706), .D(n_707), .Y(n_703) );
NAND4xp25_ASAP7_75t_L g708 ( .A(n_709), .B(n_710), .C(n_711), .D(n_712), .Y(n_708) );
INVx2_ASAP7_75t_L g713 ( .A(n_714), .Y(n_713) );
AO22x2_ASAP7_75t_L g714 ( .A1(n_715), .A2(n_751), .B1(n_752), .B2(n_769), .Y(n_714) );
INVx2_ASAP7_75t_L g769 ( .A(n_715), .Y(n_769) );
XOR2x1_ASAP7_75t_SL g715 ( .A(n_716), .B(n_733), .Y(n_715) );
NAND2xp5_ASAP7_75t_SL g717 ( .A(n_718), .B(n_726), .Y(n_717) );
NOR2xp33_ASAP7_75t_L g718 ( .A(n_719), .B(n_723), .Y(n_718) );
OAI21xp5_ASAP7_75t_SL g719 ( .A1(n_720), .A2(n_721), .B(n_722), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_724), .B(n_725), .Y(n_723) );
NOR2xp33_ASAP7_75t_L g726 ( .A(n_727), .B(n_730), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g727 ( .A(n_728), .B(n_729), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g730 ( .A(n_731), .B(n_732), .Y(n_730) );
XNOR2x1_ASAP7_75t_L g733 ( .A(n_734), .B(n_750), .Y(n_733) );
OR2x2_ASAP7_75t_L g734 ( .A(n_735), .B(n_742), .Y(n_734) );
NAND4xp25_ASAP7_75t_L g735 ( .A(n_736), .B(n_738), .C(n_740), .D(n_741), .Y(n_735) );
NAND4xp25_ASAP7_75t_L g742 ( .A(n_743), .B(n_746), .C(n_748), .D(n_749), .Y(n_742) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
XOR2x2_ASAP7_75t_L g752 ( .A(n_753), .B(n_768), .Y(n_752) );
NAND2x1_ASAP7_75t_L g753 ( .A(n_754), .B(n_761), .Y(n_753) );
NOR2x1_ASAP7_75t_L g754 ( .A(n_755), .B(n_758), .Y(n_754) );
NAND2xp5_ASAP7_75t_L g755 ( .A(n_756), .B(n_757), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g758 ( .A(n_759), .B(n_760), .Y(n_758) );
NOR2x1_ASAP7_75t_L g761 ( .A(n_762), .B(n_765), .Y(n_761) );
NAND2xp5_ASAP7_75t_L g762 ( .A(n_763), .B(n_764), .Y(n_762) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_766), .B(n_767), .Y(n_765) );
INVx1_ASAP7_75t_L g892 ( .A(n_771), .Y(n_892) );
OAI22xp5_ASAP7_75t_L g771 ( .A1(n_772), .A2(n_773), .B1(n_853), .B2(n_891), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
INVx1_ASAP7_75t_L g773 ( .A(n_774), .Y(n_773) );
AO22x2_ASAP7_75t_L g774 ( .A1(n_775), .A2(n_831), .B1(n_832), .B2(n_852), .Y(n_774) );
INVx1_ASAP7_75t_L g852 ( .A(n_775), .Y(n_852) );
XNOR2xp5_ASAP7_75t_L g775 ( .A(n_776), .B(n_803), .Y(n_775) );
OAI21x1_ASAP7_75t_L g776 ( .A1(n_777), .A2(n_778), .B(n_802), .Y(n_776) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_777), .B(n_780), .Y(n_802) );
INVx1_ASAP7_75t_L g778 ( .A(n_779), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
NAND2xp5_ASAP7_75t_L g780 ( .A(n_781), .B(n_795), .Y(n_780) );
NOR4xp75_ASAP7_75t_L g781 ( .A(n_782), .B(n_785), .C(n_787), .D(n_791), .Y(n_781) );
INVx2_ASAP7_75t_SL g783 ( .A(n_784), .Y(n_783) );
OAI21xp5_ASAP7_75t_SL g836 ( .A1(n_784), .A2(n_837), .B(n_838), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g795 ( .A(n_796), .B(n_799), .Y(n_795) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_797), .B(n_798), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_800), .B(n_801), .Y(n_799) );
INVx2_ASAP7_75t_SL g829 ( .A(n_804), .Y(n_829) );
AND2x2_ASAP7_75t_L g804 ( .A(n_805), .B(n_815), .Y(n_804) );
NOR2xp33_ASAP7_75t_L g805 ( .A(n_806), .B(n_811), .Y(n_805) );
OAI21xp33_ASAP7_75t_SL g806 ( .A1(n_807), .A2(n_808), .B(n_809), .Y(n_806) );
NAND2xp5_ASAP7_75t_L g811 ( .A(n_812), .B(n_813), .Y(n_811) );
NOR2xp33_ASAP7_75t_L g815 ( .A(n_816), .B(n_822), .Y(n_815) );
NAND2xp5_ASAP7_75t_L g816 ( .A(n_817), .B(n_819), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g822 ( .A(n_823), .B(n_827), .Y(n_822) );
INVx2_ASAP7_75t_SL g825 ( .A(n_826), .Y(n_825) );
INVx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx2_ASAP7_75t_L g851 ( .A(n_833), .Y(n_851) );
NAND2x1_ASAP7_75t_SL g834 ( .A(n_835), .B(n_842), .Y(n_834) );
NOR2x1_ASAP7_75t_L g835 ( .A(n_836), .B(n_839), .Y(n_835) );
NAND2xp5_ASAP7_75t_L g839 ( .A(n_840), .B(n_841), .Y(n_839) );
NOR2x1_ASAP7_75t_L g842 ( .A(n_843), .B(n_847), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_848), .B(n_850), .Y(n_847) );
INVx1_ASAP7_75t_L g891 ( .A(n_853), .Y(n_891) );
OAI22xp5_ASAP7_75t_SL g853 ( .A1(n_854), .A2(n_870), .B1(n_889), .B2(n_890), .Y(n_853) );
INVx3_ASAP7_75t_L g889 ( .A(n_854), .Y(n_889) );
INVx5_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
NOR2x1_ASAP7_75t_L g856 ( .A(n_857), .B(n_865), .Y(n_856) );
NAND4xp25_ASAP7_75t_L g857 ( .A(n_858), .B(n_859), .C(n_860), .D(n_864), .Y(n_857) );
BUFx6f_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
NAND4xp25_ASAP7_75t_L g865 ( .A(n_866), .B(n_867), .C(n_868), .D(n_869), .Y(n_865) );
INVx1_ASAP7_75t_L g890 ( .A(n_870), .Y(n_890) );
BUFx2_ASAP7_75t_L g870 ( .A(n_871), .Y(n_870) );
INVx1_ASAP7_75t_L g871 ( .A(n_872), .Y(n_871) );
INVx1_ASAP7_75t_L g888 ( .A(n_873), .Y(n_888) );
NOR2x1_ASAP7_75t_L g873 ( .A(n_874), .B(n_879), .Y(n_873) );
NAND4xp25_ASAP7_75t_L g874 ( .A(n_875), .B(n_876), .C(n_877), .D(n_878), .Y(n_874) );
NAND4xp25_ASAP7_75t_L g879 ( .A(n_880), .B(n_883), .C(n_885), .D(n_886), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx3_ASAP7_75t_SL g895 ( .A(n_896), .Y(n_895) );
AND2x2_ASAP7_75t_L g896 ( .A(n_897), .B(n_899), .Y(n_896) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_897), .B(n_900), .Y(n_935) );
INVx1_ASAP7_75t_L g899 ( .A(n_900), .Y(n_899) );
NAND2xp5_ASAP7_75t_L g901 ( .A(n_902), .B(n_903), .Y(n_901) );
OAI222xp33_ASAP7_75t_L g904 ( .A1(n_905), .A2(n_927), .B1(n_929), .B2(n_933), .C1(n_936), .C2(n_937), .Y(n_904) );
CKINVDCx20_ASAP7_75t_R g906 ( .A(n_907), .Y(n_906) );
HB1xp67_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
NAND2x1_ASAP7_75t_L g908 ( .A(n_909), .B(n_918), .Y(n_908) );
NOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_914), .Y(n_909) );
OAI21xp5_ASAP7_75t_SL g910 ( .A1(n_911), .A2(n_912), .B(n_913), .Y(n_910) );
NAND2xp5_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
NOR2x1_ASAP7_75t_L g918 ( .A(n_919), .B(n_923), .Y(n_918) );
NAND2xp5_ASAP7_75t_L g919 ( .A(n_920), .B(n_921), .Y(n_919) );
NAND2xp5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
INVx1_ASAP7_75t_SL g927 ( .A(n_928), .Y(n_927) );
INVx3_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx2_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g931 ( .A(n_932), .Y(n_931) );
CKINVDCx20_ASAP7_75t_R g933 ( .A(n_934), .Y(n_933) );
CKINVDCx6p67_ASAP7_75t_R g934 ( .A(n_935), .Y(n_934) );
endmodule