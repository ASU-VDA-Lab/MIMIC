module real_aes_12836_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_222;
wire n_750;
wire n_631;
wire n_943;
wire n_287;
wire n_357;
wire n_905;
wire n_503;
wire n_386;
wire n_673;
wire n_635;
wire n_518;
wire n_254;
wire n_792;
wire n_207;
wire n_878;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_132;
wire n_857;
wire n_919;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_379;
wire n_374;
wire n_453;
wire n_932;
wire n_235;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_870;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_883;
wire n_356;
wire n_478;
wire n_918;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_121;
wire n_352;
wire n_935;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_263;
wire n_906;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_104;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_860;
wire n_298;
wire n_523;
wire n_909;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_649;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_455;
wire n_310;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_903;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_936;
wire n_610;
wire n_581;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_722;
wire n_745;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_879;
wire n_331;
wire n_182;
wire n_449;
wire n_363;
wire n_417;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_947;
wire n_142;
wire n_561;
wire n_876;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_502;
wire n_434;
wire n_505;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_880;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_869;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_945;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_898;
wire n_848;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_756;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_749;
wire n_663;
wire n_588;
wire n_109;
wire n_914;
wire n_203;
wire n_536;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_133;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_939;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_155;
wire n_653;
wire n_243;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_679;
wire n_633;
wire n_520;
wire n_926;
wire n_922;
wire n_149;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_861;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_639;
wire n_151;
wire n_546;
wire n_587;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_888;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_911;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_170;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_849;
wire n_192;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_237;
wire n_668;
wire n_797;
wire n_862;
INVx2_ASAP7_75t_SL g293 ( .A(n_0), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_1), .Y(n_146) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_2), .A2(n_49), .B(n_132), .Y(n_131) );
INVx1_ASAP7_75t_L g192 ( .A(n_2), .Y(n_192) );
NAND2xp5_ASAP7_75t_SL g240 ( .A(n_3), .B(n_182), .Y(n_240) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_4), .B(n_304), .Y(n_303) );
NAND2xp5_ASAP7_75t_SL g569 ( .A(n_5), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g644 ( .A(n_6), .B(n_329), .Y(n_644) );
AND2x2_ASAP7_75t_L g197 ( .A(n_7), .B(n_161), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g327 ( .A(n_8), .B(n_328), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_9), .B(n_270), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g634 ( .A(n_10), .B(n_270), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g683 ( .A(n_11), .B(n_583), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_12), .B(n_173), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_13), .B(n_154), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_14), .B(n_292), .Y(n_568) );
CKINVDCx5p33_ASAP7_75t_R g618 ( .A(n_15), .Y(n_618) );
BUFx3_ASAP7_75t_L g138 ( .A(n_16), .Y(n_138) );
INVx1_ASAP7_75t_L g152 ( .A(n_16), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_17), .B(n_160), .Y(n_244) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_18), .B(n_169), .Y(n_598) );
CKINVDCx5p33_ASAP7_75t_R g641 ( .A(n_19), .Y(n_641) );
BUFx10_ASAP7_75t_L g113 ( .A(n_20), .Y(n_113) );
NAND2xp5_ASAP7_75t_SL g593 ( .A(n_21), .B(n_210), .Y(n_593) );
CKINVDCx5p33_ASAP7_75t_R g611 ( .A(n_22), .Y(n_611) );
CKINVDCx5p33_ASAP7_75t_R g227 ( .A(n_23), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g627 ( .A(n_24), .B(n_570), .Y(n_627) );
NAND3xp33_ASAP7_75t_L g309 ( .A(n_25), .B(n_136), .C(n_307), .Y(n_309) );
NAND2xp5_ASAP7_75t_SL g597 ( .A(n_26), .B(n_210), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_27), .B(n_270), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g662 ( .A(n_28), .B(n_169), .Y(n_662) );
NAND2xp33_ASAP7_75t_L g573 ( .A(n_29), .B(n_141), .Y(n_573) );
INVx1_ASAP7_75t_L g158 ( .A(n_30), .Y(n_158) );
A2O1A1Ixp33_ASAP7_75t_L g609 ( .A1(n_31), .A2(n_153), .B(n_171), .C(n_610), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g286 ( .A(n_32), .B(n_287), .Y(n_286) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_33), .A2(n_104), .B1(n_937), .B2(n_947), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_34), .B(n_148), .Y(n_594) );
NAND2xp5_ASAP7_75t_SL g682 ( .A(n_35), .B(n_182), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g633 ( .A(n_36), .B(n_238), .Y(n_633) );
INVx1_ASAP7_75t_L g556 ( .A(n_37), .Y(n_556) );
AND3x2_ASAP7_75t_L g936 ( .A(n_37), .B(n_108), .C(n_110), .Y(n_936) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_38), .B(n_272), .Y(n_271) );
AO221x1_ASAP7_75t_L g580 ( .A1(n_39), .A2(n_85), .B1(n_210), .B2(n_237), .C(n_284), .Y(n_580) );
NAND2xp5_ASAP7_75t_SL g642 ( .A(n_40), .B(n_630), .Y(n_642) );
NAND2xp5_ASAP7_75t_SL g149 ( .A(n_41), .B(n_150), .Y(n_149) );
AND2x4_ASAP7_75t_L g157 ( .A(n_42), .B(n_158), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_43), .B(n_160), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g289 ( .A(n_44), .B(n_261), .Y(n_289) );
NAND3xp33_ASAP7_75t_L g665 ( .A(n_45), .B(n_150), .C(n_153), .Y(n_665) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_46), .B(n_160), .Y(n_323) );
AOI21xp33_ASAP7_75t_L g931 ( .A1(n_47), .A2(n_926), .B(n_932), .Y(n_931) );
OAI22x1_ASAP7_75t_L g899 ( .A1(n_48), .A2(n_53), .B1(n_900), .B2(n_901), .Y(n_899) );
CKINVDCx5p33_ASAP7_75t_R g900 ( .A(n_48), .Y(n_900) );
INVx1_ASAP7_75t_L g191 ( .A(n_49), .Y(n_191) );
AND2x2_ASAP7_75t_L g926 ( .A(n_50), .B(n_927), .Y(n_926) );
CKINVDCx5p33_ASAP7_75t_R g180 ( .A(n_51), .Y(n_180) );
A2O1A1Ixp33_ASAP7_75t_L g290 ( .A1(n_52), .A2(n_181), .B(n_291), .C(n_294), .Y(n_290) );
INVx1_ASAP7_75t_L g901 ( .A(n_53), .Y(n_901) );
INVx1_ASAP7_75t_L g132 ( .A(n_54), .Y(n_132) );
CKINVDCx5p33_ASAP7_75t_R g615 ( .A(n_55), .Y(n_615) );
A2O1A1Ixp33_ASAP7_75t_L g675 ( .A1(n_56), .A2(n_676), .B(n_677), .C(n_679), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_57), .B(n_160), .Y(n_159) );
AOI22xp5_ASAP7_75t_L g116 ( .A1(n_58), .A2(n_117), .B1(n_903), .B2(n_904), .Y(n_116) );
CKINVDCx5p33_ASAP7_75t_R g903 ( .A(n_58), .Y(n_903) );
INVx2_ASAP7_75t_L g678 ( .A(n_59), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_60), .B(n_261), .Y(n_646) );
AND2x4_ASAP7_75t_L g945 ( .A(n_61), .B(n_946), .Y(n_945) );
INVx3_ASAP7_75t_L g224 ( .A(n_62), .Y(n_224) );
NOR2xp67_ASAP7_75t_L g109 ( .A(n_63), .B(n_77), .Y(n_109) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_64), .B(n_629), .Y(n_628) );
INVx1_ASAP7_75t_L g946 ( .A(n_65), .Y(n_946) );
NAND2xp5_ASAP7_75t_SL g334 ( .A(n_66), .B(n_220), .Y(n_334) );
INVx1_ASAP7_75t_L g236 ( .A(n_67), .Y(n_236) );
AND2x2_ASAP7_75t_L g635 ( .A(n_68), .B(n_261), .Y(n_635) );
INVx1_ASAP7_75t_L g586 ( .A(n_69), .Y(n_586) );
OAI22xp5_ASAP7_75t_L g912 ( .A1(n_70), .A2(n_75), .B1(n_913), .B2(n_914), .Y(n_912) );
INVx1_ASAP7_75t_L g914 ( .A(n_70), .Y(n_914) );
INVx2_ASAP7_75t_L g111 ( .A(n_71), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g170 ( .A(n_72), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_73), .B(n_140), .Y(n_302) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_74), .B(n_136), .Y(n_135) );
INVxp67_ASAP7_75t_SL g913 ( .A(n_75), .Y(n_913) );
OAI22xp33_ASAP7_75t_L g582 ( .A1(n_76), .A2(n_79), .B1(n_570), .B2(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g664 ( .A(n_78), .B(n_153), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_80), .B(n_277), .Y(n_276) );
INVx1_ASAP7_75t_L g285 ( .A(n_81), .Y(n_285) );
CKINVDCx5p33_ASAP7_75t_R g183 ( .A(n_82), .Y(n_183) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_83), .B(n_242), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_84), .B(n_307), .Y(n_306) );
AND2x2_ASAP7_75t_L g685 ( .A(n_86), .B(n_161), .Y(n_685) );
INVx1_ASAP7_75t_L g144 ( .A(n_87), .Y(n_144) );
BUFx3_ASAP7_75t_L g154 ( .A(n_87), .Y(n_154) );
INVx1_ASAP7_75t_L g187 ( .A(n_87), .Y(n_187) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_88), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g222 ( .A(n_89), .Y(n_222) );
NAND2xp5_ASAP7_75t_SL g588 ( .A(n_90), .B(n_589), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_91), .B(n_189), .Y(n_619) );
OAI22xp5_ASAP7_75t_L g909 ( .A1(n_92), .A2(n_910), .B1(n_911), .B2(n_917), .Y(n_909) );
INVx1_ASAP7_75t_L g910 ( .A(n_92), .Y(n_910) );
NAND2xp5_ASAP7_75t_SL g275 ( .A(n_93), .B(n_172), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_94), .B(n_161), .Y(n_278) );
NAND2xp5_ASAP7_75t_SL g661 ( .A(n_95), .B(n_630), .Y(n_661) );
NAND2xp5_ASAP7_75t_L g575 ( .A(n_96), .B(n_261), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g331 ( .A(n_97), .B(n_332), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_98), .Y(n_214) );
INVx1_ASAP7_75t_L g209 ( .A(n_99), .Y(n_209) );
CKINVDCx5p33_ASAP7_75t_R g667 ( .A(n_100), .Y(n_667) );
CKINVDCx5p33_ASAP7_75t_R g175 ( .A(n_101), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_102), .B(n_220), .Y(n_326) );
AO21x2_ASAP7_75t_L g104 ( .A1(n_105), .A2(n_114), .B(n_905), .Y(n_104) );
INVx6_ASAP7_75t_L g105 ( .A(n_106), .Y(n_105) );
OR2x6_ASAP7_75t_L g106 ( .A(n_107), .B(n_112), .Y(n_106) );
AND2x2_ASAP7_75t_L g107 ( .A(n_108), .B(n_110), .Y(n_107) );
HB1xp67_ASAP7_75t_L g108 ( .A(n_109), .Y(n_108) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_109), .B(n_556), .Y(n_925) );
BUFx2_ASAP7_75t_L g110 ( .A(n_111), .Y(n_110) );
INVx1_ASAP7_75t_L g924 ( .A(n_111), .Y(n_924) );
BUFx3_ASAP7_75t_L g907 ( .A(n_112), .Y(n_907) );
INVx3_ASAP7_75t_L g112 ( .A(n_113), .Y(n_112) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_113), .B(n_936), .Y(n_935) );
HB1xp67_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
OAI22xp5_ASAP7_75t_L g117 ( .A1(n_118), .A2(n_119), .B1(n_899), .B2(n_902), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_119), .Y(n_118) );
XNOR2xp5_ASAP7_75t_L g904 ( .A(n_119), .B(n_899), .Y(n_904) );
OAI22x1_ASAP7_75t_L g119 ( .A1(n_120), .A2(n_551), .B1(n_552), .B2(n_557), .Y(n_119) );
AO22x2_ASAP7_75t_L g911 ( .A1(n_120), .A2(n_912), .B1(n_915), .B2(n_916), .Y(n_911) );
INVx1_ASAP7_75t_L g916 ( .A(n_120), .Y(n_916) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_449), .Y(n_120) );
NOR3xp33_ASAP7_75t_L g121 ( .A(n_122), .B(n_371), .C(n_422), .Y(n_121) );
OAI221xp5_ASAP7_75t_SL g122 ( .A1(n_123), .A2(n_263), .B1(n_311), .B2(n_316), .C(n_340), .Y(n_122) );
AOI211xp5_ASAP7_75t_L g123 ( .A1(n_124), .A2(n_198), .B(n_245), .C(n_253), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
AND2x4_ASAP7_75t_L g546 ( .A(n_125), .B(n_249), .Y(n_546) );
AND2x2_ASAP7_75t_L g125 ( .A(n_126), .B(n_163), .Y(n_125) );
INVx1_ASAP7_75t_L g247 ( .A(n_126), .Y(n_247) );
AND2x2_ASAP7_75t_L g401 ( .A(n_126), .B(n_347), .Y(n_401) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_126), .Y(n_446) );
INVx1_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
INVx2_ASAP7_75t_L g256 ( .A(n_127), .Y(n_256) );
INVx3_ASAP7_75t_L g349 ( .A(n_127), .Y(n_349) );
AND2x2_ASAP7_75t_L g377 ( .A(n_127), .B(n_258), .Y(n_377) );
AND2x2_ASAP7_75t_L g384 ( .A(n_127), .B(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g127 ( .A(n_128), .Y(n_127) );
OAI21x1_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_133), .B(n_159), .Y(n_128) );
OAI21x1_ASAP7_75t_L g229 ( .A1(n_129), .A2(n_230), .B(n_244), .Y(n_229) );
OAI21x1_ASAP7_75t_L g638 ( .A1(n_129), .A2(n_639), .B(n_646), .Y(n_638) );
BUFx3_ASAP7_75t_L g129 ( .A(n_130), .Y(n_129) );
INVxp67_ASAP7_75t_L g668 ( .A(n_130), .Y(n_668) );
BUFx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g162 ( .A(n_131), .Y(n_162) );
BUFx6f_ASAP7_75t_L g261 ( .A(n_131), .Y(n_261) );
INVx1_ASAP7_75t_L g193 ( .A(n_132), .Y(n_193) );
OAI21xp5_ASAP7_75t_L g133 ( .A1(n_134), .A2(n_145), .B(n_155), .Y(n_133) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_139), .B(n_142), .Y(n_134) );
INVx1_ASAP7_75t_L g136 ( .A(n_137), .Y(n_136) );
INVx2_ASAP7_75t_L g238 ( .A(n_137), .Y(n_238) );
INVx2_ASAP7_75t_L g570 ( .A(n_137), .Y(n_570) );
INVx2_ASAP7_75t_L g630 ( .A(n_137), .Y(n_630) );
INVx2_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_138), .Y(n_141) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_138), .Y(n_216) );
INVx2_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx2_ASAP7_75t_L g148 ( .A(n_141), .Y(n_148) );
INVx3_ASAP7_75t_L g169 ( .A(n_141), .Y(n_169) );
INVx2_ASAP7_75t_L g179 ( .A(n_141), .Y(n_179) );
INVx2_ASAP7_75t_L g270 ( .A(n_141), .Y(n_270) );
INVx3_ASAP7_75t_L g284 ( .A(n_141), .Y(n_284) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_142), .A2(n_240), .B(n_241), .Y(n_239) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_142), .A2(n_275), .B(n_276), .Y(n_274) );
AOI21xp5_ASAP7_75t_L g632 ( .A1(n_142), .A2(n_633), .B(n_634), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g643 ( .A1(n_142), .A2(n_644), .B(n_645), .Y(n_643) );
INVx1_ASAP7_75t_L g684 ( .A(n_142), .Y(n_684) );
BUFx10_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
INVx1_ASAP7_75t_L g307 ( .A(n_143), .Y(n_307) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
BUFx3_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
O2A1O1Ixp5_ASAP7_75t_L g145 ( .A1(n_146), .A2(n_147), .B(n_149), .C(n_153), .Y(n_145) );
OAI21xp5_ASAP7_75t_L g663 ( .A1(n_147), .A2(n_664), .B(n_665), .Y(n_663) );
INVx2_ASAP7_75t_L g147 ( .A(n_148), .Y(n_147) );
INVx2_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
INVx2_ASAP7_75t_L g182 ( .A(n_151), .Y(n_182) );
INVx2_ASAP7_75t_L g329 ( .A(n_151), .Y(n_329) );
INVx1_ASAP7_75t_L g333 ( .A(n_151), .Y(n_333) );
INVx1_ASAP7_75t_L g616 ( .A(n_151), .Y(n_616) );
BUFx6f_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
INVx2_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
NOR2xp33_ASAP7_75t_L g211 ( .A(n_154), .B(n_212), .Y(n_211) );
NOR3xp33_ASAP7_75t_L g221 ( .A(n_154), .B(n_212), .C(n_222), .Y(n_221) );
INVx2_ASAP7_75t_L g237 ( .A(n_154), .Y(n_237) );
INVx1_ASAP7_75t_L g599 ( .A(n_154), .Y(n_599) );
OAI21x1_ASAP7_75t_L g300 ( .A1(n_155), .A2(n_301), .B(n_305), .Y(n_300) );
INVx1_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx2_ASAP7_75t_SL g338 ( .A(n_156), .Y(n_338) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
INVx1_ASAP7_75t_L g196 ( .A(n_157), .Y(n_196) );
INVx3_ASAP7_75t_L g212 ( .A(n_157), .Y(n_212) );
BUFx6f_ASAP7_75t_SL g243 ( .A(n_157), .Y(n_243) );
HB1xp67_ASAP7_75t_L g299 ( .A(n_160), .Y(n_299) );
BUFx6f_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_162), .Y(n_161) );
INVx1_ASAP7_75t_L g163 ( .A(n_164), .Y(n_163) );
OR2x2_ASAP7_75t_L g358 ( .A(n_164), .B(n_315), .Y(n_358) );
AO31x2_ASAP7_75t_L g164 ( .A1(n_165), .A2(n_188), .A3(n_194), .B(n_197), .Y(n_164) );
AO31x2_ASAP7_75t_L g369 ( .A1(n_165), .A2(n_188), .A3(n_194), .B(n_197), .Y(n_369) );
INVx2_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OAI21x1_ASAP7_75t_L g258 ( .A1(n_166), .A2(n_259), .B(n_262), .Y(n_258) );
AOI22x1_ASAP7_75t_L g166 ( .A1(n_167), .A2(n_176), .B1(n_177), .B2(n_184), .Y(n_166) );
OAI22x1_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_170), .B1(n_171), .B2(n_175), .Y(n_167) );
INVxp67_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_173), .Y(n_172) );
INVx2_ASAP7_75t_L g272 ( .A(n_173), .Y(n_272) );
HB1xp67_ASAP7_75t_L g287 ( .A(n_173), .Y(n_287) );
INVx2_ASAP7_75t_L g304 ( .A(n_173), .Y(n_304) );
NOR2xp33_ASAP7_75t_L g617 ( .A(n_173), .B(n_618), .Y(n_617) );
INVx3_ASAP7_75t_L g173 ( .A(n_174), .Y(n_173) );
BUFx6f_ASAP7_75t_L g210 ( .A(n_174), .Y(n_210) );
INVx1_ASAP7_75t_L g294 ( .A(n_176), .Y(n_294) );
AOI21x1_ASAP7_75t_L g301 ( .A1(n_176), .A2(n_302), .B(n_303), .Y(n_301) );
AOI21xp5_ASAP7_75t_SL g626 ( .A1(n_176), .A2(n_627), .B(n_628), .Y(n_626) );
OAI22xp5_ASAP7_75t_L g177 ( .A1(n_178), .A2(n_180), .B1(n_181), .B2(n_183), .Y(n_177) );
INVxp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVxp67_ASAP7_75t_L g232 ( .A(n_179), .Y(n_232) );
INVx2_ASAP7_75t_L g181 ( .A(n_182), .Y(n_181) );
AOI21x1_ASAP7_75t_SL g282 ( .A1(n_184), .A2(n_283), .B(n_286), .Y(n_282) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
AOI21xp5_ASAP7_75t_L g325 ( .A1(n_185), .A2(n_326), .B(n_327), .Y(n_325) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_185), .B(n_582), .Y(n_581) );
INVx2_ASAP7_75t_L g185 ( .A(n_186), .Y(n_185) );
INVx2_ASAP7_75t_L g218 ( .A(n_186), .Y(n_218) );
AOI21xp5_ASAP7_75t_L g567 ( .A1(n_186), .A2(n_568), .B(n_569), .Y(n_567) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
BUFx3_ASAP7_75t_L g273 ( .A(n_187), .Y(n_273) );
INVxp67_ASAP7_75t_L g188 ( .A(n_189), .Y(n_188) );
OAI21xp33_ASAP7_75t_L g295 ( .A1(n_189), .A2(n_196), .B(n_289), .Y(n_295) );
INVx2_ASAP7_75t_L g189 ( .A(n_190), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g607 ( .A(n_190), .B(n_338), .Y(n_607) );
AO21x2_ASAP7_75t_L g190 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_190) );
AOI21x1_ASAP7_75t_L g205 ( .A1(n_191), .A2(n_192), .B(n_193), .Y(n_205) );
BUFx2_ASAP7_75t_L g194 ( .A(n_195), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_196), .Y(n_195) );
INVx1_ASAP7_75t_L g262 ( .A(n_197), .Y(n_262) );
INVx1_ASAP7_75t_L g198 ( .A(n_199), .Y(n_198) );
AOI322xp5_ASAP7_75t_L g372 ( .A1(n_199), .A2(n_373), .A3(n_377), .B1(n_378), .B2(n_381), .C1(n_388), .C2(n_396), .Y(n_372) );
INVx1_ASAP7_75t_L g199 ( .A(n_200), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
AND2x2_ASAP7_75t_L g396 ( .A(n_201), .B(n_348), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_201), .B(n_348), .Y(n_411) );
AND2x2_ASAP7_75t_L g464 ( .A(n_201), .B(n_377), .Y(n_464) );
AND2x2_ASAP7_75t_L g201 ( .A(n_202), .B(n_228), .Y(n_201) );
INVx3_ASAP7_75t_L g251 ( .A(n_202), .Y(n_251) );
AO21x2_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_206), .B(n_226), .Y(n_202) );
AO21x1_ASAP7_75t_L g386 ( .A1(n_203), .A2(n_206), .B(n_226), .Y(n_386) );
HB1xp67_ASAP7_75t_L g203 ( .A(n_204), .Y(n_203) );
NOR2xp33_ASAP7_75t_SL g226 ( .A(n_204), .B(n_227), .Y(n_226) );
NOR2xp33_ASAP7_75t_L g585 ( .A(n_204), .B(n_586), .Y(n_585) );
INVx2_ASAP7_75t_L g204 ( .A(n_205), .Y(n_204) );
NOR2xp33_ASAP7_75t_R g584 ( .A(n_205), .B(n_212), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_207), .B(n_219), .Y(n_206) );
AOI22xp5_ASAP7_75t_L g207 ( .A1(n_208), .A2(n_211), .B1(n_213), .B2(n_217), .Y(n_207) );
NOR2xp33_ASAP7_75t_L g208 ( .A(n_209), .B(n_210), .Y(n_208) );
INVx1_ASAP7_75t_L g225 ( .A(n_210), .Y(n_225) );
INVx2_ASAP7_75t_L g277 ( .A(n_210), .Y(n_277) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_212), .B(n_218), .Y(n_217) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_212), .B(n_218), .C(n_224), .Y(n_223) );
INVx2_ASAP7_75t_L g574 ( .A(n_212), .Y(n_574) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_212), .B(n_261), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_214), .B(n_215), .Y(n_213) );
INVx2_ASAP7_75t_L g220 ( .A(n_215), .Y(n_220) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
INVx1_ASAP7_75t_L g242 ( .A(n_216), .Y(n_242) );
INVx2_ASAP7_75t_L g292 ( .A(n_216), .Y(n_292) );
INVx2_ASAP7_75t_L g583 ( .A(n_216), .Y(n_583) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_220), .A2(n_221), .B1(n_223), .B2(n_225), .Y(n_219) );
INVx1_ASAP7_75t_L g252 ( .A(n_228), .Y(n_252) );
AND2x2_ASAP7_75t_L g257 ( .A(n_228), .B(n_258), .Y(n_257) );
INVx3_ASAP7_75t_L g315 ( .A(n_228), .Y(n_315) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_228), .Y(n_406) );
INVx2_ASAP7_75t_L g419 ( .A(n_228), .Y(n_419) );
AND2x2_ASAP7_75t_L g429 ( .A(n_228), .B(n_251), .Y(n_429) );
INVx1_ASAP7_75t_L g490 ( .A(n_228), .Y(n_490) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_229), .Y(n_228) );
OAI21x1_ASAP7_75t_L g230 ( .A1(n_231), .A2(n_239), .B(n_243), .Y(n_230) );
OAI21xp5_ASAP7_75t_L g231 ( .A1(n_232), .A2(n_233), .B(n_234), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_235), .B(n_238), .Y(n_234) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_236), .B(n_237), .Y(n_235) );
INVx1_ASAP7_75t_L g595 ( .A(n_237), .Y(n_595) );
OAI21x1_ASAP7_75t_L g267 ( .A1(n_243), .A2(n_268), .B(n_274), .Y(n_267) );
OAI21x1_ASAP7_75t_L g639 ( .A1(n_243), .A2(n_640), .B(n_643), .Y(n_639) );
NOR2xp67_ASAP7_75t_L g245 ( .A(n_246), .B(n_248), .Y(n_245) );
HB1xp67_ASAP7_75t_L g246 ( .A(n_247), .Y(n_246) );
INVx2_ASAP7_75t_L g507 ( .A(n_247), .Y(n_507) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_250), .Y(n_249) );
OR2x2_ASAP7_75t_L g533 ( .A(n_250), .B(n_368), .Y(n_533) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g347 ( .A(n_251), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_251), .B(n_349), .Y(n_370) );
INVx1_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
NAND2xp5_ASAP7_75t_SL g254 ( .A(n_255), .B(n_257), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_255), .B(n_455), .Y(n_479) );
INVx1_ASAP7_75t_L g255 ( .A(n_256), .Y(n_255) );
NOR2xp67_ASAP7_75t_L g313 ( .A(n_256), .B(n_314), .Y(n_313) );
AND2x4_ASAP7_75t_L g438 ( .A(n_257), .B(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_L g348 ( .A(n_258), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g457 ( .A(n_258), .Y(n_457) );
OAI21x1_ASAP7_75t_L g266 ( .A1(n_259), .A2(n_267), .B(n_278), .Y(n_266) );
OAI21x1_ASAP7_75t_L g319 ( .A1(n_259), .A2(n_267), .B(n_278), .Y(n_319) );
BUFx6f_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
NOR2x1_ASAP7_75t_SL g336 ( .A(n_260), .B(n_337), .Y(n_336) );
BUFx6f_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g356 ( .A(n_261), .Y(n_356) );
INVxp67_ASAP7_75t_SL g590 ( .A(n_261), .Y(n_590) );
INVx2_ASAP7_75t_L g625 ( .A(n_261), .Y(n_625) );
OR2x2_ASAP7_75t_L g263 ( .A(n_264), .B(n_279), .Y(n_263) );
AND2x2_ASAP7_75t_L g363 ( .A(n_264), .B(n_321), .Y(n_363) );
OR2x2_ASAP7_75t_L g530 ( .A(n_264), .B(n_361), .Y(n_530) );
INVx1_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g343 ( .A(n_265), .B(n_344), .Y(n_343) );
BUFx3_ASAP7_75t_L g375 ( .A(n_265), .Y(n_375) );
AND2x2_ASAP7_75t_L g502 ( .A(n_265), .B(n_280), .Y(n_502) );
AND2x4_ASAP7_75t_L g518 ( .A(n_265), .B(n_415), .Y(n_518) );
INVx2_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g462 ( .A(n_266), .Y(n_462) );
AOI21xp5_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_271), .B(n_273), .Y(n_268) );
INVx2_ASAP7_75t_L g335 ( .A(n_273), .Y(n_335) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_273), .A2(n_572), .B(n_573), .Y(n_571) );
INVx1_ASAP7_75t_L g679 ( .A(n_273), .Y(n_679) );
INVxp67_ASAP7_75t_L g308 ( .A(n_277), .Y(n_308) );
OR2x2_ASAP7_75t_L g379 ( .A(n_279), .B(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g426 ( .A(n_279), .Y(n_426) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_296), .Y(n_279) );
AND2x4_ASAP7_75t_L g318 ( .A(n_280), .B(n_319), .Y(n_318) );
HB1xp67_ASAP7_75t_L g365 ( .A(n_280), .Y(n_365) );
INVx1_ASAP7_75t_L g391 ( .A(n_280), .Y(n_391) );
AND2x2_ASAP7_75t_L g434 ( .A(n_280), .B(n_354), .Y(n_434) );
INVx2_ASAP7_75t_L g280 ( .A(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g353 ( .A(n_281), .Y(n_353) );
OAI21x1_ASAP7_75t_L g281 ( .A1(n_282), .A2(n_288), .B(n_295), .Y(n_281) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
NOR2xp33_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
AND2x4_ASAP7_75t_L g395 ( .A(n_296), .B(n_321), .Y(n_395) );
INVx1_ASAP7_75t_L g409 ( .A(n_296), .Y(n_409) );
INVx2_ASAP7_75t_L g296 ( .A(n_297), .Y(n_296) );
INVxp67_ASAP7_75t_SL g339 ( .A(n_297), .Y(n_339) );
INVx2_ASAP7_75t_L g362 ( .A(n_297), .Y(n_362) );
INVx2_ASAP7_75t_L g297 ( .A(n_298), .Y(n_297) );
OAI21x1_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_300), .B(n_310), .Y(n_298) );
OA21x2_ASAP7_75t_L g354 ( .A1(n_300), .A2(n_310), .B(n_355), .Y(n_354) );
O2A1O1Ixp5_ASAP7_75t_L g640 ( .A1(n_304), .A2(n_599), .B(n_641), .C(n_642), .Y(n_640) );
OAI21xp5_ASAP7_75t_L g305 ( .A1(n_306), .A2(n_308), .B(n_309), .Y(n_305) );
INVxp67_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
HB1xp67_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
OR2x2_ASAP7_75t_L g476 ( .A(n_314), .B(n_477), .Y(n_476) );
BUFx2_ASAP7_75t_L g497 ( .A(n_314), .Y(n_497) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_315), .B(n_486), .Y(n_500) );
OR2x2_ASAP7_75t_L g316 ( .A(n_317), .B(n_320), .Y(n_316) );
INVx2_ASAP7_75t_L g317 ( .A(n_318), .Y(n_317) );
AND2x2_ASAP7_75t_L g407 ( .A(n_318), .B(n_408), .Y(n_407) );
AND2x2_ASAP7_75t_L g470 ( .A(n_318), .B(n_471), .Y(n_470) );
AND2x2_ASAP7_75t_L g495 ( .A(n_318), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g539 ( .A(n_318), .Y(n_539) );
AND2x2_ASAP7_75t_L g392 ( .A(n_319), .B(n_362), .Y(n_392) );
AND2x4_ASAP7_75t_L g394 ( .A(n_319), .B(n_395), .Y(n_394) );
OR2x2_ASAP7_75t_L g399 ( .A(n_319), .B(n_352), .Y(n_399) );
AND2x4_ASAP7_75t_L g414 ( .A(n_319), .B(n_415), .Y(n_414) );
OR2x2_ASAP7_75t_L g320 ( .A(n_321), .B(n_339), .Y(n_320) );
INVx2_ASAP7_75t_L g344 ( .A(n_321), .Y(n_344) );
INVx2_ASAP7_75t_L g366 ( .A(n_321), .Y(n_366) );
BUFx2_ASAP7_75t_L g380 ( .A(n_321), .Y(n_380) );
INVx1_ASAP7_75t_L g436 ( .A(n_321), .Y(n_436) );
AND2x2_ASAP7_75t_L g496 ( .A(n_321), .B(n_354), .Y(n_496) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
NAND2x1_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
OAI21x1_ASAP7_75t_SL g324 ( .A1(n_325), .A2(n_330), .B(n_336), .Y(n_324) );
INVx2_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AOI21xp5_ASAP7_75t_L g330 ( .A1(n_331), .A2(n_334), .B(n_335), .Y(n_330) );
INVx1_ASAP7_75t_L g332 ( .A(n_333), .Y(n_332) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
AND2x2_ASAP7_75t_L g376 ( .A(n_339), .B(n_344), .Y(n_376) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_350), .B(n_357), .Y(n_340) );
INVxp67_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_343), .B(n_345), .Y(n_342) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_343), .B(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g519 ( .A(n_343), .Y(n_519) );
AND2x2_ASAP7_75t_L g531 ( .A(n_343), .B(n_351), .Y(n_531) );
BUFx2_ASAP7_75t_L g471 ( .A(n_344), .Y(n_471) );
INVx1_ASAP7_75t_L g545 ( .A(n_344), .Y(n_545) );
INVx1_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
NAND2xp5_ASAP7_75t_L g346 ( .A(n_347), .B(n_348), .Y(n_346) );
NAND2xp5_ASAP7_75t_L g404 ( .A(n_348), .B(n_405), .Y(n_404) );
INVx2_ASAP7_75t_L g420 ( .A(n_348), .Y(n_420) );
INVx2_ASAP7_75t_SL g350 ( .A(n_351), .Y(n_350) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_351), .A2(n_542), .B1(n_544), .B2(n_546), .Y(n_541) );
INVx2_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
OR2x2_ASAP7_75t_SL g352 ( .A(n_353), .B(n_354), .Y(n_352) );
OR2x6_ASAP7_75t_L g361 ( .A(n_353), .B(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g415 ( .A(n_353), .Y(n_415) );
OA21x2_ASAP7_75t_L g565 ( .A1(n_355), .A2(n_566), .B(n_575), .Y(n_565) );
INVx1_ASAP7_75t_SL g355 ( .A(n_356), .Y(n_355) );
OAI22xp5_ASAP7_75t_L g357 ( .A1(n_358), .A2(n_359), .B1(n_364), .B2(n_367), .Y(n_357) );
INVx2_ASAP7_75t_SL g402 ( .A(n_358), .Y(n_402) );
OR2x2_ASAP7_75t_L g431 ( .A(n_358), .B(n_370), .Y(n_431) );
INVx2_ASAP7_75t_L g468 ( .A(n_359), .Y(n_468) );
NAND2x1p5_ASAP7_75t_L g359 ( .A(n_360), .B(n_363), .Y(n_359) );
INVx2_ASAP7_75t_SL g360 ( .A(n_361), .Y(n_360) );
OR2x2_ASAP7_75t_L g516 ( .A(n_361), .B(n_366), .Y(n_516) );
OR2x2_ASAP7_75t_L g549 ( .A(n_361), .B(n_375), .Y(n_549) );
NAND2xp5_ASAP7_75t_L g364 ( .A(n_365), .B(n_366), .Y(n_364) );
AND2x2_ASAP7_75t_L g437 ( .A(n_365), .B(n_392), .Y(n_437) );
INVx1_ASAP7_75t_L g413 ( .A(n_366), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_366), .B(n_390), .Y(n_453) );
OR2x2_ASAP7_75t_L g489 ( .A(n_366), .B(n_490), .Y(n_489) );
OR2x2_ASAP7_75t_L g367 ( .A(n_368), .B(n_370), .Y(n_367) );
INVx1_ASAP7_75t_L g486 ( .A(n_368), .Y(n_486) );
BUFx3_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
INVx2_ASAP7_75t_L g387 ( .A(n_369), .Y(n_387) );
INVx1_ASAP7_75t_L g439 ( .A(n_370), .Y(n_439) );
HB1xp67_ASAP7_75t_L g473 ( .A(n_370), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g371 ( .A(n_372), .B(n_397), .Y(n_371) );
INVx2_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_375), .B(n_376), .Y(n_374) );
INVx2_ASAP7_75t_L g443 ( .A(n_375), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_375), .B(n_395), .Y(n_448) );
AND2x2_ASAP7_75t_L g461 ( .A(n_376), .B(n_462), .Y(n_461) );
BUFx3_ASAP7_75t_L g521 ( .A(n_376), .Y(n_521) );
INVx1_ASAP7_75t_L g523 ( .A(n_377), .Y(n_523) );
INVx1_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
AND2x2_ASAP7_75t_L g501 ( .A(n_380), .B(n_502), .Y(n_501) );
NAND2x1_ASAP7_75t_L g487 ( .A(n_381), .B(n_488), .Y(n_487) );
INVx3_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
INVx2_ASAP7_75t_L g514 ( .A(n_382), .Y(n_514) );
OR2x6_ASAP7_75t_L g382 ( .A(n_383), .B(n_387), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g477 ( .A(n_384), .Y(n_477) );
AND2x2_ASAP7_75t_L g537 ( .A(n_384), .B(n_387), .Y(n_537) );
INVx1_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g418 ( .A(n_386), .B(n_419), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_386), .B(n_457), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_387), .B(n_429), .Y(n_428) );
INVx2_ASAP7_75t_L g528 ( .A(n_387), .Y(n_528) );
NAND2x1_ASAP7_75t_L g388 ( .A(n_389), .B(n_393), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
HB1xp67_ASAP7_75t_L g491 ( .A(n_390), .Y(n_491) );
AND2x2_ASAP7_75t_L g390 ( .A(n_391), .B(n_392), .Y(n_390) );
INVx2_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
AOI221x1_ASAP7_75t_L g397 ( .A1(n_398), .A2(n_400), .B1(n_403), .B2(n_407), .C(n_410), .Y(n_397) );
INVx3_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
AOI22xp5_ASAP7_75t_L g432 ( .A1(n_400), .A2(n_433), .B1(n_437), .B2(n_438), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g440 ( .A1(n_400), .A2(n_441), .B1(n_444), .B2(n_447), .Y(n_440) );
INVxp67_ASAP7_75t_SL g538 ( .A(n_400), .Y(n_538) );
AND2x4_ASAP7_75t_L g400 ( .A(n_401), .B(n_402), .Y(n_400) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OR2x2_ASAP7_75t_L g478 ( .A(n_405), .B(n_479), .Y(n_478) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_408), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g442 ( .A(n_408), .B(n_443), .Y(n_442) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
OAI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B1(n_416), .B2(n_421), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_413), .B(n_414), .Y(n_412) );
AND2x4_ASAP7_75t_L g481 ( .A(n_413), .B(n_426), .Y(n_481) );
AOI22xp5_ASAP7_75t_L g423 ( .A1(n_414), .A2(n_424), .B1(n_427), .B2(n_430), .Y(n_423) );
AND2x2_ASAP7_75t_L g504 ( .A(n_414), .B(n_471), .Y(n_504) );
OR2x2_ASAP7_75t_L g416 ( .A(n_417), .B(n_420), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
AND2x2_ASAP7_75t_L g485 ( .A(n_418), .B(n_486), .Y(n_485) );
INVx1_ASAP7_75t_L g506 ( .A(n_418), .Y(n_506) );
AND2x2_ASAP7_75t_L g527 ( .A(n_418), .B(n_528), .Y(n_527) );
AND2x2_ASAP7_75t_L g544 ( .A(n_418), .B(n_545), .Y(n_544) );
NAND3xp33_ASAP7_75t_SL g422 ( .A(n_423), .B(n_432), .C(n_440), .Y(n_422) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVx1_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_429), .B(n_446), .Y(n_445) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
AND2x2_ASAP7_75t_L g433 ( .A(n_434), .B(n_435), .Y(n_433) );
INVx2_ASAP7_75t_L g435 ( .A(n_436), .Y(n_435) );
INVxp67_ASAP7_75t_L g475 ( .A(n_437), .Y(n_475) );
OAI21xp5_ASAP7_75t_L g498 ( .A1(n_438), .A2(n_499), .B(n_501), .Y(n_498) );
INVx1_ASAP7_75t_L g441 ( .A(n_442), .Y(n_441) );
INVxp67_ASAP7_75t_SL g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g543 ( .A(n_446), .Y(n_543) );
INVx1_ASAP7_75t_L g459 ( .A(n_447), .Y(n_459) );
INVx2_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
NOR2x1_ASAP7_75t_L g449 ( .A(n_450), .B(n_508), .Y(n_449) );
NAND3xp33_ASAP7_75t_SL g450 ( .A(n_451), .B(n_465), .C(n_482), .Y(n_450) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_452), .A2(n_454), .B(n_458), .Y(n_451) );
INVx1_ASAP7_75t_L g452 ( .A(n_453), .Y(n_452) );
HB1xp67_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
AOI21xp5_ASAP7_75t_L g458 ( .A1(n_459), .A2(n_460), .B(n_463), .Y(n_458) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
OAI22xp5_ASAP7_75t_SL g542 ( .A1(n_462), .A2(n_517), .B1(n_528), .B2(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g550 ( .A(n_462), .Y(n_550) );
INVx2_ASAP7_75t_L g463 ( .A(n_464), .Y(n_463) );
AOI21xp5_ASAP7_75t_L g465 ( .A1(n_466), .A2(n_472), .B(n_474), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_467), .B(n_469), .Y(n_466) );
INVx2_ASAP7_75t_SL g467 ( .A(n_468), .Y(n_467) );
INVx1_ASAP7_75t_L g469 ( .A(n_470), .Y(n_469) );
INVx1_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
OAI22xp5_ASAP7_75t_L g474 ( .A1(n_475), .A2(n_476), .B1(n_478), .B2(n_480), .Y(n_474) );
INVx1_ASAP7_75t_L g494 ( .A(n_477), .Y(n_494) );
INVx2_ASAP7_75t_L g480 ( .A(n_481), .Y(n_480) );
AOI21xp5_ASAP7_75t_L g524 ( .A1(n_481), .A2(n_505), .B(n_525), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g482 ( .A1(n_483), .A2(n_491), .B(n_492), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_484), .B(n_487), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_488), .B(n_537), .Y(n_536) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx2_ASAP7_75t_L g513 ( .A(n_490), .Y(n_513) );
NAND3xp33_ASAP7_75t_SL g492 ( .A(n_493), .B(n_498), .C(n_503), .Y(n_492) );
NAND3xp33_ASAP7_75t_SL g493 ( .A(n_494), .B(n_495), .C(n_497), .Y(n_493) );
AND2x2_ASAP7_75t_L g525 ( .A(n_496), .B(n_518), .Y(n_525) );
INVx1_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
NAND3xp33_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .C(n_507), .Y(n_503) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_509), .B(n_534), .Y(n_508) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_510), .A2(n_515), .B(n_522), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_512), .B(n_514), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_513), .Y(n_512) );
NAND4xp25_ASAP7_75t_SL g515 ( .A(n_516), .B(n_517), .C(n_519), .D(n_520), .Y(n_515) );
INVx3_ASAP7_75t_R g517 ( .A(n_518), .Y(n_517) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI21xp5_ASAP7_75t_SL g522 ( .A1(n_523), .A2(n_524), .B(n_526), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g526 ( .A1(n_527), .A2(n_529), .B1(n_531), .B2(n_532), .Y(n_526) );
INVx2_ASAP7_75t_L g529 ( .A(n_530), .Y(n_529) );
INVx2_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
NOR2xp33_ASAP7_75t_L g534 ( .A(n_535), .B(n_540), .Y(n_534) );
AOI21xp5_ASAP7_75t_SL g535 ( .A1(n_536), .A2(n_538), .B(n_539), .Y(n_535) );
AOI22xp5_ASAP7_75t_L g547 ( .A1(n_537), .A2(n_546), .B1(n_548), .B2(n_550), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g540 ( .A(n_541), .B(n_547), .Y(n_540) );
INVx2_ASAP7_75t_SL g548 ( .A(n_549), .Y(n_548) );
CKINVDCx5p33_ASAP7_75t_R g551 ( .A(n_552), .Y(n_551) );
CKINVDCx10_ASAP7_75t_R g552 ( .A(n_553), .Y(n_552) );
BUFx6f_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
BUFx2_ASAP7_75t_L g555 ( .A(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
NAND4xp75_ASAP7_75t_L g558 ( .A(n_559), .B(n_750), .C(n_817), .D(n_859), .Y(n_558) );
NOR3x1_ASAP7_75t_L g559 ( .A(n_560), .B(n_703), .C(n_744), .Y(n_559) );
INVx1_ASAP7_75t_L g560 ( .A(n_561), .Y(n_560) );
AOI211x1_ASAP7_75t_L g561 ( .A1(n_562), .A2(n_601), .B(n_647), .C(n_687), .Y(n_561) );
NOR2xp33_ASAP7_75t_L g562 ( .A(n_563), .B(n_576), .Y(n_562) );
OAI32xp33_ASAP7_75t_L g647 ( .A1(n_563), .A2(n_648), .A3(n_652), .B1(n_655), .B2(n_670), .Y(n_647) );
INVx2_ASAP7_75t_SL g857 ( .A(n_563), .Y(n_857) );
AND2x4_ASAP7_75t_L g874 ( .A(n_563), .B(n_746), .Y(n_874) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
INVx1_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
AND2x2_ASAP7_75t_L g669 ( .A(n_565), .B(n_587), .Y(n_669) );
HB1xp67_ASAP7_75t_L g702 ( .A(n_565), .Y(n_702) );
INVx1_ASAP7_75t_L g708 ( .A(n_565), .Y(n_708) );
INVx1_ASAP7_75t_L g724 ( .A(n_565), .Y(n_724) );
AND2x2_ASAP7_75t_L g732 ( .A(n_565), .B(n_658), .Y(n_732) );
NOR2xp33_ASAP7_75t_L g739 ( .A(n_565), .B(n_587), .Y(n_739) );
OAI21xp5_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B(n_574), .Y(n_566) );
AND2x4_ASAP7_75t_L g624 ( .A(n_574), .B(n_625), .Y(n_624) );
AOI21xp33_ASAP7_75t_L g686 ( .A1(n_574), .A2(n_668), .B(n_685), .Y(n_686) );
O2A1O1Ixp33_ASAP7_75t_L g811 ( .A1(n_576), .A2(n_731), .B(n_812), .C(n_816), .Y(n_811) );
INVx1_ASAP7_75t_L g576 ( .A(n_577), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g654 ( .A(n_578), .Y(n_654) );
OR2x2_ASAP7_75t_L g722 ( .A(n_578), .B(n_723), .Y(n_722) );
NOR2x1_ASAP7_75t_L g778 ( .A(n_578), .B(n_657), .Y(n_778) );
OR2x2_ASAP7_75t_L g578 ( .A(n_579), .B(n_587), .Y(n_578) );
INVx2_ASAP7_75t_SL g696 ( .A(n_579), .Y(n_696) );
AND2x2_ASAP7_75t_L g709 ( .A(n_579), .B(n_700), .Y(n_709) );
AND2x2_ASAP7_75t_L g718 ( .A(n_579), .B(n_701), .Y(n_718) );
AND2x2_ASAP7_75t_L g735 ( .A(n_579), .B(n_698), .Y(n_735) );
BUFx3_ASAP7_75t_L g763 ( .A(n_579), .Y(n_763) );
AND2x2_ASAP7_75t_L g858 ( .A(n_579), .B(n_697), .Y(n_858) );
OR2x2_ASAP7_75t_L g891 ( .A(n_579), .B(n_708), .Y(n_891) );
AO31x2_ASAP7_75t_L g579 ( .A1(n_580), .A2(n_581), .A3(n_584), .B(n_585), .Y(n_579) );
NOR2xp33_ASAP7_75t_L g610 ( .A(n_583), .B(n_611), .Y(n_610) );
INVx3_ASAP7_75t_L g698 ( .A(n_587), .Y(n_698) );
AND2x2_ASAP7_75t_L g707 ( .A(n_587), .B(n_708), .Y(n_707) );
AND2x4_ASAP7_75t_L g587 ( .A(n_588), .B(n_591), .Y(n_587) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI21xp5_ASAP7_75t_L g591 ( .A1(n_592), .A2(n_596), .B(n_600), .Y(n_591) );
AOI21xp5_ASAP7_75t_L g592 ( .A1(n_593), .A2(n_594), .B(n_595), .Y(n_592) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_595), .A2(n_614), .B(n_617), .Y(n_613) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_597), .A2(n_598), .B(n_599), .Y(n_596) );
AOI21xp5_ASAP7_75t_L g660 ( .A1(n_599), .A2(n_661), .B(n_662), .Y(n_660) );
INVxp67_ASAP7_75t_L g601 ( .A(n_602), .Y(n_601) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_620), .Y(n_602) );
AND2x4_ASAP7_75t_L g728 ( .A(n_603), .B(n_729), .Y(n_728) );
AND2x4_ASAP7_75t_L g748 ( .A(n_603), .B(n_749), .Y(n_748) );
NAND2x1_ASAP7_75t_L g827 ( .A(n_603), .B(n_764), .Y(n_827) );
INVx5_ASAP7_75t_L g603 ( .A(n_604), .Y(n_603) );
AND2x4_ASAP7_75t_SL g653 ( .A(n_604), .B(n_654), .Y(n_653) );
AND2x2_ASAP7_75t_L g768 ( .A(n_604), .B(n_763), .Y(n_768) );
AND2x4_ASAP7_75t_L g772 ( .A(n_604), .B(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g797 ( .A(n_604), .B(n_673), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g888 ( .A(n_604), .B(n_620), .Y(n_888) );
BUFx6f_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
INVxp67_ASAP7_75t_L g743 ( .A(n_605), .Y(n_743) );
AO21x1_ASAP7_75t_SL g605 ( .A1(n_606), .A2(n_608), .B(n_612), .Y(n_605) );
AO21x2_ASAP7_75t_L g757 ( .A1(n_606), .A2(n_608), .B(n_612), .Y(n_757) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_607), .Y(n_606) );
OAI21x1_ASAP7_75t_SL g612 ( .A1(n_607), .A2(n_613), .B(n_619), .Y(n_612) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_615), .B(n_616), .Y(n_614) );
INVx1_ASAP7_75t_L g676 ( .A(n_616), .Y(n_676) );
INVx1_ASAP7_75t_L g715 ( .A(n_620), .Y(n_715) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_636), .Y(n_620) );
INVx3_ASAP7_75t_L g712 ( .A(n_621), .Y(n_712) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
INVx2_ASAP7_75t_L g650 ( .A(n_622), .Y(n_650) );
OR2x2_ASAP7_75t_L g690 ( .A(n_622), .B(n_674), .Y(n_690) );
AND2x2_ASAP7_75t_L g766 ( .A(n_622), .B(n_638), .Y(n_766) );
AND2x2_ASAP7_75t_L g884 ( .A(n_622), .B(n_637), .Y(n_884) );
NAND2x1p5_ASAP7_75t_L g622 ( .A(n_623), .B(n_631), .Y(n_622) );
NAND2x1_ASAP7_75t_L g623 ( .A(n_624), .B(n_626), .Y(n_623) );
AOI21x1_ASAP7_75t_L g631 ( .A1(n_624), .A2(n_632), .B(n_635), .Y(n_631) );
O2A1O1Ixp5_ASAP7_75t_L g659 ( .A1(n_624), .A2(n_660), .B(n_663), .C(n_666), .Y(n_659) );
INVx2_ASAP7_75t_SL g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_L g671 ( .A(n_636), .Y(n_671) );
OR2x2_ASAP7_75t_L g736 ( .A(n_636), .B(n_690), .Y(n_736) );
INVx1_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g651 ( .A(n_637), .Y(n_651) );
INVx1_ASAP7_75t_L g692 ( .A(n_637), .Y(n_692) );
INVx2_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
INVxp33_ASAP7_75t_L g730 ( .A(n_638), .Y(n_730) );
OR2x2_ASAP7_75t_L g816 ( .A(n_648), .B(n_810), .Y(n_816) );
INVx1_ASAP7_75t_L g849 ( .A(n_648), .Y(n_849) );
OR2x2_ASAP7_75t_L g648 ( .A(n_649), .B(n_651), .Y(n_648) );
AND2x2_ASAP7_75t_L g773 ( .A(n_649), .B(n_674), .Y(n_773) );
NAND2xp5_ASAP7_75t_L g815 ( .A(n_649), .B(n_714), .Y(n_815) );
INVx2_ASAP7_75t_L g649 ( .A(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g673 ( .A(n_650), .B(n_674), .Y(n_673) );
AND2x2_ASAP7_75t_L g713 ( .A(n_651), .B(n_714), .Y(n_713) );
AND2x2_ASAP7_75t_L g830 ( .A(n_651), .B(n_757), .Y(n_830) );
INVx2_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
AND2x2_ASAP7_75t_L g822 ( .A(n_653), .B(n_823), .Y(n_822) );
AND2x2_ASAP7_75t_L g877 ( .A(n_654), .B(n_657), .Y(n_877) );
INVx1_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g767 ( .A(n_656), .B(n_768), .Y(n_767) );
AND2x2_ASAP7_75t_L g656 ( .A(n_657), .B(n_669), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g761 ( .A(n_657), .B(n_762), .Y(n_761) );
INVx2_ASAP7_75t_L g821 ( .A(n_657), .Y(n_821) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
INVx2_ASAP7_75t_L g701 ( .A(n_658), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g723 ( .A(n_658), .B(n_724), .Y(n_723) );
BUFx2_ASAP7_75t_SL g835 ( .A(n_658), .Y(n_835) );
INVx2_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
NOR2xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .Y(n_666) );
AND2x4_ASAP7_75t_SL g780 ( .A(n_669), .B(n_696), .Y(n_780) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_669), .B(n_763), .Y(n_806) );
AND2x2_ASAP7_75t_L g834 ( .A(n_669), .B(n_835), .Y(n_834) );
OR2x2_ASAP7_75t_L g670 ( .A(n_671), .B(n_672), .Y(n_670) );
AND2x2_ASAP7_75t_L g776 ( .A(n_671), .B(n_673), .Y(n_776) );
AND2x2_ASAP7_75t_L g784 ( .A(n_671), .B(n_785), .Y(n_784) );
INVx1_ASAP7_75t_L g824 ( .A(n_671), .Y(n_824) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
NAND2xp5_ASAP7_75t_L g829 ( .A(n_673), .B(n_830), .Y(n_829) );
INVx1_ASAP7_75t_L g714 ( .A(n_674), .Y(n_714) );
INVx2_ASAP7_75t_L g721 ( .A(n_674), .Y(n_721) );
INVx1_ASAP7_75t_L g787 ( .A(n_674), .Y(n_787) );
AND2x2_ASAP7_75t_L g893 ( .A(n_674), .B(n_756), .Y(n_893) );
AO21x2_ASAP7_75t_L g674 ( .A1(n_675), .A2(n_680), .B(n_686), .Y(n_674) );
NOR2xp67_ASAP7_75t_L g677 ( .A(n_676), .B(n_678), .Y(n_677) );
AOI21xp5_ASAP7_75t_L g680 ( .A1(n_681), .A2(n_684), .B(n_685), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_682), .B(n_683), .Y(n_681) );
AOI21x1_ASAP7_75t_L g687 ( .A1(n_688), .A2(n_691), .B(n_693), .Y(n_687) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
AND2x4_ASAP7_75t_SL g749 ( .A(n_689), .B(n_692), .Y(n_749) );
INVx1_ASAP7_75t_L g689 ( .A(n_690), .Y(n_689) );
INVx2_ASAP7_75t_L g754 ( .A(n_690), .Y(n_754) );
BUFx2_ASAP7_75t_L g691 ( .A(n_692), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_692), .B(n_789), .Y(n_788) );
INVx2_ASAP7_75t_L g845 ( .A(n_692), .Y(n_845) );
OR2x2_ASAP7_75t_L g868 ( .A(n_692), .B(n_815), .Y(n_868) );
OR2x6_ASAP7_75t_L g693 ( .A(n_694), .B(n_699), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g861 ( .A(n_695), .Y(n_861) );
AND2x2_ASAP7_75t_L g695 ( .A(n_696), .B(n_697), .Y(n_695) );
AND2x2_ASAP7_75t_L g840 ( .A(n_696), .B(n_803), .Y(n_840) );
INVx1_ASAP7_75t_L g760 ( .A(n_697), .Y(n_760) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_698), .B(n_701), .Y(n_747) );
INVx1_ASAP7_75t_L g863 ( .A(n_699), .Y(n_863) );
OR2x2_ASAP7_75t_L g699 ( .A(n_700), .B(n_702), .Y(n_699) );
INVx1_ASAP7_75t_L g741 ( .A(n_700), .Y(n_741) );
AND2x2_ASAP7_75t_L g793 ( .A(n_700), .B(n_780), .Y(n_793) );
INVx2_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
NAND2x1_ASAP7_75t_L g703 ( .A(n_704), .B(n_725), .Y(n_703) );
OA222x2_ASAP7_75t_L g704 ( .A1(n_705), .A2(n_710), .B1(n_715), .B2(n_716), .C1(n_719), .C2(n_722), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
OAI21xp33_ASAP7_75t_L g878 ( .A1(n_706), .A2(n_879), .B(n_881), .Y(n_878) );
AND2x4_ASAP7_75t_L g706 ( .A(n_707), .B(n_709), .Y(n_706) );
AND2x4_ASAP7_75t_L g717 ( .A(n_707), .B(n_718), .Y(n_717) );
NAND2x1_ASAP7_75t_L g740 ( .A(n_707), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_L g825 ( .A1(n_707), .A2(n_826), .B(n_828), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g774 ( .A1(n_710), .A2(n_775), .B1(n_777), .B2(n_779), .Y(n_774) );
INVx2_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_712), .B(n_713), .Y(n_711) );
NAND2x1p5_ASAP7_75t_L g742 ( .A(n_712), .B(n_743), .Y(n_742) );
INVx4_ASAP7_75t_L g716 ( .A(n_717), .Y(n_716) );
AND2x4_ASAP7_75t_L g738 ( .A(n_718), .B(n_739), .Y(n_738) );
AOI22xp5_ASAP7_75t_L g894 ( .A1(n_718), .A2(n_828), .B1(n_895), .B2(n_896), .Y(n_894) );
NOR2xp33_ASAP7_75t_SL g854 ( .A(n_719), .B(n_845), .Y(n_854) );
INVx1_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2x1_ASAP7_75t_L g838 ( .A(n_720), .B(n_764), .Y(n_838) );
INVx1_ASAP7_75t_L g720 ( .A(n_721), .Y(n_720) );
AND2x2_ASAP7_75t_L g729 ( .A(n_721), .B(n_730), .Y(n_729) );
AND2x2_ASAP7_75t_L g789 ( .A(n_721), .B(n_756), .Y(n_789) );
OR2x2_ASAP7_75t_L g810 ( .A(n_721), .B(n_756), .Y(n_810) );
INVx2_ASAP7_75t_L g803 ( .A(n_723), .Y(n_803) );
INVx1_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
OAI322xp33_ASAP7_75t_L g726 ( .A1(n_727), .A2(n_731), .A3(n_733), .B1(n_736), .B2(n_737), .C1(n_740), .C2(n_742), .Y(n_726) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
AND2x2_ASAP7_75t_L g755 ( .A(n_730), .B(n_756), .Y(n_755) );
OR2x2_ASAP7_75t_L g865 ( .A(n_731), .B(n_866), .Y(n_865) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
AND2x4_ASAP7_75t_L g791 ( .A(n_732), .B(n_735), .Y(n_791) );
AO221x1_ASAP7_75t_L g860 ( .A1(n_733), .A2(n_857), .B1(n_861), .B2(n_862), .C(n_864), .Y(n_860) );
INVx1_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
AND2x2_ASAP7_75t_L g846 ( .A(n_735), .B(n_803), .Y(n_846) );
AOI21xp5_ASAP7_75t_SL g770 ( .A1(n_737), .A2(n_765), .B(n_771), .Y(n_770) );
INVx4_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
AOI22xp5_ASAP7_75t_L g853 ( .A1(n_738), .A2(n_784), .B1(n_854), .B2(n_855), .Y(n_853) );
AND2x2_ASAP7_75t_L g895 ( .A(n_741), .B(n_858), .Y(n_895) );
AND2x2_ASAP7_75t_L g744 ( .A(n_745), .B(n_748), .Y(n_744) );
HB1xp67_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx2_ASAP7_75t_L g746 ( .A(n_747), .Y(n_746) );
OAI21xp5_ASAP7_75t_L g841 ( .A1(n_749), .A2(n_842), .B(n_846), .Y(n_841) );
INVx2_ASAP7_75t_L g851 ( .A(n_749), .Y(n_851) );
AOI22xp5_ASAP7_75t_L g870 ( .A1(n_749), .A2(n_871), .B1(n_872), .B2(n_875), .Y(n_870) );
NOR3x1_ASAP7_75t_L g750 ( .A(n_751), .B(n_781), .C(n_804), .Y(n_750) );
NAND2xp5_ASAP7_75t_L g751 ( .A(n_752), .B(n_769), .Y(n_751) );
AOI22xp5_ASAP7_75t_L g752 ( .A1(n_753), .A2(n_758), .B1(n_764), .B2(n_767), .Y(n_752) );
AND2x2_ASAP7_75t_L g753 ( .A(n_754), .B(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g800 ( .A(n_754), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g799 ( .A(n_755), .B(n_800), .Y(n_799) );
NOR2xp33_ASAP7_75t_L g848 ( .A(n_755), .B(n_849), .Y(n_848) );
NAND2xp5_ASAP7_75t_L g897 ( .A(n_755), .B(n_898), .Y(n_897) );
INVx2_ASAP7_75t_L g814 ( .A(n_756), .Y(n_814) );
INVx3_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_757), .B(n_787), .Y(n_786) );
INVx2_ASAP7_75t_SL g758 ( .A(n_759), .Y(n_758) );
OR2x2_ASAP7_75t_L g759 ( .A(n_760), .B(n_761), .Y(n_759) );
NAND2xp5_ASAP7_75t_L g802 ( .A(n_760), .B(n_803), .Y(n_802) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_761), .Y(n_880) );
INVx2_ASAP7_75t_L g762 ( .A(n_763), .Y(n_762) );
INVx1_ASAP7_75t_L g866 ( .A(n_763), .Y(n_866) );
HB1xp67_ASAP7_75t_L g873 ( .A(n_763), .Y(n_873) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_764), .B(n_809), .Y(n_808) );
INVx6_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
INVx4_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
AND2x2_ASAP7_75t_L g892 ( .A(n_766), .B(n_893), .Y(n_892) );
NAND2xp5_ASAP7_75t_L g852 ( .A(n_768), .B(n_834), .Y(n_852) );
NOR2xp67_ASAP7_75t_SL g769 ( .A(n_770), .B(n_774), .Y(n_769) );
INVx2_ASAP7_75t_L g771 ( .A(n_772), .Y(n_771) );
INVx2_ASAP7_75t_SL g775 ( .A(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g777 ( .A(n_778), .Y(n_777) );
INVx2_ASAP7_75t_L g779 ( .A(n_780), .Y(n_779) );
OAI21xp5_ASAP7_75t_L g781 ( .A1(n_782), .A2(n_790), .B(n_792), .Y(n_781) );
AND2x2_ASAP7_75t_L g782 ( .A(n_783), .B(n_788), .Y(n_782) );
INVx1_ASAP7_75t_L g783 ( .A(n_784), .Y(n_783) );
INVx1_ASAP7_75t_L g844 ( .A(n_785), .Y(n_844) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
INVx1_ASAP7_75t_L g795 ( .A(n_789), .Y(n_795) );
INVxp67_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
AOI22xp5_ASAP7_75t_L g792 ( .A1(n_793), .A2(n_794), .B1(n_798), .B2(n_801), .Y(n_792) );
INVx2_ASAP7_75t_L g850 ( .A(n_793), .Y(n_850) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_795), .B(n_796), .Y(n_794) );
INVx2_ASAP7_75t_SL g796 ( .A(n_797), .Y(n_796) );
INVxp67_ASAP7_75t_SL g798 ( .A(n_799), .Y(n_798) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
AO21x1_ASAP7_75t_L g804 ( .A1(n_805), .A2(n_807), .B(n_811), .Y(n_804) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVxp67_ASAP7_75t_SL g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g809 ( .A(n_810), .Y(n_809) );
INVx1_ASAP7_75t_L g871 ( .A(n_812), .Y(n_871) );
OR2x2_ASAP7_75t_L g812 ( .A(n_813), .B(n_815), .Y(n_812) );
OR2x2_ASAP7_75t_L g882 ( .A(n_813), .B(n_883), .Y(n_882) );
INVx2_ASAP7_75t_L g813 ( .A(n_814), .Y(n_813) );
BUFx2_ASAP7_75t_SL g837 ( .A(n_814), .Y(n_837) );
OR2x2_ASAP7_75t_L g836 ( .A(n_815), .B(n_837), .Y(n_836) );
INVx1_ASAP7_75t_L g898 ( .A(n_815), .Y(n_898) );
NOR2x1_ASAP7_75t_L g817 ( .A(n_818), .B(n_847), .Y(n_817) );
NAND4xp75_ASAP7_75t_L g818 ( .A(n_819), .B(n_825), .C(n_831), .D(n_841), .Y(n_818) );
NAND2xp5_ASAP7_75t_L g819 ( .A(n_820), .B(n_822), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g823 ( .A(n_824), .Y(n_823) );
INVx1_ASAP7_75t_L g826 ( .A(n_827), .Y(n_826) );
INVx1_ASAP7_75t_L g828 ( .A(n_829), .Y(n_828) );
INVx1_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_836), .B1(n_838), .B2(n_839), .Y(n_832) );
INVx2_ASAP7_75t_L g833 ( .A(n_834), .Y(n_833) );
INVx2_ASAP7_75t_L g839 ( .A(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g842 ( .A(n_843), .Y(n_842) );
OR2x2_ASAP7_75t_L g843 ( .A(n_844), .B(n_845), .Y(n_843) );
AOI22xp5_ASAP7_75t_L g886 ( .A1(n_846), .A2(n_887), .B1(n_889), .B2(n_892), .Y(n_886) );
OAI221xp5_ASAP7_75t_L g847 ( .A1(n_848), .A2(n_850), .B1(n_851), .B2(n_852), .C(n_853), .Y(n_847) );
INVx1_ASAP7_75t_L g855 ( .A(n_856), .Y(n_855) );
NAND2xp5_ASAP7_75t_L g856 ( .A(n_857), .B(n_858), .Y(n_856) );
AOI211x1_ASAP7_75t_L g859 ( .A1(n_860), .A2(n_867), .B(n_869), .C(n_885), .Y(n_859) );
INVx1_ASAP7_75t_L g862 ( .A(n_863), .Y(n_862) );
INVx2_ASAP7_75t_L g864 ( .A(n_865), .Y(n_864) );
INVx1_ASAP7_75t_L g867 ( .A(n_868), .Y(n_867) );
NAND2xp5_ASAP7_75t_SL g869 ( .A(n_870), .B(n_878), .Y(n_869) );
AND2x4_ASAP7_75t_L g872 ( .A(n_873), .B(n_874), .Y(n_872) );
INVx1_ASAP7_75t_L g875 ( .A(n_876), .Y(n_875) );
INVx2_ASAP7_75t_SL g876 ( .A(n_877), .Y(n_876) );
INVxp67_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g881 ( .A(n_882), .Y(n_881) );
INVx1_ASAP7_75t_L g883 ( .A(n_884), .Y(n_883) );
NAND2xp5_ASAP7_75t_SL g885 ( .A(n_886), .B(n_894), .Y(n_885) );
INVx2_ASAP7_75t_L g887 ( .A(n_888), .Y(n_887) );
INVx1_ASAP7_75t_L g889 ( .A(n_890), .Y(n_889) );
HB1xp67_ASAP7_75t_L g890 ( .A(n_891), .Y(n_890) );
INVxp67_ASAP7_75t_SL g896 ( .A(n_897), .Y(n_896) );
INVxp67_ASAP7_75t_L g902 ( .A(n_899), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g905 ( .A1(n_906), .A2(n_908), .B(n_931), .Y(n_905) );
INVx3_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
AOI21xp5_ASAP7_75t_L g908 ( .A1(n_909), .A2(n_918), .B(n_926), .Y(n_908) );
INVxp67_ASAP7_75t_L g917 ( .A(n_911), .Y(n_917) );
CKINVDCx5p33_ASAP7_75t_R g915 ( .A(n_912), .Y(n_915) );
INVx1_ASAP7_75t_L g918 ( .A(n_919), .Y(n_918) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
INVx2_ASAP7_75t_SL g920 ( .A(n_921), .Y(n_920) );
INVx2_ASAP7_75t_L g921 ( .A(n_922), .Y(n_921) );
INVx2_ASAP7_75t_SL g922 ( .A(n_923), .Y(n_922) );
INVx2_ASAP7_75t_L g930 ( .A(n_923), .Y(n_930) );
NOR2x1p5_ASAP7_75t_L g923 ( .A(n_924), .B(n_925), .Y(n_923) );
CKINVDCx8_ASAP7_75t_R g927 ( .A(n_928), .Y(n_927) );
BUFx6f_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
BUFx3_ASAP7_75t_L g929 ( .A(n_930), .Y(n_929) );
INVx1_ASAP7_75t_L g932 ( .A(n_933), .Y(n_932) );
BUFx3_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
BUFx3_ASAP7_75t_L g934 ( .A(n_935), .Y(n_934) );
AND2x2_ASAP7_75t_L g940 ( .A(n_936), .B(n_941), .Y(n_940) );
INVx1_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
INVx4_ASAP7_75t_SL g938 ( .A(n_939), .Y(n_938) );
BUFx6f_ASAP7_75t_L g939 ( .A(n_940), .Y(n_939) );
BUFx6f_ASAP7_75t_L g948 ( .A(n_940), .Y(n_948) );
INVx1_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx1_ASAP7_75t_L g942 ( .A(n_943), .Y(n_942) );
INVx1_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
INVx1_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
CKINVDCx5p33_ASAP7_75t_R g947 ( .A(n_948), .Y(n_947) );
endmodule