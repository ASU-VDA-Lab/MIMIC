module fake_jpeg_19770_n_94 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_94);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_94;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx13_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_1),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_4),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_2),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_18),
.B(n_12),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_23),
.B(n_21),
.Y(n_38)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_18),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_26),
.B(n_28),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g27 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_27),
.A2(n_12),
.B1(n_21),
.B2(n_20),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_6),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_SL g29 ( 
.A(n_20),
.B(n_0),
.Y(n_29)
);

AND2x2_ASAP7_75t_L g36 ( 
.A(n_29),
.B(n_21),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g31 ( 
.A(n_23),
.B(n_22),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_31),
.B(n_36),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_32),
.A2(n_33),
.B1(n_13),
.B2(n_14),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g33 ( 
.A(n_24),
.B(n_14),
.C(n_13),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_30),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g40 ( 
.A(n_38),
.B(n_16),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_47),
.C(n_17),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_31),
.B(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_42),
.B(n_45),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_39),
.A2(n_13),
.B1(n_26),
.B2(n_25),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_43),
.A2(n_50),
.B1(n_16),
.B2(n_11),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_49),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_31),
.B(n_15),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_35),
.Y(n_46)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_L g47 ( 
.A1(n_36),
.A2(n_19),
.B(n_16),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_39),
.A2(n_33),
.B1(n_34),
.B2(n_25),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g54 ( 
.A1(n_48),
.A2(n_34),
.B1(n_37),
.B2(n_16),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_30),
.B1(n_26),
.B2(n_17),
.Y(n_50)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_37),
.Y(n_51)
);

NAND3xp33_ASAP7_75t_L g59 ( 
.A(n_51),
.B(n_5),
.C(n_7),
.Y(n_59)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_35),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_52),
.B(n_3),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_53),
.B(n_45),
.C(n_42),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_54),
.A2(n_61),
.B1(n_63),
.B2(n_9),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_62),
.Y(n_67)
);

NOR2x1_ASAP7_75t_L g56 ( 
.A(n_41),
.B(n_11),
.Y(n_56)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_56),
.A2(n_59),
.B(n_44),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_49),
.A2(n_11),
.B1(n_3),
.B2(n_1),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_63)
);

MAJx2_ASAP7_75t_L g64 ( 
.A(n_53),
.B(n_40),
.C(n_47),
.Y(n_64)
);

XNOR2xp5_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_71),
.Y(n_77)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_66),
.B(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_58),
.B(n_41),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_69),
.B(n_70),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_58),
.A2(n_50),
.B(n_52),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_46),
.C(n_8),
.Y(n_71)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_68),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_74),
.B(n_60),
.Y(n_81)
);

BUFx2_ASAP7_75t_L g76 ( 
.A(n_67),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_75),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_63),
.B1(n_54),
.B2(n_64),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_80),
.B(n_81),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_56),
.B1(n_62),
.B2(n_57),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g86 ( 
.A(n_82),
.B(n_83),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_77),
.B(n_78),
.Y(n_84)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_84),
.B(n_77),
.C(n_79),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g90 ( 
.A(n_85),
.B(n_86),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g88 ( 
.A1(n_87),
.A2(n_82),
.B(n_84),
.Y(n_88)
);

BUFx24_ASAP7_75t_SL g91 ( 
.A(n_88),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_76),
.Y(n_89)
);

BUFx2_ASAP7_75t_L g92 ( 
.A(n_89),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g93 ( 
.A1(n_91),
.A2(n_90),
.B(n_92),
.Y(n_93)
);

BUFx24_ASAP7_75t_SL g94 ( 
.A(n_93),
.Y(n_94)
);


endmodule