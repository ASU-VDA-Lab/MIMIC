module fake_jpeg_26583_n_116 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_116);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_10;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_L g9 ( 
.A(n_0),
.Y(n_9)
);

INVx1_ASAP7_75t_L g10 ( 
.A(n_8),
.Y(n_10)
);

BUFx12f_ASAP7_75t_L g11 ( 
.A(n_6),
.Y(n_11)
);

BUFx5_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx16_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVx11_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_11),
.Y(n_18)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_19),
.B(n_20),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_15),
.B(n_0),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_21),
.B(n_17),
.Y(n_33)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_22),
.B(n_17),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_11),
.Y(n_23)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

INVx8_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_24),
.Y(n_26)
);

AOI22xp33_ASAP7_75t_SL g25 ( 
.A1(n_18),
.A2(n_15),
.B1(n_9),
.B2(n_10),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_25),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g27 ( 
.A1(n_22),
.A2(n_16),
.B1(n_17),
.B2(n_14),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_27),
.A2(n_32),
.B1(n_24),
.B2(n_13),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g42 ( 
.A1(n_28),
.A2(n_33),
.B(n_13),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g32 ( 
.A1(n_22),
.A2(n_18),
.B1(n_24),
.B2(n_16),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_29),
.B(n_20),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_34),
.B(n_41),
.Y(n_44)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_36),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_25),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_37),
.A2(n_30),
.B1(n_26),
.B2(n_9),
.Y(n_53)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_39),
.Y(n_50)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_26),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_29),
.B(n_20),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_42),
.A2(n_28),
.B(n_9),
.Y(n_47)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_23),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_36),
.A2(n_32),
.B1(n_28),
.B2(n_31),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_45),
.A2(n_48),
.B1(n_51),
.B2(n_53),
.Y(n_55)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

MAJx2_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_52),
.C(n_51),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_40),
.A2(n_32),
.B1(n_37),
.B2(n_41),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_34),
.A2(n_26),
.B1(n_24),
.B2(n_27),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_SL g52 ( 
.A(n_42),
.B(n_33),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_50),
.Y(n_56)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_56),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_46),
.Y(n_58)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_58),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_44),
.B(n_10),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_59),
.B(n_1),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_60),
.A2(n_63),
.B1(n_45),
.B2(n_52),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_53),
.Y(n_62)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_62),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_48),
.A2(n_38),
.B1(n_35),
.B2(n_39),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g82 ( 
.A(n_65),
.B(n_1),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_SL g80 ( 
.A1(n_67),
.A2(n_21),
.B(n_23),
.Y(n_80)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_68),
.B(n_70),
.Y(n_77)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_57),
.Y(n_70)
);

AO22x1_ASAP7_75t_SL g73 ( 
.A1(n_55),
.A2(n_43),
.B1(n_38),
.B2(n_35),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_55),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_71),
.B(n_56),
.Y(n_74)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_74),
.Y(n_87)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_75),
.B(n_79),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_67),
.B(n_60),
.C(n_54),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_64),
.C(n_69),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_78),
.A2(n_80),
.B(n_81),
.Y(n_90)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

XNOR2x1_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_21),
.Y(n_81)
);

NAND3xp33_ASAP7_75t_L g84 ( 
.A(n_82),
.B(n_1),
.C(n_2),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_66),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_83),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g96 ( 
.A1(n_84),
.A2(n_88),
.B(n_89),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_86),
.B(n_87),
.C(n_85),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_80),
.A2(n_68),
.B1(n_72),
.B2(n_39),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g89 ( 
.A1(n_77),
.A2(n_26),
.B1(n_43),
.B2(n_30),
.Y(n_89)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_76),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_23),
.C(n_12),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_93),
.B(n_94),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_81),
.C(n_30),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_23),
.C(n_19),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_95),
.B(n_19),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_14),
.B1(n_12),
.B2(n_4),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g100 ( 
.A1(n_97),
.A2(n_14),
.B1(n_12),
.B2(n_5),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g98 ( 
.A1(n_91),
.A2(n_2),
.B(n_3),
.Y(n_98)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_98),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_100),
.A2(n_3),
.B1(n_5),
.B2(n_7),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_101),
.B(n_23),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_92),
.C(n_96),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_104),
.B(n_105),
.C(n_102),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_99),
.A2(n_3),
.B(n_4),
.Y(n_105)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_106),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_107),
.B(n_103),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_108),
.B(n_109),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g111 ( 
.A1(n_110),
.A2(n_7),
.B(n_8),
.Y(n_111)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_111),
.Y(n_113)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_113),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_L g115 ( 
.A1(n_114),
.A2(n_112),
.B(n_7),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_8),
.Y(n_116)
);


endmodule