module fake_jpeg_28375_n_355 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_355);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_355;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_SL g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx12f_ASAP7_75t_L g22 ( 
.A(n_14),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_1),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx2_ASAP7_75t_SL g26 ( 
.A(n_0),
.Y(n_26)
);

INVx11_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx16_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_1),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_4),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_22),
.Y(n_38)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_38),
.Y(n_68)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_39),
.Y(n_81)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g71 ( 
.A(n_40),
.Y(n_71)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_22),
.Y(n_41)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_22),
.B(n_12),
.Y(n_42)
);

NOR3xp33_ASAP7_75t_L g77 ( 
.A(n_42),
.B(n_30),
.C(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_16),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_44),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_23),
.Y(n_45)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_45),
.Y(n_79)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_46),
.Y(n_91)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_34),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_27),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_48),
.B(n_18),
.Y(n_93)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_34),
.Y(n_49)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_49),
.Y(n_60)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_50),
.Y(n_80)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_27),
.Y(n_51)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_51),
.Y(n_69)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_53),
.B(n_30),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_23),
.Y(n_54)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_54),
.Y(n_66)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_23),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_23),
.Y(n_56)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_56),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_45),
.A2(n_56),
.B1(n_55),
.B2(n_26),
.Y(n_57)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_57),
.A2(n_59),
.B1(n_61),
.B2(n_74),
.Y(n_125)
);

INVx4_ASAP7_75t_SL g58 ( 
.A(n_46),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_58),
.B(n_77),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_45),
.A2(n_26),
.B1(n_17),
.B2(n_35),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_38),
.A2(n_26),
.B1(n_17),
.B2(n_35),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_40),
.A2(n_26),
.B1(n_17),
.B2(n_25),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_62),
.Y(n_95)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_63),
.B(n_31),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_39),
.A2(n_17),
.B1(n_37),
.B2(n_25),
.Y(n_65)
);

CKINVDCx14_ASAP7_75t_R g102 ( 
.A(n_65),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_41),
.A2(n_37),
.B1(n_33),
.B2(n_24),
.Y(n_67)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_67),
.Y(n_123)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_70),
.Y(n_96)
);

NAND2xp33_ASAP7_75t_SL g73 ( 
.A(n_49),
.B(n_29),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g114 ( 
.A1(n_73),
.A2(n_78),
.B(n_71),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_44),
.A2(n_33),
.B1(n_19),
.B2(n_20),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_19),
.B1(n_20),
.B2(n_18),
.Y(n_75)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_75),
.Y(n_133)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_82),
.Y(n_104)
);

INVx6_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

BUFx2_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_50),
.A2(n_18),
.B1(n_28),
.B2(n_29),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g98 ( 
.A(n_84),
.Y(n_98)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_49),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_86),
.B(n_87),
.Y(n_110)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_52),
.Y(n_88)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_88),
.Y(n_122)
);

INVx3_ASAP7_75t_L g90 ( 
.A(n_54),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_90),
.B(n_92),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_53),
.B(n_28),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_93),
.B(n_21),
.Y(n_124)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_97),
.Y(n_137)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_60),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_108),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_61),
.B(n_42),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_100),
.B(n_116),
.Y(n_134)
);

BUFx24_ASAP7_75t_L g101 ( 
.A(n_68),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_101),
.Y(n_141)
);

AO22x1_ASAP7_75t_SL g103 ( 
.A1(n_73),
.A2(n_31),
.B1(n_29),
.B2(n_28),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_103),
.A2(n_111),
.B1(n_91),
.B2(n_82),
.Y(n_146)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_57),
.Y(n_105)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_105),
.Y(n_142)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_59),
.Y(n_106)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_106),
.Y(n_143)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_88),
.Y(n_107)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_68),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_64),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_109),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_L g111 ( 
.A1(n_66),
.A2(n_48),
.B1(n_31),
.B2(n_36),
.Y(n_111)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_58),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_112),
.B(n_119),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_64),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_113),
.Y(n_152)
);

AOI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_114),
.A2(n_79),
.B(n_89),
.Y(n_139)
);

OR2x2_ASAP7_75t_L g115 ( 
.A(n_76),
.B(n_36),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g149 ( 
.A1(n_115),
.A2(n_91),
.B(n_69),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_76),
.B(n_81),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_88),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

INVx13_ASAP7_75t_L g119 ( 
.A(n_60),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_81),
.B(n_31),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_120),
.B(n_130),
.Y(n_150)
);

CKINVDCx14_ASAP7_75t_R g155 ( 
.A(n_124),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_72),
.B(n_36),
.Y(n_126)
);

XNOR2xp5_ASAP7_75t_L g138 ( 
.A(n_126),
.B(n_21),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_66),
.A2(n_83),
.B1(n_79),
.B2(n_90),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_127),
.A2(n_69),
.B1(n_86),
.B2(n_3),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g128 ( 
.A(n_60),
.Y(n_128)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_128),
.Y(n_164)
);

INVx4_ASAP7_75t_L g129 ( 
.A(n_80),
.Y(n_129)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_129),
.Y(n_165)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_70),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_131),
.B(n_132),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_71),
.B(n_21),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_126),
.B(n_85),
.C(n_63),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_140),
.C(n_144),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_138),
.B(n_115),
.Y(n_177)
);

OAI21xp5_ASAP7_75t_SL g185 ( 
.A1(n_139),
.A2(n_151),
.B(n_96),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_114),
.B(n_85),
.C(n_89),
.Y(n_140)
);

MAJx2_ASAP7_75t_L g144 ( 
.A(n_100),
.B(n_94),
.C(n_102),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_146),
.A2(n_161),
.B1(n_129),
.B2(n_109),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_149),
.A2(n_157),
.B(n_115),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_95),
.A2(n_0),
.B(n_1),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_125),
.B(n_80),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_153),
.B(n_138),
.C(n_140),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_154),
.A2(n_159),
.B1(n_122),
.B2(n_99),
.Y(n_195)
);

AND2x6_ASAP7_75t_L g156 ( 
.A(n_123),
.B(n_9),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_156),
.B(n_103),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g157 ( 
.A1(n_95),
.A2(n_133),
.B(n_98),
.C(n_106),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_105),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_98),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_125),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_161)
);

OA22x2_ASAP7_75t_L g162 ( 
.A1(n_133),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_162),
.B(n_2),
.Y(n_189)
);

BUFx5_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_166),
.B(n_175),
.Y(n_210)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_150),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_167),
.B(n_173),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_134),
.B(n_116),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_168),
.B(n_171),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_169),
.A2(n_170),
.B1(n_188),
.B2(n_16),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_161),
.A2(n_103),
.B1(n_113),
.B2(n_121),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_134),
.B(n_137),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_172),
.A2(n_189),
.B(n_143),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_137),
.B(n_110),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_150),
.B(n_97),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_174),
.B(n_176),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_153),
.B(n_120),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_177),
.B(n_198),
.C(n_142),
.Y(n_204)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_157),
.A2(n_131),
.B(n_130),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g223 ( 
.A1(n_178),
.A2(n_179),
.B(n_185),
.Y(n_223)
);

AOI21xp5_ASAP7_75t_L g179 ( 
.A1(n_149),
.A2(n_96),
.B(n_112),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_155),
.B(n_101),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_180),
.B(n_181),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_163),
.B(n_101),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_135),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_182),
.B(n_186),
.Y(n_227)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_163),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_108),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_187),
.B(n_190),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_146),
.A2(n_111),
.B1(n_122),
.B2(n_118),
.Y(n_188)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_145),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_147),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_191),
.B(n_193),
.Y(n_202)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_164),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_200),
.Y(n_230)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_152),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_159),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g234 ( 
.A(n_194),
.B(n_197),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_143),
.B1(n_165),
.B2(n_158),
.Y(n_208)
);

OAI21xp33_ASAP7_75t_L g196 ( 
.A1(n_151),
.A2(n_144),
.B(n_139),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g203 ( 
.A(n_196),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_154),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_148),
.B(n_101),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g224 ( 
.A(n_199),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_142),
.B(n_11),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_141),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g218 ( 
.A(n_201),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_204),
.B(n_215),
.C(n_228),
.Y(n_236)
);

OAI21xp5_ASAP7_75t_L g261 ( 
.A1(n_206),
.A2(n_8),
.B(n_229),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_208),
.A2(n_193),
.B1(n_191),
.B2(n_182),
.Y(n_246)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_199),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_209),
.B(n_213),
.Y(n_235)
);

OAI32xp33_ASAP7_75t_L g211 ( 
.A1(n_171),
.A2(n_176),
.A3(n_167),
.B1(n_187),
.B2(n_168),
.Y(n_211)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

AND2x2_ASAP7_75t_SL g212 ( 
.A(n_178),
.B(n_158),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_212),
.A2(n_6),
.B(n_7),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_180),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_183),
.B(n_148),
.C(n_165),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_197),
.A2(n_156),
.B1(n_162),
.B2(n_141),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_216),
.A2(n_221),
.B1(n_222),
.B2(n_225),
.Y(n_247)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_181),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_217),
.B(n_219),
.Y(n_240)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_174),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_162),
.B1(n_104),
.B2(n_118),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g243 ( 
.A1(n_220),
.A2(n_226),
.B1(n_189),
.B2(n_184),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_194),
.A2(n_162),
.B1(n_118),
.B2(n_104),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_195),
.A2(n_119),
.B1(n_128),
.B2(n_10),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_170),
.A2(n_189),
.B1(n_188),
.B2(n_186),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_13),
.C(n_12),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_198),
.B(n_13),
.C(n_11),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_184),
.C(n_200),
.Y(n_244)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_173),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_232),
.B(n_190),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_204),
.B(n_177),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_237),
.B(n_255),
.Y(n_283)
);

AOI21xp5_ASAP7_75t_L g239 ( 
.A1(n_223),
.A2(n_185),
.B(n_172),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_239),
.A2(n_253),
.B(n_256),
.Y(n_262)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_202),
.Y(n_241)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_241),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_202),
.Y(n_242)
);

CKINVDCx16_ASAP7_75t_R g272 ( 
.A(n_242),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g271 ( 
.A1(n_243),
.A2(n_251),
.B1(n_259),
.B2(n_222),
.Y(n_271)
);

MAJx2_ASAP7_75t_L g278 ( 
.A(n_244),
.B(n_228),
.C(n_231),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_166),
.Y(n_245)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_245),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_246),
.A2(n_212),
.B1(n_217),
.B2(n_224),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_230),
.B(n_192),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_248),
.B(n_252),
.Y(n_263)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_250),
.Y(n_269)
);

AOI22xp33_ASAP7_75t_SL g251 ( 
.A1(n_209),
.A2(n_201),
.B1(n_179),
.B2(n_5),
.Y(n_251)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_210),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_223),
.A2(n_2),
.B(n_3),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_205),
.B(n_6),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_254),
.B(n_258),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_215),
.B(n_11),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_13),
.C(n_7),
.Y(n_257)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_257),
.B(n_253),
.Y(n_268)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_234),
.Y(n_258)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_208),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_226),
.A2(n_8),
.B1(n_220),
.B2(n_212),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_260),
.A2(n_218),
.B1(n_207),
.B2(n_8),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g276 ( 
.A1(n_261),
.A2(n_256),
.B(n_229),
.Y(n_276)
);

OAI22x1_ASAP7_75t_L g264 ( 
.A1(n_243),
.A2(n_212),
.B1(n_216),
.B2(n_221),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g286 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_277),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_247),
.A2(n_233),
.B1(n_203),
.B2(n_219),
.Y(n_266)
);

AOI21xp33_ASAP7_75t_L g267 ( 
.A1(n_252),
.A2(n_232),
.B(n_206),
.Y(n_267)
);

BUFx12f_ASAP7_75t_SL g300 ( 
.A(n_267),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_268),
.B(n_282),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_237),
.B(n_211),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_270),
.B(n_236),
.Y(n_284)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_271),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g296 ( 
.A1(n_276),
.A2(n_261),
.B(n_258),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_247),
.A2(n_225),
.B1(n_214),
.B2(n_227),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_278),
.B(n_236),
.C(n_283),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g279 ( 
.A(n_239),
.B(n_207),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_SL g301 ( 
.A(n_279),
.B(n_240),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_214),
.B1(n_227),
.B2(n_205),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_280),
.B(n_249),
.Y(n_288)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_281),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_250),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_289),
.Y(n_314)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_287),
.B(n_288),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_283),
.B(n_255),
.C(n_238),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_290),
.B(n_291),
.C(n_268),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_270),
.B(n_278),
.C(n_279),
.Y(n_291)
);

XNOR2xp5_ASAP7_75t_L g293 ( 
.A(n_266),
.B(n_238),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_296),
.Y(n_317)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_269),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_297),
.Y(n_315)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_269),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_263),
.Y(n_298)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_298),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g299 ( 
.A(n_265),
.Y(n_299)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_299),
.Y(n_312)
);

XNOR2x1_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_264),
.Y(n_304)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_274),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_302),
.B(n_235),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_307),
.Y(n_323)
);

INVx2_ASAP7_75t_L g306 ( 
.A(n_300),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_306),
.B(n_313),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_275),
.C(n_273),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_314),
.C(n_307),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_299),
.A2(n_246),
.B1(n_281),
.B2(n_277),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_309),
.B(n_292),
.Y(n_321)
);

INVxp33_ASAP7_75t_L g310 ( 
.A(n_287),
.Y(n_310)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_310),
.Y(n_330)
);

NOR2xp67_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_262),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_311),
.B(n_262),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g316 ( 
.A(n_288),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g325 ( 
.A(n_316),
.B(n_241),
.Y(n_325)
);

A2O1A1Ixp33_ASAP7_75t_L g318 ( 
.A1(n_312),
.A2(n_240),
.B(n_294),
.C(n_285),
.Y(n_318)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_318),
.Y(n_336)
);

A2O1A1Ixp33_ASAP7_75t_L g319 ( 
.A1(n_304),
.A2(n_294),
.B(n_293),
.C(n_301),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_319),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_308),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_320),
.B(n_325),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_321),
.A2(n_315),
.B1(n_290),
.B2(n_276),
.Y(n_335)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_322),
.B(n_327),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_305),
.B(n_280),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_326),
.B(n_328),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_314),
.B(n_284),
.C(n_306),
.Y(n_328)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_291),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_329),
.B(n_317),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g333 ( 
.A1(n_330),
.A2(n_292),
.B1(n_303),
.B2(n_310),
.Y(n_333)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_333),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g334 ( 
.A1(n_324),
.A2(n_309),
.B1(n_260),
.B2(n_296),
.Y(n_334)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_334),
.Y(n_342)
);

AOI21xp5_ASAP7_75t_L g343 ( 
.A1(n_335),
.A2(n_319),
.B(n_323),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g346 ( 
.A(n_339),
.B(n_244),
.Y(n_346)
);

NOR4xp25_ASAP7_75t_L g340 ( 
.A(n_337),
.B(n_286),
.C(n_328),
.D(n_318),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g348 ( 
.A1(n_340),
.A2(n_345),
.B(n_346),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_343),
.B(n_335),
.C(n_336),
.Y(n_349)
);

OAI21x1_ASAP7_75t_L g344 ( 
.A1(n_332),
.A2(n_327),
.B(n_323),
.Y(n_344)
);

INVxp33_ASAP7_75t_L g347 ( 
.A(n_344),
.Y(n_347)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_331),
.A2(n_254),
.B(n_257),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_349),
.B(n_332),
.C(n_333),
.Y(n_352)
);

HB1xp67_ASAP7_75t_L g350 ( 
.A(n_341),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_350),
.A2(n_338),
.B(n_342),
.Y(n_351)
);

BUFx24_ASAP7_75t_SL g353 ( 
.A(n_351),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_SL g354 ( 
.A1(n_353),
.A2(n_352),
.B1(n_348),
.B2(n_347),
.Y(n_354)
);

XOR2xp5_ASAP7_75t_L g355 ( 
.A(n_354),
.B(n_8),
.Y(n_355)
);


endmodule