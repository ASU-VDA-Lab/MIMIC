module fake_netlist_5_1829_n_2311 (n_137, n_210, n_168, n_164, n_191, n_91, n_208, n_82, n_122, n_194, n_142, n_176, n_10, n_214, n_140, n_24, n_124, n_86, n_136, n_146, n_182, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_180, n_184, n_65, n_78, n_74, n_144, n_207, n_114, n_57, n_96, n_37, n_189, n_165, n_111, n_108, n_213, n_129, n_31, n_13, n_66, n_98, n_177, n_60, n_155, n_152, n_197, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_195, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_203, n_205, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_179, n_125, n_35, n_167, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_202, n_130, n_157, n_29, n_79, n_193, n_131, n_151, n_47, n_173, n_192, n_25, n_53, n_160, n_198, n_188, n_190, n_8, n_201, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_212, n_85, n_159, n_163, n_95, n_119, n_183, n_185, n_175, n_169, n_59, n_26, n_133, n_215, n_55, n_196, n_99, n_2, n_211, n_218, n_181, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_178, n_12, n_67, n_121, n_36, n_76, n_200, n_87, n_150, n_162, n_27, n_170, n_64, n_77, n_102, n_106, n_161, n_209, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_174, n_186, n_199, n_134, n_187, n_32, n_41, n_104, n_172, n_103, n_56, n_51, n_63, n_97, n_141, n_166, n_11, n_206, n_217, n_171, n_153, n_7, n_15, n_145, n_48, n_204, n_50, n_52, n_88, n_110, n_216, n_2311);

input n_137;
input n_210;
input n_168;
input n_164;
input n_191;
input n_91;
input n_208;
input n_82;
input n_122;
input n_194;
input n_142;
input n_176;
input n_10;
input n_214;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_182;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_180;
input n_184;
input n_65;
input n_78;
input n_74;
input n_144;
input n_207;
input n_114;
input n_57;
input n_96;
input n_37;
input n_189;
input n_165;
input n_111;
input n_108;
input n_213;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_177;
input n_60;
input n_155;
input n_152;
input n_197;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_195;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_203;
input n_205;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_179;
input n_125;
input n_35;
input n_167;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_202;
input n_130;
input n_157;
input n_29;
input n_79;
input n_193;
input n_131;
input n_151;
input n_47;
input n_173;
input n_192;
input n_25;
input n_53;
input n_160;
input n_198;
input n_188;
input n_190;
input n_8;
input n_201;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_212;
input n_85;
input n_159;
input n_163;
input n_95;
input n_119;
input n_183;
input n_185;
input n_175;
input n_169;
input n_59;
input n_26;
input n_133;
input n_215;
input n_55;
input n_196;
input n_99;
input n_2;
input n_211;
input n_218;
input n_181;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_178;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_200;
input n_87;
input n_150;
input n_162;
input n_27;
input n_170;
input n_64;
input n_77;
input n_102;
input n_106;
input n_161;
input n_209;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_174;
input n_186;
input n_199;
input n_134;
input n_187;
input n_32;
input n_41;
input n_104;
input n_172;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_166;
input n_11;
input n_206;
input n_217;
input n_171;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_204;
input n_50;
input n_52;
input n_88;
input n_110;
input n_216;

output n_2311;

wire n_924;
wire n_1263;
wire n_977;
wire n_1378;
wire n_2253;
wire n_611;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_1166;
wire n_1751;
wire n_469;
wire n_1508;
wire n_785;
wire n_549;
wire n_2200;
wire n_532;
wire n_1161;
wire n_1859;
wire n_1677;
wire n_1150;
wire n_226;
wire n_1780;
wire n_1488;
wire n_667;
wire n_790;
wire n_1055;
wire n_1501;
wire n_880;
wire n_544;
wire n_1007;
wire n_552;
wire n_1528;
wire n_1370;
wire n_1292;
wire n_1198;
wire n_1360;
wire n_1099;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_1021;
wire n_1960;
wire n_2185;
wire n_551;
wire n_2143;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_1353;
wire n_800;
wire n_1347;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_864;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_275;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2024;
wire n_1696;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_1359;
wire n_530;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_2031;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_1896;
wire n_2165;
wire n_2147;
wire n_929;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_1104;
wire n_1294;
wire n_659;
wire n_1705;
wire n_1257;
wire n_1182;
wire n_579;
wire n_1698;
wire n_1261;
wire n_938;
wire n_1098;
wire n_2142;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_1135;
wire n_519;
wire n_406;
wire n_2203;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2047;
wire n_1280;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2058;
wire n_291;
wire n_231;
wire n_257;
wire n_731;
wire n_371;
wire n_1483;
wire n_1314;
wire n_1512;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_569;
wire n_2144;
wire n_1778;
wire n_227;
wire n_2306;
wire n_920;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_335;
wire n_2085;
wire n_1669;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2149;
wire n_1078;
wire n_1670;
wire n_775;
wire n_219;
wire n_600;
wire n_1484;
wire n_2071;
wire n_1374;
wire n_1328;
wire n_223;
wire n_2141;
wire n_1948;
wire n_1984;
wire n_2099;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_1723;
wire n_955;
wire n_1850;
wire n_339;
wire n_1146;
wire n_882;
wire n_243;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_550;
wire n_696;
wire n_897;
wire n_350;
wire n_798;
wire n_646;
wire n_1428;
wire n_436;
wire n_1394;
wire n_1414;
wire n_1216;
wire n_580;
wire n_290;
wire n_1040;
wire n_2202;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_926;
wire n_2180;
wire n_2249;
wire n_344;
wire n_1218;
wire n_1931;
wire n_2276;
wire n_475;
wire n_422;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_1755;
wire n_415;
wire n_1071;
wire n_485;
wire n_1165;
wire n_1267;
wire n_1561;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_528;
wire n_2300;
wire n_1796;
wire n_680;
wire n_1473;
wire n_1587;
wire n_395;
wire n_553;
wire n_901;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_2174;
wire n_1748;
wire n_1672;
wire n_675;
wire n_888;
wire n_1880;
wire n_1167;
wire n_1626;
wire n_637;
wire n_1384;
wire n_1556;
wire n_446;
wire n_1863;
wire n_1064;
wire n_858;
wire n_2079;
wire n_2238;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_881;
wire n_1405;
wire n_1706;
wire n_468;
wire n_342;
wire n_464;
wire n_363;
wire n_1582;
wire n_1069;
wire n_1784;
wire n_1075;
wire n_1836;
wire n_1450;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2072;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_973;
wire n_1700;
wire n_477;
wire n_571;
wire n_1585;
wire n_461;
wire n_1971;
wire n_1599;
wire n_2275;
wire n_1211;
wire n_1197;
wire n_1523;
wire n_1950;
wire n_907;
wire n_1447;
wire n_2251;
wire n_1377;
wire n_989;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_1403;
wire n_2248;
wire n_488;
wire n_736;
wire n_892;
wire n_1000;
wire n_1202;
wire n_1278;
wire n_2062;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_332;
wire n_1053;
wire n_1224;
wire n_349;
wire n_1926;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_2150;
wire n_2241;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2140;
wire n_1819;
wire n_2139;
wire n_476;
wire n_1527;
wire n_2042;
wire n_534;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2175;
wire n_1854;
wire n_1565;
wire n_1809;
wire n_1856;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_561;
wire n_1319;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_1532;
wire n_2271;
wire n_1027;
wire n_971;
wire n_1156;
wire n_326;
wire n_794;
wire n_404;
wire n_2293;
wire n_686;
wire n_847;
wire n_1393;
wire n_596;
wire n_1775;
wire n_2028;
wire n_1368;
wire n_558;
wire n_702;
wire n_1276;
wire n_822;
wire n_1412;
wire n_1709;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_352;
wire n_1884;
wire n_1038;
wire n_520;
wire n_1369;
wire n_409;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2195;
wire n_300;
wire n_809;
wire n_931;
wire n_870;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_868;
wire n_639;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_1629;
wire n_1293;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_1175;
wire n_360;
wire n_1479;
wire n_1810;
wire n_1888;
wire n_2009;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_1997;
wire n_1766;
wire n_1477;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_1189;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_747;
wire n_2064;
wire n_784;
wire n_1733;
wire n_1244;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_697;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_1415;
wire n_367;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_1829;
wire n_1464;
wire n_649;
wire n_547;
wire n_1444;
wire n_1191;
wire n_1674;
wire n_1833;
wire n_1830;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_1734;
wire n_744;
wire n_629;
wire n_590;
wire n_1308;
wire n_2178;
wire n_1767;
wire n_254;
wire n_1680;
wire n_1233;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_293;
wire n_677;
wire n_372;
wire n_244;
wire n_1333;
wire n_1121;
wire n_314;
wire n_433;
wire n_604;
wire n_368;
wire n_2007;
wire n_949;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_738;
wire n_1624;
wire n_640;
wire n_1510;
wire n_624;
wire n_252;
wire n_1380;
wire n_1744;
wire n_1617;
wire n_295;
wire n_1010;
wire n_1994;
wire n_1231;
wire n_739;
wire n_1279;
wire n_1406;
wire n_1195;
wire n_1837;
wire n_1839;
wire n_610;
wire n_1760;
wire n_936;
wire n_568;
wire n_1500;
wire n_1090;
wire n_757;
wire n_633;
wire n_439;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_2046;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_1158;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_1987;
wire n_1145;
wire n_878;
wire n_524;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_1871;
wire n_1964;
wire n_331;
wire n_906;
wire n_1163;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2035;
wire n_658;
wire n_2061;
wire n_1740;
wire n_1362;
wire n_1586;
wire n_456;
wire n_959;
wire n_535;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_1923;
wire n_1773;
wire n_592;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_1017;
wire n_2171;
wire n_978;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2137;
wire n_603;
wire n_1431;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_1148;
wire n_2051;
wire n_750;
wire n_742;
wire n_2029;
wire n_995;
wire n_454;
wire n_2168;
wire n_1609;
wire n_374;
wire n_1989;
wire n_396;
wire n_1887;
wire n_1383;
wire n_1073;
wire n_255;
wire n_662;
wire n_459;
wire n_962;
wire n_1215;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_1336;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_1574;
wire n_473;
wire n_2048;
wire n_2133;
wire n_1921;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_355;
wire n_486;
wire n_1800;
wire n_1548;
wire n_614;
wire n_337;
wire n_1421;
wire n_1286;
wire n_1177;
wire n_1355;
wire n_974;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_2124;
wire n_743;
wire n_2081;
wire n_299;
wire n_303;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2261;
wire n_1820;
wire n_829;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_1724;
wire n_2111;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_1420;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_1127;
wire n_2277;
wire n_761;
wire n_1785;
wire n_1568;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2090;
wire n_1870;
wire n_309;
wire n_512;
wire n_1591;
wire n_2033;
wire n_322;
wire n_1682;
wire n_1980;
wire n_1249;
wire n_652;
wire n_1111;
wire n_1365;
wire n_1927;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_1909;
wire n_224;
wire n_1562;
wire n_383;
wire n_834;
wire n_765;
wire n_2255;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_1913;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_358;
wire n_1101;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_1324;
wire n_987;
wire n_1846;
wire n_261;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_1903;
wire n_1407;
wire n_1551;
wire n_545;
wire n_441;
wire n_860;
wire n_450;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_628;
wire n_365;
wire n_1849;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_1430;
wire n_513;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_1044;
wire n_1205;
wire n_346;
wire n_1209;
wire n_1552;
wire n_495;
wire n_602;
wire n_574;
wire n_1435;
wire n_879;
wire n_623;
wire n_2088;
wire n_405;
wire n_824;
wire n_359;
wire n_1645;
wire n_490;
wire n_1327;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_1717;
wire n_572;
wire n_366;
wire n_815;
wire n_1795;
wire n_2128;
wire n_1821;
wire n_327;
wire n_1381;
wire n_1611;
wire n_1037;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_1316;
wire n_1708;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2092;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2281;
wire n_2131;
wire n_2216;
wire n_531;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_960;
wire n_2308;
wire n_1893;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_1311;
wire n_2191;
wire n_1519;
wire n_256;
wire n_950;
wire n_1553;
wire n_1811;
wire n_380;
wire n_419;
wire n_1346;
wire n_444;
wire n_1299;
wire n_2158;
wire n_1808;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_418;
wire n_248;
wire n_912;
wire n_968;
wire n_315;
wire n_451;
wire n_619;
wire n_408;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_1139;
wire n_515;
wire n_351;
wire n_885;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_1157;
wire n_841;
wire n_1050;
wire n_802;
wire n_1954;
wire n_2265;
wire n_1608;
wire n_983;
wire n_1844;
wire n_280;
wire n_1305;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_2304;
wire n_762;
wire n_1283;
wire n_1644;
wire n_690;
wire n_1974;
wire n_583;
wire n_2086;
wire n_2289;
wire n_302;
wire n_1343;
wire n_2263;
wire n_1203;
wire n_1631;
wire n_821;
wire n_1763;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_753;
wire n_621;
wire n_455;
wire n_1048;
wire n_1719;
wire n_1288;
wire n_385;
wire n_507;
wire n_2269;
wire n_2309;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2123;
wire n_972;
wire n_692;
wire n_2037;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_1911;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_1688;
wire n_945;
wire n_492;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_1932;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_2082;
wire n_286;
wire n_1992;
wire n_1643;
wire n_883;
wire n_1983;
wire n_470;
wire n_449;
wire n_325;
wire n_1594;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_856;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_540;
wire n_618;
wire n_896;
wire n_2310;
wire n_323;
wire n_2287;
wire n_356;
wire n_2291;
wire n_894;
wire n_1636;
wire n_2056;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_234;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_833;
wire n_2020;
wire n_1646;
wire n_225;
wire n_1307;
wire n_1881;
wire n_988;
wire n_2043;
wire n_1940;
wire n_814;
wire n_1549;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_387;
wire n_1149;
wire n_398;
wire n_1671;
wire n_635;
wire n_763;
wire n_1020;
wire n_1062;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_1814;
wire n_1035;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_1188;
wire n_1722;
wire n_661;
wire n_1802;
wire n_849;
wire n_584;
wire n_681;
wire n_336;
wire n_1638;
wire n_1786;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_311;
wire n_830;
wire n_2098;
wire n_1296;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_749;
wire n_1895;
wire n_1134;
wire n_1358;
wire n_717;
wire n_939;
wire n_482;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_866;
wire n_969;
wire n_1401;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_338;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_836;
wire n_990;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_567;
wire n_1465;
wire n_778;
wire n_1122;
wire n_306;
wire n_458;
wire n_770;
wire n_1375;
wire n_1102;
wire n_1843;
wire n_711;
wire n_1499;
wire n_1187;
wire n_1441;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_489;
wire n_1174;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_1572;
wire n_1968;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_726;
wire n_982;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_1658;
wire n_899;
wire n_1253;
wire n_1737;
wire n_2201;
wire n_2117;
wire n_1904;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2205;
wire n_1335;
wire n_1514;
wire n_1777;
wire n_1957;
wire n_1059;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_2067;
wire n_527;
wire n_707;
wire n_1168;
wire n_2219;
wire n_2148;
wire n_937;
wire n_1427;
wire n_393;
wire n_487;
wire n_1584;
wire n_665;
wire n_1726;
wire n_1835;
wire n_1440;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_1787;
wire n_910;
wire n_2232;
wire n_2212;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_1496;
wire n_1125;
wire n_410;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_232;
wire n_1915;
wire n_1109;
wire n_895;
wire n_1310;
wire n_2121;
wire n_1803;
wire n_427;
wire n_1399;
wire n_1543;
wire n_1991;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_808;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_500;
wire n_1067;
wire n_1720;
wire n_435;
wire n_2003;
wire n_766;
wire n_1457;
wire n_541;
wire n_538;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_869;
wire n_810;
wire n_416;
wire n_827;
wire n_401;
wire n_1703;
wire n_1352;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_2211;
wire n_2095;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_1602;
wire n_855;
wire n_1178;
wire n_1461;
wire n_850;
wire n_684;
wire n_268;
wire n_2286;
wire n_664;
wire n_1999;
wire n_503;
wire n_2065;
wire n_2136;
wire n_235;
wire n_1372;
wire n_605;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_916;
wire n_1081;
wire n_493;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_998;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_725;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_672;
wire n_1985;
wire n_1898;
wire n_2107;
wire n_581;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_265;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_714;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_997;
wire n_932;
wire n_612;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_1268;
wire n_559;
wire n_825;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_509;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_1376;
wire n_941;
wire n_981;
wire n_1569;
wire n_2188;
wire n_867;
wire n_2239;
wire n_587;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_548;
wire n_812;
wire n_298;
wire n_2104;
wire n_518;
wire n_505;
wire n_2057;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_782;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_1900;
wire n_1620;
wire n_381;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_481;
wire n_1675;
wire n_1924;
wire n_1727;
wire n_1554;
wire n_1745;
wire n_769;
wire n_2006;
wire n_1995;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_1813;
wire n_886;
wire n_2014;
wire n_1221;
wire n_654;
wire n_1172;
wire n_379;
wire n_428;
wire n_1341;
wire n_570;
wire n_1641;
wire n_1361;
wire n_1707;
wire n_853;
wire n_377;
wire n_751;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_1129;
wire n_392;
wire n_704;
wire n_787;
wire n_1770;
wire n_961;
wire n_2250;
wire n_1756;
wire n_771;
wire n_276;
wire n_1716;
wire n_1225;
wire n_1520;
wire n_522;
wire n_1287;
wire n_1262;
wire n_400;
wire n_930;
wire n_1873;
wire n_1411;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_1087;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_1498;
wire n_2167;
wire n_1223;
wire n_1272;
wire n_682;
wire n_1567;
wire n_1247;
wire n_922;
wire n_816;
wire n_1648;
wire n_591;
wire n_1536;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_839;
wire n_1210;
wire n_1364;
wire n_2183;
wire n_328;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_1555;
wire n_499;
wire n_1589;
wire n_517;
wire n_413;
wire n_402;
wire n_1086;
wire n_796;
wire n_1858;
wire n_1619;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_1348;
wire n_2030;
wire n_903;
wire n_1525;
wire n_1752;
wire n_740;
wire n_384;
wire n_2208;
wire n_1404;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_1910;
wire n_333;
wire n_1298;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_1193;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2146;
wire n_844;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_1627;
wire n_1245;
wire n_846;
wire n_1673;
wire n_465;
wire n_362;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_1739;
wire n_270;
wire n_616;
wire n_2278;
wire n_1914;
wire n_2135;
wire n_745;
wire n_1654;
wire n_1103;
wire n_648;
wire n_1379;
wire n_312;
wire n_2196;
wire n_2170;
wire n_1076;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_730;
wire n_2036;
wire n_1325;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2083;
wire n_695;
wire n_656;
wire n_1606;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_229;
wire n_1936;
wire n_1956;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2027;
wire n_453;
wire n_403;
wire n_1130;
wire n_720;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_1604;
wire n_1275;
wire n_1764;
wire n_712;
wire n_246;
wire n_1583;
wire n_1042;
wire n_1402;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_1621;
wire n_2113;
wire n_251;
wire n_566;
wire n_565;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2274;
wire n_811;
wire n_334;
wire n_1558;
wire n_807;
wire n_2166;
wire n_835;
wire n_666;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_2044;
wire n_1990;
wire n_1004;
wire n_1186;
wire n_1032;
wire n_242;
wire n_1681;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_1693;
wire n_438;
wire n_713;
wire n_904;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_1180;
wire n_1827;
wire n_1271;
wire n_533;
wire n_1542;
wire n_1251;
wire n_278;
wire n_2268;

INVx1_ASAP7_75t_L g219 ( 
.A(n_55),
.Y(n_219)
);

INVx1_ASAP7_75t_SL g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_92),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_189),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_170),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_32),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_49),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_25),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_43),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_205),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_143),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_69),
.Y(n_230)
);

BUFx10_ASAP7_75t_L g231 ( 
.A(n_92),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_49),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_80),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_25),
.Y(n_234)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_11),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_171),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_105),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_145),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_115),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_16),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_195),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_198),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_83),
.Y(n_243)
);

BUFx10_ASAP7_75t_L g244 ( 
.A(n_165),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_67),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_93),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_14),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_113),
.Y(n_248)
);

BUFx10_ASAP7_75t_L g249 ( 
.A(n_72),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_75),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_38),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_35),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_156),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_65),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_73),
.Y(n_255)
);

INVx2_ASAP7_75t_L g256 ( 
.A(n_147),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_33),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_117),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_160),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_42),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_150),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_26),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_192),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_46),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_207),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_212),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_127),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_44),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_216),
.Y(n_269)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_123),
.Y(n_270)
);

BUFx6f_ASAP7_75t_L g271 ( 
.A(n_132),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_179),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_169),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_135),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_110),
.Y(n_275)
);

CKINVDCx5p33_ASAP7_75t_R g276 ( 
.A(n_125),
.Y(n_276)
);

CKINVDCx16_ASAP7_75t_R g277 ( 
.A(n_121),
.Y(n_277)
);

CKINVDCx5p33_ASAP7_75t_R g278 ( 
.A(n_78),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_193),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_122),
.Y(n_280)
);

BUFx6f_ASAP7_75t_L g281 ( 
.A(n_157),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g282 ( 
.A(n_111),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_17),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_130),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_118),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_5),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_186),
.Y(n_287)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_196),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_154),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_28),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_148),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_53),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_66),
.Y(n_293)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_11),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_14),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_213),
.Y(n_296)
);

BUFx2_ASAP7_75t_L g297 ( 
.A(n_43),
.Y(n_297)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_103),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_73),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_102),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_159),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_8),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_50),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_52),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_218),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_10),
.Y(n_306)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_60),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_138),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_129),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_194),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_191),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_178),
.Y(n_312)
);

BUFx3_ASAP7_75t_L g313 ( 
.A(n_183),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_141),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_163),
.Y(n_315)
);

INVx1_ASAP7_75t_SL g316 ( 
.A(n_1),
.Y(n_316)
);

BUFx5_ASAP7_75t_L g317 ( 
.A(n_162),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_153),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_48),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_124),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_204),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_13),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_199),
.Y(n_323)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_44),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_60),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_119),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_61),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_70),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_36),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_106),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_131),
.Y(n_331)
);

INVx2_ASAP7_75t_L g332 ( 
.A(n_36),
.Y(n_332)
);

CKINVDCx5p33_ASAP7_75t_R g333 ( 
.A(n_176),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_95),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_7),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_6),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_151),
.Y(n_337)
);

BUFx10_ASAP7_75t_L g338 ( 
.A(n_34),
.Y(n_338)
);

CKINVDCx14_ASAP7_75t_R g339 ( 
.A(n_149),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_99),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_167),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_70),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_74),
.Y(n_343)
);

INVx1_ASAP7_75t_SL g344 ( 
.A(n_72),
.Y(n_344)
);

CKINVDCx5p33_ASAP7_75t_R g345 ( 
.A(n_142),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_214),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_15),
.Y(n_347)
);

INVx2_ASAP7_75t_L g348 ( 
.A(n_175),
.Y(n_348)
);

INVx1_ASAP7_75t_SL g349 ( 
.A(n_56),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_59),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_76),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_109),
.Y(n_352)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_83),
.Y(n_353)
);

CKINVDCx5p33_ASAP7_75t_R g354 ( 
.A(n_37),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_208),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_203),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_97),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_66),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_8),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_177),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_23),
.Y(n_361)
);

CKINVDCx5p33_ASAP7_75t_R g362 ( 
.A(n_76),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_17),
.Y(n_363)
);

CKINVDCx5p33_ASAP7_75t_R g364 ( 
.A(n_40),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_168),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_20),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_108),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_98),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_23),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_137),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_126),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_100),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_12),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_200),
.Y(n_374)
);

CKINVDCx5p33_ASAP7_75t_R g375 ( 
.A(n_6),
.Y(n_375)
);

BUFx5_ASAP7_75t_L g376 ( 
.A(n_91),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_42),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_24),
.Y(n_378)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_197),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_27),
.Y(n_380)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_139),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_34),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_15),
.Y(n_383)
);

CKINVDCx20_ASAP7_75t_R g384 ( 
.A(n_10),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_55),
.Y(n_385)
);

CKINVDCx5p33_ASAP7_75t_R g386 ( 
.A(n_77),
.Y(n_386)
);

CKINVDCx16_ASAP7_75t_R g387 ( 
.A(n_93),
.Y(n_387)
);

CKINVDCx20_ASAP7_75t_R g388 ( 
.A(n_107),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_152),
.Y(n_389)
);

CKINVDCx5p33_ASAP7_75t_R g390 ( 
.A(n_77),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_53),
.Y(n_391)
);

INVx2_ASAP7_75t_SL g392 ( 
.A(n_22),
.Y(n_392)
);

CKINVDCx5p33_ASAP7_75t_R g393 ( 
.A(n_12),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g394 ( 
.A(n_65),
.Y(n_394)
);

INVx2_ASAP7_75t_L g395 ( 
.A(n_50),
.Y(n_395)
);

CKINVDCx5p33_ASAP7_75t_R g396 ( 
.A(n_114),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_21),
.Y(n_397)
);

CKINVDCx5p33_ASAP7_75t_R g398 ( 
.A(n_19),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_166),
.Y(n_399)
);

CKINVDCx5p33_ASAP7_75t_R g400 ( 
.A(n_38),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_202),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_2),
.Y(n_402)
);

CKINVDCx5p33_ASAP7_75t_R g403 ( 
.A(n_161),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g404 ( 
.A(n_210),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_64),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_5),
.Y(n_406)
);

CKINVDCx16_ASAP7_75t_R g407 ( 
.A(n_158),
.Y(n_407)
);

CKINVDCx5p33_ASAP7_75t_R g408 ( 
.A(n_81),
.Y(n_408)
);

CKINVDCx5p33_ASAP7_75t_R g409 ( 
.A(n_85),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_54),
.Y(n_410)
);

CKINVDCx16_ASAP7_75t_R g411 ( 
.A(n_209),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_89),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_30),
.Y(n_413)
);

CKINVDCx5p33_ASAP7_75t_R g414 ( 
.A(n_85),
.Y(n_414)
);

CKINVDCx5p33_ASAP7_75t_R g415 ( 
.A(n_155),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_24),
.Y(n_416)
);

CKINVDCx5p33_ASAP7_75t_R g417 ( 
.A(n_29),
.Y(n_417)
);

CKINVDCx5p33_ASAP7_75t_R g418 ( 
.A(n_81),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_79),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_78),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_30),
.Y(n_421)
);

CKINVDCx5p33_ASAP7_75t_R g422 ( 
.A(n_174),
.Y(n_422)
);

CKINVDCx5p33_ASAP7_75t_R g423 ( 
.A(n_215),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_9),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_211),
.Y(n_425)
);

CKINVDCx5p33_ASAP7_75t_R g426 ( 
.A(n_13),
.Y(n_426)
);

INVx2_ASAP7_75t_SL g427 ( 
.A(n_79),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_48),
.Y(n_428)
);

CKINVDCx5p33_ASAP7_75t_R g429 ( 
.A(n_69),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_67),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_128),
.Y(n_431)
);

CKINVDCx20_ASAP7_75t_R g432 ( 
.A(n_253),
.Y(n_432)
);

INVx2_ASAP7_75t_L g433 ( 
.A(n_376),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_376),
.Y(n_434)
);

CKINVDCx5p33_ASAP7_75t_R g435 ( 
.A(n_222),
.Y(n_435)
);

INVxp67_ASAP7_75t_SL g436 ( 
.A(n_282),
.Y(n_436)
);

CKINVDCx20_ASAP7_75t_R g437 ( 
.A(n_270),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_376),
.Y(n_438)
);

CKINVDCx5p33_ASAP7_75t_R g439 ( 
.A(n_228),
.Y(n_439)
);

HB1xp67_ASAP7_75t_L g440 ( 
.A(n_297),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_376),
.Y(n_441)
);

HB1xp67_ASAP7_75t_L g442 ( 
.A(n_297),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_229),
.Y(n_443)
);

CKINVDCx5p33_ASAP7_75t_R g444 ( 
.A(n_236),
.Y(n_444)
);

INVxp67_ASAP7_75t_SL g445 ( 
.A(n_282),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_309),
.B(n_0),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_376),
.Y(n_447)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_376),
.B(n_0),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_237),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_238),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_376),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_376),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_239),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_376),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_308),
.Y(n_455)
);

INVxp67_ASAP7_75t_L g456 ( 
.A(n_219),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_283),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_283),
.Y(n_458)
);

CKINVDCx16_ASAP7_75t_R g459 ( 
.A(n_268),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_332),
.Y(n_460)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_320),
.Y(n_461)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_332),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_241),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_395),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_395),
.Y(n_465)
);

BUFx3_ASAP7_75t_L g466 ( 
.A(n_313),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_416),
.Y(n_467)
);

CKINVDCx20_ASAP7_75t_R g468 ( 
.A(n_388),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_416),
.Y(n_469)
);

BUFx2_ASAP7_75t_L g470 ( 
.A(n_268),
.Y(n_470)
);

CKINVDCx5p33_ASAP7_75t_R g471 ( 
.A(n_242),
.Y(n_471)
);

CKINVDCx20_ASAP7_75t_R g472 ( 
.A(n_277),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_219),
.Y(n_473)
);

NOR2xp67_ASAP7_75t_L g474 ( 
.A(n_392),
.B(n_1),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_313),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_225),
.Y(n_476)
);

CKINVDCx5p33_ASAP7_75t_R g477 ( 
.A(n_248),
.Y(n_477)
);

CKINVDCx5p33_ASAP7_75t_R g478 ( 
.A(n_258),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_317),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_225),
.Y(n_480)
);

INVxp33_ASAP7_75t_SL g481 ( 
.A(n_221),
.Y(n_481)
);

INVxp67_ASAP7_75t_L g482 ( 
.A(n_227),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_227),
.Y(n_483)
);

CKINVDCx20_ASAP7_75t_R g484 ( 
.A(n_277),
.Y(n_484)
);

CKINVDCx5p33_ASAP7_75t_R g485 ( 
.A(n_259),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_240),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_240),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g488 ( 
.A(n_407),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_261),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_263),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_317),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_257),
.Y(n_492)
);

CKINVDCx5p33_ASAP7_75t_R g493 ( 
.A(n_266),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_257),
.Y(n_494)
);

CKINVDCx5p33_ASAP7_75t_R g495 ( 
.A(n_267),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g496 ( 
.A(n_407),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_269),
.Y(n_497)
);

NOR2xp67_ASAP7_75t_L g498 ( 
.A(n_392),
.B(n_2),
.Y(n_498)
);

CKINVDCx5p33_ASAP7_75t_R g499 ( 
.A(n_273),
.Y(n_499)
);

CKINVDCx5p33_ASAP7_75t_R g500 ( 
.A(n_274),
.Y(n_500)
);

CKINVDCx5p33_ASAP7_75t_R g501 ( 
.A(n_275),
.Y(n_501)
);

CKINVDCx20_ASAP7_75t_R g502 ( 
.A(n_411),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_276),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_307),
.Y(n_504)
);

CKINVDCx20_ASAP7_75t_R g505 ( 
.A(n_411),
.Y(n_505)
);

AND2x2_ASAP7_75t_L g506 ( 
.A(n_387),
.B(n_3),
.Y(n_506)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_307),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_279),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_309),
.B(n_3),
.Y(n_509)
);

CKINVDCx20_ASAP7_75t_R g510 ( 
.A(n_339),
.Y(n_510)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_319),
.Y(n_511)
);

CKINVDCx20_ASAP7_75t_R g512 ( 
.A(n_280),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_319),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_328),
.Y(n_514)
);

CKINVDCx5p33_ASAP7_75t_R g515 ( 
.A(n_284),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_289),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_223),
.B(n_4),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_328),
.Y(n_518)
);

INVxp67_ASAP7_75t_L g519 ( 
.A(n_350),
.Y(n_519)
);

CKINVDCx20_ASAP7_75t_R g520 ( 
.A(n_291),
.Y(n_520)
);

CKINVDCx20_ASAP7_75t_R g521 ( 
.A(n_305),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_350),
.Y(n_522)
);

CKINVDCx20_ASAP7_75t_R g523 ( 
.A(n_311),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_256),
.B(n_4),
.Y(n_524)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_314),
.Y(n_525)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_353),
.Y(n_526)
);

CKINVDCx16_ASAP7_75t_R g527 ( 
.A(n_387),
.Y(n_527)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_353),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_315),
.Y(n_529)
);

NOR2xp67_ASAP7_75t_L g530 ( 
.A(n_427),
.B(n_7),
.Y(n_530)
);

INVx2_ASAP7_75t_L g531 ( 
.A(n_317),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g532 ( 
.A(n_318),
.Y(n_532)
);

CKINVDCx20_ASAP7_75t_R g533 ( 
.A(n_321),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_358),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_323),
.Y(n_535)
);

CKINVDCx20_ASAP7_75t_R g536 ( 
.A(n_333),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_358),
.Y(n_537)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_337),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_359),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_340),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_345),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_359),
.Y(n_542)
);

CKINVDCx20_ASAP7_75t_R g543 ( 
.A(n_346),
.Y(n_543)
);

CKINVDCx5p33_ASAP7_75t_R g544 ( 
.A(n_352),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_377),
.Y(n_545)
);

BUFx6f_ASAP7_75t_L g546 ( 
.A(n_433),
.Y(n_546)
);

CKINVDCx5p33_ASAP7_75t_R g547 ( 
.A(n_435),
.Y(n_547)
);

NOR2xp67_ASAP7_75t_L g548 ( 
.A(n_434),
.B(n_256),
.Y(n_548)
);

CKINVDCx5p33_ASAP7_75t_R g549 ( 
.A(n_439),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g550 ( 
.A(n_470),
.Y(n_550)
);

HB1xp67_ASAP7_75t_L g551 ( 
.A(n_459),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_473),
.Y(n_552)
);

AND2x6_ASAP7_75t_L g553 ( 
.A(n_434),
.B(n_271),
.Y(n_553)
);

AND2x2_ASAP7_75t_SL g554 ( 
.A(n_506),
.B(n_265),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_475),
.B(n_427),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_L g556 ( 
.A(n_446),
.B(n_357),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_473),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_433),
.Y(n_558)
);

INVx3_ASAP7_75t_L g559 ( 
.A(n_438),
.Y(n_559)
);

CKINVDCx5p33_ASAP7_75t_R g560 ( 
.A(n_443),
.Y(n_560)
);

INVx3_ASAP7_75t_L g561 ( 
.A(n_438),
.Y(n_561)
);

HB1xp67_ASAP7_75t_L g562 ( 
.A(n_459),
.Y(n_562)
);

CKINVDCx5p33_ASAP7_75t_R g563 ( 
.A(n_444),
.Y(n_563)
);

BUFx2_ASAP7_75t_L g564 ( 
.A(n_472),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_L g565 ( 
.A(n_481),
.B(n_288),
.Y(n_565)
);

CKINVDCx5p33_ASAP7_75t_R g566 ( 
.A(n_449),
.Y(n_566)
);

NOR2xp33_ASAP7_75t_L g567 ( 
.A(n_436),
.B(n_301),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_441),
.Y(n_568)
);

BUFx2_ASAP7_75t_L g569 ( 
.A(n_484),
.Y(n_569)
);

INVx1_ASAP7_75t_L g570 ( 
.A(n_476),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_441),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_476),
.Y(n_572)
);

BUFx3_ASAP7_75t_L g573 ( 
.A(n_466),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_480),
.Y(n_574)
);

INVxp67_ASAP7_75t_L g575 ( 
.A(n_470),
.Y(n_575)
);

CKINVDCx20_ASAP7_75t_R g576 ( 
.A(n_432),
.Y(n_576)
);

INVx2_ASAP7_75t_L g577 ( 
.A(n_447),
.Y(n_577)
);

CKINVDCx20_ASAP7_75t_R g578 ( 
.A(n_437),
.Y(n_578)
);

CKINVDCx5p33_ASAP7_75t_R g579 ( 
.A(n_450),
.Y(n_579)
);

INVx1_ASAP7_75t_L g580 ( 
.A(n_480),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_483),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_447),
.Y(n_582)
);

CKINVDCx5p33_ASAP7_75t_R g583 ( 
.A(n_453),
.Y(n_583)
);

CKINVDCx5p33_ASAP7_75t_R g584 ( 
.A(n_463),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_483),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_486),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_486),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_487),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_487),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_492),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_451),
.B(n_404),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_492),
.Y(n_592)
);

INVx2_ASAP7_75t_L g593 ( 
.A(n_451),
.Y(n_593)
);

INVx1_ASAP7_75t_L g594 ( 
.A(n_494),
.Y(n_594)
);

BUFx6f_ASAP7_75t_L g595 ( 
.A(n_452),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_452),
.Y(n_596)
);

AND2x2_ASAP7_75t_L g597 ( 
.A(n_466),
.B(n_404),
.Y(n_597)
);

HB1xp67_ASAP7_75t_L g598 ( 
.A(n_527),
.Y(n_598)
);

INVx5_ASAP7_75t_L g599 ( 
.A(n_479),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_471),
.B(n_477),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_478),
.B(n_265),
.Y(n_601)
);

INVx1_ASAP7_75t_L g602 ( 
.A(n_494),
.Y(n_602)
);

INVx3_ASAP7_75t_L g603 ( 
.A(n_454),
.Y(n_603)
);

BUFx2_ASAP7_75t_L g604 ( 
.A(n_488),
.Y(n_604)
);

INVx1_ASAP7_75t_L g605 ( 
.A(n_504),
.Y(n_605)
);

INVx1_ASAP7_75t_L g606 ( 
.A(n_504),
.Y(n_606)
);

BUFx2_ASAP7_75t_L g607 ( 
.A(n_496),
.Y(n_607)
);

AND2x6_ASAP7_75t_L g608 ( 
.A(n_454),
.B(n_271),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_507),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_507),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_448),
.Y(n_611)
);

CKINVDCx5p33_ASAP7_75t_R g612 ( 
.A(n_485),
.Y(n_612)
);

CKINVDCx5p33_ASAP7_75t_R g613 ( 
.A(n_489),
.Y(n_613)
);

INVx3_ASAP7_75t_L g614 ( 
.A(n_479),
.Y(n_614)
);

CKINVDCx20_ASAP7_75t_R g615 ( 
.A(n_455),
.Y(n_615)
);

AND2x4_ASAP7_75t_L g616 ( 
.A(n_524),
.B(n_348),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_511),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_511),
.Y(n_618)
);

CKINVDCx5p33_ASAP7_75t_R g619 ( 
.A(n_490),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_SL g620 ( 
.A(n_527),
.B(n_244),
.Y(n_620)
);

INVx1_ASAP7_75t_L g621 ( 
.A(n_513),
.Y(n_621)
);

INVx5_ASAP7_75t_L g622 ( 
.A(n_491),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_513),
.Y(n_623)
);

CKINVDCx16_ASAP7_75t_R g624 ( 
.A(n_502),
.Y(n_624)
);

AOI22xp5_ASAP7_75t_L g625 ( 
.A1(n_506),
.A2(n_293),
.B1(n_369),
.B2(n_299),
.Y(n_625)
);

HB1xp67_ASAP7_75t_L g626 ( 
.A(n_493),
.Y(n_626)
);

AND2x4_ASAP7_75t_L g627 ( 
.A(n_491),
.B(n_348),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_514),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_531),
.Y(n_629)
);

INVx1_ASAP7_75t_L g630 ( 
.A(n_514),
.Y(n_630)
);

INVx1_ASAP7_75t_L g631 ( 
.A(n_518),
.Y(n_631)
);

CKINVDCx20_ASAP7_75t_R g632 ( 
.A(n_461),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_518),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_522),
.Y(n_634)
);

CKINVDCx20_ASAP7_75t_R g635 ( 
.A(n_468),
.Y(n_635)
);

NAND2xp5_ASAP7_75t_SL g636 ( 
.A(n_565),
.B(n_495),
.Y(n_636)
);

AND2x6_ASAP7_75t_L g637 ( 
.A(n_611),
.B(n_223),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_L g638 ( 
.A(n_554),
.B(n_497),
.Y(n_638)
);

INVx2_ASAP7_75t_L g639 ( 
.A(n_558),
.Y(n_639)
);

INVx4_ASAP7_75t_L g640 ( 
.A(n_571),
.Y(n_640)
);

NAND2x1p5_ASAP7_75t_L g641 ( 
.A(n_554),
.B(n_272),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_559),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_550),
.B(n_445),
.Y(n_643)
);

INVx4_ASAP7_75t_SL g644 ( 
.A(n_553),
.Y(n_644)
);

INVx1_ASAP7_75t_L g645 ( 
.A(n_559),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_554),
.B(n_499),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_568),
.Y(n_647)
);

INVx5_ASAP7_75t_L g648 ( 
.A(n_553),
.Y(n_648)
);

AND2x2_ASAP7_75t_L g649 ( 
.A(n_555),
.B(n_457),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_568),
.Y(n_650)
);

BUFx3_ASAP7_75t_L g651 ( 
.A(n_573),
.Y(n_651)
);

INVx3_ASAP7_75t_L g652 ( 
.A(n_546),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_555),
.B(n_457),
.Y(n_653)
);

OAI22xp33_ASAP7_75t_L g654 ( 
.A1(n_625),
.A2(n_509),
.B1(n_304),
.B2(n_316),
.Y(n_654)
);

AND2x2_ASAP7_75t_L g655 ( 
.A(n_597),
.B(n_458),
.Y(n_655)
);

INVx1_ASAP7_75t_L g656 ( 
.A(n_559),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_558),
.Y(n_657)
);

INVx5_ASAP7_75t_L g658 ( 
.A(n_553),
.Y(n_658)
);

AND2x6_ASAP7_75t_L g659 ( 
.A(n_611),
.B(n_272),
.Y(n_659)
);

INVx2_ASAP7_75t_L g660 ( 
.A(n_558),
.Y(n_660)
);

INVx4_ASAP7_75t_L g661 ( 
.A(n_571),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_611),
.B(n_500),
.Y(n_662)
);

AOI22xp33_ASAP7_75t_L g663 ( 
.A1(n_616),
.A2(n_517),
.B1(n_442),
.B2(n_440),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_611),
.B(n_501),
.Y(n_664)
);

NAND2xp33_ASAP7_75t_L g665 ( 
.A(n_611),
.B(n_317),
.Y(n_665)
);

BUFx6f_ASAP7_75t_L g666 ( 
.A(n_546),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_611),
.B(n_503),
.Y(n_667)
);

INVx1_ASAP7_75t_SL g668 ( 
.A(n_576),
.Y(n_668)
);

CKINVDCx20_ASAP7_75t_R g669 ( 
.A(n_578),
.Y(n_669)
);

INVx2_ASAP7_75t_L g670 ( 
.A(n_629),
.Y(n_670)
);

INVx4_ASAP7_75t_L g671 ( 
.A(n_571),
.Y(n_671)
);

BUFx3_ASAP7_75t_L g672 ( 
.A(n_573),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_556),
.B(n_601),
.Y(n_673)
);

INVx1_ASAP7_75t_L g674 ( 
.A(n_568),
.Y(n_674)
);

OR2x2_ASAP7_75t_L g675 ( 
.A(n_575),
.B(n_508),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_559),
.Y(n_676)
);

NAND2xp33_ASAP7_75t_L g677 ( 
.A(n_556),
.B(n_317),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_591),
.B(n_515),
.Y(n_678)
);

INVx1_ASAP7_75t_L g679 ( 
.A(n_577),
.Y(n_679)
);

INVx1_ASAP7_75t_L g680 ( 
.A(n_577),
.Y(n_680)
);

INVx3_ASAP7_75t_L g681 ( 
.A(n_546),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_SL g682 ( 
.A(n_567),
.B(n_516),
.Y(n_682)
);

BUFx6f_ASAP7_75t_L g683 ( 
.A(n_546),
.Y(n_683)
);

NOR2xp33_ASAP7_75t_L g684 ( 
.A(n_600),
.B(n_529),
.Y(n_684)
);

CKINVDCx16_ASAP7_75t_R g685 ( 
.A(n_624),
.Y(n_685)
);

INVx2_ASAP7_75t_L g686 ( 
.A(n_629),
.Y(n_686)
);

INVx4_ASAP7_75t_L g687 ( 
.A(n_571),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_577),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_629),
.Y(n_689)
);

OR2x2_ASAP7_75t_L g690 ( 
.A(n_597),
.B(n_540),
.Y(n_690)
);

OR2x2_ASAP7_75t_L g691 ( 
.A(n_551),
.B(n_544),
.Y(n_691)
);

AND2x6_ASAP7_75t_L g692 ( 
.A(n_616),
.B(n_285),
.Y(n_692)
);

INVx2_ASAP7_75t_L g693 ( 
.A(n_593),
.Y(n_693)
);

INVx2_ASAP7_75t_SL g694 ( 
.A(n_573),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_593),
.Y(n_695)
);

INVx2_ASAP7_75t_SL g696 ( 
.A(n_591),
.Y(n_696)
);

INVx1_ASAP7_75t_SL g697 ( 
.A(n_615),
.Y(n_697)
);

BUFx10_ASAP7_75t_L g698 ( 
.A(n_547),
.Y(n_698)
);

NAND2xp5_ASAP7_75t_SL g699 ( 
.A(n_549),
.B(n_510),
.Y(n_699)
);

BUFx6f_ASAP7_75t_L g700 ( 
.A(n_546),
.Y(n_700)
);

INVx4_ASAP7_75t_L g701 ( 
.A(n_571),
.Y(n_701)
);

CKINVDCx5p33_ASAP7_75t_R g702 ( 
.A(n_632),
.Y(n_702)
);

AND2x4_ASAP7_75t_L g703 ( 
.A(n_591),
.B(n_285),
.Y(n_703)
);

BUFx3_ASAP7_75t_L g704 ( 
.A(n_591),
.Y(n_704)
);

INVx1_ASAP7_75t_SL g705 ( 
.A(n_635),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_560),
.B(n_512),
.Y(n_706)
);

BUFx6f_ASAP7_75t_L g707 ( 
.A(n_546),
.Y(n_707)
);

INVx2_ASAP7_75t_SL g708 ( 
.A(n_616),
.Y(n_708)
);

AND2x4_ASAP7_75t_L g709 ( 
.A(n_616),
.B(n_287),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_563),
.B(n_520),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_L g711 ( 
.A(n_566),
.B(n_521),
.Y(n_711)
);

INVx2_ASAP7_75t_SL g712 ( 
.A(n_562),
.Y(n_712)
);

AOI22xp33_ASAP7_75t_L g713 ( 
.A1(n_627),
.A2(n_498),
.B1(n_530),
.B2(n_474),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_579),
.B(n_523),
.Y(n_714)
);

INVxp67_ASAP7_75t_L g715 ( 
.A(n_598),
.Y(n_715)
);

BUFx6f_ASAP7_75t_L g716 ( 
.A(n_571),
.Y(n_716)
);

OAI22xp5_ASAP7_75t_L g717 ( 
.A1(n_620),
.A2(n_532),
.B1(n_533),
.B2(n_525),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_561),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_583),
.Y(n_719)
);

AND2x4_ASAP7_75t_L g720 ( 
.A(n_552),
.B(n_287),
.Y(n_720)
);

INVx1_ASAP7_75t_L g721 ( 
.A(n_561),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_SL g722 ( 
.A(n_584),
.B(n_535),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_561),
.B(n_365),
.Y(n_723)
);

AND2x4_ASAP7_75t_L g724 ( 
.A(n_552),
.B(n_296),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_561),
.Y(n_725)
);

INVx4_ASAP7_75t_L g726 ( 
.A(n_582),
.Y(n_726)
);

INVx2_ASAP7_75t_SL g727 ( 
.A(n_627),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_593),
.Y(n_728)
);

NAND2xp5_ASAP7_75t_L g729 ( 
.A(n_603),
.B(n_381),
.Y(n_729)
);

INVx3_ASAP7_75t_L g730 ( 
.A(n_614),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_582),
.Y(n_731)
);

INVx1_ASAP7_75t_SL g732 ( 
.A(n_564),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_L g733 ( 
.A(n_603),
.B(n_396),
.Y(n_733)
);

BUFx10_ASAP7_75t_L g734 ( 
.A(n_612),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_596),
.Y(n_735)
);

AOI22xp33_ASAP7_75t_L g736 ( 
.A1(n_627),
.A2(n_498),
.B1(n_530),
.B2(n_474),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_596),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_596),
.Y(n_738)
);

AOI22xp5_ASAP7_75t_L g739 ( 
.A1(n_613),
.A2(n_536),
.B1(n_541),
.B2(n_538),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_603),
.Y(n_740)
);

NAND2xp33_ASAP7_75t_L g741 ( 
.A(n_553),
.B(n_317),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_SL g742 ( 
.A(n_619),
.B(n_543),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_557),
.B(n_570),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_626),
.B(n_505),
.Y(n_744)
);

NOR2xp33_ASAP7_75t_L g745 ( 
.A(n_557),
.B(n_456),
.Y(n_745)
);

INVx6_ASAP7_75t_L g746 ( 
.A(n_582),
.Y(n_746)
);

BUFx6f_ASAP7_75t_L g747 ( 
.A(n_582),
.Y(n_747)
);

AND2x4_ASAP7_75t_L g748 ( 
.A(n_570),
.B(n_296),
.Y(n_748)
);

AND2x4_ASAP7_75t_L g749 ( 
.A(n_572),
.B(n_300),
.Y(n_749)
);

INVx3_ASAP7_75t_L g750 ( 
.A(n_614),
.Y(n_750)
);

INVx2_ASAP7_75t_L g751 ( 
.A(n_614),
.Y(n_751)
);

BUFx6f_ASAP7_75t_L g752 ( 
.A(n_582),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_603),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_582),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_614),
.Y(n_755)
);

AND2x2_ASAP7_75t_SL g756 ( 
.A(n_625),
.B(n_300),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_595),
.B(n_403),
.Y(n_757)
);

INVx1_ASAP7_75t_L g758 ( 
.A(n_627),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_572),
.B(n_458),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_595),
.Y(n_760)
);

INVx3_ASAP7_75t_L g761 ( 
.A(n_595),
.Y(n_761)
);

CKINVDCx5p33_ASAP7_75t_R g762 ( 
.A(n_624),
.Y(n_762)
);

INVx1_ASAP7_75t_L g763 ( 
.A(n_595),
.Y(n_763)
);

INVx2_ASAP7_75t_SL g764 ( 
.A(n_574),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_574),
.B(n_460),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_595),
.B(n_415),
.Y(n_766)
);

AND2x6_ASAP7_75t_L g767 ( 
.A(n_595),
.B(n_310),
.Y(n_767)
);

INVx1_ASAP7_75t_L g768 ( 
.A(n_580),
.Y(n_768)
);

AND2x2_ASAP7_75t_L g769 ( 
.A(n_580),
.B(n_460),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_581),
.B(n_244),
.Y(n_770)
);

INVx2_ASAP7_75t_L g771 ( 
.A(n_581),
.Y(n_771)
);

INVx1_ASAP7_75t_L g772 ( 
.A(n_585),
.Y(n_772)
);

BUFx6f_ASAP7_75t_L g773 ( 
.A(n_599),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_548),
.B(n_422),
.Y(n_774)
);

CKINVDCx5p33_ASAP7_75t_R g775 ( 
.A(n_564),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_585),
.B(n_462),
.Y(n_776)
);

AND2x2_ASAP7_75t_L g777 ( 
.A(n_586),
.B(n_587),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_586),
.Y(n_778)
);

HB1xp67_ASAP7_75t_L g779 ( 
.A(n_569),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_587),
.B(n_462),
.Y(n_780)
);

NOR2xp33_ASAP7_75t_L g781 ( 
.A(n_588),
.B(n_482),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_588),
.B(n_464),
.Y(n_782)
);

INVx3_ASAP7_75t_L g783 ( 
.A(n_599),
.Y(n_783)
);

INVx1_ASAP7_75t_L g784 ( 
.A(n_589),
.Y(n_784)
);

CKINVDCx5p33_ASAP7_75t_R g785 ( 
.A(n_569),
.Y(n_785)
);

INVx1_ASAP7_75t_L g786 ( 
.A(n_589),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_590),
.B(n_464),
.Y(n_787)
);

BUFx6f_ASAP7_75t_L g788 ( 
.A(n_599),
.Y(n_788)
);

AND2x4_ASAP7_75t_L g789 ( 
.A(n_590),
.B(n_310),
.Y(n_789)
);

AND2x4_ASAP7_75t_L g790 ( 
.A(n_592),
.B(n_312),
.Y(n_790)
);

AOI22xp33_ASAP7_75t_L g791 ( 
.A1(n_708),
.A2(n_548),
.B1(n_312),
.B2(n_330),
.Y(n_791)
);

AOI22xp33_ASAP7_75t_L g792 ( 
.A1(n_708),
.A2(n_326),
.B1(n_331),
.B2(n_330),
.Y(n_792)
);

NOR2xp33_ASAP7_75t_L g793 ( 
.A(n_673),
.B(n_604),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_704),
.Y(n_794)
);

HB1xp67_ASAP7_75t_L g795 ( 
.A(n_779),
.Y(n_795)
);

AOI22xp33_ASAP7_75t_L g796 ( 
.A1(n_709),
.A2(n_326),
.B1(n_341),
.B2(n_331),
.Y(n_796)
);

AND2x6_ASAP7_75t_SL g797 ( 
.A(n_744),
.B(n_377),
.Y(n_797)
);

INVx8_ASAP7_75t_L g798 ( 
.A(n_692),
.Y(n_798)
);

NOR2xp33_ASAP7_75t_L g799 ( 
.A(n_684),
.B(n_604),
.Y(n_799)
);

CKINVDCx16_ASAP7_75t_R g800 ( 
.A(n_685),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_727),
.B(n_553),
.Y(n_801)
);

AOI22xp33_ASAP7_75t_L g802 ( 
.A1(n_709),
.A2(n_341),
.B1(n_356),
.B2(n_355),
.Y(n_802)
);

NOR2xp33_ASAP7_75t_L g803 ( 
.A(n_636),
.B(n_607),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_758),
.Y(n_804)
);

AND2x4_ASAP7_75t_L g805 ( 
.A(n_694),
.B(n_592),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_727),
.B(n_553),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_758),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_709),
.A2(n_355),
.B1(n_360),
.B2(n_356),
.Y(n_808)
);

AND2x6_ASAP7_75t_SL g809 ( 
.A(n_706),
.B(n_710),
.Y(n_809)
);

INVx2_ASAP7_75t_L g810 ( 
.A(n_771),
.Y(n_810)
);

INVx2_ASAP7_75t_L g811 ( 
.A(n_771),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_704),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_639),
.Y(n_813)
);

INVx1_ASAP7_75t_L g814 ( 
.A(n_743),
.Y(n_814)
);

INVx1_ASAP7_75t_L g815 ( 
.A(n_743),
.Y(n_815)
);

NOR2xp33_ASAP7_75t_L g816 ( 
.A(n_638),
.B(n_607),
.Y(n_816)
);

INVx1_ASAP7_75t_L g817 ( 
.A(n_777),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_777),
.Y(n_818)
);

INVx2_ASAP7_75t_L g819 ( 
.A(n_639),
.Y(n_819)
);

OR2x2_ASAP7_75t_L g820 ( 
.A(n_643),
.B(n_220),
.Y(n_820)
);

INVx2_ASAP7_75t_L g821 ( 
.A(n_657),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_SL g822 ( 
.A(n_696),
.B(n_271),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_SL g823 ( 
.A(n_696),
.B(n_271),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_662),
.B(n_553),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_768),
.Y(n_825)
);

AND2x2_ASAP7_75t_L g826 ( 
.A(n_649),
.B(n_594),
.Y(n_826)
);

INVx1_ASAP7_75t_L g827 ( 
.A(n_768),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_L g828 ( 
.A(n_646),
.B(n_344),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_664),
.B(n_553),
.Y(n_829)
);

AOI22xp33_ASAP7_75t_L g830 ( 
.A1(n_641),
.A2(n_360),
.B1(n_368),
.B2(n_367),
.Y(n_830)
);

INVx3_ASAP7_75t_L g831 ( 
.A(n_730),
.Y(n_831)
);

AOI22xp5_ASAP7_75t_L g832 ( 
.A1(n_667),
.A2(n_425),
.B1(n_423),
.B2(n_368),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_SL g833 ( 
.A(n_641),
.B(n_271),
.Y(n_833)
);

INVx4_ASAP7_75t_L g834 ( 
.A(n_716),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_764),
.B(n_608),
.Y(n_835)
);

NOR2xp33_ASAP7_75t_L g836 ( 
.A(n_682),
.B(n_349),
.Y(n_836)
);

INVx2_ASAP7_75t_L g837 ( 
.A(n_657),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_L g838 ( 
.A(n_764),
.B(n_608),
.Y(n_838)
);

A2O1A1Ixp33_ASAP7_75t_SL g839 ( 
.A1(n_677),
.A2(n_370),
.B(n_371),
.C(n_367),
.Y(n_839)
);

OAI22xp5_ASAP7_75t_L g840 ( 
.A1(n_641),
.A2(n_371),
.B1(n_372),
.B2(n_370),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_713),
.B(n_608),
.Y(n_841)
);

OAI21xp5_ASAP7_75t_L g842 ( 
.A1(n_642),
.A2(n_608),
.B(n_374),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_655),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_675),
.B(n_224),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_772),
.Y(n_845)
);

AND2x2_ASAP7_75t_L g846 ( 
.A(n_649),
.B(n_594),
.Y(n_846)
);

NOR2xp33_ASAP7_75t_L g847 ( 
.A(n_675),
.B(n_226),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_736),
.B(n_608),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_772),
.B(n_778),
.Y(n_849)
);

OAI22xp5_ASAP7_75t_L g850 ( 
.A1(n_678),
.A2(n_374),
.B1(n_379),
.B2(n_372),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_778),
.Y(n_851)
);

INVx3_ASAP7_75t_L g852 ( 
.A(n_730),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_660),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_SL g854 ( 
.A(n_703),
.B(n_281),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_692),
.A2(n_756),
.B1(n_703),
.B2(n_677),
.Y(n_855)
);

AOI22xp5_ASAP7_75t_L g856 ( 
.A1(n_692),
.A2(n_389),
.B1(n_399),
.B2(n_379),
.Y(n_856)
);

AND2x4_ASAP7_75t_L g857 ( 
.A(n_694),
.B(n_602),
.Y(n_857)
);

NOR2xp33_ASAP7_75t_L g858 ( 
.A(n_690),
.B(n_230),
.Y(n_858)
);

AOI22xp5_ASAP7_75t_L g859 ( 
.A1(n_692),
.A2(n_399),
.B1(n_401),
.B2(n_389),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_651),
.B(n_602),
.Y(n_860)
);

NAND2xp5_ASAP7_75t_L g861 ( 
.A(n_784),
.B(n_608),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_653),
.B(n_519),
.Y(n_862)
);

AOI22xp33_ASAP7_75t_L g863 ( 
.A1(n_692),
.A2(n_756),
.B1(n_703),
.B2(n_659),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_786),
.B(n_608),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_660),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_L g866 ( 
.A(n_653),
.B(n_608),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_SL g867 ( 
.A(n_648),
.B(n_281),
.Y(n_867)
);

AOI22xp33_ASAP7_75t_L g868 ( 
.A1(n_692),
.A2(n_431),
.B1(n_401),
.B2(n_294),
.Y(n_868)
);

BUFx6f_ASAP7_75t_L g869 ( 
.A(n_651),
.Y(n_869)
);

BUFx6f_ASAP7_75t_L g870 ( 
.A(n_672),
.Y(n_870)
);

BUFx6f_ASAP7_75t_SL g871 ( 
.A(n_698),
.Y(n_871)
);

AND2x6_ASAP7_75t_SL g872 ( 
.A(n_711),
.B(n_382),
.Y(n_872)
);

AOI22xp5_ASAP7_75t_L g873 ( 
.A1(n_654),
.A2(n_655),
.B1(n_729),
.B2(n_723),
.Y(n_873)
);

INVx2_ASAP7_75t_SL g874 ( 
.A(n_690),
.Y(n_874)
);

NAND2xp33_ASAP7_75t_L g875 ( 
.A(n_637),
.B(n_317),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_645),
.B(n_431),
.Y(n_876)
);

INVx5_ASAP7_75t_L g877 ( 
.A(n_773),
.Y(n_877)
);

NAND2xp5_ASAP7_75t_L g878 ( 
.A(n_656),
.B(n_605),
.Y(n_878)
);

AOI22xp33_ASAP7_75t_L g879 ( 
.A1(n_637),
.A2(n_298),
.B1(n_281),
.B2(n_317),
.Y(n_879)
);

NAND2xp5_ASAP7_75t_L g880 ( 
.A(n_676),
.B(n_605),
.Y(n_880)
);

NOR2xp33_ASAP7_75t_L g881 ( 
.A(n_643),
.B(n_232),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_670),
.Y(n_882)
);

NOR2xp33_ASAP7_75t_L g883 ( 
.A(n_715),
.B(n_691),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_L g884 ( 
.A(n_718),
.B(n_721),
.Y(n_884)
);

INVx2_ASAP7_75t_L g885 ( 
.A(n_670),
.Y(n_885)
);

BUFx3_ASAP7_75t_L g886 ( 
.A(n_672),
.Y(n_886)
);

INVx2_ASAP7_75t_SL g887 ( 
.A(n_720),
.Y(n_887)
);

BUFx6f_ASAP7_75t_L g888 ( 
.A(n_716),
.Y(n_888)
);

NAND2xp5_ASAP7_75t_L g889 ( 
.A(n_725),
.B(n_606),
.Y(n_889)
);

INVx8_ASAP7_75t_L g890 ( 
.A(n_637),
.Y(n_890)
);

OAI22xp5_ASAP7_75t_L g891 ( 
.A1(n_663),
.A2(n_324),
.B1(n_281),
.B2(n_298),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_759),
.Y(n_892)
);

AOI22xp5_ASAP7_75t_L g893 ( 
.A1(n_733),
.A2(n_634),
.B1(n_633),
.B2(n_631),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_L g894 ( 
.A(n_740),
.B(n_606),
.Y(n_894)
);

NOR2xp33_ASAP7_75t_L g895 ( 
.A(n_691),
.B(n_233),
.Y(n_895)
);

INVx4_ASAP7_75t_L g896 ( 
.A(n_716),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_SL g897 ( 
.A(n_648),
.B(n_281),
.Y(n_897)
);

AOI21xp5_ASAP7_75t_L g898 ( 
.A1(n_757),
.A2(n_766),
.B(n_665),
.Y(n_898)
);

OAI22xp5_ASAP7_75t_SL g899 ( 
.A1(n_669),
.A2(n_384),
.B1(n_380),
.B2(n_378),
.Y(n_899)
);

HB1xp67_ASAP7_75t_L g900 ( 
.A(n_712),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_753),
.B(n_609),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_730),
.B(n_609),
.Y(n_902)
);

OAI22xp33_ASAP7_75t_L g903 ( 
.A1(n_712),
.A2(n_382),
.B1(n_430),
.B2(n_383),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_750),
.B(n_610),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_665),
.A2(n_634),
.B(n_633),
.C(n_631),
.Y(n_905)
);

AOI22xp33_ASAP7_75t_L g906 ( 
.A1(n_637),
.A2(n_298),
.B1(n_317),
.B2(n_412),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_750),
.B(n_610),
.Y(n_907)
);

AOI22xp33_ASAP7_75t_L g908 ( 
.A1(n_637),
.A2(n_298),
.B1(n_430),
.B2(n_413),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_750),
.B(n_617),
.Y(n_909)
);

A2O1A1Ixp33_ASAP7_75t_L g910 ( 
.A1(n_745),
.A2(n_383),
.B(n_385),
.C(n_391),
.Y(n_910)
);

CKINVDCx5p33_ASAP7_75t_R g911 ( 
.A(n_719),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_763),
.B(n_617),
.Y(n_912)
);

INVx1_ASAP7_75t_L g913 ( 
.A(n_759),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_763),
.B(n_618),
.Y(n_914)
);

OR2x2_ASAP7_75t_L g915 ( 
.A(n_732),
.B(n_618),
.Y(n_915)
);

O2A1O1Ixp33_ASAP7_75t_L g916 ( 
.A1(n_741),
.A2(n_630),
.B(n_628),
.C(n_623),
.Y(n_916)
);

AOI22xp33_ASAP7_75t_L g917 ( 
.A1(n_637),
.A2(n_298),
.B1(n_421),
.B2(n_412),
.Y(n_917)
);

INVx2_ASAP7_75t_SL g918 ( 
.A(n_790),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_719),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_SL g920 ( 
.A(n_648),
.B(n_531),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_760),
.B(n_761),
.Y(n_921)
);

INVx2_ASAP7_75t_L g922 ( 
.A(n_686),
.Y(n_922)
);

INVx2_ASAP7_75t_L g923 ( 
.A(n_686),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_SL g924 ( 
.A(n_648),
.B(n_599),
.Y(n_924)
);

BUFx6f_ASAP7_75t_L g925 ( 
.A(n_716),
.Y(n_925)
);

BUFx3_ASAP7_75t_L g926 ( 
.A(n_698),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_659),
.A2(n_630),
.B1(n_628),
.B2(n_623),
.Y(n_927)
);

BUFx5_ASAP7_75t_L g928 ( 
.A(n_659),
.Y(n_928)
);

NAND2xp5_ASAP7_75t_L g929 ( 
.A(n_760),
.B(n_621),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_L g930 ( 
.A(n_781),
.B(n_243),
.C(n_234),
.Y(n_930)
);

NAND2xp5_ASAP7_75t_L g931 ( 
.A(n_761),
.B(n_621),
.Y(n_931)
);

AOI22xp33_ASAP7_75t_L g932 ( 
.A1(n_659),
.A2(n_391),
.B1(n_421),
.B2(n_420),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_761),
.B(n_622),
.Y(n_933)
);

AND2x2_ASAP7_75t_L g934 ( 
.A(n_720),
.B(n_724),
.Y(n_934)
);

NOR2xp67_ASAP7_75t_L g935 ( 
.A(n_739),
.B(n_96),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_652),
.B(n_599),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_652),
.B(n_599),
.Y(n_937)
);

INVx2_ASAP7_75t_L g938 ( 
.A(n_689),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_652),
.B(n_599),
.Y(n_939)
);

OAI22xp5_ASAP7_75t_L g940 ( 
.A1(n_720),
.A2(n_245),
.B1(n_246),
.B2(n_247),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_681),
.B(n_622),
.Y(n_941)
);

AOI22xp5_ASAP7_75t_L g942 ( 
.A1(n_659),
.A2(n_244),
.B1(n_373),
.B2(n_366),
.Y(n_942)
);

AOI22xp33_ASAP7_75t_L g943 ( 
.A1(n_659),
.A2(n_385),
.B1(n_410),
.B2(n_413),
.Y(n_943)
);

AOI22xp5_ASAP7_75t_L g944 ( 
.A1(n_724),
.A2(n_244),
.B1(n_386),
.B2(n_375),
.Y(n_944)
);

INVx1_ASAP7_75t_L g945 ( 
.A(n_765),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_L g946 ( 
.A(n_681),
.B(n_622),
.Y(n_946)
);

INVx1_ASAP7_75t_L g947 ( 
.A(n_765),
.Y(n_947)
);

NAND2xp5_ASAP7_75t_SL g948 ( 
.A(n_648),
.B(n_622),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_681),
.B(n_622),
.Y(n_949)
);

AND2x2_ASAP7_75t_L g950 ( 
.A(n_698),
.B(n_231),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_769),
.Y(n_951)
);

AOI22xp33_ASAP7_75t_L g952 ( 
.A1(n_724),
.A2(n_410),
.B1(n_420),
.B2(n_419),
.Y(n_952)
);

AOI22xp5_ASAP7_75t_L g953 ( 
.A1(n_790),
.A2(n_362),
.B1(n_252),
.B2(n_254),
.Y(n_953)
);

NAND2x1p5_ASAP7_75t_L g954 ( 
.A(n_658),
.B(n_622),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_658),
.B(n_622),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_754),
.B(n_790),
.Y(n_956)
);

NOR2xp33_ASAP7_75t_L g957 ( 
.A(n_770),
.B(n_250),
.Y(n_957)
);

NAND2xp5_ASAP7_75t_SL g958 ( 
.A(n_658),
.B(n_251),
.Y(n_958)
);

OR2x6_ASAP7_75t_L g959 ( 
.A(n_714),
.B(n_419),
.Y(n_959)
);

AND2x4_ASAP7_75t_L g960 ( 
.A(n_748),
.B(n_522),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_SL g961 ( 
.A(n_658),
.B(n_255),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_L g962 ( 
.A(n_789),
.B(n_526),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_804),
.Y(n_963)
);

INVx5_ASAP7_75t_L g964 ( 
.A(n_798),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_804),
.Y(n_965)
);

NOR2xp33_ASAP7_75t_R g966 ( 
.A(n_911),
.B(n_669),
.Y(n_966)
);

AND2x4_ASAP7_75t_L g967 ( 
.A(n_886),
.B(n_748),
.Y(n_967)
);

OR2x2_ASAP7_75t_L g968 ( 
.A(n_820),
.B(n_668),
.Y(n_968)
);

CKINVDCx5p33_ASAP7_75t_R g969 ( 
.A(n_911),
.Y(n_969)
);

INVx2_ASAP7_75t_L g970 ( 
.A(n_807),
.Y(n_970)
);

NAND2xp5_ASAP7_75t_L g971 ( 
.A(n_828),
.B(n_748),
.Y(n_971)
);

NOR3xp33_ASAP7_75t_SL g972 ( 
.A(n_899),
.B(n_785),
.C(n_775),
.Y(n_972)
);

NOR3xp33_ASAP7_75t_SL g973 ( 
.A(n_903),
.B(n_785),
.C(n_775),
.Y(n_973)
);

BUFx12f_ASAP7_75t_L g974 ( 
.A(n_919),
.Y(n_974)
);

NAND2xp5_ASAP7_75t_SL g975 ( 
.A(n_863),
.B(n_855),
.Y(n_975)
);

AND2x4_ASAP7_75t_L g976 ( 
.A(n_886),
.B(n_749),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_805),
.B(n_857),
.Y(n_977)
);

INVx2_ASAP7_75t_L g978 ( 
.A(n_807),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_805),
.B(n_749),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_810),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_L g981 ( 
.A(n_805),
.B(n_749),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_857),
.B(n_789),
.Y(n_982)
);

HB1xp67_ASAP7_75t_L g983 ( 
.A(n_900),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_810),
.Y(n_984)
);

NAND2xp33_ASAP7_75t_R g985 ( 
.A(n_919),
.B(n_762),
.Y(n_985)
);

NAND3xp33_ASAP7_75t_L g986 ( 
.A(n_836),
.B(n_717),
.C(n_722),
.Y(n_986)
);

AND2x2_ASAP7_75t_L g987 ( 
.A(n_826),
.B(n_789),
.Y(n_987)
);

AOI22xp33_ASAP7_75t_L g988 ( 
.A1(n_934),
.A2(n_830),
.B1(n_815),
.B2(n_817),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_811),
.Y(n_989)
);

AOI22xp33_ASAP7_75t_L g990 ( 
.A1(n_934),
.A2(n_650),
.B1(n_674),
.B2(n_679),
.Y(n_990)
);

NAND2xp5_ASAP7_75t_SL g991 ( 
.A(n_873),
.B(n_734),
.Y(n_991)
);

NAND2xp5_ASAP7_75t_L g992 ( 
.A(n_857),
.B(n_647),
.Y(n_992)
);

INVx2_ASAP7_75t_SL g993 ( 
.A(n_915),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_826),
.B(n_647),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_811),
.Y(n_995)
);

INVx2_ASAP7_75t_SL g996 ( 
.A(n_846),
.Y(n_996)
);

BUFx6f_ASAP7_75t_L g997 ( 
.A(n_888),
.Y(n_997)
);

BUFx6f_ASAP7_75t_L g998 ( 
.A(n_888),
.Y(n_998)
);

INVx5_ASAP7_75t_L g999 ( 
.A(n_798),
.Y(n_999)
);

NOR2xp33_ASAP7_75t_L g1000 ( 
.A(n_793),
.B(n_697),
.Y(n_1000)
);

BUFx6f_ASAP7_75t_L g1001 ( 
.A(n_888),
.Y(n_1001)
);

INVx2_ASAP7_75t_L g1002 ( 
.A(n_813),
.Y(n_1002)
);

NAND2xp5_ASAP7_75t_L g1003 ( 
.A(n_846),
.B(n_825),
.Y(n_1003)
);

AOI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_887),
.A2(n_742),
.B1(n_774),
.B2(n_699),
.Y(n_1004)
);

INVx2_ASAP7_75t_SL g1005 ( 
.A(n_860),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_827),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_813),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_845),
.Y(n_1008)
);

INVx2_ASAP7_75t_L g1009 ( 
.A(n_819),
.Y(n_1009)
);

INVx2_ASAP7_75t_L g1010 ( 
.A(n_819),
.Y(n_1010)
);

NAND2xp5_ASAP7_75t_L g1011 ( 
.A(n_851),
.B(n_843),
.Y(n_1011)
);

INVx3_ASAP7_75t_L g1012 ( 
.A(n_831),
.Y(n_1012)
);

HB1xp67_ASAP7_75t_L g1013 ( 
.A(n_795),
.Y(n_1013)
);

INVx2_ASAP7_75t_L g1014 ( 
.A(n_821),
.Y(n_1014)
);

HB1xp67_ASAP7_75t_L g1015 ( 
.A(n_874),
.Y(n_1015)
);

INVx1_ASAP7_75t_L g1016 ( 
.A(n_929),
.Y(n_1016)
);

BUFx5_ASAP7_75t_L g1017 ( 
.A(n_794),
.Y(n_1017)
);

INVx4_ASAP7_75t_L g1018 ( 
.A(n_888),
.Y(n_1018)
);

BUFx3_ASAP7_75t_L g1019 ( 
.A(n_869),
.Y(n_1019)
);

OR2x6_ASAP7_75t_L g1020 ( 
.A(n_798),
.B(n_769),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_884),
.Y(n_1021)
);

CKINVDCx14_ASAP7_75t_R g1022 ( 
.A(n_926),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_931),
.Y(n_1023)
);

INVx1_ASAP7_75t_L g1024 ( 
.A(n_912),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_869),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_874),
.Y(n_1026)
);

INVx2_ASAP7_75t_L g1027 ( 
.A(n_821),
.Y(n_1027)
);

NOR2xp33_ASAP7_75t_R g1028 ( 
.A(n_800),
.B(n_702),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_914),
.Y(n_1029)
);

AND2x4_ASAP7_75t_L g1030 ( 
.A(n_860),
.B(n_776),
.Y(n_1030)
);

BUFx12f_ASAP7_75t_L g1031 ( 
.A(n_872),
.Y(n_1031)
);

CKINVDCx20_ASAP7_75t_R g1032 ( 
.A(n_926),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_843),
.B(n_650),
.Y(n_1033)
);

NAND2xp33_ASAP7_75t_L g1034 ( 
.A(n_928),
.B(n_658),
.Y(n_1034)
);

NOR2xp33_ASAP7_75t_R g1035 ( 
.A(n_809),
.B(n_702),
.Y(n_1035)
);

INVx3_ASAP7_75t_SL g1036 ( 
.A(n_959),
.Y(n_1036)
);

INVx3_ASAP7_75t_L g1037 ( 
.A(n_831),
.Y(n_1037)
);

INVx2_ASAP7_75t_L g1038 ( 
.A(n_837),
.Y(n_1038)
);

NAND3xp33_ASAP7_75t_SL g1039 ( 
.A(n_799),
.B(n_762),
.C(n_705),
.Y(n_1039)
);

NOR3xp33_ASAP7_75t_SL g1040 ( 
.A(n_816),
.B(n_262),
.C(n_260),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_849),
.B(n_814),
.Y(n_1041)
);

BUFx6f_ASAP7_75t_L g1042 ( 
.A(n_925),
.Y(n_1042)
);

INVx2_ASAP7_75t_L g1043 ( 
.A(n_837),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_853),
.Y(n_1044)
);

INVx2_ASAP7_75t_L g1045 ( 
.A(n_853),
.Y(n_1045)
);

INVx2_ASAP7_75t_L g1046 ( 
.A(n_865),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_812),
.Y(n_1047)
);

NAND2xp5_ASAP7_75t_L g1048 ( 
.A(n_818),
.B(n_674),
.Y(n_1048)
);

BUFx4_ASAP7_75t_SL g1049 ( 
.A(n_797),
.Y(n_1049)
);

HB1xp67_ASAP7_75t_L g1050 ( 
.A(n_860),
.Y(n_1050)
);

INVx3_ASAP7_75t_L g1051 ( 
.A(n_831),
.Y(n_1051)
);

INVx3_ASAP7_75t_L g1052 ( 
.A(n_852),
.Y(n_1052)
);

INVx1_ASAP7_75t_L g1053 ( 
.A(n_902),
.Y(n_1053)
);

BUFx4f_ASAP7_75t_L g1054 ( 
.A(n_869),
.Y(n_1054)
);

BUFx6f_ASAP7_75t_SL g1055 ( 
.A(n_959),
.Y(n_1055)
);

BUFx6f_ASAP7_75t_L g1056 ( 
.A(n_925),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_862),
.B(n_776),
.Y(n_1057)
);

OR2x4_ASAP7_75t_L g1058 ( 
.A(n_803),
.B(n_883),
.Y(n_1058)
);

INVx4_ASAP7_75t_L g1059 ( 
.A(n_925),
.Y(n_1059)
);

HB1xp67_ASAP7_75t_L g1060 ( 
.A(n_959),
.Y(n_1060)
);

HB1xp67_ASAP7_75t_L g1061 ( 
.A(n_959),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_887),
.B(n_679),
.Y(n_1062)
);

AND2x4_ASAP7_75t_L g1063 ( 
.A(n_918),
.B(n_780),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_918),
.B(n_680),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_844),
.B(n_734),
.Y(n_1065)
);

INVx2_ASAP7_75t_L g1066 ( 
.A(n_865),
.Y(n_1066)
);

INVx2_ASAP7_75t_L g1067 ( 
.A(n_882),
.Y(n_1067)
);

AND2x4_ASAP7_75t_L g1068 ( 
.A(n_869),
.B(n_780),
.Y(n_1068)
);

OAI21xp5_ASAP7_75t_L g1069 ( 
.A1(n_833),
.A2(n_688),
.B(n_680),
.Y(n_1069)
);

AOI22xp33_ASAP7_75t_L g1070 ( 
.A1(n_840),
.A2(n_738),
.B1(n_735),
.B2(n_688),
.Y(n_1070)
);

NOR3xp33_ASAP7_75t_SL g1071 ( 
.A(n_930),
.B(n_278),
.C(n_264),
.Y(n_1071)
);

AND2x6_ASAP7_75t_L g1072 ( 
.A(n_824),
.B(n_695),
.Y(n_1072)
);

BUFx2_ASAP7_75t_L g1073 ( 
.A(n_870),
.Y(n_1073)
);

INVx2_ASAP7_75t_L g1074 ( 
.A(n_882),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_885),
.Y(n_1075)
);

AOI22xp5_ASAP7_75t_L g1076 ( 
.A1(n_847),
.A2(n_746),
.B1(n_767),
.B2(n_782),
.Y(n_1076)
);

AOI22xp5_ASAP7_75t_L g1077 ( 
.A1(n_858),
.A2(n_881),
.B1(n_913),
.B2(n_892),
.Y(n_1077)
);

HB1xp67_ASAP7_75t_L g1078 ( 
.A(n_870),
.Y(n_1078)
);

NAND2xp5_ASAP7_75t_L g1079 ( 
.A(n_945),
.B(n_695),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_904),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_907),
.Y(n_1081)
);

NAND2xp5_ASAP7_75t_L g1082 ( 
.A(n_947),
.B(n_735),
.Y(n_1082)
);

INVx1_ASAP7_75t_SL g1083 ( 
.A(n_950),
.Y(n_1083)
);

INVx5_ASAP7_75t_L g1084 ( 
.A(n_798),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_909),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_951),
.B(n_737),
.Y(n_1086)
);

INVx2_ASAP7_75t_L g1087 ( 
.A(n_885),
.Y(n_1087)
);

INVx1_ASAP7_75t_L g1088 ( 
.A(n_852),
.Y(n_1088)
);

NOR2xp67_ASAP7_75t_L g1089 ( 
.A(n_957),
.B(n_782),
.Y(n_1089)
);

INVx4_ASAP7_75t_L g1090 ( 
.A(n_925),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_852),
.Y(n_1091)
);

INVx3_ASAP7_75t_L g1092 ( 
.A(n_834),
.Y(n_1092)
);

BUFx6f_ASAP7_75t_L g1093 ( 
.A(n_890),
.Y(n_1093)
);

INVx3_ASAP7_75t_L g1094 ( 
.A(n_834),
.Y(n_1094)
);

NOR2xp33_ASAP7_75t_L g1095 ( 
.A(n_895),
.B(n_734),
.Y(n_1095)
);

AOI22xp33_ASAP7_75t_L g1096 ( 
.A1(n_960),
.A2(n_738),
.B1(n_737),
.B2(n_767),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_871),
.Y(n_1097)
);

NOR3xp33_ASAP7_75t_SL g1098 ( 
.A(n_940),
.B(n_290),
.C(n_286),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_878),
.Y(n_1099)
);

INVx3_ASAP7_75t_L g1100 ( 
.A(n_834),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_880),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_889),
.Y(n_1102)
);

INVx2_ASAP7_75t_L g1103 ( 
.A(n_922),
.Y(n_1103)
);

NAND2xp5_ASAP7_75t_L g1104 ( 
.A(n_960),
.B(n_693),
.Y(n_1104)
);

NAND2x1p5_ASAP7_75t_L g1105 ( 
.A(n_896),
.B(n_640),
.Y(n_1105)
);

INVx3_ASAP7_75t_L g1106 ( 
.A(n_896),
.Y(n_1106)
);

O2A1O1Ixp33_ASAP7_75t_L g1107 ( 
.A1(n_891),
.A2(n_741),
.B(n_787),
.C(n_693),
.Y(n_1107)
);

INVx5_ASAP7_75t_L g1108 ( 
.A(n_890),
.Y(n_1108)
);

NOR2xp33_ASAP7_75t_R g1109 ( 
.A(n_871),
.B(n_292),
.Y(n_1109)
);

AND2x2_ASAP7_75t_L g1110 ( 
.A(n_960),
.B(n_787),
.Y(n_1110)
);

INVx2_ASAP7_75t_L g1111 ( 
.A(n_922),
.Y(n_1111)
);

AND2x4_ASAP7_75t_L g1112 ( 
.A(n_870),
.B(n_644),
.Y(n_1112)
);

BUFx6f_ASAP7_75t_L g1113 ( 
.A(n_890),
.Y(n_1113)
);

AND2x4_ASAP7_75t_L g1114 ( 
.A(n_870),
.B(n_644),
.Y(n_1114)
);

INVx3_ASAP7_75t_SL g1115 ( 
.A(n_958),
.Y(n_1115)
);

NAND2xp5_ASAP7_75t_L g1116 ( 
.A(n_893),
.B(n_728),
.Y(n_1116)
);

NAND2xp33_ASAP7_75t_SL g1117 ( 
.A(n_871),
.B(n_716),
.Y(n_1117)
);

NAND2xp33_ASAP7_75t_SL g1118 ( 
.A(n_841),
.B(n_731),
.Y(n_1118)
);

INVx3_ASAP7_75t_L g1119 ( 
.A(n_896),
.Y(n_1119)
);

HB1xp67_ASAP7_75t_L g1120 ( 
.A(n_962),
.Y(n_1120)
);

INVx1_ASAP7_75t_L g1121 ( 
.A(n_894),
.Y(n_1121)
);

BUFx2_ASAP7_75t_L g1122 ( 
.A(n_866),
.Y(n_1122)
);

HB1xp67_ASAP7_75t_L g1123 ( 
.A(n_935),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_901),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_923),
.Y(n_1125)
);

AND2x2_ASAP7_75t_L g1126 ( 
.A(n_952),
.B(n_728),
.Y(n_1126)
);

NAND2xp5_ASAP7_75t_L g1127 ( 
.A(n_796),
.B(n_689),
.Y(n_1127)
);

BUFx12f_ASAP7_75t_L g1128 ( 
.A(n_910),
.Y(n_1128)
);

AND2x4_ASAP7_75t_L g1129 ( 
.A(n_956),
.B(n_644),
.Y(n_1129)
);

NOR3xp33_ASAP7_75t_SL g1130 ( 
.A(n_910),
.B(n_302),
.C(n_295),
.Y(n_1130)
);

INVx2_ASAP7_75t_L g1131 ( 
.A(n_923),
.Y(n_1131)
);

AOI22xp5_ASAP7_75t_L g1132 ( 
.A1(n_832),
.A2(n_746),
.B1(n_767),
.B2(n_661),
.Y(n_1132)
);

INVx1_ASAP7_75t_L g1133 ( 
.A(n_938),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_802),
.B(n_751),
.Y(n_1134)
);

OR2x2_ASAP7_75t_L g1135 ( 
.A(n_953),
.B(n_526),
.Y(n_1135)
);

OR2x6_ASAP7_75t_L g1136 ( 
.A(n_890),
.B(n_746),
.Y(n_1136)
);

AOI22xp5_ASAP7_75t_L g1137 ( 
.A1(n_833),
.A2(n_746),
.B1(n_767),
.B2(n_661),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_938),
.Y(n_1138)
);

INVx1_ASAP7_75t_L g1139 ( 
.A(n_905),
.Y(n_1139)
);

AND2x2_ASAP7_75t_L g1140 ( 
.A(n_848),
.B(n_944),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_928),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_808),
.B(n_751),
.Y(n_1142)
);

AND2x4_ASAP7_75t_L g1143 ( 
.A(n_927),
.B(n_644),
.Y(n_1143)
);

INVx2_ASAP7_75t_L g1144 ( 
.A(n_921),
.Y(n_1144)
);

NOR3xp33_ASAP7_75t_SL g1145 ( 
.A(n_850),
.B(n_306),
.C(n_303),
.Y(n_1145)
);

BUFx6f_ASAP7_75t_L g1146 ( 
.A(n_801),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_916),
.Y(n_1147)
);

NAND2xp5_ASAP7_75t_L g1148 ( 
.A(n_792),
.B(n_755),
.Y(n_1148)
);

NOR3xp33_ASAP7_75t_L g1149 ( 
.A(n_961),
.B(n_325),
.C(n_322),
.Y(n_1149)
);

BUFx6f_ASAP7_75t_L g1150 ( 
.A(n_806),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_876),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_856),
.Y(n_1152)
);

NAND2xp5_ASAP7_75t_SL g1153 ( 
.A(n_928),
.B(n_731),
.Y(n_1153)
);

BUFx2_ASAP7_75t_L g1154 ( 
.A(n_859),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_942),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_861),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_965),
.Y(n_1157)
);

AOI31xp67_ASAP7_75t_L g1158 ( 
.A1(n_991),
.A2(n_970),
.A3(n_978),
.B(n_965),
.Y(n_1158)
);

AO21x1_ASAP7_75t_L g1159 ( 
.A1(n_1118),
.A2(n_898),
.B(n_823),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_SL g1160 ( 
.A(n_1089),
.B(n_928),
.Y(n_1160)
);

BUFx6f_ASAP7_75t_L g1161 ( 
.A(n_997),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1099),
.B(n_868),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_970),
.Y(n_1163)
);

BUFx4f_ASAP7_75t_SL g1164 ( 
.A(n_974),
.Y(n_1164)
);

OAI21x1_ASAP7_75t_L g1165 ( 
.A1(n_1153),
.A2(n_937),
.B(n_936),
.Y(n_1165)
);

OR2x2_ASAP7_75t_L g1166 ( 
.A(n_968),
.B(n_854),
.Y(n_1166)
);

INVx1_ASAP7_75t_L g1167 ( 
.A(n_978),
.Y(n_1167)
);

OAI21x1_ASAP7_75t_L g1168 ( 
.A1(n_1069),
.A2(n_941),
.B(n_939),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1101),
.B(n_1102),
.Y(n_1169)
);

OAI22xp5_ASAP7_75t_L g1170 ( 
.A1(n_975),
.A2(n_791),
.B1(n_829),
.B2(n_838),
.Y(n_1170)
);

AO31x2_ASAP7_75t_L g1171 ( 
.A1(n_1147),
.A2(n_864),
.A3(n_835),
.B(n_424),
.Y(n_1171)
);

A2O1A1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_975),
.A2(n_943),
.B(n_932),
.C(n_879),
.Y(n_1172)
);

AND2x4_ASAP7_75t_L g1173 ( 
.A(n_1030),
.B(n_854),
.Y(n_1173)
);

AOI221xp5_ASAP7_75t_L g1174 ( 
.A1(n_986),
.A2(n_335),
.B1(n_327),
.B2(n_329),
.C(n_334),
.Y(n_1174)
);

AO31x2_ASAP7_75t_L g1175 ( 
.A1(n_1139),
.A2(n_424),
.A3(n_755),
.B(n_671),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1121),
.B(n_822),
.Y(n_1176)
);

OAI21x1_ASAP7_75t_L g1177 ( 
.A1(n_1153),
.A2(n_949),
.B(n_946),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_1065),
.A2(n_875),
.B(n_906),
.C(n_908),
.Y(n_1178)
);

CKINVDCx8_ASAP7_75t_R g1179 ( 
.A(n_969),
.Y(n_1179)
);

OAI21x1_ASAP7_75t_L g1180 ( 
.A1(n_1105),
.A2(n_933),
.B(n_823),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_963),
.Y(n_1181)
);

OAI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_971),
.A2(n_822),
.B(n_920),
.Y(n_1182)
);

INVx1_ASAP7_75t_SL g1183 ( 
.A(n_1013),
.Y(n_1183)
);

BUFx8_ASAP7_75t_L g1184 ( 
.A(n_1055),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_SL g1185 ( 
.A(n_1077),
.B(n_928),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_1006),
.Y(n_1186)
);

OAI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1140),
.A2(n_920),
.B(n_842),
.Y(n_1187)
);

AND2x2_ASAP7_75t_L g1188 ( 
.A(n_1057),
.B(n_231),
.Y(n_1188)
);

BUFx3_ASAP7_75t_L g1189 ( 
.A(n_974),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_1008),
.Y(n_1190)
);

OAI21x1_ASAP7_75t_L g1191 ( 
.A1(n_1105),
.A2(n_958),
.B(n_961),
.Y(n_1191)
);

OAI21x1_ASAP7_75t_L g1192 ( 
.A1(n_1105),
.A2(n_1037),
.B(n_1012),
.Y(n_1192)
);

OAI21x1_ASAP7_75t_L g1193 ( 
.A1(n_1012),
.A2(n_948),
.B(n_924),
.Y(n_1193)
);

BUFx6f_ASAP7_75t_L g1194 ( 
.A(n_997),
.Y(n_1194)
);

AOI21xp5_ASAP7_75t_L g1195 ( 
.A1(n_1034),
.A2(n_661),
.B(n_640),
.Y(n_1195)
);

AND2x2_ASAP7_75t_L g1196 ( 
.A(n_1057),
.B(n_231),
.Y(n_1196)
);

OAI21x1_ASAP7_75t_L g1197 ( 
.A1(n_1012),
.A2(n_948),
.B(n_924),
.Y(n_1197)
);

INVx2_ASAP7_75t_L g1198 ( 
.A(n_1002),
.Y(n_1198)
);

NOR2x1_ASAP7_75t_SL g1199 ( 
.A(n_1136),
.B(n_867),
.Y(n_1199)
);

OAI21x1_ASAP7_75t_L g1200 ( 
.A1(n_1037),
.A2(n_955),
.B(n_897),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1002),
.Y(n_1201)
);

OAI21x1_ASAP7_75t_L g1202 ( 
.A1(n_1037),
.A2(n_955),
.B(n_897),
.Y(n_1202)
);

BUFx2_ASAP7_75t_L g1203 ( 
.A(n_1026),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_984),
.Y(n_1204)
);

OAI21x1_ASAP7_75t_L g1205 ( 
.A1(n_1051),
.A2(n_867),
.B(n_954),
.Y(n_1205)
);

OAI21x1_ASAP7_75t_SL g1206 ( 
.A1(n_977),
.A2(n_917),
.B(n_671),
.Y(n_1206)
);

AOI21xp5_ASAP7_75t_L g1207 ( 
.A1(n_1034),
.A2(n_671),
.B(n_640),
.Y(n_1207)
);

A2O1A1Ixp33_ASAP7_75t_L g1208 ( 
.A1(n_1095),
.A2(n_875),
.B(n_839),
.C(n_534),
.Y(n_1208)
);

OAI22xp5_ASAP7_75t_L g1209 ( 
.A1(n_988),
.A2(n_979),
.B1(n_982),
.B2(n_981),
.Y(n_1209)
);

NOR2x1_ASAP7_75t_SL g1210 ( 
.A(n_1136),
.B(n_731),
.Y(n_1210)
);

AO31x2_ASAP7_75t_L g1211 ( 
.A1(n_1122),
.A2(n_726),
.A3(n_701),
.B(n_687),
.Y(n_1211)
);

OAI21x1_ASAP7_75t_L g1212 ( 
.A1(n_1051),
.A2(n_954),
.B(n_783),
.Y(n_1212)
);

OAI21x1_ASAP7_75t_L g1213 ( 
.A1(n_1051),
.A2(n_783),
.B(n_928),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_995),
.Y(n_1214)
);

AOI22xp5_ASAP7_75t_SL g1215 ( 
.A1(n_1000),
.A2(n_406),
.B1(n_405),
.B2(n_402),
.Y(n_1215)
);

AO31x2_ASAP7_75t_L g1216 ( 
.A1(n_1122),
.A2(n_687),
.A3(n_701),
.B(n_726),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1141),
.A2(n_701),
.B(n_726),
.Y(n_1217)
);

OAI21x1_ASAP7_75t_L g1218 ( 
.A1(n_1052),
.A2(n_783),
.B(n_928),
.Y(n_1218)
);

BUFx6f_ASAP7_75t_L g1219 ( 
.A(n_997),
.Y(n_1219)
);

A2O1A1Ixp33_ASAP7_75t_L g1220 ( 
.A1(n_996),
.A2(n_839),
.B(n_545),
.C(n_542),
.Y(n_1220)
);

OAI22xp5_ASAP7_75t_L g1221 ( 
.A1(n_1058),
.A2(n_700),
.B1(n_666),
.B2(n_683),
.Y(n_1221)
);

AOI221x1_ASAP7_75t_L g1222 ( 
.A1(n_1118),
.A2(n_1149),
.B1(n_1117),
.B2(n_1039),
.C(n_1140),
.Y(n_1222)
);

OR2x2_ASAP7_75t_L g1223 ( 
.A(n_968),
.B(n_528),
.Y(n_1223)
);

OAI21xp5_ASAP7_75t_L g1224 ( 
.A1(n_1107),
.A2(n_687),
.B(n_767),
.Y(n_1224)
);

NOR2xp33_ASAP7_75t_L g1225 ( 
.A(n_1058),
.B(n_336),
.Y(n_1225)
);

BUFx3_ASAP7_75t_L g1226 ( 
.A(n_1032),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1052),
.A2(n_545),
.B(n_528),
.Y(n_1227)
);

AOI21xp5_ASAP7_75t_SL g1228 ( 
.A1(n_1141),
.A2(n_747),
.B(n_731),
.Y(n_1228)
);

OAI21x1_ASAP7_75t_L g1229 ( 
.A1(n_1052),
.A2(n_534),
.B(n_537),
.Y(n_1229)
);

NOR2x1_ASAP7_75t_L g1230 ( 
.A(n_1019),
.B(n_537),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1124),
.B(n_666),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_1141),
.A2(n_877),
.B(n_700),
.Y(n_1232)
);

AOI21xp33_ASAP7_75t_L g1233 ( 
.A1(n_993),
.A2(n_354),
.B(n_351),
.Y(n_1233)
);

NAND2xp33_ASAP7_75t_L g1234 ( 
.A(n_964),
.B(n_767),
.Y(n_1234)
);

OAI22xp5_ASAP7_75t_L g1235 ( 
.A1(n_1041),
.A2(n_700),
.B1(n_666),
.B2(n_683),
.Y(n_1235)
);

AND2x2_ASAP7_75t_L g1236 ( 
.A(n_993),
.B(n_231),
.Y(n_1236)
);

OAI22xp5_ASAP7_75t_L g1237 ( 
.A1(n_1024),
.A2(n_700),
.B1(n_666),
.B2(n_683),
.Y(n_1237)
);

OA21x2_ASAP7_75t_L g1238 ( 
.A1(n_1156),
.A2(n_539),
.B(n_542),
.Y(n_1238)
);

AO31x2_ASAP7_75t_L g1239 ( 
.A1(n_1116),
.A2(n_539),
.A3(n_467),
.B(n_469),
.Y(n_1239)
);

OAI21x1_ASAP7_75t_L g1240 ( 
.A1(n_1144),
.A2(n_465),
.B(n_467),
.Y(n_1240)
);

AOI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1083),
.A2(n_342),
.B(n_343),
.Y(n_1241)
);

OR2x6_ASAP7_75t_L g1242 ( 
.A(n_1020),
.B(n_1005),
.Y(n_1242)
);

OAI22xp5_ASAP7_75t_L g1243 ( 
.A1(n_1029),
.A2(n_700),
.B1(n_666),
.B2(n_683),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1144),
.A2(n_465),
.B(n_469),
.Y(n_1244)
);

INVx5_ASAP7_75t_L g1245 ( 
.A(n_1136),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1104),
.A2(n_877),
.B(n_409),
.Y(n_1246)
);

AO32x2_ASAP7_75t_L g1247 ( 
.A1(n_996),
.A2(n_235),
.A3(n_249),
.B1(n_338),
.B2(n_19),
.Y(n_1247)
);

NAND3x1_ASAP7_75t_L g1248 ( 
.A(n_1004),
.B(n_235),
.C(n_249),
.Y(n_1248)
);

A2O1A1Ixp33_ASAP7_75t_L g1249 ( 
.A1(n_1003),
.A2(n_400),
.B(n_429),
.C(n_428),
.Y(n_1249)
);

BUFx10_ASAP7_75t_L g1250 ( 
.A(n_969),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_980),
.Y(n_1251)
);

AOI21xp5_ASAP7_75t_L g1252 ( 
.A1(n_1092),
.A2(n_877),
.B(n_683),
.Y(n_1252)
);

OAI21x1_ASAP7_75t_L g1253 ( 
.A1(n_980),
.A2(n_877),
.B(n_752),
.Y(n_1253)
);

AOI21xp5_ASAP7_75t_L g1254 ( 
.A1(n_1092),
.A2(n_877),
.B(n_707),
.Y(n_1254)
);

BUFx3_ASAP7_75t_L g1255 ( 
.A(n_1032),
.Y(n_1255)
);

BUFx8_ASAP7_75t_L g1256 ( 
.A(n_1055),
.Y(n_1256)
);

OAI21xp5_ASAP7_75t_L g1257 ( 
.A1(n_1053),
.A2(n_347),
.B(n_361),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1021),
.B(n_707),
.Y(n_1258)
);

BUFx6f_ASAP7_75t_L g1259 ( 
.A(n_997),
.Y(n_1259)
);

AOI21xp5_ASAP7_75t_L g1260 ( 
.A1(n_1092),
.A2(n_1100),
.B(n_1094),
.Y(n_1260)
);

NAND3xp33_ASAP7_75t_L g1261 ( 
.A(n_1040),
.B(n_398),
.C(n_426),
.Y(n_1261)
);

NOR2xp67_ASAP7_75t_SL g1262 ( 
.A(n_1108),
.B(n_731),
.Y(n_1262)
);

NAND2xp5_ASAP7_75t_L g1263 ( 
.A(n_987),
.B(n_707),
.Y(n_1263)
);

OAI21x1_ASAP7_75t_L g1264 ( 
.A1(n_989),
.A2(n_747),
.B(n_752),
.Y(n_1264)
);

OAI21x1_ASAP7_75t_L g1265 ( 
.A1(n_989),
.A2(n_747),
.B(n_752),
.Y(n_1265)
);

AND2x2_ASAP7_75t_L g1266 ( 
.A(n_1110),
.B(n_235),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1007),
.A2(n_747),
.B(n_752),
.Y(n_1267)
);

AOI21xp5_ASAP7_75t_L g1268 ( 
.A1(n_1094),
.A2(n_707),
.B(n_752),
.Y(n_1268)
);

NAND2xp5_ASAP7_75t_L g1269 ( 
.A(n_987),
.B(n_707),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1005),
.A2(n_1080),
.B1(n_1085),
.B2(n_1081),
.Y(n_1270)
);

AO31x2_ASAP7_75t_L g1271 ( 
.A1(n_1023),
.A2(n_1151),
.A3(n_1016),
.B(n_994),
.Y(n_1271)
);

OAI21x1_ASAP7_75t_L g1272 ( 
.A1(n_1007),
.A2(n_747),
.B(n_101),
.Y(n_1272)
);

AND2x2_ASAP7_75t_L g1273 ( 
.A(n_1110),
.B(n_235),
.Y(n_1273)
);

NAND2xp5_ASAP7_75t_SL g1274 ( 
.A(n_1068),
.B(n_363),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_1125),
.Y(n_1275)
);

OAI21xp5_ASAP7_75t_L g1276 ( 
.A1(n_992),
.A2(n_364),
.B(n_390),
.Y(n_1276)
);

OAI22x1_ASAP7_75t_L g1277 ( 
.A1(n_1036),
.A2(n_418),
.B1(n_417),
.B2(n_414),
.Y(n_1277)
);

OAI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1148),
.A2(n_393),
.B(n_394),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1120),
.B(n_397),
.Y(n_1279)
);

NAND2xp5_ASAP7_75t_L g1280 ( 
.A(n_1063),
.B(n_408),
.Y(n_1280)
);

A2O1A1Ixp33_ASAP7_75t_L g1281 ( 
.A1(n_991),
.A2(n_338),
.B(n_249),
.C(n_18),
.Y(n_1281)
);

AOI21xp5_ASAP7_75t_L g1282 ( 
.A1(n_1094),
.A2(n_1106),
.B(n_1100),
.Y(n_1282)
);

OAI21xp5_ASAP7_75t_L g1283 ( 
.A1(n_1134),
.A2(n_180),
.B(n_112),
.Y(n_1283)
);

INVxp67_ASAP7_75t_SL g1284 ( 
.A(n_1100),
.Y(n_1284)
);

OAI21x1_ASAP7_75t_L g1285 ( 
.A1(n_1009),
.A2(n_173),
.B(n_116),
.Y(n_1285)
);

AOI21xp5_ASAP7_75t_L g1286 ( 
.A1(n_1106),
.A2(n_1119),
.B(n_1108),
.Y(n_1286)
);

NAND2xp33_ASAP7_75t_L g1287 ( 
.A(n_964),
.B(n_773),
.Y(n_1287)
);

AOI31xp67_ASAP7_75t_L g1288 ( 
.A1(n_1076),
.A2(n_181),
.A3(n_120),
.B(n_217),
.Y(n_1288)
);

AOI21xp5_ASAP7_75t_L g1289 ( 
.A1(n_1106),
.A2(n_788),
.B(n_773),
.Y(n_1289)
);

AOI21xp5_ASAP7_75t_L g1290 ( 
.A1(n_1119),
.A2(n_788),
.B(n_773),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1133),
.Y(n_1291)
);

INVx4_ASAP7_75t_SL g1292 ( 
.A(n_997),
.Y(n_1292)
);

NAND2xp5_ASAP7_75t_L g1293 ( 
.A(n_1063),
.B(n_249),
.Y(n_1293)
);

NAND2xp5_ASAP7_75t_L g1294 ( 
.A(n_1063),
.B(n_338),
.Y(n_1294)
);

INVx1_ASAP7_75t_L g1295 ( 
.A(n_1009),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1030),
.B(n_338),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1030),
.B(n_9),
.Y(n_1297)
);

INVx4_ASAP7_75t_L g1298 ( 
.A(n_1054),
.Y(n_1298)
);

OAI21x1_ASAP7_75t_L g1299 ( 
.A1(n_1010),
.A2(n_182),
.B(n_133),
.Y(n_1299)
);

OAI21x1_ASAP7_75t_L g1300 ( 
.A1(n_1119),
.A2(n_184),
.B(n_134),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_L g1301 ( 
.A1(n_1142),
.A2(n_185),
.B(n_136),
.Y(n_1301)
);

OAI21x1_ASAP7_75t_L g1302 ( 
.A1(n_1010),
.A2(n_1027),
.B(n_1014),
.Y(n_1302)
);

NAND2xp5_ASAP7_75t_L g1303 ( 
.A(n_1151),
.B(n_16),
.Y(n_1303)
);

BUFx3_ASAP7_75t_L g1304 ( 
.A(n_1026),
.Y(n_1304)
);

OAI21x1_ASAP7_75t_L g1305 ( 
.A1(n_1014),
.A2(n_187),
.B(n_140),
.Y(n_1305)
);

AOI21xp5_ASAP7_75t_L g1306 ( 
.A1(n_1108),
.A2(n_788),
.B(n_773),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1015),
.B(n_18),
.Y(n_1307)
);

BUFx6f_ASAP7_75t_L g1308 ( 
.A(n_998),
.Y(n_1308)
);

OAI21xp5_ASAP7_75t_L g1309 ( 
.A1(n_1127),
.A2(n_172),
.B(n_206),
.Y(n_1309)
);

AOI21xp5_ASAP7_75t_SL g1310 ( 
.A1(n_1093),
.A2(n_788),
.B(n_201),
.Y(n_1310)
);

AOI21xp5_ASAP7_75t_L g1311 ( 
.A1(n_1108),
.A2(n_788),
.B(n_190),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_983),
.B(n_20),
.Y(n_1312)
);

AND2x2_ASAP7_75t_L g1313 ( 
.A(n_1050),
.B(n_21),
.Y(n_1313)
);

AOI21xp5_ASAP7_75t_L g1314 ( 
.A1(n_1108),
.A2(n_188),
.B(n_164),
.Y(n_1314)
);

OAI21x1_ASAP7_75t_L g1315 ( 
.A1(n_1027),
.A2(n_146),
.B(n_144),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1071),
.B(n_22),
.C(n_27),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1068),
.B(n_104),
.Y(n_1317)
);

AND2x4_ASAP7_75t_L g1318 ( 
.A(n_1068),
.B(n_28),
.Y(n_1318)
);

OAI21x1_ASAP7_75t_L g1319 ( 
.A1(n_1038),
.A2(n_29),
.B(n_31),
.Y(n_1319)
);

OAI21x1_ASAP7_75t_L g1320 ( 
.A1(n_1038),
.A2(n_31),
.B(n_32),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1043),
.A2(n_33),
.B(n_35),
.Y(n_1321)
);

NAND2xp5_ASAP7_75t_L g1322 ( 
.A(n_1011),
.B(n_37),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_SL g1323 ( 
.A(n_1146),
.B(n_39),
.Y(n_1323)
);

INVx3_ASAP7_75t_L g1324 ( 
.A(n_1245),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1264),
.A2(n_1064),
.B(n_1062),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1265),
.A2(n_1070),
.B(n_1046),
.Y(n_1326)
);

OAI22xp5_ASAP7_75t_L g1327 ( 
.A1(n_1169),
.A2(n_1155),
.B1(n_1123),
.B2(n_1152),
.Y(n_1327)
);

OAI21x1_ASAP7_75t_SL g1328 ( 
.A1(n_1199),
.A2(n_1048),
.B(n_1086),
.Y(n_1328)
);

INVx2_ASAP7_75t_L g1329 ( 
.A(n_1163),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_L g1330 ( 
.A1(n_1225),
.A2(n_1155),
.B1(n_1154),
.B2(n_1152),
.Y(n_1330)
);

NAND2x1p5_ASAP7_75t_L g1331 ( 
.A(n_1245),
.B(n_964),
.Y(n_1331)
);

A2O1A1Ixp33_ASAP7_75t_L g1332 ( 
.A1(n_1178),
.A2(n_1098),
.B(n_1145),
.C(n_1135),
.Y(n_1332)
);

AO21x2_ASAP7_75t_L g1333 ( 
.A1(n_1224),
.A2(n_1132),
.B(n_1137),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_1163),
.Y(n_1334)
);

NAND2xp5_ASAP7_75t_L g1335 ( 
.A(n_1188),
.B(n_1135),
.Y(n_1335)
);

AND2x4_ASAP7_75t_L g1336 ( 
.A(n_1245),
.B(n_967),
.Y(n_1336)
);

INVx4_ASAP7_75t_L g1337 ( 
.A(n_1245),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1228),
.A2(n_964),
.B(n_1084),
.Y(n_1338)
);

NAND3xp33_ASAP7_75t_L g1339 ( 
.A(n_1215),
.B(n_973),
.C(n_985),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_SL g1340 ( 
.A1(n_1159),
.A2(n_1079),
.B(n_1082),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1186),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1190),
.Y(n_1342)
);

HB1xp67_ASAP7_75t_L g1343 ( 
.A(n_1203),
.Y(n_1343)
);

AO21x2_ASAP7_75t_L g1344 ( 
.A1(n_1208),
.A2(n_1033),
.B(n_1130),
.Y(n_1344)
);

AND2x2_ASAP7_75t_L g1345 ( 
.A(n_1318),
.B(n_1126),
.Y(n_1345)
);

OAI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1267),
.A2(n_1067),
.B(n_1111),
.Y(n_1346)
);

AO21x2_ASAP7_75t_L g1347 ( 
.A1(n_1208),
.A2(n_1088),
.B(n_1091),
.Y(n_1347)
);

OAI21xp5_ASAP7_75t_L g1348 ( 
.A1(n_1209),
.A2(n_990),
.B(n_1126),
.Y(n_1348)
);

CKINVDCx11_ASAP7_75t_R g1349 ( 
.A(n_1179),
.Y(n_1349)
);

AND2x4_ASAP7_75t_L g1350 ( 
.A(n_1242),
.B(n_967),
.Y(n_1350)
);

INVxp67_ASAP7_75t_L g1351 ( 
.A(n_1183),
.Y(n_1351)
);

AO21x1_ASAP7_75t_L g1352 ( 
.A1(n_1309),
.A2(n_1117),
.B(n_1047),
.Y(n_1352)
);

AND2x4_ASAP7_75t_L g1353 ( 
.A(n_1242),
.B(n_967),
.Y(n_1353)
);

OAI22xp5_ASAP7_75t_L g1354 ( 
.A1(n_1284),
.A2(n_1154),
.B1(n_1054),
.B2(n_976),
.Y(n_1354)
);

AO21x2_ASAP7_75t_L g1355 ( 
.A1(n_1246),
.A2(n_1067),
.B(n_1046),
.Y(n_1355)
);

AO21x2_ASAP7_75t_L g1356 ( 
.A1(n_1206),
.A2(n_1066),
.B(n_1044),
.Y(n_1356)
);

OAI21x1_ASAP7_75t_SL g1357 ( 
.A1(n_1210),
.A2(n_1018),
.B(n_1059),
.Y(n_1357)
);

NOR2xp33_ASAP7_75t_L g1358 ( 
.A(n_1233),
.B(n_1036),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1198),
.Y(n_1359)
);

INVx3_ASAP7_75t_L g1360 ( 
.A(n_1192),
.Y(n_1360)
);

AO31x2_ASAP7_75t_L g1361 ( 
.A1(n_1220),
.A2(n_1087),
.A3(n_1045),
.B(n_1066),
.Y(n_1361)
);

OAI21x1_ASAP7_75t_L g1362 ( 
.A1(n_1272),
.A2(n_1075),
.B(n_1138),
.Y(n_1362)
);

BUFx10_ASAP7_75t_L g1363 ( 
.A(n_1225),
.Y(n_1363)
);

INVxp67_ASAP7_75t_L g1364 ( 
.A(n_1223),
.Y(n_1364)
);

INVx2_ASAP7_75t_L g1365 ( 
.A(n_1198),
.Y(n_1365)
);

AOI22xp33_ASAP7_75t_L g1366 ( 
.A1(n_1173),
.A2(n_1128),
.B1(n_1061),
.B2(n_1060),
.Y(n_1366)
);

NAND2xp5_ASAP7_75t_SL g1367 ( 
.A(n_1304),
.B(n_966),
.Y(n_1367)
);

AOI22xp33_ASAP7_75t_L g1368 ( 
.A1(n_1173),
.A2(n_1128),
.B1(n_1055),
.B2(n_976),
.Y(n_1368)
);

OAI21x1_ASAP7_75t_L g1369 ( 
.A1(n_1177),
.A2(n_1074),
.B(n_1075),
.Y(n_1369)
);

BUFx3_ASAP7_75t_L g1370 ( 
.A(n_1304),
.Y(n_1370)
);

AND2x2_ASAP7_75t_L g1371 ( 
.A(n_1318),
.B(n_976),
.Y(n_1371)
);

OA21x2_ASAP7_75t_L g1372 ( 
.A1(n_1240),
.A2(n_1045),
.B(n_1074),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1204),
.Y(n_1373)
);

AOI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1185),
.A2(n_1087),
.B(n_1043),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1214),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1201),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1250),
.Y(n_1377)
);

OA21x2_ASAP7_75t_L g1378 ( 
.A1(n_1240),
.A2(n_1111),
.B(n_1103),
.Y(n_1378)
);

AOI221xp5_ASAP7_75t_L g1379 ( 
.A1(n_1174),
.A2(n_972),
.B1(n_1035),
.B2(n_1109),
.C(n_1028),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1275),
.Y(n_1380)
);

OA21x2_ASAP7_75t_L g1381 ( 
.A1(n_1244),
.A2(n_1103),
.B(n_1138),
.Y(n_1381)
);

OAI22xp5_ASAP7_75t_L g1382 ( 
.A1(n_1284),
.A2(n_1054),
.B1(n_964),
.B2(n_999),
.Y(n_1382)
);

AOI22xp33_ASAP7_75t_SL g1383 ( 
.A1(n_1184),
.A2(n_1022),
.B1(n_1097),
.B2(n_1031),
.Y(n_1383)
);

OAI21xp5_ASAP7_75t_L g1384 ( 
.A1(n_1178),
.A2(n_1096),
.B(n_1072),
.Y(n_1384)
);

OAI21x1_ASAP7_75t_L g1385 ( 
.A1(n_1177),
.A2(n_1131),
.B(n_1044),
.Y(n_1385)
);

AND2x4_ASAP7_75t_L g1386 ( 
.A(n_1242),
.B(n_1114),
.Y(n_1386)
);

NAND2x1p5_ASAP7_75t_L g1387 ( 
.A(n_1192),
.B(n_1084),
.Y(n_1387)
);

OAI21x1_ASAP7_75t_L g1388 ( 
.A1(n_1302),
.A2(n_1131),
.B(n_1078),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1196),
.B(n_1073),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1291),
.Y(n_1390)
);

INVx2_ASAP7_75t_L g1391 ( 
.A(n_1201),
.Y(n_1391)
);

OAI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1302),
.A2(n_1072),
.B(n_1017),
.Y(n_1392)
);

OR2x2_ASAP7_75t_L g1393 ( 
.A(n_1271),
.B(n_1115),
.Y(n_1393)
);

OAI21x1_ASAP7_75t_L g1394 ( 
.A1(n_1165),
.A2(n_1072),
.B(n_1017),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1180),
.A2(n_1072),
.B(n_1017),
.Y(n_1395)
);

AND2x4_ASAP7_75t_L g1396 ( 
.A(n_1173),
.B(n_1114),
.Y(n_1396)
);

OR2x6_ASAP7_75t_L g1397 ( 
.A(n_1298),
.B(n_1020),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_SL g1398 ( 
.A1(n_1283),
.A2(n_1059),
.B(n_1090),
.Y(n_1398)
);

BUFx10_ASAP7_75t_L g1399 ( 
.A(n_1318),
.Y(n_1399)
);

NOR2xp33_ASAP7_75t_L g1400 ( 
.A(n_1166),
.B(n_1022),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_1181),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1226),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1251),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1157),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1253),
.A2(n_1229),
.B(n_1227),
.Y(n_1405)
);

OAI221xp5_ASAP7_75t_L g1406 ( 
.A1(n_1257),
.A2(n_1115),
.B1(n_1097),
.B2(n_1073),
.C(n_1020),
.Y(n_1406)
);

NAND2x1p5_ASAP7_75t_L g1407 ( 
.A(n_1262),
.B(n_999),
.Y(n_1407)
);

INVx2_ASAP7_75t_L g1408 ( 
.A(n_1295),
.Y(n_1408)
);

OR2x6_ASAP7_75t_L g1409 ( 
.A(n_1298),
.B(n_1020),
.Y(n_1409)
);

BUFx6f_ASAP7_75t_L g1410 ( 
.A(n_1161),
.Y(n_1410)
);

BUFx3_ASAP7_75t_L g1411 ( 
.A(n_1226),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1167),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_1303),
.Y(n_1413)
);

AOI22xp5_ASAP7_75t_L g1414 ( 
.A1(n_1274),
.A2(n_1031),
.B1(n_1017),
.B2(n_1025),
.Y(n_1414)
);

OAI21x1_ASAP7_75t_L g1415 ( 
.A1(n_1213),
.A2(n_1072),
.B(n_1017),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1230),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1158),
.Y(n_1417)
);

A2O1A1Ixp33_ASAP7_75t_L g1418 ( 
.A1(n_1301),
.A2(n_1129),
.B(n_1025),
.C(n_1019),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1241),
.B(n_1150),
.Y(n_1419)
);

INVx1_ASAP7_75t_L g1420 ( 
.A(n_1271),
.Y(n_1420)
);

O2A1O1Ixp33_ASAP7_75t_SL g1421 ( 
.A1(n_1185),
.A2(n_1017),
.B(n_1072),
.C(n_1146),
.Y(n_1421)
);

CKINVDCx12_ASAP7_75t_R g1422 ( 
.A(n_1312),
.Y(n_1422)
);

AOI222xp33_ASAP7_75t_L g1423 ( 
.A1(n_1281),
.A2(n_1049),
.B1(n_1146),
.B2(n_1150),
.C1(n_1129),
.C2(n_1143),
.Y(n_1423)
);

BUFx2_ASAP7_75t_SL g1424 ( 
.A(n_1255),
.Y(n_1424)
);

INVx1_ASAP7_75t_L g1425 ( 
.A(n_1271),
.Y(n_1425)
);

AOI22xp33_ASAP7_75t_L g1426 ( 
.A1(n_1274),
.A2(n_1150),
.B1(n_1146),
.B2(n_1017),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_L g1427 ( 
.A(n_1162),
.B(n_1266),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1238),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1161),
.Y(n_1429)
);

OA21x2_ASAP7_75t_L g1430 ( 
.A1(n_1319),
.A2(n_1129),
.B(n_1143),
.Y(n_1430)
);

NAND3xp33_ASAP7_75t_L g1431 ( 
.A(n_1316),
.B(n_1150),
.C(n_1146),
.Y(n_1431)
);

INVx3_ASAP7_75t_L g1432 ( 
.A(n_1161),
.Y(n_1432)
);

BUFx4_ASAP7_75t_R g1433 ( 
.A(n_1250),
.Y(n_1433)
);

AOI22xp33_ASAP7_75t_L g1434 ( 
.A1(n_1278),
.A2(n_1150),
.B1(n_1143),
.B2(n_1114),
.Y(n_1434)
);

AND2x4_ASAP7_75t_L g1435 ( 
.A(n_1292),
.B(n_1112),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1271),
.Y(n_1436)
);

INVxp33_ASAP7_75t_L g1437 ( 
.A(n_1236),
.Y(n_1437)
);

INVx2_ASAP7_75t_L g1438 ( 
.A(n_1238),
.Y(n_1438)
);

NAND2x1p5_ASAP7_75t_L g1439 ( 
.A(n_1317),
.B(n_999),
.Y(n_1439)
);

AND2x4_ASAP7_75t_L g1440 ( 
.A(n_1292),
.B(n_1112),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1273),
.B(n_1112),
.Y(n_1441)
);

OAI22xp5_ASAP7_75t_L g1442 ( 
.A1(n_1270),
.A2(n_1084),
.B1(n_999),
.B2(n_1136),
.Y(n_1442)
);

OAI21x1_ASAP7_75t_L g1443 ( 
.A1(n_1218),
.A2(n_999),
.B(n_1084),
.Y(n_1443)
);

INVx3_ASAP7_75t_SL g1444 ( 
.A(n_1250),
.Y(n_1444)
);

OR2x2_ASAP7_75t_L g1445 ( 
.A(n_1176),
.B(n_1018),
.Y(n_1445)
);

O2A1O1Ixp33_ASAP7_75t_SL g1446 ( 
.A1(n_1317),
.A2(n_1056),
.B(n_1001),
.C(n_1042),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1168),
.A2(n_1191),
.B(n_1299),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1238),
.Y(n_1448)
);

OAI21x1_ASAP7_75t_L g1449 ( 
.A1(n_1168),
.A2(n_1084),
.B(n_1113),
.Y(n_1449)
);

BUFx3_ASAP7_75t_L g1450 ( 
.A(n_1255),
.Y(n_1450)
);

OAI21x1_ASAP7_75t_SL g1451 ( 
.A1(n_1286),
.A2(n_1090),
.B(n_1059),
.Y(n_1451)
);

BUFx2_ASAP7_75t_L g1452 ( 
.A(n_1292),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_SL g1453 ( 
.A1(n_1281),
.A2(n_1042),
.B(n_1001),
.C(n_998),
.Y(n_1453)
);

AOI22xp33_ASAP7_75t_L g1454 ( 
.A1(n_1297),
.A2(n_1018),
.B1(n_1090),
.B2(n_998),
.Y(n_1454)
);

NOR2x1_ASAP7_75t_SL g1455 ( 
.A(n_1161),
.B(n_1113),
.Y(n_1455)
);

AOI22xp33_ASAP7_75t_L g1456 ( 
.A1(n_1313),
.A2(n_1056),
.B1(n_1042),
.B2(n_1001),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1175),
.Y(n_1457)
);

AO21x2_ASAP7_75t_L g1458 ( 
.A1(n_1220),
.A2(n_1056),
.B(n_1042),
.Y(n_1458)
);

INVx6_ASAP7_75t_SL g1459 ( 
.A(n_1164),
.Y(n_1459)
);

INVx2_ASAP7_75t_L g1460 ( 
.A(n_1171),
.Y(n_1460)
);

INVx2_ASAP7_75t_L g1461 ( 
.A(n_1171),
.Y(n_1461)
);

OAI22xp5_ASAP7_75t_L g1462 ( 
.A1(n_1258),
.A2(n_1113),
.B1(n_1093),
.B2(n_1056),
.Y(n_1462)
);

INVx6_ASAP7_75t_L g1463 ( 
.A(n_1194),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1191),
.A2(n_1285),
.B(n_1305),
.Y(n_1464)
);

INVx2_ASAP7_75t_SL g1465 ( 
.A(n_1194),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1164),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1307),
.B(n_1056),
.Y(n_1467)
);

A2O1A1Ixp33_ASAP7_75t_L g1468 ( 
.A1(n_1249),
.A2(n_1113),
.B(n_1093),
.C(n_1042),
.Y(n_1468)
);

O2A1O1Ixp33_ASAP7_75t_SL g1469 ( 
.A1(n_1323),
.A2(n_1001),
.B(n_998),
.C(n_1113),
.Y(n_1469)
);

OAI21xp5_ASAP7_75t_L g1470 ( 
.A1(n_1187),
.A2(n_1001),
.B(n_998),
.Y(n_1470)
);

AND2x4_ASAP7_75t_L g1471 ( 
.A(n_1222),
.B(n_1093),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1305),
.A2(n_1315),
.B(n_1200),
.Y(n_1472)
);

OAI21x1_ASAP7_75t_L g1473 ( 
.A1(n_1315),
.A2(n_1093),
.B(n_40),
.Y(n_1473)
);

OAI21x1_ASAP7_75t_L g1474 ( 
.A1(n_1200),
.A2(n_39),
.B(n_41),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_1194),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1175),
.Y(n_1476)
);

OR2x6_ASAP7_75t_L g1477 ( 
.A(n_1323),
.B(n_41),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1175),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1194),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1219),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1175),
.Y(n_1481)
);

INVx2_ASAP7_75t_L g1482 ( 
.A(n_1171),
.Y(n_1482)
);

AND2x4_ASAP7_75t_L g1483 ( 
.A(n_1263),
.B(n_1269),
.Y(n_1483)
);

AO21x2_ASAP7_75t_L g1484 ( 
.A1(n_1182),
.A2(n_45),
.B(n_46),
.Y(n_1484)
);

O2A1O1Ixp33_ASAP7_75t_L g1485 ( 
.A1(n_1249),
.A2(n_45),
.B(n_47),
.C(n_51),
.Y(n_1485)
);

INVx2_ASAP7_75t_SL g1486 ( 
.A(n_1219),
.Y(n_1486)
);

BUFx2_ASAP7_75t_SL g1487 ( 
.A(n_1219),
.Y(n_1487)
);

OR2x2_ASAP7_75t_L g1488 ( 
.A(n_1322),
.B(n_47),
.Y(n_1488)
);

OAI21x1_ASAP7_75t_L g1489 ( 
.A1(n_1202),
.A2(n_51),
.B(n_52),
.Y(n_1489)
);

BUFx2_ASAP7_75t_L g1490 ( 
.A(n_1219),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1231),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1172),
.A2(n_54),
.B1(n_56),
.B2(n_57),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1293),
.Y(n_1493)
);

OAI21x1_ASAP7_75t_L g1494 ( 
.A1(n_1202),
.A2(n_57),
.B(n_58),
.Y(n_1494)
);

HB1xp67_ASAP7_75t_L g1495 ( 
.A(n_1296),
.Y(n_1495)
);

AO31x2_ASAP7_75t_L g1496 ( 
.A1(n_1170),
.A2(n_58),
.A3(n_59),
.B(n_61),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1184),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1294),
.Y(n_1498)
);

OA21x2_ASAP7_75t_L g1499 ( 
.A1(n_1319),
.A2(n_1321),
.B(n_1320),
.Y(n_1499)
);

OAI21x1_ASAP7_75t_L g1500 ( 
.A1(n_1300),
.A2(n_62),
.B(n_63),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1171),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1280),
.Y(n_1502)
);

HB1xp67_ASAP7_75t_L g1503 ( 
.A(n_1393),
.Y(n_1503)
);

OA21x2_ASAP7_75t_L g1504 ( 
.A1(n_1472),
.A2(n_1321),
.B(n_1320),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1492),
.A2(n_1276),
.B1(n_1277),
.B2(n_1261),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1341),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1329),
.Y(n_1507)
);

O2A1O1Ixp33_ASAP7_75t_SL g1508 ( 
.A1(n_1332),
.A2(n_1468),
.B(n_1418),
.C(n_1384),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1345),
.B(n_1279),
.Y(n_1509)
);

HB1xp67_ASAP7_75t_L g1510 ( 
.A(n_1393),
.Y(n_1510)
);

OR2x2_ASAP7_75t_L g1511 ( 
.A(n_1364),
.B(n_1189),
.Y(n_1511)
);

AND2x2_ASAP7_75t_L g1512 ( 
.A(n_1345),
.B(n_1247),
.Y(n_1512)
);

AOI22xp33_ASAP7_75t_SL g1513 ( 
.A1(n_1358),
.A2(n_1256),
.B1(n_1184),
.B2(n_1189),
.Y(n_1513)
);

AND2x2_ASAP7_75t_L g1514 ( 
.A(n_1330),
.B(n_1247),
.Y(n_1514)
);

AOI221xp5_ASAP7_75t_SL g1515 ( 
.A1(n_1485),
.A2(n_1221),
.B1(n_1248),
.B2(n_1243),
.C(n_1237),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1327),
.B(n_1256),
.Y(n_1516)
);

AOI22xp5_ASAP7_75t_L g1517 ( 
.A1(n_1339),
.A2(n_1248),
.B1(n_1256),
.B2(n_1160),
.Y(n_1517)
);

INVxp67_ASAP7_75t_SL g1518 ( 
.A(n_1470),
.Y(n_1518)
);

BUFx6f_ASAP7_75t_L g1519 ( 
.A(n_1435),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1467),
.B(n_1247),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1467),
.B(n_1247),
.Y(n_1521)
);

OR2x2_ASAP7_75t_L g1522 ( 
.A(n_1335),
.B(n_1239),
.Y(n_1522)
);

OAI22xp5_ASAP7_75t_L g1523 ( 
.A1(n_1437),
.A2(n_1172),
.B1(n_1282),
.B2(n_1260),
.Y(n_1523)
);

BUFx6f_ASAP7_75t_L g1524 ( 
.A(n_1435),
.Y(n_1524)
);

INVx1_ASAP7_75t_L g1525 ( 
.A(n_1342),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1334),
.Y(n_1526)
);

BUFx3_ASAP7_75t_L g1527 ( 
.A(n_1370),
.Y(n_1527)
);

INVx4_ASAP7_75t_L g1528 ( 
.A(n_1435),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1373),
.Y(n_1529)
);

BUFx12f_ASAP7_75t_L g1530 ( 
.A(n_1349),
.Y(n_1530)
);

NAND2x1_ASAP7_75t_L g1531 ( 
.A(n_1337),
.B(n_1310),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1359),
.Y(n_1532)
);

INVx1_ASAP7_75t_L g1533 ( 
.A(n_1375),
.Y(n_1533)
);

AOI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1502),
.A2(n_1160),
.B1(n_1234),
.B2(n_1314),
.Y(n_1534)
);

AND2x4_ASAP7_75t_L g1535 ( 
.A(n_1350),
.B(n_1308),
.Y(n_1535)
);

AOI22xp33_ASAP7_75t_L g1536 ( 
.A1(n_1477),
.A2(n_1300),
.B1(n_1311),
.B2(n_1235),
.Y(n_1536)
);

AOI22xp33_ASAP7_75t_L g1537 ( 
.A1(n_1477),
.A2(n_1234),
.B1(n_1308),
.B2(n_1259),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1380),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1371),
.B(n_1239),
.Y(n_1539)
);

BUFx6f_ASAP7_75t_L g1540 ( 
.A(n_1440),
.Y(n_1540)
);

OAI22xp33_ASAP7_75t_L g1541 ( 
.A1(n_1477),
.A2(n_1308),
.B1(n_1259),
.B2(n_1195),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1390),
.Y(n_1542)
);

INVx3_ASAP7_75t_L g1543 ( 
.A(n_1440),
.Y(n_1543)
);

AOI22xp33_ASAP7_75t_L g1544 ( 
.A1(n_1477),
.A2(n_1308),
.B1(n_1259),
.B2(n_1197),
.Y(n_1544)
);

OR2x2_ASAP7_75t_L g1545 ( 
.A(n_1402),
.B(n_1239),
.Y(n_1545)
);

OR2x6_ASAP7_75t_L g1546 ( 
.A(n_1397),
.B(n_1409),
.Y(n_1546)
);

AOI22xp33_ASAP7_75t_L g1547 ( 
.A1(n_1348),
.A2(n_1259),
.B1(n_1197),
.B2(n_1193),
.Y(n_1547)
);

OR2x2_ASAP7_75t_L g1548 ( 
.A(n_1427),
.B(n_1239),
.Y(n_1548)
);

A2O1A1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1488),
.A2(n_1287),
.B(n_1207),
.C(n_1268),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1413),
.A2(n_1193),
.B1(n_1287),
.B2(n_1205),
.Y(n_1550)
);

AOI22xp33_ASAP7_75t_L g1551 ( 
.A1(n_1488),
.A2(n_1288),
.B1(n_1254),
.B2(n_1252),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1371),
.B(n_1216),
.Y(n_1552)
);

OAI21xp5_ASAP7_75t_L g1553 ( 
.A1(n_1431),
.A2(n_1217),
.B(n_1212),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1493),
.B(n_1216),
.Y(n_1554)
);

BUFx4f_ASAP7_75t_L g1555 ( 
.A(n_1444),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_1349),
.Y(n_1556)
);

AOI22xp33_ASAP7_75t_SL g1557 ( 
.A1(n_1424),
.A2(n_1232),
.B1(n_63),
.B2(n_64),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1401),
.Y(n_1558)
);

CKINVDCx14_ASAP7_75t_R g1559 ( 
.A(n_1497),
.Y(n_1559)
);

AND2x2_ASAP7_75t_L g1560 ( 
.A(n_1437),
.B(n_1216),
.Y(n_1560)
);

OAI22xp5_ASAP7_75t_L g1561 ( 
.A1(n_1366),
.A2(n_1290),
.B1(n_1289),
.B2(n_1306),
.Y(n_1561)
);

AND2x2_ASAP7_75t_SL g1562 ( 
.A(n_1471),
.B(n_1216),
.Y(n_1562)
);

INVx6_ASAP7_75t_L g1563 ( 
.A(n_1399),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1498),
.B(n_1211),
.Y(n_1564)
);

AOI22xp33_ASAP7_75t_L g1565 ( 
.A1(n_1423),
.A2(n_62),
.B1(n_68),
.B2(n_71),
.Y(n_1565)
);

NAND3x1_ASAP7_75t_L g1566 ( 
.A(n_1379),
.B(n_68),
.C(n_71),
.Y(n_1566)
);

CKINVDCx8_ASAP7_75t_R g1567 ( 
.A(n_1466),
.Y(n_1567)
);

OAI22xp5_ASAP7_75t_L g1568 ( 
.A1(n_1434),
.A2(n_1211),
.B1(n_75),
.B2(n_80),
.Y(n_1568)
);

OAI21x1_ASAP7_75t_L g1569 ( 
.A1(n_1464),
.A2(n_1211),
.B(n_82),
.Y(n_1569)
);

INVx1_ASAP7_75t_L g1570 ( 
.A(n_1404),
.Y(n_1570)
);

AND2x2_ASAP7_75t_L g1571 ( 
.A(n_1495),
.B(n_1211),
.Y(n_1571)
);

OR2x6_ASAP7_75t_L g1572 ( 
.A(n_1397),
.B(n_74),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1343),
.Y(n_1573)
);

AOI211xp5_ASAP7_75t_L g1574 ( 
.A1(n_1406),
.A2(n_82),
.B(n_84),
.C(n_86),
.Y(n_1574)
);

CKINVDCx8_ASAP7_75t_R g1575 ( 
.A(n_1466),
.Y(n_1575)
);

NAND3xp33_ASAP7_75t_SL g1576 ( 
.A(n_1414),
.B(n_84),
.C(n_86),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1412),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1365),
.Y(n_1578)
);

OAI22xp5_ASAP7_75t_L g1579 ( 
.A1(n_1400),
.A2(n_87),
.B1(n_88),
.B2(n_89),
.Y(n_1579)
);

OR2x2_ASAP7_75t_L g1580 ( 
.A(n_1411),
.B(n_87),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1365),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1403),
.Y(n_1582)
);

OAI22xp5_ASAP7_75t_L g1583 ( 
.A1(n_1368),
.A2(n_88),
.B1(n_90),
.B2(n_91),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1403),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1376),
.Y(n_1585)
);

OR2x2_ASAP7_75t_L g1586 ( 
.A(n_1411),
.B(n_95),
.Y(n_1586)
);

OAI21x1_ASAP7_75t_L g1587 ( 
.A1(n_1464),
.A2(n_1472),
.B(n_1449),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1441),
.B(n_1396),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1408),
.Y(n_1589)
);

AOI221xp5_ASAP7_75t_L g1590 ( 
.A1(n_1453),
.A2(n_90),
.B1(n_94),
.B2(n_1351),
.C(n_1389),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1408),
.Y(n_1591)
);

OAI22xp33_ASAP7_75t_L g1592 ( 
.A1(n_1377),
.A2(n_94),
.B1(n_1444),
.B2(n_1450),
.Y(n_1592)
);

OAI22xp5_ASAP7_75t_L g1593 ( 
.A1(n_1377),
.A2(n_1426),
.B1(n_1419),
.B2(n_1456),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1441),
.B(n_1396),
.Y(n_1594)
);

BUFx3_ASAP7_75t_L g1595 ( 
.A(n_1370),
.Y(n_1595)
);

BUFx2_ASAP7_75t_L g1596 ( 
.A(n_1450),
.Y(n_1596)
);

AND2x4_ASAP7_75t_L g1597 ( 
.A(n_1350),
.B(n_1353),
.Y(n_1597)
);

AND2x2_ASAP7_75t_L g1598 ( 
.A(n_1396),
.B(n_1350),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1491),
.B(n_1483),
.Y(n_1599)
);

NOR2xp67_ASAP7_75t_R g1600 ( 
.A(n_1337),
.B(n_1452),
.Y(n_1600)
);

CKINVDCx11_ASAP7_75t_R g1601 ( 
.A(n_1497),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1353),
.B(n_1386),
.Y(n_1602)
);

OAI22xp5_ASAP7_75t_L g1603 ( 
.A1(n_1416),
.A2(n_1367),
.B1(n_1439),
.B2(n_1354),
.Y(n_1603)
);

AOI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1422),
.A2(n_1353),
.B1(n_1363),
.B2(n_1386),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1340),
.A2(n_1484),
.B1(n_1352),
.B2(n_1328),
.C(n_1483),
.Y(n_1605)
);

INVx4_ASAP7_75t_L g1606 ( 
.A(n_1440),
.Y(n_1606)
);

OAI22xp33_ASAP7_75t_L g1607 ( 
.A1(n_1445),
.A2(n_1409),
.B1(n_1397),
.B2(n_1439),
.Y(n_1607)
);

OAI222xp33_ASAP7_75t_L g1608 ( 
.A1(n_1439),
.A2(n_1445),
.B1(n_1409),
.B2(n_1397),
.C1(n_1383),
.C2(n_1483),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1386),
.B(n_1391),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1457),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1372),
.Y(n_1611)
);

OAI21x1_ASAP7_75t_L g1612 ( 
.A1(n_1449),
.A2(n_1405),
.B(n_1447),
.Y(n_1612)
);

INVx2_ASAP7_75t_L g1613 ( 
.A(n_1372),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1476),
.Y(n_1614)
);

OA21x2_ASAP7_75t_L g1615 ( 
.A1(n_1478),
.A2(n_1481),
.B(n_1447),
.Y(n_1615)
);

AND2x4_ASAP7_75t_L g1616 ( 
.A(n_1336),
.B(n_1409),
.Y(n_1616)
);

INVx1_ASAP7_75t_L g1617 ( 
.A(n_1420),
.Y(n_1617)
);

AOI221xp5_ASAP7_75t_L g1618 ( 
.A1(n_1340),
.A2(n_1484),
.B1(n_1352),
.B2(n_1328),
.C(n_1421),
.Y(n_1618)
);

NAND2xp33_ASAP7_75t_R g1619 ( 
.A(n_1471),
.B(n_1324),
.Y(n_1619)
);

OAI22xp33_ASAP7_75t_L g1620 ( 
.A1(n_1337),
.A2(n_1324),
.B1(n_1452),
.B2(n_1433),
.Y(n_1620)
);

OR2x6_ASAP7_75t_L g1621 ( 
.A(n_1331),
.B(n_1324),
.Y(n_1621)
);

AOI22xp33_ASAP7_75t_L g1622 ( 
.A1(n_1484),
.A2(n_1333),
.B1(n_1363),
.B2(n_1344),
.Y(n_1622)
);

O2A1O1Ixp33_ASAP7_75t_SL g1623 ( 
.A1(n_1425),
.A2(n_1436),
.B(n_1462),
.C(n_1465),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1454),
.A2(n_1471),
.B1(n_1336),
.B2(n_1407),
.Y(n_1624)
);

AND2x2_ASAP7_75t_L g1625 ( 
.A(n_1363),
.B(n_1399),
.Y(n_1625)
);

A2O1A1Ixp33_ASAP7_75t_L g1626 ( 
.A1(n_1338),
.A2(n_1474),
.B(n_1494),
.C(n_1489),
.Y(n_1626)
);

NAND3xp33_ASAP7_75t_L g1627 ( 
.A(n_1469),
.B(n_1446),
.C(n_1336),
.Y(n_1627)
);

AND2x4_ASAP7_75t_L g1628 ( 
.A(n_1490),
.B(n_1432),
.Y(n_1628)
);

HB1xp67_ASAP7_75t_L g1629 ( 
.A(n_1347),
.Y(n_1629)
);

NAND2xp33_ASAP7_75t_SL g1630 ( 
.A(n_1433),
.B(n_1459),
.Y(n_1630)
);

NAND2x1_ASAP7_75t_L g1631 ( 
.A(n_1357),
.B(n_1451),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1407),
.A2(n_1442),
.B1(n_1331),
.B2(n_1487),
.Y(n_1632)
);

OAI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1407),
.A2(n_1331),
.B1(n_1487),
.B2(n_1382),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1333),
.A2(n_1344),
.B1(n_1399),
.B2(n_1501),
.Y(n_1634)
);

CKINVDCx5p33_ASAP7_75t_R g1635 ( 
.A(n_1459),
.Y(n_1635)
);

NAND3xp33_ASAP7_75t_SL g1636 ( 
.A(n_1422),
.B(n_1490),
.C(n_1459),
.Y(n_1636)
);

INVx2_ASAP7_75t_L g1637 ( 
.A(n_1378),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1496),
.Y(n_1638)
);

A2O1A1Ixp33_ASAP7_75t_L g1639 ( 
.A1(n_1474),
.A2(n_1494),
.B(n_1489),
.C(n_1500),
.Y(n_1639)
);

AND2x2_ASAP7_75t_L g1640 ( 
.A(n_1432),
.B(n_1486),
.Y(n_1640)
);

BUFx12f_ASAP7_75t_L g1641 ( 
.A(n_1410),
.Y(n_1641)
);

AOI22xp5_ASAP7_75t_L g1642 ( 
.A1(n_1344),
.A2(n_1333),
.B1(n_1355),
.B2(n_1356),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1496),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1463),
.Y(n_1644)
);

OAI22xp33_ASAP7_75t_L g1645 ( 
.A1(n_1460),
.A2(n_1501),
.B1(n_1461),
.B2(n_1482),
.Y(n_1645)
);

BUFx3_ASAP7_75t_L g1646 ( 
.A(n_1463),
.Y(n_1646)
);

AOI22xp33_ASAP7_75t_L g1647 ( 
.A1(n_1460),
.A2(n_1461),
.B1(n_1482),
.B2(n_1347),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1496),
.Y(n_1648)
);

CKINVDCx11_ASAP7_75t_R g1649 ( 
.A(n_1410),
.Y(n_1649)
);

AND2x4_ASAP7_75t_L g1650 ( 
.A(n_1432),
.B(n_1479),
.Y(n_1650)
);

INVx2_ASAP7_75t_L g1651 ( 
.A(n_1378),
.Y(n_1651)
);

AOI22xp33_ASAP7_75t_SL g1652 ( 
.A1(n_1398),
.A2(n_1455),
.B1(n_1500),
.B2(n_1355),
.Y(n_1652)
);

AND2x4_ASAP7_75t_L g1653 ( 
.A(n_1465),
.B(n_1479),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1496),
.Y(n_1654)
);

AOI22xp33_ASAP7_75t_L g1655 ( 
.A1(n_1347),
.A2(n_1355),
.B1(n_1356),
.B2(n_1398),
.Y(n_1655)
);

BUFx12f_ASAP7_75t_L g1656 ( 
.A(n_1410),
.Y(n_1656)
);

NAND3xp33_ASAP7_75t_L g1657 ( 
.A(n_1430),
.B(n_1499),
.C(n_1429),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1361),
.Y(n_1658)
);

OAI22xp5_ASAP7_75t_L g1659 ( 
.A1(n_1463),
.A2(n_1486),
.B1(n_1430),
.B2(n_1387),
.Y(n_1659)
);

OAI22xp5_ASAP7_75t_L g1660 ( 
.A1(n_1463),
.A2(n_1430),
.B1(n_1387),
.B2(n_1475),
.Y(n_1660)
);

OAI22xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1410),
.A2(n_1429),
.B1(n_1480),
.B2(n_1475),
.Y(n_1661)
);

NAND2xp33_ASAP7_75t_L g1662 ( 
.A(n_1410),
.B(n_1429),
.Y(n_1662)
);

BUFx2_ASAP7_75t_L g1663 ( 
.A(n_1429),
.Y(n_1663)
);

INVx6_ASAP7_75t_L g1664 ( 
.A(n_1429),
.Y(n_1664)
);

HB1xp67_ASAP7_75t_L g1665 ( 
.A(n_1361),
.Y(n_1665)
);

OAI22xp5_ASAP7_75t_L g1666 ( 
.A1(n_1387),
.A2(n_1480),
.B1(n_1475),
.B2(n_1374),
.Y(n_1666)
);

AOI221xp5_ASAP7_75t_L g1667 ( 
.A1(n_1356),
.A2(n_1438),
.B1(n_1448),
.B2(n_1428),
.C(n_1417),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1496),
.B(n_1480),
.Y(n_1668)
);

NAND2xp5_ASAP7_75t_L g1669 ( 
.A(n_1475),
.B(n_1480),
.Y(n_1669)
);

AOI22xp33_ASAP7_75t_L g1670 ( 
.A1(n_1428),
.A2(n_1438),
.B1(n_1448),
.B2(n_1458),
.Y(n_1670)
);

INVx8_ASAP7_75t_L g1671 ( 
.A(n_1475),
.Y(n_1671)
);

INVx3_ASAP7_75t_L g1672 ( 
.A(n_1480),
.Y(n_1672)
);

AOI21xp33_ASAP7_75t_L g1673 ( 
.A1(n_1458),
.A2(n_1325),
.B(n_1451),
.Y(n_1673)
);

INVx6_ASAP7_75t_L g1674 ( 
.A(n_1357),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1361),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1361),
.B(n_1473),
.Y(n_1676)
);

CKINVDCx5p33_ASAP7_75t_R g1677 ( 
.A(n_1360),
.Y(n_1677)
);

BUFx2_ASAP7_75t_L g1678 ( 
.A(n_1458),
.Y(n_1678)
);

AOI22xp33_ASAP7_75t_SL g1679 ( 
.A1(n_1473),
.A2(n_1394),
.B1(n_1499),
.B2(n_1395),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1443),
.A2(n_1392),
.B(n_1395),
.Y(n_1680)
);

AOI22xp33_ASAP7_75t_L g1681 ( 
.A1(n_1417),
.A2(n_1381),
.B1(n_1499),
.B2(n_1385),
.Y(n_1681)
);

NOR2xp33_ASAP7_75t_L g1682 ( 
.A(n_1374),
.B(n_1381),
.Y(n_1682)
);

OR2x2_ASAP7_75t_L g1683 ( 
.A(n_1361),
.B(n_1385),
.Y(n_1683)
);

BUFx2_ASAP7_75t_L g1684 ( 
.A(n_1360),
.Y(n_1684)
);

A2O1A1Ixp33_ASAP7_75t_L g1685 ( 
.A1(n_1574),
.A2(n_1392),
.B(n_1394),
.C(n_1415),
.Y(n_1685)
);

INVx3_ASAP7_75t_L g1686 ( 
.A(n_1674),
.Y(n_1686)
);

AOI21xp5_ASAP7_75t_L g1687 ( 
.A1(n_1508),
.A2(n_1443),
.B(n_1415),
.Y(n_1687)
);

AND2x6_ASAP7_75t_SL g1688 ( 
.A(n_1516),
.B(n_1369),
.Y(n_1688)
);

AOI321xp33_ASAP7_75t_L g1689 ( 
.A1(n_1565),
.A2(n_1360),
.A3(n_1369),
.B1(n_1388),
.B2(n_1325),
.C(n_1362),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1611),
.Y(n_1690)
);

AO21x2_ASAP7_75t_L g1691 ( 
.A1(n_1626),
.A2(n_1388),
.B(n_1405),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1545),
.B(n_1381),
.Y(n_1692)
);

AND2x4_ASAP7_75t_L g1693 ( 
.A(n_1546),
.B(n_1362),
.Y(n_1693)
);

OAI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1565),
.A2(n_1326),
.B1(n_1346),
.B2(n_1505),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1516),
.A2(n_1326),
.B1(n_1346),
.B2(n_1505),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1613),
.Y(n_1696)
);

OAI22xp33_ASAP7_75t_L g1697 ( 
.A1(n_1592),
.A2(n_1572),
.B1(n_1517),
.B2(n_1604),
.Y(n_1697)
);

AOI222xp33_ASAP7_75t_L g1698 ( 
.A1(n_1590),
.A2(n_1576),
.B1(n_1579),
.B2(n_1583),
.C1(n_1514),
.C2(n_1592),
.Y(n_1698)
);

OAI221xp5_ASAP7_75t_L g1699 ( 
.A1(n_1513),
.A2(n_1557),
.B1(n_1536),
.B2(n_1515),
.C(n_1572),
.Y(n_1699)
);

OAI22xp33_ASAP7_75t_L g1700 ( 
.A1(n_1572),
.A2(n_1586),
.B1(n_1580),
.B2(n_1511),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1568),
.A2(n_1630),
.B1(n_1559),
.B2(n_1522),
.Y(n_1701)
);

AOI22xp33_ASAP7_75t_L g1702 ( 
.A1(n_1559),
.A2(n_1599),
.B1(n_1601),
.B2(n_1636),
.Y(n_1702)
);

AOI22xp33_ASAP7_75t_L g1703 ( 
.A1(n_1601),
.A2(n_1593),
.B1(n_1539),
.B2(n_1560),
.Y(n_1703)
);

OAI211xp5_ASAP7_75t_L g1704 ( 
.A1(n_1508),
.A2(n_1622),
.B(n_1536),
.C(n_1605),
.Y(n_1704)
);

AOI22xp33_ASAP7_75t_L g1705 ( 
.A1(n_1506),
.A2(n_1538),
.B1(n_1558),
.B2(n_1529),
.Y(n_1705)
);

OAI22xp33_ASAP7_75t_L g1706 ( 
.A1(n_1546),
.A2(n_1555),
.B1(n_1619),
.B2(n_1573),
.Y(n_1706)
);

HB1xp67_ASAP7_75t_L g1707 ( 
.A(n_1609),
.Y(n_1707)
);

OAI22xp5_ASAP7_75t_L g1708 ( 
.A1(n_1537),
.A2(n_1555),
.B1(n_1566),
.B2(n_1596),
.Y(n_1708)
);

NAND3xp33_ASAP7_75t_L g1709 ( 
.A(n_1622),
.B(n_1603),
.C(n_1618),
.Y(n_1709)
);

OAI221xp5_ASAP7_75t_L g1710 ( 
.A1(n_1534),
.A2(n_1549),
.B1(n_1537),
.B2(n_1523),
.C(n_1551),
.Y(n_1710)
);

OAI22xp5_ASAP7_75t_L g1711 ( 
.A1(n_1620),
.A2(n_1544),
.B1(n_1595),
.B2(n_1527),
.Y(n_1711)
);

AOI221xp5_ASAP7_75t_L g1712 ( 
.A1(n_1638),
.A2(n_1648),
.B1(n_1643),
.B2(n_1654),
.C(n_1518),
.Y(n_1712)
);

OAI211xp5_ASAP7_75t_L g1713 ( 
.A1(n_1554),
.A2(n_1564),
.B(n_1548),
.C(n_1642),
.Y(n_1713)
);

OAI22xp5_ASAP7_75t_L g1714 ( 
.A1(n_1620),
.A2(n_1544),
.B1(n_1595),
.B2(n_1527),
.Y(n_1714)
);

AOI22xp33_ASAP7_75t_SL g1715 ( 
.A1(n_1624),
.A2(n_1661),
.B1(n_1602),
.B2(n_1616),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1617),
.Y(n_1716)
);

AOI221xp5_ASAP7_75t_L g1717 ( 
.A1(n_1518),
.A2(n_1607),
.B1(n_1634),
.B2(n_1571),
.C(n_1525),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1546),
.B(n_1616),
.Y(n_1718)
);

AND2x2_ASAP7_75t_L g1719 ( 
.A(n_1594),
.B(n_1598),
.Y(n_1719)
);

AOI222xp33_ASAP7_75t_L g1720 ( 
.A1(n_1512),
.A2(n_1608),
.B1(n_1530),
.B2(n_1520),
.C1(n_1521),
.C2(n_1533),
.Y(n_1720)
);

OAI221xp5_ASAP7_75t_L g1721 ( 
.A1(n_1549),
.A2(n_1551),
.B1(n_1561),
.B2(n_1531),
.C(n_1634),
.Y(n_1721)
);

INVx2_ASAP7_75t_L g1722 ( 
.A(n_1637),
.Y(n_1722)
);

AOI21xp5_ASAP7_75t_L g1723 ( 
.A1(n_1541),
.A2(n_1662),
.B(n_1623),
.Y(n_1723)
);

AND2x4_ASAP7_75t_L g1724 ( 
.A(n_1597),
.B(n_1621),
.Y(n_1724)
);

INVx1_ASAP7_75t_L g1725 ( 
.A(n_1542),
.Y(n_1725)
);

OAI21xp5_ASAP7_75t_L g1726 ( 
.A1(n_1553),
.A2(n_1550),
.B(n_1569),
.Y(n_1726)
);

AND2x2_ASAP7_75t_L g1727 ( 
.A(n_1597),
.B(n_1552),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1570),
.Y(n_1728)
);

AND2x2_ASAP7_75t_L g1729 ( 
.A(n_1628),
.B(n_1625),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1628),
.B(n_1640),
.Y(n_1730)
);

AOI22xp33_ASAP7_75t_L g1731 ( 
.A1(n_1577),
.A2(n_1591),
.B1(n_1589),
.B2(n_1584),
.Y(n_1731)
);

AND2x4_ASAP7_75t_L g1732 ( 
.A(n_1621),
.B(n_1535),
.Y(n_1732)
);

INVx3_ASAP7_75t_L g1733 ( 
.A(n_1674),
.Y(n_1733)
);

INVx4_ASAP7_75t_L g1734 ( 
.A(n_1649),
.Y(n_1734)
);

CKINVDCx5p33_ASAP7_75t_R g1735 ( 
.A(n_1556),
.Y(n_1735)
);

AND2x2_ASAP7_75t_L g1736 ( 
.A(n_1535),
.B(n_1543),
.Y(n_1736)
);

BUFx2_ASAP7_75t_L g1737 ( 
.A(n_1646),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1610),
.Y(n_1738)
);

INVx1_ASAP7_75t_L g1739 ( 
.A(n_1614),
.Y(n_1739)
);

AOI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1582),
.A2(n_1503),
.B1(n_1510),
.B2(n_1607),
.Y(n_1740)
);

NAND2xp5_ASAP7_75t_L g1741 ( 
.A(n_1503),
.B(n_1510),
.Y(n_1741)
);

OAI22xp5_ASAP7_75t_L g1742 ( 
.A1(n_1567),
.A2(n_1575),
.B1(n_1543),
.B2(n_1606),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1650),
.B(n_1519),
.Y(n_1743)
);

AND2x2_ASAP7_75t_L g1744 ( 
.A(n_1650),
.B(n_1519),
.Y(n_1744)
);

OAI211xp5_ASAP7_75t_L g1745 ( 
.A1(n_1668),
.A2(n_1639),
.B(n_1655),
.C(n_1652),
.Y(n_1745)
);

AOI22xp33_ASAP7_75t_L g1746 ( 
.A1(n_1541),
.A2(n_1606),
.B1(n_1528),
.B2(n_1540),
.Y(n_1746)
);

INVx2_ASAP7_75t_SL g1747 ( 
.A(n_1635),
.Y(n_1747)
);

AND2x2_ASAP7_75t_L g1748 ( 
.A(n_1519),
.B(n_1524),
.Y(n_1748)
);

OAI211xp5_ASAP7_75t_SL g1749 ( 
.A1(n_1655),
.A2(n_1639),
.B(n_1673),
.C(n_1626),
.Y(n_1749)
);

AOI221xp5_ASAP7_75t_L g1750 ( 
.A1(n_1623),
.A2(n_1645),
.B1(n_1647),
.B2(n_1629),
.C(n_1665),
.Y(n_1750)
);

NOR2x1_ASAP7_75t_SL g1751 ( 
.A(n_1627),
.B(n_1621),
.Y(n_1751)
);

AND2x2_ASAP7_75t_L g1752 ( 
.A(n_1519),
.B(n_1524),
.Y(n_1752)
);

AOI22xp33_ASAP7_75t_L g1753 ( 
.A1(n_1528),
.A2(n_1540),
.B1(n_1524),
.B2(n_1507),
.Y(n_1753)
);

OAI22xp5_ASAP7_75t_L g1754 ( 
.A1(n_1563),
.A2(n_1677),
.B1(n_1550),
.B2(n_1547),
.Y(n_1754)
);

NAND2xp5_ASAP7_75t_L g1755 ( 
.A(n_1526),
.B(n_1581),
.Y(n_1755)
);

OAI221xp5_ASAP7_75t_L g1756 ( 
.A1(n_1547),
.A2(n_1632),
.B1(n_1633),
.B2(n_1679),
.C(n_1563),
.Y(n_1756)
);

OAI22xp5_ASAP7_75t_L g1757 ( 
.A1(n_1563),
.A2(n_1524),
.B1(n_1540),
.B2(n_1562),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1562),
.A2(n_1674),
.B1(n_1619),
.B2(n_1678),
.Y(n_1758)
);

OAI22xp33_ASAP7_75t_L g1759 ( 
.A1(n_1540),
.A2(n_1646),
.B1(n_1644),
.B2(n_1659),
.Y(n_1759)
);

NAND3xp33_ASAP7_75t_L g1760 ( 
.A(n_1647),
.B(n_1660),
.C(n_1629),
.Y(n_1760)
);

OAI22xp5_ASAP7_75t_L g1761 ( 
.A1(n_1670),
.A2(n_1669),
.B1(n_1664),
.B2(n_1653),
.Y(n_1761)
);

BUFx5_ASAP7_75t_L g1762 ( 
.A(n_1676),
.Y(n_1762)
);

OAI22xp5_ASAP7_75t_L g1763 ( 
.A1(n_1670),
.A2(n_1664),
.B1(n_1653),
.B2(n_1663),
.Y(n_1763)
);

A2O1A1Ixp33_ASAP7_75t_L g1764 ( 
.A1(n_1682),
.A2(n_1657),
.B(n_1665),
.C(n_1667),
.Y(n_1764)
);

CKINVDCx5p33_ASAP7_75t_R g1765 ( 
.A(n_1649),
.Y(n_1765)
);

OAI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1664),
.A2(n_1672),
.B1(n_1641),
.B2(n_1656),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1631),
.A2(n_1666),
.B1(n_1672),
.B2(n_1671),
.Y(n_1767)
);

AOI22xp33_ASAP7_75t_L g1768 ( 
.A1(n_1532),
.A2(n_1578),
.B1(n_1585),
.B2(n_1658),
.Y(n_1768)
);

AOI222xp33_ASAP7_75t_L g1769 ( 
.A1(n_1585),
.A2(n_1600),
.B1(n_1658),
.B2(n_1675),
.C1(n_1645),
.C2(n_1684),
.Y(n_1769)
);

OR2x2_ASAP7_75t_L g1770 ( 
.A(n_1675),
.B(n_1683),
.Y(n_1770)
);

AOI21xp33_ASAP7_75t_L g1771 ( 
.A1(n_1504),
.A2(n_1682),
.B(n_1615),
.Y(n_1771)
);

AND2x4_ASAP7_75t_L g1772 ( 
.A(n_1587),
.B(n_1612),
.Y(n_1772)
);

INVxp67_ASAP7_75t_L g1773 ( 
.A(n_1615),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_SL g1774 ( 
.A(n_1671),
.B(n_1680),
.Y(n_1774)
);

OA21x2_ASAP7_75t_L g1775 ( 
.A1(n_1681),
.A2(n_1651),
.B(n_1504),
.Y(n_1775)
);

NAND3xp33_ASAP7_75t_L g1776 ( 
.A(n_1504),
.B(n_1615),
.C(n_1681),
.Y(n_1776)
);

OAI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1671),
.A2(n_1565),
.B1(n_1330),
.B2(n_1095),
.Y(n_1777)
);

OAI22xp5_ASAP7_75t_SL g1778 ( 
.A1(n_1516),
.A2(n_1095),
.B1(n_986),
.B2(n_1065),
.Y(n_1778)
);

AOI22xp33_ASAP7_75t_L g1779 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1779)
);

BUFx2_ASAP7_75t_L g1780 ( 
.A(n_1527),
.Y(n_1780)
);

OAI211xp5_ASAP7_75t_L g1781 ( 
.A1(n_1574),
.A2(n_1565),
.B(n_986),
.C(n_836),
.Y(n_1781)
);

AO21x2_ASAP7_75t_L g1782 ( 
.A1(n_1626),
.A2(n_1673),
.B(n_1639),
.Y(n_1782)
);

OAI21xp33_ASAP7_75t_L g1783 ( 
.A1(n_1505),
.A2(n_1095),
.B(n_1065),
.Y(n_1783)
);

AND2x2_ASAP7_75t_L g1784 ( 
.A(n_1509),
.B(n_1588),
.Y(n_1784)
);

INVx1_ASAP7_75t_L g1785 ( 
.A(n_1617),
.Y(n_1785)
);

AND2x2_ASAP7_75t_L g1786 ( 
.A(n_1509),
.B(n_1588),
.Y(n_1786)
);

AOI22xp33_ASAP7_75t_L g1787 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1787)
);

HB1xp67_ASAP7_75t_L g1788 ( 
.A(n_1609),
.Y(n_1788)
);

AOI221xp5_ASAP7_75t_L g1789 ( 
.A1(n_1565),
.A2(n_654),
.B1(n_986),
.B2(n_836),
.C(n_1492),
.Y(n_1789)
);

OAI22xp5_ASAP7_75t_L g1790 ( 
.A1(n_1565),
.A2(n_1330),
.B1(n_1095),
.B2(n_1065),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1546),
.B(n_1616),
.Y(n_1791)
);

AOI22xp5_ASAP7_75t_L g1792 ( 
.A1(n_1516),
.A2(n_1095),
.B1(n_1065),
.B2(n_799),
.Y(n_1792)
);

NAND2xp5_ASAP7_75t_L g1793 ( 
.A(n_1509),
.B(n_1413),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1509),
.B(n_1413),
.Y(n_1794)
);

OR2x2_ASAP7_75t_L g1795 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1795)
);

OAI22xp33_ASAP7_75t_L g1796 ( 
.A1(n_1592),
.A2(n_986),
.B1(n_1058),
.B2(n_1065),
.Y(n_1796)
);

AOI22xp33_ASAP7_75t_SL g1797 ( 
.A1(n_1516),
.A2(n_1095),
.B1(n_1065),
.B2(n_986),
.Y(n_1797)
);

AOI22xp33_ASAP7_75t_L g1798 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1509),
.B(n_1327),
.Y(n_1799)
);

CKINVDCx6p67_ASAP7_75t_R g1800 ( 
.A(n_1530),
.Y(n_1800)
);

BUFx2_ASAP7_75t_L g1801 ( 
.A(n_1527),
.Y(n_1801)
);

OAI322xp33_ASAP7_75t_L g1802 ( 
.A1(n_1592),
.A2(n_654),
.A3(n_625),
.B1(n_387),
.B2(n_268),
.C1(n_1215),
.C2(n_517),
.Y(n_1802)
);

AOI22xp33_ASAP7_75t_L g1803 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1803)
);

NOR2x1_ASAP7_75t_SL g1804 ( 
.A(n_1546),
.B(n_1627),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1509),
.B(n_1413),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1617),
.Y(n_1806)
);

BUFx3_ASAP7_75t_L g1807 ( 
.A(n_1527),
.Y(n_1807)
);

AOI22xp33_ASAP7_75t_L g1808 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1808)
);

BUFx3_ASAP7_75t_L g1809 ( 
.A(n_1527),
.Y(n_1809)
);

AOI22xp33_ASAP7_75t_L g1810 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1810)
);

OAI211xp5_ASAP7_75t_L g1811 ( 
.A1(n_1574),
.A2(n_1565),
.B(n_986),
.C(n_836),
.Y(n_1811)
);

CKINVDCx20_ASAP7_75t_R g1812 ( 
.A(n_1601),
.Y(n_1812)
);

OAI22xp33_ASAP7_75t_L g1813 ( 
.A1(n_1592),
.A2(n_986),
.B1(n_1058),
.B2(n_1065),
.Y(n_1813)
);

AOI21xp5_ASAP7_75t_L g1814 ( 
.A1(n_1508),
.A2(n_1338),
.B(n_975),
.Y(n_1814)
);

OR2x2_ASAP7_75t_L g1815 ( 
.A(n_1545),
.B(n_1522),
.Y(n_1815)
);

INVx3_ASAP7_75t_L g1816 ( 
.A(n_1674),
.Y(n_1816)
);

OAI21x1_ASAP7_75t_L g1817 ( 
.A1(n_1680),
.A2(n_1612),
.B(n_1587),
.Y(n_1817)
);

OAI22xp33_ASAP7_75t_L g1818 ( 
.A1(n_1592),
.A2(n_986),
.B1(n_1058),
.B2(n_1065),
.Y(n_1818)
);

OAI22xp5_ASAP7_75t_L g1819 ( 
.A1(n_1565),
.A2(n_1330),
.B1(n_1095),
.B2(n_1065),
.Y(n_1819)
);

INVx3_ASAP7_75t_SL g1820 ( 
.A(n_1556),
.Y(n_1820)
);

AOI22xp33_ASAP7_75t_L g1821 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1574),
.A2(n_986),
.B1(n_799),
.B2(n_1095),
.C(n_1065),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_SL g1823 ( 
.A1(n_1516),
.A2(n_1095),
.B1(n_1065),
.B2(n_986),
.Y(n_1823)
);

AOI22xp33_ASAP7_75t_L g1824 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1824)
);

AOI22xp33_ASAP7_75t_L g1825 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1509),
.B(n_1413),
.Y(n_1826)
);

INVx2_ASAP7_75t_L g1827 ( 
.A(n_1611),
.Y(n_1827)
);

AOI22xp33_ASAP7_75t_SL g1828 ( 
.A1(n_1516),
.A2(n_1095),
.B1(n_1065),
.B2(n_986),
.Y(n_1828)
);

OAI22xp33_ASAP7_75t_L g1829 ( 
.A1(n_1592),
.A2(n_986),
.B1(n_1058),
.B2(n_1065),
.Y(n_1829)
);

INVx3_ASAP7_75t_L g1830 ( 
.A(n_1674),
.Y(n_1830)
);

OAI22xp5_ASAP7_75t_SL g1831 ( 
.A1(n_1516),
.A2(n_1095),
.B1(n_986),
.B2(n_1065),
.Y(n_1831)
);

AOI22xp33_ASAP7_75t_L g1832 ( 
.A1(n_1565),
.A2(n_986),
.B1(n_1590),
.B2(n_1492),
.Y(n_1832)
);

AND2x4_ASAP7_75t_L g1833 ( 
.A(n_1693),
.B(n_1772),
.Y(n_1833)
);

AND2x4_ASAP7_75t_L g1834 ( 
.A(n_1693),
.B(n_1772),
.Y(n_1834)
);

BUFx2_ASAP7_75t_L g1835 ( 
.A(n_1693),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1716),
.Y(n_1836)
);

NAND2xp5_ASAP7_75t_L g1837 ( 
.A(n_1741),
.B(n_1795),
.Y(n_1837)
);

HB1xp67_ASAP7_75t_L g1838 ( 
.A(n_1773),
.Y(n_1838)
);

AND2x2_ASAP7_75t_L g1839 ( 
.A(n_1762),
.B(n_1690),
.Y(n_1839)
);

INVx2_ASAP7_75t_L g1840 ( 
.A(n_1775),
.Y(n_1840)
);

AOI22xp5_ASAP7_75t_L g1841 ( 
.A1(n_1790),
.A2(n_1819),
.B1(n_1811),
.B2(n_1781),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1738),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1815),
.B(n_1739),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1785),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1806),
.Y(n_1845)
);

CKINVDCx20_ASAP7_75t_R g1846 ( 
.A(n_1812),
.Y(n_1846)
);

INVx2_ASAP7_75t_L g1847 ( 
.A(n_1775),
.Y(n_1847)
);

INVx2_ASAP7_75t_L g1848 ( 
.A(n_1775),
.Y(n_1848)
);

AO21x2_ASAP7_75t_L g1849 ( 
.A1(n_1726),
.A2(n_1771),
.B(n_1776),
.Y(n_1849)
);

INVx2_ASAP7_75t_L g1850 ( 
.A(n_1696),
.Y(n_1850)
);

NOR2xp67_ASAP7_75t_L g1851 ( 
.A(n_1713),
.B(n_1709),
.Y(n_1851)
);

AND2x4_ASAP7_75t_L g1852 ( 
.A(n_1772),
.B(n_1718),
.Y(n_1852)
);

INVx1_ASAP7_75t_L g1853 ( 
.A(n_1722),
.Y(n_1853)
);

BUFx2_ASAP7_75t_L g1854 ( 
.A(n_1770),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1725),
.B(n_1728),
.Y(n_1855)
);

AND4x1_ASAP7_75t_L g1856 ( 
.A(n_1792),
.B(n_1783),
.C(n_1789),
.D(n_1824),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1827),
.B(n_1764),
.Y(n_1857)
);

INVx3_ASAP7_75t_L g1858 ( 
.A(n_1817),
.Y(n_1858)
);

AOI22xp5_ASAP7_75t_L g1859 ( 
.A1(n_1822),
.A2(n_1778),
.B1(n_1831),
.B2(n_1832),
.Y(n_1859)
);

NOR2x1_ASAP7_75t_L g1860 ( 
.A(n_1686),
.B(n_1733),
.Y(n_1860)
);

AND2x2_ASAP7_75t_L g1861 ( 
.A(n_1764),
.B(n_1692),
.Y(n_1861)
);

OR2x2_ASAP7_75t_L g1862 ( 
.A(n_1760),
.B(n_1782),
.Y(n_1862)
);

AND2x2_ASAP7_75t_L g1863 ( 
.A(n_1782),
.B(n_1758),
.Y(n_1863)
);

OR2x2_ASAP7_75t_L g1864 ( 
.A(n_1745),
.B(n_1740),
.Y(n_1864)
);

OAI22xp5_ASAP7_75t_L g1865 ( 
.A1(n_1779),
.A2(n_1832),
.B1(n_1787),
.B2(n_1808),
.Y(n_1865)
);

AND2x4_ASAP7_75t_L g1866 ( 
.A(n_1718),
.B(n_1791),
.Y(n_1866)
);

BUFx2_ASAP7_75t_L g1867 ( 
.A(n_1691),
.Y(n_1867)
);

INVx2_ASAP7_75t_L g1868 ( 
.A(n_1817),
.Y(n_1868)
);

AND2x2_ASAP7_75t_L g1869 ( 
.A(n_1691),
.B(n_1750),
.Y(n_1869)
);

AND2x2_ASAP7_75t_L g1870 ( 
.A(n_1712),
.B(n_1740),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1717),
.B(n_1705),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1695),
.B(n_1768),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1768),
.B(n_1727),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1755),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1705),
.B(n_1799),
.Y(n_1875)
);

AND2x2_ASAP7_75t_L g1876 ( 
.A(n_1704),
.B(n_1720),
.Y(n_1876)
);

INVx4_ASAP7_75t_L g1877 ( 
.A(n_1686),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1686),
.Y(n_1878)
);

OR2x2_ASAP7_75t_L g1879 ( 
.A(n_1707),
.B(n_1788),
.Y(n_1879)
);

HB1xp67_ASAP7_75t_L g1880 ( 
.A(n_1763),
.Y(n_1880)
);

AND2x4_ASAP7_75t_L g1881 ( 
.A(n_1732),
.B(n_1724),
.Y(n_1881)
);

AND2x2_ASAP7_75t_L g1882 ( 
.A(n_1784),
.B(n_1786),
.Y(n_1882)
);

OR2x2_ASAP7_75t_L g1883 ( 
.A(n_1761),
.B(n_1721),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1731),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1731),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1774),
.Y(n_1886)
);

INVx1_ASAP7_75t_L g1887 ( 
.A(n_1723),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1689),
.Y(n_1888)
);

INVx1_ASAP7_75t_L g1889 ( 
.A(n_1749),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1754),
.B(n_1710),
.Y(n_1890)
);

BUFx2_ASAP7_75t_L g1891 ( 
.A(n_1688),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1816),
.Y(n_1892)
);

INVx1_ASAP7_75t_L g1893 ( 
.A(n_1816),
.Y(n_1893)
);

HB1xp67_ASAP7_75t_L g1894 ( 
.A(n_1756),
.Y(n_1894)
);

BUFx3_ASAP7_75t_L g1895 ( 
.A(n_1816),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1799),
.B(n_1730),
.Y(n_1896)
);

OR2x2_ASAP7_75t_L g1897 ( 
.A(n_1694),
.B(n_1711),
.Y(n_1897)
);

OR2x6_ASAP7_75t_L g1898 ( 
.A(n_1687),
.B(n_1814),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1769),
.B(n_1703),
.Y(n_1899)
);

AND2x2_ASAP7_75t_L g1900 ( 
.A(n_1703),
.B(n_1685),
.Y(n_1900)
);

AND2x2_ASAP7_75t_L g1901 ( 
.A(n_1685),
.B(n_1729),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1804),
.B(n_1751),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1830),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1767),
.Y(n_1904)
);

INVx1_ASAP7_75t_L g1905 ( 
.A(n_1757),
.Y(n_1905)
);

OAI211xp5_ASAP7_75t_L g1906 ( 
.A1(n_1779),
.A2(n_1787),
.B(n_1808),
.C(n_1810),
.Y(n_1906)
);

INVx1_ASAP7_75t_L g1907 ( 
.A(n_1759),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_R g1908 ( 
.A(n_1846),
.B(n_1812),
.Y(n_1908)
);

INVx1_ASAP7_75t_L g1909 ( 
.A(n_1836),
.Y(n_1909)
);

HB1xp67_ASAP7_75t_L g1910 ( 
.A(n_1854),
.Y(n_1910)
);

INVx1_ASAP7_75t_L g1911 ( 
.A(n_1836),
.Y(n_1911)
);

BUFx3_ASAP7_75t_L g1912 ( 
.A(n_1895),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1840),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1865),
.A2(n_1798),
.B1(n_1803),
.B2(n_1810),
.Y(n_1914)
);

NAND2xp5_ASAP7_75t_L g1915 ( 
.A(n_1837),
.B(n_1794),
.Y(n_1915)
);

OAI211xp5_ASAP7_75t_L g1916 ( 
.A1(n_1859),
.A2(n_1797),
.B(n_1823),
.C(n_1828),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1842),
.Y(n_1917)
);

AOI22xp33_ASAP7_75t_L g1918 ( 
.A1(n_1865),
.A2(n_1821),
.B1(n_1803),
.B2(n_1798),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1842),
.Y(n_1919)
);

CKINVDCx5p33_ASAP7_75t_R g1920 ( 
.A(n_1846),
.Y(n_1920)
);

AND2x2_ASAP7_75t_L g1921 ( 
.A(n_1835),
.B(n_1715),
.Y(n_1921)
);

HB1xp67_ASAP7_75t_L g1922 ( 
.A(n_1854),
.Y(n_1922)
);

INVx1_ASAP7_75t_L g1923 ( 
.A(n_1844),
.Y(n_1923)
);

AOI22xp33_ASAP7_75t_L g1924 ( 
.A1(n_1859),
.A2(n_1824),
.B1(n_1825),
.B2(n_1821),
.Y(n_1924)
);

AOI21x1_ASAP7_75t_L g1925 ( 
.A1(n_1851),
.A2(n_1742),
.B(n_1766),
.Y(n_1925)
);

NAND3xp33_ASAP7_75t_L g1926 ( 
.A(n_1856),
.B(n_1825),
.C(n_1698),
.Y(n_1926)
);

AOI22xp33_ASAP7_75t_L g1927 ( 
.A1(n_1894),
.A2(n_1802),
.B1(n_1699),
.B2(n_1777),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1844),
.Y(n_1928)
);

OAI221xp5_ASAP7_75t_L g1929 ( 
.A1(n_1856),
.A2(n_1702),
.B1(n_1701),
.B2(n_1826),
.C(n_1793),
.Y(n_1929)
);

BUFx10_ASAP7_75t_L g1930 ( 
.A(n_1886),
.Y(n_1930)
);

OR2x2_ASAP7_75t_L g1931 ( 
.A(n_1854),
.B(n_1805),
.Y(n_1931)
);

OR2x2_ASAP7_75t_L g1932 ( 
.A(n_1837),
.B(n_1801),
.Y(n_1932)
);

OAI21x1_ASAP7_75t_L g1933 ( 
.A1(n_1858),
.A2(n_1714),
.B(n_1746),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1875),
.B(n_1879),
.Y(n_1934)
);

AOI22xp33_ASAP7_75t_L g1935 ( 
.A1(n_1894),
.A2(n_1697),
.B1(n_1829),
.B2(n_1796),
.Y(n_1935)
);

AOI22xp33_ASAP7_75t_L g1936 ( 
.A1(n_1876),
.A2(n_1841),
.B1(n_1851),
.B2(n_1899),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1845),
.Y(n_1937)
);

BUFx2_ASAP7_75t_L g1938 ( 
.A(n_1833),
.Y(n_1938)
);

INVx2_ASAP7_75t_L g1939 ( 
.A(n_1840),
.Y(n_1939)
);

OAI31xp33_ASAP7_75t_L g1940 ( 
.A1(n_1906),
.A2(n_1813),
.A3(n_1818),
.B(n_1700),
.Y(n_1940)
);

HB1xp67_ASAP7_75t_L g1941 ( 
.A(n_1879),
.Y(n_1941)
);

OAI211xp5_ASAP7_75t_L g1942 ( 
.A1(n_1841),
.A2(n_1701),
.B(n_1702),
.C(n_1734),
.Y(n_1942)
);

AO21x2_ASAP7_75t_L g1943 ( 
.A1(n_1868),
.A2(n_1706),
.B(n_1708),
.Y(n_1943)
);

NAND3xp33_ASAP7_75t_L g1944 ( 
.A(n_1889),
.B(n_1753),
.C(n_1746),
.Y(n_1944)
);

INVx2_ASAP7_75t_L g1945 ( 
.A(n_1847),
.Y(n_1945)
);

AOI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1889),
.A2(n_1719),
.B1(n_1780),
.B2(n_1737),
.C(n_1736),
.Y(n_1946)
);

AOI221xp5_ASAP7_75t_L g1947 ( 
.A1(n_1888),
.A2(n_1807),
.B1(n_1809),
.B2(n_1734),
.C(n_1753),
.Y(n_1947)
);

OAI22xp5_ASAP7_75t_L g1948 ( 
.A1(n_1906),
.A2(n_1765),
.B1(n_1734),
.B2(n_1807),
.Y(n_1948)
);

OAI221xp5_ASAP7_75t_L g1949 ( 
.A1(n_1891),
.A2(n_1747),
.B1(n_1820),
.B2(n_1809),
.C(n_1765),
.Y(n_1949)
);

AOI22xp33_ASAP7_75t_L g1950 ( 
.A1(n_1876),
.A2(n_1800),
.B1(n_1743),
.B2(n_1744),
.Y(n_1950)
);

NOR2x1_ASAP7_75t_L g1951 ( 
.A(n_1891),
.B(n_1748),
.Y(n_1951)
);

NOR2xp33_ASAP7_75t_L g1952 ( 
.A(n_1896),
.B(n_1820),
.Y(n_1952)
);

NOR2xp33_ASAP7_75t_SL g1953 ( 
.A(n_1877),
.B(n_1735),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1876),
.A2(n_1735),
.B1(n_1752),
.B2(n_1899),
.Y(n_1954)
);

INVx2_ASAP7_75t_L g1955 ( 
.A(n_1847),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_L g1956 ( 
.A(n_1875),
.B(n_1879),
.Y(n_1956)
);

INVx2_ASAP7_75t_L g1957 ( 
.A(n_1847),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1848),
.Y(n_1958)
);

AO22x1_ASAP7_75t_L g1959 ( 
.A1(n_1891),
.A2(n_1899),
.B1(n_1902),
.B2(n_1870),
.Y(n_1959)
);

INVx2_ASAP7_75t_L g1960 ( 
.A(n_1848),
.Y(n_1960)
);

INVx2_ASAP7_75t_L g1961 ( 
.A(n_1848),
.Y(n_1961)
);

NAND3xp33_ASAP7_75t_L g1962 ( 
.A(n_1862),
.B(n_1888),
.C(n_1890),
.Y(n_1962)
);

INVx1_ASAP7_75t_SL g1963 ( 
.A(n_1882),
.Y(n_1963)
);

AOI21xp5_ASAP7_75t_L g1964 ( 
.A1(n_1898),
.A2(n_1871),
.B(n_1890),
.Y(n_1964)
);

AND2x2_ASAP7_75t_L g1965 ( 
.A(n_1835),
.B(n_1839),
.Y(n_1965)
);

BUFx2_ASAP7_75t_L g1966 ( 
.A(n_1833),
.Y(n_1966)
);

NOR2xp67_ASAP7_75t_L g1967 ( 
.A(n_1838),
.B(n_1833),
.Y(n_1967)
);

AND2x2_ASAP7_75t_L g1968 ( 
.A(n_1835),
.B(n_1839),
.Y(n_1968)
);

INVx1_ASAP7_75t_L g1969 ( 
.A(n_1838),
.Y(n_1969)
);

INVx2_ASAP7_75t_L g1970 ( 
.A(n_1850),
.Y(n_1970)
);

INVx5_ASAP7_75t_SL g1971 ( 
.A(n_1898),
.Y(n_1971)
);

AOI221xp5_ASAP7_75t_L g1972 ( 
.A1(n_1900),
.A2(n_1871),
.B1(n_1869),
.B2(n_1870),
.C(n_1907),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1853),
.Y(n_1973)
);

AOI22xp33_ASAP7_75t_L g1974 ( 
.A1(n_1900),
.A2(n_1890),
.B1(n_1897),
.B2(n_1864),
.Y(n_1974)
);

INVx1_ASAP7_75t_L g1975 ( 
.A(n_1853),
.Y(n_1975)
);

AOI22xp33_ASAP7_75t_L g1976 ( 
.A1(n_1900),
.A2(n_1897),
.B1(n_1864),
.B2(n_1883),
.Y(n_1976)
);

AOI221xp5_ASAP7_75t_L g1977 ( 
.A1(n_1869),
.A2(n_1870),
.B1(n_1907),
.B2(n_1885),
.C(n_1884),
.Y(n_1977)
);

NOR4xp25_ASAP7_75t_SL g1978 ( 
.A(n_1887),
.B(n_1886),
.C(n_1904),
.D(n_1867),
.Y(n_1978)
);

NOR2x1_ASAP7_75t_L g1979 ( 
.A(n_1887),
.B(n_1860),
.Y(n_1979)
);

INVx1_ASAP7_75t_L g1980 ( 
.A(n_1909),
.Y(n_1980)
);

OR2x2_ASAP7_75t_L g1981 ( 
.A(n_1910),
.B(n_1862),
.Y(n_1981)
);

INVxp67_ASAP7_75t_L g1982 ( 
.A(n_1962),
.Y(n_1982)
);

INVx1_ASAP7_75t_L g1983 ( 
.A(n_1909),
.Y(n_1983)
);

AND3x1_ASAP7_75t_L g1984 ( 
.A(n_1936),
.B(n_1902),
.C(n_1863),
.Y(n_1984)
);

INVx1_ASAP7_75t_L g1985 ( 
.A(n_1911),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_L g1986 ( 
.A(n_1949),
.B(n_1896),
.Y(n_1986)
);

AND2x2_ASAP7_75t_L g1987 ( 
.A(n_1965),
.B(n_1863),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1934),
.B(n_1861),
.Y(n_1988)
);

INVx1_ASAP7_75t_L g1989 ( 
.A(n_1911),
.Y(n_1989)
);

AND2x2_ASAP7_75t_L g1990 ( 
.A(n_1938),
.B(n_1833),
.Y(n_1990)
);

OR2x2_ASAP7_75t_L g1991 ( 
.A(n_1922),
.B(n_1862),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_L g1992 ( 
.A(n_1956),
.B(n_1861),
.Y(n_1992)
);

NOR2x1_ASAP7_75t_L g1993 ( 
.A(n_1951),
.B(n_1860),
.Y(n_1993)
);

INVx3_ASAP7_75t_L g1994 ( 
.A(n_1913),
.Y(n_1994)
);

INVx1_ASAP7_75t_L g1995 ( 
.A(n_1917),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1965),
.B(n_1863),
.Y(n_1996)
);

OR2x2_ASAP7_75t_L g1997 ( 
.A(n_1941),
.B(n_1931),
.Y(n_1997)
);

AND2x2_ASAP7_75t_L g1998 ( 
.A(n_1968),
.B(n_1869),
.Y(n_1998)
);

AND2x2_ASAP7_75t_L g1999 ( 
.A(n_1938),
.B(n_1833),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1969),
.B(n_1861),
.Y(n_2000)
);

INVx1_ASAP7_75t_L g2001 ( 
.A(n_1917),
.Y(n_2001)
);

INVx2_ASAP7_75t_SL g2002 ( 
.A(n_1913),
.Y(n_2002)
);

OR2x2_ASAP7_75t_L g2003 ( 
.A(n_1931),
.B(n_1843),
.Y(n_2003)
);

INVx1_ASAP7_75t_L g2004 ( 
.A(n_1919),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1966),
.B(n_1834),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1969),
.B(n_1843),
.Y(n_2006)
);

INVx1_ASAP7_75t_SL g2007 ( 
.A(n_1951),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1919),
.Y(n_2008)
);

AND2x2_ASAP7_75t_L g2009 ( 
.A(n_1968),
.B(n_1834),
.Y(n_2009)
);

INVx2_ASAP7_75t_SL g2010 ( 
.A(n_1939),
.Y(n_2010)
);

AND2x2_ASAP7_75t_L g2011 ( 
.A(n_1966),
.B(n_1834),
.Y(n_2011)
);

HB1xp67_ASAP7_75t_L g2012 ( 
.A(n_1970),
.Y(n_2012)
);

OR2x2_ASAP7_75t_L g2013 ( 
.A(n_1932),
.B(n_1849),
.Y(n_2013)
);

HB1xp67_ASAP7_75t_L g2014 ( 
.A(n_1970),
.Y(n_2014)
);

INVx2_ASAP7_75t_L g2015 ( 
.A(n_1945),
.Y(n_2015)
);

NOR2xp33_ASAP7_75t_L g2016 ( 
.A(n_1952),
.B(n_1896),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1945),
.B(n_1834),
.Y(n_2017)
);

AND2x2_ASAP7_75t_L g2018 ( 
.A(n_1955),
.B(n_1834),
.Y(n_2018)
);

INVx1_ASAP7_75t_SL g2019 ( 
.A(n_1930),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_L g2020 ( 
.A(n_1964),
.B(n_1857),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1967),
.B(n_1852),
.Y(n_2021)
);

AND2x2_ASAP7_75t_L g2022 ( 
.A(n_1963),
.B(n_1852),
.Y(n_2022)
);

OR2x2_ASAP7_75t_L g2023 ( 
.A(n_1932),
.B(n_1849),
.Y(n_2023)
);

NOR2xp33_ASAP7_75t_R g2024 ( 
.A(n_1920),
.B(n_1904),
.Y(n_2024)
);

OR2x2_ASAP7_75t_L g2025 ( 
.A(n_1955),
.B(n_1849),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1967),
.B(n_1852),
.Y(n_2026)
);

AOI22xp33_ASAP7_75t_L g2027 ( 
.A1(n_1926),
.A2(n_1897),
.B1(n_1883),
.B2(n_1864),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_L g2028 ( 
.A(n_1973),
.B(n_1857),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1923),
.Y(n_2029)
);

INVx2_ASAP7_75t_L g2030 ( 
.A(n_1957),
.Y(n_2030)
);

INVx1_ASAP7_75t_L g2031 ( 
.A(n_1923),
.Y(n_2031)
);

AND2x2_ASAP7_75t_L g2032 ( 
.A(n_1912),
.B(n_1852),
.Y(n_2032)
);

INVx1_ASAP7_75t_L g2033 ( 
.A(n_1928),
.Y(n_2033)
);

OR2x2_ASAP7_75t_L g2034 ( 
.A(n_1958),
.B(n_1849),
.Y(n_2034)
);

INVx1_ASAP7_75t_L g2035 ( 
.A(n_1928),
.Y(n_2035)
);

INVx1_ASAP7_75t_L g2036 ( 
.A(n_1937),
.Y(n_2036)
);

AND2x2_ASAP7_75t_L g2037 ( 
.A(n_1912),
.B(n_1852),
.Y(n_2037)
);

AND2x2_ASAP7_75t_L g2038 ( 
.A(n_1921),
.B(n_1901),
.Y(n_2038)
);

NAND2xp5_ASAP7_75t_L g2039 ( 
.A(n_1973),
.B(n_1857),
.Y(n_2039)
);

AND2x2_ASAP7_75t_L g2040 ( 
.A(n_1958),
.B(n_1867),
.Y(n_2040)
);

AND2x2_ASAP7_75t_L g2041 ( 
.A(n_1960),
.B(n_1867),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_L g2042 ( 
.A(n_1975),
.B(n_1874),
.Y(n_2042)
);

OR2x2_ASAP7_75t_L g2043 ( 
.A(n_2013),
.B(n_1915),
.Y(n_2043)
);

AND2x2_ASAP7_75t_L g2044 ( 
.A(n_1987),
.B(n_1971),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1994),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1980),
.Y(n_2046)
);

INVx2_ASAP7_75t_L g2047 ( 
.A(n_1994),
.Y(n_2047)
);

AOI22xp33_ASAP7_75t_L g2048 ( 
.A1(n_1982),
.A2(n_1918),
.B1(n_1914),
.B2(n_1927),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1980),
.Y(n_2049)
);

INVx1_ASAP7_75t_L g2050 ( 
.A(n_1983),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_2028),
.Y(n_2051)
);

NOR2xp33_ASAP7_75t_L g2052 ( 
.A(n_1986),
.B(n_1920),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1983),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1982),
.B(n_1972),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_L g2055 ( 
.A(n_1988),
.B(n_1992),
.Y(n_2055)
);

INVx1_ASAP7_75t_L g2056 ( 
.A(n_1985),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1987),
.B(n_1971),
.Y(n_2057)
);

INVx1_ASAP7_75t_L g2058 ( 
.A(n_1985),
.Y(n_2058)
);

NAND2x1p5_ASAP7_75t_L g2059 ( 
.A(n_1993),
.B(n_1979),
.Y(n_2059)
);

INVx2_ASAP7_75t_L g2060 ( 
.A(n_1994),
.Y(n_2060)
);

OR2x2_ASAP7_75t_L g2061 ( 
.A(n_2013),
.B(n_1961),
.Y(n_2061)
);

INVx2_ASAP7_75t_L g2062 ( 
.A(n_1994),
.Y(n_2062)
);

INVx2_ASAP7_75t_L g2063 ( 
.A(n_2002),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1989),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1987),
.B(n_1971),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_L g2066 ( 
.A(n_1988),
.B(n_1977),
.Y(n_2066)
);

HB1xp67_ASAP7_75t_L g2067 ( 
.A(n_2028),
.Y(n_2067)
);

AND2x2_ASAP7_75t_L g2068 ( 
.A(n_1996),
.B(n_1971),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1989),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1996),
.B(n_1921),
.Y(n_2070)
);

NOR2xp33_ASAP7_75t_L g2071 ( 
.A(n_2016),
.B(n_1954),
.Y(n_2071)
);

AND2x2_ASAP7_75t_L g2072 ( 
.A(n_1996),
.B(n_1901),
.Y(n_2072)
);

NAND2xp5_ASAP7_75t_L g2073 ( 
.A(n_1992),
.B(n_1959),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_2020),
.B(n_1959),
.Y(n_2074)
);

AOI31xp33_ASAP7_75t_L g2075 ( 
.A1(n_1984),
.A2(n_1916),
.A3(n_1935),
.B(n_1942),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_2020),
.B(n_1976),
.Y(n_2076)
);

INVx1_ASAP7_75t_L g2077 ( 
.A(n_1995),
.Y(n_2077)
);

AND2x2_ASAP7_75t_L g2078 ( 
.A(n_1998),
.B(n_2021),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1995),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_2001),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_L g2081 ( 
.A(n_2038),
.B(n_1974),
.Y(n_2081)
);

INVx1_ASAP7_75t_L g2082 ( 
.A(n_2001),
.Y(n_2082)
);

OR2x2_ASAP7_75t_L g2083 ( 
.A(n_2023),
.B(n_1961),
.Y(n_2083)
);

NOR2x1_ASAP7_75t_L g2084 ( 
.A(n_1993),
.B(n_1979),
.Y(n_2084)
);

INVx1_ASAP7_75t_L g2085 ( 
.A(n_2004),
.Y(n_2085)
);

OR2x6_ASAP7_75t_L g2086 ( 
.A(n_2023),
.B(n_1898),
.Y(n_2086)
);

AND2x2_ASAP7_75t_L g2087 ( 
.A(n_1998),
.B(n_1901),
.Y(n_2087)
);

INVx2_ASAP7_75t_L g2088 ( 
.A(n_2002),
.Y(n_2088)
);

NAND2xp5_ASAP7_75t_L g2089 ( 
.A(n_2000),
.B(n_1937),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_L g2090 ( 
.A(n_2038),
.B(n_1880),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_2004),
.Y(n_2091)
);

NAND2x1_ASAP7_75t_L g2092 ( 
.A(n_2021),
.B(n_1898),
.Y(n_2092)
);

HB1xp67_ASAP7_75t_L g2093 ( 
.A(n_2039),
.Y(n_2093)
);

OR2x2_ASAP7_75t_L g2094 ( 
.A(n_2000),
.B(n_1975),
.Y(n_2094)
);

AOI21xp33_ASAP7_75t_SL g2095 ( 
.A1(n_2027),
.A2(n_1940),
.B(n_1948),
.Y(n_2095)
);

INVx2_ASAP7_75t_SL g2096 ( 
.A(n_2021),
.Y(n_2096)
);

INVx1_ASAP7_75t_L g2097 ( 
.A(n_2046),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_L g2098 ( 
.A(n_2054),
.B(n_2039),
.Y(n_2098)
);

OR2x2_ASAP7_75t_L g2099 ( 
.A(n_2055),
.B(n_1981),
.Y(n_2099)
);

BUFx2_ASAP7_75t_L g2100 ( 
.A(n_2084),
.Y(n_2100)
);

AND2x2_ASAP7_75t_L g2101 ( 
.A(n_2078),
.B(n_1998),
.Y(n_2101)
);

NOR2xp33_ASAP7_75t_R g2102 ( 
.A(n_2052),
.B(n_1925),
.Y(n_2102)
);

NOR3xp33_ASAP7_75t_L g2103 ( 
.A(n_2095),
.B(n_1929),
.C(n_1944),
.Y(n_2103)
);

NAND2x1_ASAP7_75t_L g2104 ( 
.A(n_2084),
.B(n_2021),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_2066),
.B(n_2003),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_2095),
.B(n_1984),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_2046),
.Y(n_2107)
);

AND2x4_ASAP7_75t_SL g2108 ( 
.A(n_2044),
.B(n_1930),
.Y(n_2108)
);

AND2x2_ASAP7_75t_L g2109 ( 
.A(n_2078),
.B(n_2009),
.Y(n_2109)
);

NOR2xp67_ASAP7_75t_L g2110 ( 
.A(n_2096),
.B(n_2026),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_L g2111 ( 
.A(n_2076),
.B(n_2003),
.Y(n_2111)
);

AND2x2_ASAP7_75t_L g2112 ( 
.A(n_2087),
.B(n_2009),
.Y(n_2112)
);

CKINVDCx16_ASAP7_75t_R g2113 ( 
.A(n_2070),
.Y(n_2113)
);

NAND3xp33_ASAP7_75t_L g2114 ( 
.A(n_2075),
.B(n_1924),
.C(n_1947),
.Y(n_2114)
);

NAND2xp5_ASAP7_75t_L g2115 ( 
.A(n_2081),
.B(n_2006),
.Y(n_2115)
);

INVx3_ASAP7_75t_SL g2116 ( 
.A(n_2070),
.Y(n_2116)
);

AND2x2_ASAP7_75t_L g2117 ( 
.A(n_2087),
.B(n_2009),
.Y(n_2117)
);

NOR2xp67_ASAP7_75t_SL g2118 ( 
.A(n_2074),
.B(n_1883),
.Y(n_2118)
);

INVx2_ASAP7_75t_L g2119 ( 
.A(n_2045),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2049),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_L g2121 ( 
.A(n_2090),
.B(n_2006),
.Y(n_2121)
);

O2A1O1Ixp5_ASAP7_75t_SL g2122 ( 
.A1(n_2049),
.A2(n_2008),
.B(n_2029),
.C(n_2031),
.Y(n_2122)
);

NOR2xp33_ASAP7_75t_R g2123 ( 
.A(n_2048),
.B(n_1925),
.Y(n_2123)
);

OR2x6_ASAP7_75t_L g2124 ( 
.A(n_2059),
.B(n_1902),
.Y(n_2124)
);

AND2x2_ASAP7_75t_L g2125 ( 
.A(n_2072),
.B(n_1990),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2045),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_2072),
.B(n_1990),
.Y(n_2127)
);

INVx1_ASAP7_75t_L g2128 ( 
.A(n_2050),
.Y(n_2128)
);

NOR2xp33_ASAP7_75t_SL g2129 ( 
.A(n_2071),
.B(n_1953),
.Y(n_2129)
);

NAND2xp33_ASAP7_75t_R g2130 ( 
.A(n_2073),
.B(n_1908),
.Y(n_2130)
);

AND2x2_ASAP7_75t_L g2131 ( 
.A(n_2044),
.B(n_1999),
.Y(n_2131)
);

INVx1_ASAP7_75t_L g2132 ( 
.A(n_2050),
.Y(n_2132)
);

AOI22xp5_ASAP7_75t_L g2133 ( 
.A1(n_2057),
.A2(n_1943),
.B1(n_1872),
.B2(n_1905),
.Y(n_2133)
);

INVx1_ASAP7_75t_L g2134 ( 
.A(n_2053),
.Y(n_2134)
);

INVx1_ASAP7_75t_L g2135 ( 
.A(n_2053),
.Y(n_2135)
);

INVx1_ASAP7_75t_L g2136 ( 
.A(n_2056),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_2055),
.B(n_1997),
.Y(n_2137)
);

NAND2xp33_ASAP7_75t_SL g2138 ( 
.A(n_2075),
.B(n_2024),
.Y(n_2138)
);

NOR4xp25_ASAP7_75t_SL g2139 ( 
.A(n_2059),
.B(n_2007),
.C(n_1978),
.D(n_1946),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_2056),
.Y(n_2140)
);

NAND2xp33_ASAP7_75t_R g2141 ( 
.A(n_2057),
.B(n_1981),
.Y(n_2141)
);

NOR2xp33_ASAP7_75t_R g2142 ( 
.A(n_2065),
.B(n_1950),
.Y(n_2142)
);

AND2x2_ASAP7_75t_L g2143 ( 
.A(n_2065),
.B(n_1999),
.Y(n_2143)
);

AND2x2_ASAP7_75t_L g2144 ( 
.A(n_2068),
.B(n_2005),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_2051),
.B(n_1997),
.Y(n_2145)
);

OAI22xp5_ASAP7_75t_L g2146 ( 
.A1(n_2106),
.A2(n_2007),
.B1(n_2096),
.B2(n_2059),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_2097),
.Y(n_2147)
);

NAND2xp5_ASAP7_75t_L g2148 ( 
.A(n_2103),
.B(n_2106),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_2138),
.A2(n_1872),
.B1(n_2068),
.B2(n_1880),
.Y(n_2149)
);

HB1xp67_ASAP7_75t_L g2150 ( 
.A(n_2100),
.Y(n_2150)
);

OAI21xp5_ASAP7_75t_SL g2151 ( 
.A1(n_2114),
.A2(n_2133),
.B(n_2138),
.Y(n_2151)
);

INVx2_ASAP7_75t_L g2152 ( 
.A(n_2116),
.Y(n_2152)
);

AOI22xp5_ASAP7_75t_L g2153 ( 
.A1(n_2130),
.A2(n_1943),
.B1(n_2086),
.B2(n_1905),
.Y(n_2153)
);

OAI21xp5_ASAP7_75t_L g2154 ( 
.A1(n_2122),
.A2(n_1933),
.B(n_2019),
.Y(n_2154)
);

INVx1_ASAP7_75t_L g2155 ( 
.A(n_2107),
.Y(n_2155)
);

OAI21xp33_ASAP7_75t_L g2156 ( 
.A1(n_2123),
.A2(n_2086),
.B(n_2043),
.Y(n_2156)
);

XOR2x2_ASAP7_75t_L g2157 ( 
.A(n_2116),
.B(n_1943),
.Y(n_2157)
);

INVx1_ASAP7_75t_L g2158 ( 
.A(n_2120),
.Y(n_2158)
);

NOR2xp33_ASAP7_75t_SL g2159 ( 
.A(n_2129),
.B(n_2019),
.Y(n_2159)
);

NAND3xp33_ASAP7_75t_L g2160 ( 
.A(n_2139),
.B(n_2086),
.C(n_1884),
.Y(n_2160)
);

NAND2xp33_ASAP7_75t_SL g2161 ( 
.A(n_2102),
.B(n_2092),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_SL g2162 ( 
.A1(n_2113),
.A2(n_2092),
.B1(n_2086),
.B2(n_1898),
.Y(n_2162)
);

INVx2_ASAP7_75t_L g2163 ( 
.A(n_2100),
.Y(n_2163)
);

AND2x2_ASAP7_75t_L g2164 ( 
.A(n_2109),
.B(n_2067),
.Y(n_2164)
);

AND2x2_ASAP7_75t_L g2165 ( 
.A(n_2109),
.B(n_2093),
.Y(n_2165)
);

AOI31xp33_ASAP7_75t_L g2166 ( 
.A1(n_2141),
.A2(n_2105),
.A3(n_2098),
.B(n_2111),
.Y(n_2166)
);

OAI21xp5_ASAP7_75t_L g2167 ( 
.A1(n_2122),
.A2(n_1933),
.B(n_2089),
.Y(n_2167)
);

INVx1_ASAP7_75t_L g2168 ( 
.A(n_2128),
.Y(n_2168)
);

OAI21xp33_ASAP7_75t_L g2169 ( 
.A1(n_2115),
.A2(n_2086),
.B(n_2043),
.Y(n_2169)
);

OR2x2_ASAP7_75t_L g2170 ( 
.A(n_2137),
.B(n_2094),
.Y(n_2170)
);

INVx1_ASAP7_75t_L g2171 ( 
.A(n_2132),
.Y(n_2171)
);

NAND3xp33_ASAP7_75t_L g2172 ( 
.A(n_2118),
.B(n_1885),
.C(n_2025),
.Y(n_2172)
);

NAND2xp5_ASAP7_75t_SL g2173 ( 
.A(n_2142),
.B(n_2026),
.Y(n_2173)
);

NOR2xp33_ASAP7_75t_L g2174 ( 
.A(n_2118),
.B(n_1882),
.Y(n_2174)
);

INVx2_ASAP7_75t_L g2175 ( 
.A(n_2101),
.Y(n_2175)
);

INVx1_ASAP7_75t_L g2176 ( 
.A(n_2134),
.Y(n_2176)
);

NAND2x1_ASAP7_75t_L g2177 ( 
.A(n_2124),
.B(n_2063),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_L g2178 ( 
.A(n_2125),
.B(n_2089),
.Y(n_2178)
);

INVx2_ASAP7_75t_L g2179 ( 
.A(n_2101),
.Y(n_2179)
);

INVx2_ASAP7_75t_L g2180 ( 
.A(n_2119),
.Y(n_2180)
);

AOI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_2104),
.A2(n_1849),
.B(n_1991),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_2108),
.B(n_1930),
.Y(n_2182)
);

NAND2xp33_ASAP7_75t_SL g2183 ( 
.A(n_2131),
.B(n_1991),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_2110),
.A2(n_2034),
.B(n_2025),
.Y(n_2184)
);

INVx2_ASAP7_75t_L g2185 ( 
.A(n_2177),
.Y(n_2185)
);

OAI311xp33_ASAP7_75t_L g2186 ( 
.A1(n_2151),
.A2(n_2145),
.A3(n_2099),
.B1(n_2121),
.C1(n_2140),
.Y(n_2186)
);

AND2x2_ASAP7_75t_L g2187 ( 
.A(n_2152),
.B(n_2124),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_2147),
.Y(n_2188)
);

INVx1_ASAP7_75t_SL g2189 ( 
.A(n_2152),
.Y(n_2189)
);

OAI21xp33_ASAP7_75t_SL g2190 ( 
.A1(n_2166),
.A2(n_2124),
.B(n_2112),
.Y(n_2190)
);

OAI22xp5_ASAP7_75t_L g2191 ( 
.A1(n_2160),
.A2(n_2124),
.B1(n_2108),
.B2(n_2143),
.Y(n_2191)
);

OR2x2_ASAP7_75t_L g2192 ( 
.A(n_2170),
.B(n_2099),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_2147),
.Y(n_2193)
);

O2A1O1Ixp33_ASAP7_75t_SL g2194 ( 
.A1(n_2148),
.A2(n_2136),
.B(n_2135),
.C(n_2063),
.Y(n_2194)
);

OAI222xp33_ASAP7_75t_L g2195 ( 
.A1(n_2146),
.A2(n_2144),
.B1(n_2143),
.B2(n_2131),
.C1(n_2112),
.C2(n_2117),
.Y(n_2195)
);

AND2x2_ASAP7_75t_L g2196 ( 
.A(n_2175),
.B(n_2144),
.Y(n_2196)
);

NAND2xp33_ASAP7_75t_L g2197 ( 
.A(n_2149),
.B(n_2125),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_2155),
.Y(n_2198)
);

HB1xp67_ASAP7_75t_L g2199 ( 
.A(n_2150),
.Y(n_2199)
);

INVx2_ASAP7_75t_L g2200 ( 
.A(n_2177),
.Y(n_2200)
);

NAND2xp5_ASAP7_75t_SL g2201 ( 
.A(n_2159),
.B(n_2127),
.Y(n_2201)
);

INVx1_ASAP7_75t_L g2202 ( 
.A(n_2155),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2174),
.B(n_2127),
.Y(n_2203)
);

AOI222xp33_ASAP7_75t_L g2204 ( 
.A1(n_2156),
.A2(n_1872),
.B1(n_2117),
.B2(n_2063),
.C1(n_2088),
.C2(n_2091),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2168),
.Y(n_2205)
);

NOR2xp33_ASAP7_75t_L g2206 ( 
.A(n_2173),
.B(n_2094),
.Y(n_2206)
);

OAI221xp5_ASAP7_75t_L g2207 ( 
.A1(n_2153),
.A2(n_2126),
.B1(n_2119),
.B2(n_2034),
.C(n_2080),
.Y(n_2207)
);

AOI31xp33_ASAP7_75t_L g2208 ( 
.A1(n_2182),
.A2(n_2088),
.A3(n_2126),
.B(n_2037),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2168),
.Y(n_2209)
);

OAI21xp5_ASAP7_75t_SL g2210 ( 
.A1(n_2169),
.A2(n_1866),
.B(n_1873),
.Y(n_2210)
);

OAI22xp5_ASAP7_75t_L g2211 ( 
.A1(n_2172),
.A2(n_1898),
.B1(n_2058),
.B2(n_2085),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2171),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_2171),
.Y(n_2213)
);

INVx1_ASAP7_75t_L g2214 ( 
.A(n_2199),
.Y(n_2214)
);

NAND2xp33_ASAP7_75t_SL g2215 ( 
.A(n_2201),
.B(n_2163),
.Y(n_2215)
);

OR2x2_ASAP7_75t_L g2216 ( 
.A(n_2189),
.B(n_2175),
.Y(n_2216)
);

NOR2x1_ASAP7_75t_L g2217 ( 
.A(n_2185),
.B(n_2163),
.Y(n_2217)
);

CKINVDCx20_ASAP7_75t_R g2218 ( 
.A(n_2191),
.Y(n_2218)
);

INVx2_ASAP7_75t_SL g2219 ( 
.A(n_2185),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2188),
.Y(n_2220)
);

AND2x4_ASAP7_75t_L g2221 ( 
.A(n_2200),
.B(n_2179),
.Y(n_2221)
);

NOR2xp67_ASAP7_75t_L g2222 ( 
.A(n_2190),
.B(n_2179),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_2188),
.Y(n_2223)
);

NAND2xp5_ASAP7_75t_L g2224 ( 
.A(n_2196),
.B(n_2197),
.Y(n_2224)
);

XNOR2xp5_ASAP7_75t_L g2225 ( 
.A(n_2187),
.B(n_2157),
.Y(n_2225)
);

AND2x2_ASAP7_75t_L g2226 ( 
.A(n_2187),
.B(n_2164),
.Y(n_2226)
);

XOR2x2_ASAP7_75t_L g2227 ( 
.A(n_2186),
.B(n_2157),
.Y(n_2227)
);

INVx1_ASAP7_75t_L g2228 ( 
.A(n_2193),
.Y(n_2228)
);

AND2x2_ASAP7_75t_L g2229 ( 
.A(n_2196),
.B(n_2164),
.Y(n_2229)
);

NAND2xp5_ASAP7_75t_L g2230 ( 
.A(n_2197),
.B(n_2165),
.Y(n_2230)
);

NOR2x1_ASAP7_75t_L g2231 ( 
.A(n_2200),
.B(n_2176),
.Y(n_2231)
);

INVxp67_ASAP7_75t_L g2232 ( 
.A(n_2192),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2206),
.B(n_2165),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_2193),
.Y(n_2234)
);

NOR3xp33_ASAP7_75t_SL g2235 ( 
.A(n_2195),
.B(n_2161),
.C(n_2162),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2192),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_2236),
.Y(n_2237)
);

NOR2xp33_ASAP7_75t_L g2238 ( 
.A(n_2232),
.B(n_2203),
.Y(n_2238)
);

OAI21xp5_ASAP7_75t_SL g2239 ( 
.A1(n_2230),
.A2(n_2210),
.B(n_2208),
.Y(n_2239)
);

INVx1_ASAP7_75t_L g2240 ( 
.A(n_2236),
.Y(n_2240)
);

NOR2x1_ASAP7_75t_L g2241 ( 
.A(n_2217),
.B(n_2202),
.Y(n_2241)
);

NAND3xp33_ASAP7_75t_L g2242 ( 
.A(n_2215),
.B(n_2194),
.C(n_2204),
.Y(n_2242)
);

NOR3x1_ASAP7_75t_L g2243 ( 
.A(n_2224),
.B(n_2198),
.C(n_2205),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_2226),
.B(n_2202),
.Y(n_2244)
);

INVx1_ASAP7_75t_L g2245 ( 
.A(n_2214),
.Y(n_2245)
);

AOI221xp5_ASAP7_75t_L g2246 ( 
.A1(n_2215),
.A2(n_2207),
.B1(n_2211),
.B2(n_2212),
.C(n_2209),
.Y(n_2246)
);

AOI221xp5_ASAP7_75t_L g2247 ( 
.A1(n_2235),
.A2(n_2213),
.B1(n_2212),
.B2(n_2209),
.C(n_2161),
.Y(n_2247)
);

INVx1_ASAP7_75t_L g2248 ( 
.A(n_2216),
.Y(n_2248)
);

AND3x1_ASAP7_75t_L g2249 ( 
.A(n_2235),
.B(n_2213),
.C(n_2154),
.Y(n_2249)
);

NOR3xp33_ASAP7_75t_SL g2250 ( 
.A(n_2233),
.B(n_2183),
.C(n_2181),
.Y(n_2250)
);

NAND2xp5_ASAP7_75t_L g2251 ( 
.A(n_2229),
.B(n_2158),
.Y(n_2251)
);

INVx1_ASAP7_75t_L g2252 ( 
.A(n_2241),
.Y(n_2252)
);

NAND2xp33_ASAP7_75t_L g2253 ( 
.A(n_2250),
.B(n_2225),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_R g2254 ( 
.A(n_2248),
.B(n_2218),
.Y(n_2254)
);

OAI211xp5_ASAP7_75t_SL g2255 ( 
.A1(n_2247),
.A2(n_2227),
.B(n_2231),
.C(n_2228),
.Y(n_2255)
);

OAI211xp5_ASAP7_75t_SL g2256 ( 
.A1(n_2239),
.A2(n_2227),
.B(n_2234),
.C(n_2223),
.Y(n_2256)
);

AOI21xp33_ASAP7_75t_SL g2257 ( 
.A1(n_2242),
.A2(n_2219),
.B(n_2221),
.Y(n_2257)
);

NAND2xp33_ASAP7_75t_L g2258 ( 
.A(n_2250),
.B(n_2218),
.Y(n_2258)
);

INVxp67_ASAP7_75t_L g2259 ( 
.A(n_2238),
.Y(n_2259)
);

AND2x4_ASAP7_75t_L g2260 ( 
.A(n_2237),
.B(n_2219),
.Y(n_2260)
);

OAI211xp5_ASAP7_75t_SL g2261 ( 
.A1(n_2246),
.A2(n_2220),
.B(n_2167),
.C(n_2222),
.Y(n_2261)
);

NAND4xp25_ASAP7_75t_L g2262 ( 
.A(n_2243),
.B(n_2221),
.C(n_2183),
.D(n_2176),
.Y(n_2262)
);

OAI211xp5_ASAP7_75t_L g2263 ( 
.A1(n_2244),
.A2(n_2184),
.B(n_2180),
.C(n_2170),
.Y(n_2263)
);

AOI221xp5_ASAP7_75t_L g2264 ( 
.A1(n_2249),
.A2(n_2221),
.B1(n_2180),
.B2(n_2178),
.C(n_2091),
.Y(n_2264)
);

INVx1_ASAP7_75t_L g2265 ( 
.A(n_2240),
.Y(n_2265)
);

NOR2x1_ASAP7_75t_R g2266 ( 
.A(n_2245),
.B(n_1877),
.Y(n_2266)
);

CKINVDCx16_ASAP7_75t_R g2267 ( 
.A(n_2254),
.Y(n_2267)
);

BUFx12f_ASAP7_75t_L g2268 ( 
.A(n_2260),
.Y(n_2268)
);

AOI211xp5_ASAP7_75t_L g2269 ( 
.A1(n_2255),
.A2(n_2251),
.B(n_2088),
.C(n_2085),
.Y(n_2269)
);

NAND4xp25_ASAP7_75t_L g2270 ( 
.A(n_2256),
.B(n_2032),
.C(n_2037),
.D(n_2011),
.Y(n_2270)
);

OAI22xp5_ASAP7_75t_L g2271 ( 
.A1(n_2252),
.A2(n_2045),
.B1(n_2047),
.B2(n_2060),
.Y(n_2271)
);

OAI211xp5_ASAP7_75t_L g2272 ( 
.A1(n_2257),
.A2(n_2261),
.B(n_2262),
.C(n_2259),
.Y(n_2272)
);

INVx1_ASAP7_75t_L g2273 ( 
.A(n_2260),
.Y(n_2273)
);

CKINVDCx5p33_ASAP7_75t_R g2274 ( 
.A(n_2265),
.Y(n_2274)
);

XNOR2xp5_ASAP7_75t_L g2275 ( 
.A(n_2264),
.B(n_1881),
.Y(n_2275)
);

OAI22xp5_ASAP7_75t_L g2276 ( 
.A1(n_2263),
.A2(n_2047),
.B1(n_2060),
.B2(n_2062),
.Y(n_2276)
);

O2A1O1Ixp33_ASAP7_75t_L g2277 ( 
.A1(n_2253),
.A2(n_1898),
.B(n_2082),
.C(n_2080),
.Y(n_2277)
);

AOI211xp5_ASAP7_75t_L g2278 ( 
.A1(n_2272),
.A2(n_2258),
.B(n_2266),
.C(n_2077),
.Y(n_2278)
);

NOR2x1_ASAP7_75t_L g2279 ( 
.A(n_2273),
.B(n_2058),
.Y(n_2279)
);

AOI21x1_ASAP7_75t_L g2280 ( 
.A1(n_2268),
.A2(n_2047),
.B(n_2060),
.Y(n_2280)
);

NAND3xp33_ASAP7_75t_L g2281 ( 
.A(n_2269),
.B(n_2082),
.C(n_2079),
.Y(n_2281)
);

NAND2xp5_ASAP7_75t_L g2282 ( 
.A(n_2267),
.B(n_2064),
.Y(n_2282)
);

NAND3xp33_ASAP7_75t_SL g2283 ( 
.A(n_2274),
.B(n_2083),
.C(n_2061),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_2275),
.B(n_2064),
.Y(n_2284)
);

AOI221xp5_ASAP7_75t_SL g2285 ( 
.A1(n_2270),
.A2(n_2079),
.B1(n_2077),
.B2(n_2069),
.C(n_2062),
.Y(n_2285)
);

NAND2xp5_ASAP7_75t_L g2286 ( 
.A(n_2278),
.B(n_2277),
.Y(n_2286)
);

O2A1O1Ixp33_ASAP7_75t_L g2287 ( 
.A1(n_2282),
.A2(n_2276),
.B(n_2271),
.C(n_2062),
.Y(n_2287)
);

NAND3xp33_ASAP7_75t_SL g2288 ( 
.A(n_2284),
.B(n_2083),
.C(n_2061),
.Y(n_2288)
);

AO22x2_ASAP7_75t_L g2289 ( 
.A1(n_2283),
.A2(n_2069),
.B1(n_2002),
.B2(n_2010),
.Y(n_2289)
);

NOR3xp33_ASAP7_75t_L g2290 ( 
.A(n_2279),
.B(n_1855),
.C(n_1893),
.Y(n_2290)
);

AND2x4_ASAP7_75t_L g2291 ( 
.A(n_2280),
.B(n_2281),
.Y(n_2291)
);

NOR2x2_ASAP7_75t_L g2292 ( 
.A(n_2285),
.B(n_1878),
.Y(n_2292)
);

AOI21xp5_ASAP7_75t_L g2293 ( 
.A1(n_2282),
.A2(n_1855),
.B(n_2042),
.Y(n_2293)
);

INVx1_ASAP7_75t_SL g2294 ( 
.A(n_2291),
.Y(n_2294)
);

INVx2_ASAP7_75t_L g2295 ( 
.A(n_2292),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2286),
.A2(n_2287),
.B(n_2288),
.Y(n_2296)
);

O2A1O1Ixp33_ASAP7_75t_L g2297 ( 
.A1(n_2290),
.A2(n_2010),
.B(n_2014),
.C(n_2012),
.Y(n_2297)
);

INVxp67_ASAP7_75t_SL g2298 ( 
.A(n_2295),
.Y(n_2298)
);

AOI222xp33_ASAP7_75t_L g2299 ( 
.A1(n_2294),
.A2(n_2289),
.B1(n_2293),
.B2(n_2022),
.C1(n_2005),
.C2(n_2011),
.Y(n_2299)
);

AOI22xp33_ASAP7_75t_L g2300 ( 
.A1(n_2298),
.A2(n_2296),
.B1(n_2297),
.B2(n_1893),
.Y(n_2300)
);

OAI21xp5_ASAP7_75t_L g2301 ( 
.A1(n_2299),
.A2(n_2042),
.B(n_2032),
.Y(n_2301)
);

INVx1_ASAP7_75t_L g2302 ( 
.A(n_2300),
.Y(n_2302)
);

AOI22xp33_ASAP7_75t_R g2303 ( 
.A1(n_2301),
.A2(n_2014),
.B1(n_2012),
.B2(n_2010),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2300),
.Y(n_2304)
);

AOI22xp33_ASAP7_75t_L g2305 ( 
.A1(n_2302),
.A2(n_2008),
.B1(n_2031),
.B2(n_2033),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_2304),
.B(n_1882),
.Y(n_2306)
);

AOI222xp33_ASAP7_75t_L g2307 ( 
.A1(n_2306),
.A2(n_2303),
.B1(n_2029),
.B2(n_2033),
.C1(n_2036),
.C2(n_2035),
.Y(n_2307)
);

AOI22xp33_ASAP7_75t_SL g2308 ( 
.A1(n_2305),
.A2(n_2041),
.B1(n_2040),
.B2(n_2036),
.Y(n_2308)
);

AOI322xp5_ASAP7_75t_L g2309 ( 
.A1(n_2308),
.A2(n_2041),
.A3(n_2040),
.B1(n_2022),
.B2(n_2017),
.C1(n_2018),
.C2(n_2035),
.Y(n_2309)
);

OAI221xp5_ASAP7_75t_R g2310 ( 
.A1(n_2309),
.A2(n_2307),
.B1(n_2040),
.B2(n_2041),
.C(n_2015),
.Y(n_2310)
);

AOI211xp5_ASAP7_75t_L g2311 ( 
.A1(n_2310),
.A2(n_1892),
.B(n_1903),
.C(n_2030),
.Y(n_2311)
);


endmodule