module fake_jpeg_5886_n_170 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_170);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_170;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

HB1xp67_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

BUFx12_ASAP7_75t_L g16 ( 
.A(n_13),
.Y(n_16)
);

BUFx12_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

INVx3_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_11),
.B(n_1),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_24),
.Y(n_31)
);

INVx8_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

AND2x2_ASAP7_75t_SL g33 ( 
.A(n_15),
.B(n_0),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_35),
.Y(n_39)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_24),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_19),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_38),
.Y(n_47)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_41),
.B(n_42),
.Y(n_57)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_44),
.Y(n_72)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx8_ASAP7_75t_L g54 ( 
.A(n_45),
.Y(n_54)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_40),
.B(n_32),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_53),
.B(n_56),
.Y(n_91)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_55),
.B(n_60),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_42),
.B(n_22),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_20),
.B1(n_30),
.B2(n_22),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_L g83 ( 
.A1(n_59),
.A2(n_49),
.B1(n_27),
.B2(n_25),
.Y(n_83)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_28),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_61),
.B(n_28),
.Y(n_82)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_47),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_63),
.Y(n_80)
);

BUFx12f_ASAP7_75t_L g63 ( 
.A(n_39),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_64),
.B(n_65),
.Y(n_90)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_47),
.Y(n_65)
);

O2A1O1Ixp33_ASAP7_75t_L g66 ( 
.A1(n_51),
.A2(n_18),
.B(n_15),
.C(n_34),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_66),
.B(n_67),
.Y(n_93)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_48),
.Y(n_68)
);

INVx3_ASAP7_75t_SL g94 ( 
.A(n_68),
.Y(n_94)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_50),
.Y(n_69)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

MAJx2_ASAP7_75t_L g70 ( 
.A(n_51),
.B(n_37),
.C(n_34),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_70),
.B(n_74),
.C(n_58),
.Y(n_88)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

BUFx24_ASAP7_75t_SL g79 ( 
.A(n_71),
.Y(n_79)
);

OAI22xp5_ASAP7_75t_L g73 ( 
.A1(n_46),
.A2(n_20),
.B1(n_26),
.B2(n_25),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_73),
.B(n_74),
.Y(n_81)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_46),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_57),
.B(n_26),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_70),
.A2(n_49),
.B1(n_37),
.B2(n_31),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_78),
.A2(n_85),
.B1(n_95),
.B2(n_65),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_82),
.B(n_28),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_SL g109 ( 
.A1(n_83),
.A2(n_16),
.B1(n_63),
.B2(n_28),
.Y(n_109)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_72),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_86),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_61),
.A2(n_31),
.B1(n_38),
.B2(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_87),
.B(n_89),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_88),
.B(n_82),
.C(n_78),
.Y(n_97)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g92 ( 
.A(n_62),
.B(n_29),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_17),
.B(n_16),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_69),
.A2(n_27),
.B1(n_23),
.B2(n_19),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_109),
.B1(n_77),
.B2(n_92),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_97),
.B(n_112),
.C(n_83),
.Y(n_116)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_80),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_86),
.A2(n_58),
.B1(n_54),
.B2(n_67),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_101),
.B(n_104),
.Y(n_127)
);

NOR2x1p5_ASAP7_75t_L g102 ( 
.A(n_85),
.B(n_19),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_105),
.B(n_110),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_89),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_103),
.Y(n_118)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_76),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_88),
.A2(n_93),
.B(n_81),
.Y(n_105)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_106),
.Y(n_119)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_90),
.Y(n_107)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_107),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_21),
.Y(n_108)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g111 ( 
.A(n_75),
.B(n_0),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_111),
.Y(n_114)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_84),
.B(n_63),
.C(n_16),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_81),
.Y(n_113)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_113),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g131 ( 
.A1(n_115),
.A2(n_102),
.B1(n_101),
.B2(n_98),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_116),
.B(n_120),
.C(n_122),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_97),
.B(n_77),
.C(n_87),
.Y(n_120)
);

XOR2x2_ASAP7_75t_L g121 ( 
.A(n_105),
.B(n_79),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_121),
.A2(n_1),
.B(n_3),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_106),
.B(n_95),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_L g124 ( 
.A1(n_113),
.A2(n_92),
.B(n_94),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g134 ( 
.A(n_124),
.B(n_94),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g128 ( 
.A(n_96),
.B(n_94),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_128),
.B(n_112),
.C(n_99),
.Y(n_133)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_118),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_129),
.Y(n_146)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_131),
.A2(n_136),
.B(n_137),
.Y(n_143)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_117),
.A2(n_102),
.A3(n_110),
.B1(n_108),
.B2(n_107),
.C1(n_100),
.C2(n_104),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_132),
.B(n_134),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_133),
.B(n_139),
.C(n_125),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g135 ( 
.A1(n_127),
.A2(n_17),
.B1(n_16),
.B2(n_4),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_135),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_117),
.A2(n_17),
.B1(n_12),
.B2(n_4),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_119),
.A2(n_126),
.B1(n_128),
.B2(n_124),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_116),
.A2(n_17),
.B1(n_3),
.B2(n_4),
.Y(n_138)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_122),
.Y(n_140)
);

HB1xp67_ASAP7_75t_L g148 ( 
.A(n_140),
.Y(n_148)
);

OAI321xp33_ASAP7_75t_L g141 ( 
.A1(n_137),
.A2(n_121),
.A3(n_123),
.B1(n_119),
.B2(n_120),
.C(n_114),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_131),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_142),
.B(n_149),
.C(n_1),
.Y(n_155)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_145),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_130),
.B(n_133),
.C(n_134),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_150),
.B(n_156),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_144),
.B(n_136),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_155),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_146),
.B(n_129),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_152),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_130),
.B1(n_138),
.B2(n_6),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_154),
.B(n_5),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_147),
.A2(n_148),
.B1(n_142),
.B2(n_149),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_153),
.A2(n_145),
.B1(n_144),
.B2(n_9),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_159),
.B(n_162),
.Y(n_163)
);

AOI31xp67_ASAP7_75t_L g162 ( 
.A1(n_154),
.A2(n_5),
.A3(n_8),
.B(n_9),
.Y(n_162)
);

MAJx2_ASAP7_75t_L g164 ( 
.A(n_161),
.B(n_151),
.C(n_155),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_164),
.A2(n_165),
.B(n_160),
.Y(n_166)
);

MAJx2_ASAP7_75t_L g165 ( 
.A(n_161),
.B(n_158),
.C(n_157),
.Y(n_165)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_166),
.A2(n_167),
.B1(n_10),
.B2(n_159),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_163),
.B(n_9),
.Y(n_167)
);

BUFx24_ASAP7_75t_SL g169 ( 
.A(n_168),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g170 ( 
.A(n_169),
.Y(n_170)
);


endmodule