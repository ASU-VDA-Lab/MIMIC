module fake_jpeg_11598_n_424 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_424);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_424;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx4f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_3),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_17),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_16),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_9),
.Y(n_36)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

BUFx12_ASAP7_75t_L g44 ( 
.A(n_2),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_18),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_45),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_27),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_46),
.A2(n_71),
.B1(n_28),
.B2(n_30),
.Y(n_134)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_23),
.Y(n_47)
);

INVx2_ASAP7_75t_SL g102 ( 
.A(n_47),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_44),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_48),
.B(n_53),
.Y(n_89)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_24),
.Y(n_49)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_49),
.Y(n_93)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_23),
.Y(n_50)
);

INVx3_ASAP7_75t_L g124 ( 
.A(n_50),
.Y(n_124)
);

INVx13_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_51),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_44),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_54),
.B(n_57),
.Y(n_90)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_55),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_18),
.Y(n_56)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_56),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_22),
.Y(n_57)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_24),
.Y(n_58)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_58),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_24),
.B(n_32),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g111 ( 
.A(n_59),
.B(n_63),
.Y(n_111)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

INVx4_ASAP7_75t_L g117 ( 
.A(n_60),
.Y(n_117)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_61),
.Y(n_106)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_19),
.Y(n_62)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_62),
.Y(n_91)
);

INVx4_ASAP7_75t_SL g63 ( 
.A(n_19),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_25),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_64),
.B(n_69),
.Y(n_92)
);

BUFx5_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx4_ASAP7_75t_L g123 ( 
.A(n_65),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_21),
.Y(n_66)
);

INVx6_ASAP7_75t_L g99 ( 
.A(n_66),
.Y(n_99)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_27),
.Y(n_68)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_68),
.Y(n_130)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_23),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g101 ( 
.A(n_70),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_32),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_27),
.Y(n_72)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_72),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_21),
.Y(n_73)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_74),
.Y(n_118)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_23),
.Y(n_75)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_75),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_31),
.Y(n_76)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_76),
.Y(n_133)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_23),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g120 ( 
.A(n_77),
.B(n_79),
.Y(n_120)
);

BUFx12_ASAP7_75t_L g78 ( 
.A(n_23),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_78),
.B(n_80),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_31),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_31),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_20),
.B(n_0),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_81),
.B(n_82),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_20),
.B(n_4),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

AO22x1_ASAP7_75t_L g114 ( 
.A1(n_83),
.A2(n_22),
.B1(n_42),
.B2(n_43),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_33),
.B(n_4),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g109 ( 
.A(n_84),
.B(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_31),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_86),
.B(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_59),
.B(n_32),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_59),
.B(n_38),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_49),
.B(n_35),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_96),
.B(n_108),
.Y(n_165)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_68),
.A2(n_26),
.B1(n_37),
.B2(n_42),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_L g156 ( 
.A1(n_100),
.A2(n_121),
.B1(n_122),
.B2(n_125),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_35),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_110),
.B(n_80),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_38),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_112),
.B(n_65),
.Y(n_174)
);

OA22x2_ASAP7_75t_L g177 ( 
.A1(n_114),
.A2(n_60),
.B1(n_22),
.B2(n_55),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_47),
.B(n_41),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_128),
.Y(n_147)
);

OAI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_46),
.A2(n_86),
.B1(n_85),
.B2(n_45),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_119),
.A2(n_134),
.B1(n_135),
.B2(n_56),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_72),
.A2(n_26),
.B1(n_37),
.B2(n_42),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g122 ( 
.A1(n_61),
.A2(n_37),
.B1(n_36),
.B2(n_26),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_L g125 ( 
.A1(n_67),
.A2(n_36),
.B1(n_43),
.B2(n_30),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_62),
.A2(n_42),
.B1(n_34),
.B2(n_29),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_127),
.A2(n_129),
.B1(n_132),
.B2(n_22),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_50),
.B(n_41),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g129 ( 
.A1(n_52),
.A2(n_66),
.B1(n_79),
.B2(n_76),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_73),
.A2(n_33),
.B1(n_40),
.B2(n_39),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_74),
.A2(n_42),
.B1(n_40),
.B2(n_39),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_83),
.B1(n_78),
.B2(n_63),
.Y(n_136)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_136),
.Y(n_184)
);

CKINVDCx16_ASAP7_75t_R g137 ( 
.A(n_89),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_137),
.B(n_152),
.Y(n_183)
);

OR2x2_ASAP7_75t_SL g138 ( 
.A(n_105),
.B(n_75),
.Y(n_138)
);

CKINVDCx14_ASAP7_75t_R g206 ( 
.A(n_138),
.Y(n_206)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_139),
.Y(n_188)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_93),
.Y(n_140)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_140),
.Y(n_209)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_141),
.Y(n_191)
);

INVx6_ASAP7_75t_L g143 ( 
.A(n_98),
.Y(n_143)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_143),
.Y(n_189)
);

INVx3_ASAP7_75t_L g144 ( 
.A(n_131),
.Y(n_144)
);

BUFx2_ASAP7_75t_L g212 ( 
.A(n_144),
.Y(n_212)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_130),
.Y(n_145)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_145),
.Y(n_196)
);

XNOR2x1_ASAP7_75t_L g208 ( 
.A(n_146),
.B(n_174),
.Y(n_208)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_130),
.Y(n_148)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_148),
.Y(n_207)
);

OAI22xp33_ASAP7_75t_L g149 ( 
.A1(n_122),
.A2(n_70),
.B1(n_83),
.B2(n_28),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_149),
.A2(n_125),
.B1(n_120),
.B2(n_133),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_92),
.B(n_34),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_150),
.B(n_151),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_90),
.B(n_29),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_126),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_101),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_153),
.B(n_157),
.Y(n_185)
);

INVx4_ASAP7_75t_L g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_109),
.B(n_42),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_91),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_134),
.A2(n_43),
.B1(n_28),
.B2(n_30),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_158),
.A2(n_164),
.B1(n_111),
.B2(n_123),
.Y(n_180)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_93),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_163),
.Y(n_197)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_126),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_160),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_87),
.B(n_88),
.C(n_112),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_161),
.B(n_94),
.C(n_124),
.Y(n_190)
);

A2O1A1Ixp33_ASAP7_75t_L g162 ( 
.A1(n_111),
.A2(n_51),
.B(n_78),
.C(n_55),
.Y(n_162)
);

NOR2x1_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_115),
.Y(n_194)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_95),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_166),
.A2(n_99),
.B1(n_123),
.B2(n_104),
.Y(n_203)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_95),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_168),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_120),
.Y(n_168)
);

INVx5_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_169),
.B(n_172),
.Y(n_205)
);

INVx2_ASAP7_75t_SL g170 ( 
.A(n_133),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g202 ( 
.A(n_170),
.Y(n_202)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_171),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_111),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_97),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_173),
.B(n_175),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_103),
.B(n_56),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_102),
.Y(n_176)
);

OAI21xp33_ASAP7_75t_L g181 ( 
.A1(n_176),
.A2(n_178),
.B(n_120),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_177),
.A2(n_136),
.B1(n_149),
.B2(n_162),
.Y(n_210)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_102),
.Y(n_178)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_139),
.A2(n_103),
.B1(n_135),
.B2(n_117),
.Y(n_179)
);

OAI22xp33_ASAP7_75t_SL g241 ( 
.A1(n_179),
.A2(n_203),
.B1(n_186),
.B2(n_184),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_180),
.A2(n_198),
.B1(n_201),
.B2(n_156),
.Y(n_224)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_181),
.B(n_186),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_190),
.B(n_192),
.C(n_146),
.Y(n_222)
);

XNOR2xp5_ASAP7_75t_L g192 ( 
.A(n_161),
.B(n_124),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_194),
.B(n_214),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_142),
.B(n_118),
.C(n_97),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_195),
.B(n_177),
.C(n_136),
.Y(n_237)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_164),
.A2(n_113),
.B1(n_118),
.B2(n_106),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_174),
.A2(n_113),
.B1(n_106),
.B2(n_99),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_203),
.A2(n_210),
.B1(n_170),
.B2(n_98),
.Y(n_242)
);

AOI32xp33_ASAP7_75t_L g204 ( 
.A1(n_165),
.A2(n_107),
.A3(n_91),
.B1(n_106),
.B2(n_98),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_204),
.B(n_177),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_142),
.B(n_107),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_138),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_216),
.B(n_223),
.Y(n_273)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_209),
.Y(n_217)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_217),
.Y(n_248)
);

INVxp33_ASAP7_75t_L g218 ( 
.A(n_185),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_220),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g252 ( 
.A1(n_219),
.A2(n_225),
.B(n_240),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_197),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_197),
.Y(n_221)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_221),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_222),
.B(n_199),
.C(n_213),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_188),
.B(n_147),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_224),
.A2(n_238),
.B1(n_199),
.B2(n_205),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_206),
.A2(n_146),
.B1(n_157),
.B2(n_144),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_160),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_226),
.B(n_229),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_192),
.B(n_140),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_227),
.B(n_230),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g228 ( 
.A(n_191),
.Y(n_228)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_228),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_176),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_195),
.B(n_163),
.Y(n_230)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_189),
.Y(n_231)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_183),
.B(n_171),
.Y(n_232)
);

CKINVDCx16_ASAP7_75t_R g255 ( 
.A(n_232),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_195),
.B(n_159),
.Y(n_233)
);

NOR3xp33_ASAP7_75t_SL g257 ( 
.A(n_233),
.B(n_234),
.C(n_235),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_214),
.B(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_190),
.B(n_167),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_208),
.B(n_206),
.Y(n_236)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_236),
.B(n_227),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g261 ( 
.A(n_237),
.B(n_222),
.C(n_235),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_180),
.A2(n_177),
.B1(n_170),
.B2(n_141),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_182),
.A2(n_184),
.B1(n_198),
.B2(n_194),
.Y(n_240)
);

AOI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_241),
.A2(n_194),
.B1(n_208),
.B2(n_205),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_242),
.A2(n_245),
.B1(n_201),
.B2(n_202),
.Y(n_246)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_185),
.Y(n_243)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_243),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_183),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_244),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_210),
.A2(n_104),
.B1(n_173),
.B2(n_143),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_246),
.A2(n_250),
.B1(n_259),
.B2(n_262),
.Y(n_285)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_219),
.A2(n_179),
.B1(n_208),
.B2(n_204),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_249),
.B1(n_265),
.B2(n_239),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_253),
.B(n_261),
.C(n_264),
.Y(n_297)
);

AOI21xp5_ASAP7_75t_L g254 ( 
.A1(n_239),
.A2(n_213),
.B(n_193),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g294 ( 
.A(n_254),
.B(n_169),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g259 ( 
.A1(n_241),
.A2(n_202),
.B1(n_187),
.B2(n_189),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_242),
.A2(n_212),
.B1(n_191),
.B2(n_207),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_234),
.B(n_207),
.C(n_196),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_224),
.A2(n_104),
.B1(n_212),
.B2(n_191),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_266),
.B(n_271),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_232),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_268),
.B(n_229),
.Y(n_279)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_245),
.A2(n_212),
.B1(n_196),
.B2(n_211),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_238),
.B1(n_231),
.B2(n_230),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_236),
.B(n_211),
.C(n_209),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_148),
.C(n_145),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_272),
.B(n_225),
.Y(n_286)
);

AOI32xp33_ASAP7_75t_L g275 ( 
.A1(n_268),
.A2(n_215),
.A3(n_244),
.B1(n_216),
.B2(n_223),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_275),
.B(n_280),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_247),
.A2(n_239),
.B1(n_243),
.B2(n_221),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_276),
.A2(n_278),
.B(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_258),
.B(n_220),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_277),
.B(n_279),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_249),
.A2(n_239),
.B1(n_237),
.B2(n_240),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_270),
.B(n_258),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_256),
.Y(n_281)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_281),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_283),
.A2(n_288),
.B1(n_301),
.B2(n_250),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_267),
.B(n_233),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_284),
.B(n_289),
.Y(n_313)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_272),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_L g302 ( 
.A1(n_287),
.A2(n_300),
.B1(n_255),
.B2(n_264),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_265),
.A2(n_237),
.B1(n_215),
.B2(n_231),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_267),
.B(n_226),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_256),
.B(n_217),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_290),
.B(n_291),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g291 ( 
.A(n_270),
.B(n_228),
.Y(n_291)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_248),
.Y(n_292)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_292),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_251),
.Y(n_293)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_293),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_228),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_295),
.B(n_296),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_269),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_248),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g319 ( 
.A(n_298),
.B(n_299),
.Y(n_319)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_263),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_263),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_255),
.A2(n_273),
.B1(n_253),
.B2(n_252),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_296),
.B1(n_284),
.B2(n_281),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_282),
.B(n_261),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_306),
.C(n_315),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_285),
.A2(n_261),
.B1(n_252),
.B2(n_273),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_304),
.A2(n_308),
.B1(n_298),
.B2(n_292),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_305),
.A2(n_314),
.B1(n_321),
.B2(n_5),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_282),
.B(n_266),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_287),
.A2(n_257),
.B1(n_271),
.B2(n_274),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_310),
.B(n_325),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g312 ( 
.A1(n_278),
.A2(n_254),
.B(n_259),
.Y(n_312)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_312),
.A2(n_294),
.B(n_288),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_283),
.A2(n_246),
.B1(n_262),
.B2(n_257),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_266),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g316 ( 
.A(n_297),
.B(n_274),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_316),
.B(n_320),
.C(n_289),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_301),
.B(n_257),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_276),
.A2(n_260),
.B1(n_154),
.B2(n_7),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_SL g325 ( 
.A(n_286),
.B(n_260),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_307),
.B(n_293),
.Y(n_326)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_326),
.Y(n_353)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_319),
.Y(n_328)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_328),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_324),
.B(n_277),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_329),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_330),
.B(n_336),
.Y(n_361)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_319),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g351 ( 
.A(n_331),
.B(n_333),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g362 ( 
.A(n_332),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g334 ( 
.A(n_311),
.B(n_295),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_SL g359 ( 
.A(n_334),
.B(n_339),
.Y(n_359)
);

O2A1O1Ixp33_ASAP7_75t_L g335 ( 
.A1(n_317),
.A2(n_294),
.B(n_290),
.C(n_300),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_335),
.B(n_338),
.Y(n_363)
);

CKINVDCx16_ASAP7_75t_R g337 ( 
.A(n_319),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g357 ( 
.A(n_337),
.B(n_321),
.Y(n_357)
);

CKINVDCx16_ASAP7_75t_R g338 ( 
.A(n_317),
.Y(n_338)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_316),
.B(n_299),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_303),
.B(n_5),
.C(n_6),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_341),
.B(n_322),
.C(n_309),
.Y(n_352)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_315),
.B(n_5),
.Y(n_342)
);

XOR2xp5_ASAP7_75t_L g348 ( 
.A(n_342),
.B(n_306),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_343)
);

BUFx2_ASAP7_75t_L g349 ( 
.A(n_343),
.Y(n_349)
);

OAI22xp5_ASAP7_75t_SL g360 ( 
.A1(n_344),
.A2(n_345),
.B1(n_312),
.B2(n_317),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_314),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_323),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_308),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_348),
.B(n_342),
.Y(n_372)
);

NOR3xp33_ASAP7_75t_SL g350 ( 
.A(n_329),
.B(n_313),
.C(n_326),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_SL g374 ( 
.A(n_350),
.B(n_353),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_352),
.B(n_356),
.Y(n_379)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_354),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g356 ( 
.A(n_327),
.B(n_310),
.C(n_304),
.Y(n_356)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_357),
.Y(n_373)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_327),
.B(n_325),
.C(n_320),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_358),
.B(n_364),
.C(n_340),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_360),
.B(n_344),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g364 ( 
.A(n_330),
.B(n_305),
.C(n_318),
.Y(n_364)
);

AOI21xp5_ASAP7_75t_L g366 ( 
.A1(n_363),
.A2(n_332),
.B(n_331),
.Y(n_366)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_366),
.Y(n_386)
);

OAI21xp5_ASAP7_75t_SL g367 ( 
.A1(n_362),
.A2(n_338),
.B(n_328),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_367),
.B(n_370),
.Y(n_381)
);

AOI21xp5_ASAP7_75t_SL g368 ( 
.A1(n_363),
.A2(n_318),
.B(n_334),
.Y(n_368)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_368),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_369),
.B(n_358),
.C(n_364),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_361),
.B(n_336),
.C(n_340),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_371),
.A2(n_360),
.B1(n_347),
.B2(n_351),
.Y(n_385)
);

OAI221xp5_ASAP7_75t_L g384 ( 
.A1(n_372),
.A2(n_347),
.B1(n_348),
.B2(n_351),
.C(n_352),
.Y(n_384)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_374),
.Y(n_391)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_350),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_375),
.B(n_359),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g376 ( 
.A1(n_362),
.A2(n_335),
.B(n_346),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_355),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g377 ( 
.A(n_361),
.B(n_333),
.C(n_341),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g387 ( 
.A(n_377),
.B(n_378),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g378 ( 
.A(n_356),
.B(n_345),
.C(n_343),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g399 ( 
.A(n_380),
.B(n_384),
.Y(n_399)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_382),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g398 ( 
.A1(n_383),
.A2(n_376),
.B1(n_371),
.B2(n_366),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_385),
.B(n_389),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_379),
.B(n_349),
.C(n_9),
.Y(n_389)
);

AND2x2_ASAP7_75t_L g390 ( 
.A(n_378),
.B(n_349),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g393 ( 
.A1(n_390),
.A2(n_392),
.B(n_365),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_370),
.C(n_369),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_393),
.B(n_395),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g395 ( 
.A(n_392),
.B(n_368),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_SL g396 ( 
.A(n_383),
.B(n_373),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_396),
.B(n_401),
.Y(n_407)
);

XNOR2x1_ASAP7_75t_L g408 ( 
.A(n_398),
.B(n_8),
.Y(n_408)
);

A2O1A1Ixp33_ASAP7_75t_SL g400 ( 
.A1(n_388),
.A2(n_367),
.B(n_10),
.C(n_11),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g410 ( 
.A1(n_400),
.A2(n_394),
.B(n_397),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g401 ( 
.A(n_391),
.B(n_8),
.Y(n_401)
);

AOI22xp33_ASAP7_75t_SL g402 ( 
.A1(n_386),
.A2(n_8),
.B1(n_10),
.B2(n_11),
.Y(n_402)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_402),
.A2(n_390),
.B(n_10),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_387),
.B(n_17),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g409 ( 
.A(n_403),
.B(n_10),
.Y(n_409)
);

OAI21xp5_ASAP7_75t_SL g404 ( 
.A1(n_399),
.A2(n_381),
.B(n_382),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g413 ( 
.A1(n_404),
.A2(n_411),
.B(n_12),
.Y(n_413)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_406),
.Y(n_414)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_408),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_409),
.B(n_400),
.C(n_405),
.Y(n_412)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_410),
.A2(n_407),
.B(n_13),
.Y(n_415)
);

AOI21xp33_ASAP7_75t_L g411 ( 
.A1(n_400),
.A2(n_12),
.B(n_13),
.Y(n_411)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_412),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_413),
.B(n_415),
.Y(n_419)
);

OAI321xp33_ASAP7_75t_L g417 ( 
.A1(n_414),
.A2(n_410),
.A3(n_14),
.B1(n_15),
.B2(n_17),
.C(n_12),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_417),
.B(n_14),
.Y(n_421)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_418),
.A2(n_416),
.B(n_14),
.Y(n_420)
);

OAI31xp33_ASAP7_75t_L g422 ( 
.A1(n_420),
.A2(n_421),
.A3(n_419),
.B(n_14),
.Y(n_422)
);

MAJIxp5_ASAP7_75t_L g423 ( 
.A(n_422),
.B(n_15),
.C(n_258),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_423),
.B(n_15),
.Y(n_424)
);


endmodule