module real_jpeg_4166_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_470;
wire n_219;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_323;
wire n_215;
wire n_166;
wire n_176;
wire n_286;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_450;
wire n_333;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_477;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_324;
wire n_261;
wire n_86;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_0),
.A2(n_40),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_0),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g294 ( 
.A1(n_0),
.A2(n_258),
.B1(n_295),
.B2(n_296),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_SL g349 ( 
.A1(n_0),
.A2(n_115),
.B1(n_258),
.B2(n_350),
.Y(n_349)
);

AOI22xp33_ASAP7_75t_L g442 ( 
.A1(n_0),
.A2(n_92),
.B1(n_258),
.B2(n_443),
.Y(n_442)
);

AOI22xp33_ASAP7_75t_SL g281 ( 
.A1(n_1),
.A2(n_83),
.B1(n_179),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_1),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_1),
.B(n_289),
.C(n_290),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_1),
.B(n_79),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_1),
.B(n_161),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_1),
.B(n_128),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g359 ( 
.A(n_1),
.B(n_360),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_38),
.B1(n_193),
.B2(n_194),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_2),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_2),
.A2(n_116),
.B1(n_193),
.B2(n_285),
.Y(n_284)
);

AOI22xp33_ASAP7_75t_L g302 ( 
.A1(n_2),
.A2(n_124),
.B1(n_162),
.B2(n_193),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_2),
.A2(n_193),
.B1(n_365),
.B2(n_367),
.Y(n_364)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_3),
.Y(n_161)
);

BUFx5_ASAP7_75t_L g165 ( 
.A(n_3),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_3),
.Y(n_241)
);

INVx8_ASAP7_75t_L g338 ( 
.A(n_3),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g19 ( 
.A1(n_4),
.A2(n_20),
.B1(n_23),
.B2(n_24),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_5),
.Y(n_40)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_5),
.Y(n_63)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_5),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_5),
.Y(n_190)
);

INVx6_ASAP7_75t_L g260 ( 
.A(n_5),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_6),
.A2(n_77),
.B1(n_92),
.B2(n_94),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_6),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_6),
.A2(n_62),
.B1(n_94),
.B2(n_137),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g182 ( 
.A1(n_6),
.A2(n_94),
.B1(n_109),
.B2(n_183),
.Y(n_182)
);

OAI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_6),
.A2(n_94),
.B1(n_232),
.B2(n_236),
.Y(n_231)
);

INVx3_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_7),
.Y(n_46)
);

BUFx5_ASAP7_75t_L g418 ( 
.A(n_7),
.Y(n_418)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_9),
.A2(n_179),
.B1(n_307),
.B2(n_309),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_9),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_9),
.A2(n_309),
.B1(n_323),
.B2(n_324),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g397 ( 
.A1(n_9),
.A2(n_309),
.B1(n_398),
.B2(n_399),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_9),
.A2(n_37),
.B1(n_309),
.B2(n_471),
.Y(n_470)
);

AOI22xp33_ASAP7_75t_SL g60 ( 
.A1(n_10),
.A2(n_37),
.B1(n_61),
.B2(n_64),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_10),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_10),
.A2(n_64),
.B1(n_175),
.B2(n_178),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_10),
.A2(n_64),
.B1(n_206),
.B2(n_208),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_L g428 ( 
.A1(n_10),
.A2(n_64),
.B1(n_296),
.B2(n_317),
.Y(n_428)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_11),
.Y(n_112)
);

BUFx5_ASAP7_75t_L g114 ( 
.A(n_11),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_11),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g53 ( 
.A1(n_12),
.A2(n_39),
.B1(n_54),
.B2(n_57),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g201 ( 
.A1(n_12),
.A2(n_57),
.B1(n_93),
.B2(n_202),
.Y(n_201)
);

OAI22xp33_ASAP7_75t_SL g243 ( 
.A1(n_12),
.A2(n_57),
.B1(n_244),
.B2(n_245),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_12),
.A2(n_57),
.B1(n_167),
.B2(n_296),
.Y(n_405)
);

INVx8_ASAP7_75t_L g85 ( 
.A(n_13),
.Y(n_85)
);

OAI22xp33_ASAP7_75t_L g187 ( 
.A1(n_14),
.A2(n_39),
.B1(n_188),
.B2(n_189),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_14),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_14),
.A2(n_188),
.B1(n_250),
.B2(n_254),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_14),
.A2(n_188),
.B1(n_236),
.B2(n_372),
.Y(n_371)
);

AOI22xp33_ASAP7_75t_SL g446 ( 
.A1(n_14),
.A2(n_188),
.B1(n_447),
.B2(n_450),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_15),
.Y(n_123)
);

BUFx3_ASAP7_75t_L g170 ( 
.A(n_15),
.Y(n_170)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_15),
.Y(n_235)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_16),
.Y(n_69)
);

INVx8_ASAP7_75t_L g50 ( 
.A(n_17),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_18),
.A2(n_97),
.B1(n_99),
.B2(n_102),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_18),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_18),
.A2(n_102),
.B1(n_130),
.B2(n_132),
.Y(n_129)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_18),
.A2(n_102),
.B1(n_147),
.B2(n_148),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_18),
.A2(n_102),
.B1(n_167),
.B2(n_171),
.Y(n_166)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_21),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

INVx8_ASAP7_75t_L g23 ( 
.A(n_22),
.Y(n_23)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_527),
.B(n_530),
.Y(n_24)
);

AO21x1_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_149),
.B(n_526),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g26 ( 
.A(n_27),
.B(n_145),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_L g526 ( 
.A(n_27),
.B(n_145),
.Y(n_526)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_135),
.C(n_142),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g521 ( 
.A1(n_28),
.A2(n_29),
.B1(n_522),
.B2(n_523),
.Y(n_521)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

MAJIxp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_65),
.C(n_103),
.Y(n_29)
);

XNOR2xp5_ASAP7_75t_SL g269 ( 
.A(n_30),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g30 ( 
.A1(n_31),
.A2(n_53),
.B1(n_58),
.B2(n_60),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_31),
.A2(n_58),
.B1(n_60),
.B2(n_136),
.Y(n_135)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_31),
.A2(n_58),
.B1(n_136),
.B2(n_146),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_SL g212 ( 
.A1(n_31),
.A2(n_53),
.B1(n_58),
.B2(n_213),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_31),
.A2(n_257),
.B(n_261),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_31),
.A2(n_58),
.B1(n_257),
.B2(n_470),
.Y(n_469)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_32),
.B(n_192),
.Y(n_191)
);

AOI21xp5_ASAP7_75t_L g434 ( 
.A1(n_32),
.A2(n_435),
.B(n_439),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g528 ( 
.A1(n_32),
.A2(n_59),
.B(n_529),
.Y(n_528)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_43),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g33 ( 
.A1(n_34),
.A2(n_37),
.B1(n_39),
.B2(n_41),
.Y(n_33)
);

INVx6_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_L g43 ( 
.A1(n_36),
.A2(n_44),
.B1(n_47),
.B2(n_51),
.Y(n_43)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx8_ASAP7_75t_L g147 ( 
.A(n_38),
.Y(n_147)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_43),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_45),
.B(n_356),
.Y(n_419)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g366 ( 
.A(n_48),
.Y(n_366)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_49),
.Y(n_362)
);

BUFx5_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_50),
.Y(n_52)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_50),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_50),
.Y(n_98)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_50),
.Y(n_357)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_52),
.Y(n_101)
);

INVx3_ASAP7_75t_L g204 ( 
.A(n_52),
.Y(n_204)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_52),
.Y(n_444)
);

INVx2_ASAP7_75t_SL g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g403 ( 
.A(n_58),
.B(n_282),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_L g487 ( 
.A1(n_58),
.A2(n_191),
.B(n_470),
.Y(n_487)
);

INVx1_ASAP7_75t_SL g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_59),
.B(n_187),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_59),
.B(n_192),
.Y(n_261)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_62),
.Y(n_61)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

BUFx3_ASAP7_75t_L g195 ( 
.A(n_63),
.Y(n_195)
);

INVx2_ASAP7_75t_L g472 ( 
.A(n_63),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_65),
.A2(n_103),
.B1(n_104),
.B2(n_271),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_65),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_91),
.B1(n_95),
.B2(n_96),
.Y(n_65)
);

INVx2_ASAP7_75t_SL g143 ( 
.A(n_66),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_66),
.A2(n_91),
.B1(n_95),
.B2(n_217),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_66),
.A2(n_95),
.B1(n_201),
.B2(n_249),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_66),
.A2(n_95),
.B1(n_397),
.B2(n_442),
.Y(n_441)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_67),
.B(n_79),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_68),
.A2(n_70),
.B1(n_73),
.B2(n_77),
.Y(n_67)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_69),
.Y(n_76)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_69),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_72),
.Y(n_209)
);

BUFx6f_ASAP7_75t_L g253 ( 
.A(n_72),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_72),
.Y(n_255)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx2_ASAP7_75t_L g399 ( 
.A(n_77),
.Y(n_399)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_79),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_79),
.A2(n_143),
.B(n_144),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_79),
.A2(n_143),
.B1(n_200),
.B2(n_205),
.Y(n_199)
);

AOI22x1_ASAP7_75t_L g473 ( 
.A1(n_79),
.A2(n_143),
.B1(n_401),
.B2(n_474),
.Y(n_473)
);

AO22x2_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_83),
.B1(n_86),
.B2(n_89),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_82),
.Y(n_90)
);

INVx4_ASAP7_75t_L g380 ( 
.A(n_82),
.Y(n_380)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_84),
.Y(n_116)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_85),
.Y(n_247)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_85),
.Y(n_285)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_85),
.Y(n_383)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_88),
.Y(n_109)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_88),
.Y(n_131)
);

INVx6_ASAP7_75t_L g181 ( 
.A(n_88),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g452 ( 
.A(n_88),
.Y(n_452)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

INVx6_ASAP7_75t_SL g92 ( 
.A(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_95),
.B(n_364),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g396 ( 
.A1(n_95),
.A2(n_397),
.B(n_400),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g144 ( 
.A(n_96),
.Y(n_144)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_98),
.Y(n_97)
);

INVx4_ASAP7_75t_L g207 ( 
.A(n_98),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g367 ( 
.A(n_98),
.Y(n_367)
);

INVx1_ASAP7_75t_SL g398 ( 
.A(n_99),
.Y(n_398)
);

INVx5_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g214 ( 
.A1(n_103),
.A2(n_104),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_103),
.B(n_212),
.C(n_215),
.Y(n_265)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_105),
.A2(n_127),
.B(n_129),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_SL g280 ( 
.A1(n_105),
.A2(n_281),
.B(n_283),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g348 ( 
.A1(n_105),
.A2(n_127),
.B1(n_306),
.B2(n_349),
.Y(n_348)
);

OAI21xp5_ASAP7_75t_SL g393 ( 
.A1(n_105),
.A2(n_283),
.B(n_349),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_105),
.A2(n_127),
.B1(n_446),
.B2(n_465),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_106),
.A2(n_128),
.B1(n_174),
.B2(n_182),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_106),
.A2(n_128),
.B1(n_182),
.B2(n_198),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_106),
.A2(n_128),
.B1(n_174),
.B2(n_243),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_106),
.B(n_284),
.Y(n_310)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_117),
.Y(n_106)
);

OAI22xp33_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_110),
.B1(n_113),
.B2(n_115),
.Y(n_107)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_109),
.B(n_288),
.Y(n_287)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx4_ASAP7_75t_L g289 ( 
.A(n_112),
.Y(n_289)
);

INVx4_ASAP7_75t_SL g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_114),
.Y(n_126)
);

INVx5_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_117),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g305 ( 
.A1(n_117),
.A2(n_306),
.B(n_310),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_120),
.B1(n_124),
.B2(n_126),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_123),
.Y(n_125)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_123),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g372 ( 
.A(n_123),
.Y(n_372)
);

INVx6_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g445 ( 
.A1(n_127),
.A2(n_310),
.B(n_446),
.Y(n_445)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_128),
.B(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx5_ASAP7_75t_L g177 ( 
.A(n_131),
.Y(n_177)
);

INVx1_ASAP7_75t_SL g132 ( 
.A(n_133),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_134),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g523 ( 
.A(n_135),
.B(n_142),
.Y(n_523)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx3_ASAP7_75t_L g415 ( 
.A(n_140),
.Y(n_415)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

INVx2_ASAP7_75t_L g438 ( 
.A(n_141),
.Y(n_438)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_143),
.A2(n_354),
.B(n_363),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_143),
.B(n_401),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_L g489 ( 
.A1(n_143),
.A2(n_363),
.B(n_490),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g527 ( 
.A(n_145),
.B(n_528),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_145),
.B(n_528),
.Y(n_531)
);

CKINVDCx20_ASAP7_75t_R g529 ( 
.A(n_146),
.Y(n_529)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_147),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_148),
.B(n_282),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_150),
.A2(n_520),
.B(n_525),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_273),
.B(n_517),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_262),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_153),
.B(n_219),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_153),
.B(n_219),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g532 ( 
.A(n_153),
.Y(n_532)
);

FAx1_ASAP7_75t_SL g153 ( 
.A(n_154),
.B(n_196),
.CI(n_210),
.CON(n_153),
.SN(n_153)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_154),
.B(n_196),
.C(n_210),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_155),
.A2(n_156),
.B(n_185),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_L g221 ( 
.A(n_155),
.B(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_173),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_156),
.A2(n_185),
.B1(n_223),
.B2(n_224),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_156),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g460 ( 
.A1(n_156),
.A2(n_173),
.B1(n_224),
.B2(n_461),
.Y(n_460)
);

OAI21xp5_ASAP7_75t_SL g156 ( 
.A1(n_157),
.A2(n_165),
.B(n_166),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_157),
.A2(n_166),
.B1(n_231),
.B2(n_239),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_157),
.A2(n_294),
.B(n_299),
.Y(n_293)
);

AOI21xp5_ASAP7_75t_L g319 ( 
.A1(n_157),
.A2(n_282),
.B(n_299),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g422 ( 
.A1(n_157),
.A2(n_423),
.B1(n_424),
.B2(n_427),
.Y(n_422)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_158),
.B(n_302),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g332 ( 
.A1(n_158),
.A2(n_333),
.B1(n_334),
.B2(n_335),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_158),
.A2(n_160),
.B1(n_371),
.B2(n_405),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g466 ( 
.A1(n_158),
.A2(n_300),
.B1(n_428),
.B2(n_467),
.Y(n_466)
);

OR2x2_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_162),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_161),
.Y(n_301)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx14_ASAP7_75t_R g167 ( 
.A(n_168),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_169),
.Y(n_168)
);

BUFx2_ASAP7_75t_L g295 ( 
.A(n_169),
.Y(n_295)
);

BUFx5_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

BUFx8_ASAP7_75t_L g172 ( 
.A(n_170),
.Y(n_172)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_170),
.Y(n_327)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_171),
.Y(n_317)
);

INVx8_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g461 ( 
.A(n_173),
.Y(n_461)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

AOI32xp33_ASAP7_75t_L g373 ( 
.A1(n_176),
.A2(n_359),
.A3(n_374),
.B1(n_378),
.B2(n_381),
.Y(n_373)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_177),
.Y(n_308)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

BUFx2_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx8_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

BUFx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_185),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_191),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_187),
.Y(n_213)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_196),
.A2(n_226),
.B(n_227),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g227 ( 
.A(n_197),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g226 ( 
.A(n_199),
.Y(n_226)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

OAI32xp33_ASAP7_75t_L g414 ( 
.A1(n_202),
.A2(n_415),
.A3(n_416),
.B1(n_419),
.B2(n_420),
.Y(n_414)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

INVx2_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_205),
.Y(n_217)
);

INVx6_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx3_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_214),
.B2(n_218),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_211),
.A2(n_212),
.B1(n_268),
.B2(n_269),
.Y(n_267)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_211),
.B(n_264),
.C(n_268),
.Y(n_524)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_214),
.Y(n_218)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_225),
.C(n_228),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_220),
.A2(n_221),
.B1(n_225),
.B2(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_225),
.Y(n_477)
);

XNOR2xp5_ASAP7_75t_L g475 ( 
.A(n_228),
.B(n_476),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_248),
.C(n_256),
.Y(n_228)
);

XNOR2xp5_ASAP7_75t_L g458 ( 
.A(n_229),
.B(n_459),
.Y(n_458)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_242),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_230),
.B(n_242),
.Y(n_484)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_231),
.Y(n_467)
);

INVx4_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

BUFx3_ASAP7_75t_L g234 ( 
.A(n_235),
.Y(n_234)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g291 ( 
.A(n_235),
.Y(n_291)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

INVx4_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g321 ( 
.A1(n_239),
.A2(n_322),
.B(n_328),
.Y(n_321)
);

INVx4_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

INVx4_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_243),
.Y(n_465)
);

BUFx2_ASAP7_75t_L g351 ( 
.A(n_244),
.Y(n_351)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

BUFx3_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx4_ASAP7_75t_L g449 ( 
.A(n_247),
.Y(n_449)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_248),
.B(n_256),
.Y(n_459)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_249),
.Y(n_474)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_251),
.Y(n_250)
);

INVx5_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx5_ASAP7_75t_L g377 ( 
.A(n_255),
.Y(n_377)
);

INVx8_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_261),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_262),
.A2(n_518),
.B(n_519),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_263),
.B(n_272),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_263),
.B(n_272),
.Y(n_519)
);

OAI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_269),
.Y(n_268)
);

OAI311xp33_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_455),
.A3(n_493),
.B1(n_511),
.C1(n_512),
.Y(n_273)
);

AOI21x1_ASAP7_75t_L g274 ( 
.A1(n_275),
.A2(n_408),
.B(n_454),
.Y(n_274)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_276),
.A2(n_388),
.B(n_407),
.Y(n_275)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_277),
.A2(n_343),
.B(n_387),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_313),
.B(n_342),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_279),
.B(n_292),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_279),
.B(n_292),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_280),
.B(n_286),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_280),
.A2(n_286),
.B1(n_287),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_280),
.Y(n_340)
);

OAI21xp33_ASAP7_75t_SL g354 ( 
.A1(n_282),
.A2(n_355),
.B(n_358),
.Y(n_354)
);

OAI21xp33_ASAP7_75t_SL g435 ( 
.A1(n_282),
.A2(n_420),
.B(n_436),
.Y(n_435)
);

CKINVDCx16_ASAP7_75t_R g286 ( 
.A(n_287),
.Y(n_286)
);

INVx2_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_291),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_303),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_293),
.B(n_304),
.C(n_312),
.Y(n_344)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_294),
.Y(n_334)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_297),
.Y(n_296)
);

INVx6_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_300),
.B(n_302),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g369 ( 
.A1(n_301),
.A2(n_328),
.B(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_304),
.A2(n_305),
.B1(n_311),
.B2(n_312),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_305),
.Y(n_304)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.Y(n_307)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_331),
.B(n_341),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g314 ( 
.A1(n_315),
.A2(n_320),
.B(n_330),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_319),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_321),
.B(n_329),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_321),
.B(n_329),
.Y(n_330)
);

INVxp67_ASAP7_75t_L g333 ( 
.A(n_322),
.Y(n_333)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_339),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_332),
.B(n_339),
.Y(n_341)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx8_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_344),
.B(n_345),
.Y(n_387)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_368),
.Y(n_345)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_347),
.A2(n_348),
.B1(n_352),
.B2(n_353),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_348),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g389 ( 
.A(n_348),
.B(n_352),
.C(n_368),
.Y(n_389)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_351),
.Y(n_350)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_353),
.Y(n_352)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_359),
.Y(n_358)
);

INVx2_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx4_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

INVx3_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

XOR2xp5_ASAP7_75t_L g368 ( 
.A(n_369),
.B(n_373),
.Y(n_368)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_369),
.B(n_373),
.Y(n_394)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_371),
.Y(n_370)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_375),
.Y(n_374)
);

INVx3_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

INVx6_ASAP7_75t_L g376 ( 
.A(n_377),
.Y(n_376)
);

INVx4_ASAP7_75t_L g378 ( 
.A(n_379),
.Y(n_378)
);

INVx8_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

INVx6_ASAP7_75t_L g386 ( 
.A(n_380),
.Y(n_386)
);

NAND2xp33_ASAP7_75t_SL g381 ( 
.A(n_382),
.B(n_384),
.Y(n_381)
);

INVx5_ASAP7_75t_L g382 ( 
.A(n_383),
.Y(n_382)
);

INVx2_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx3_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_390),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_SL g407 ( 
.A(n_389),
.B(n_390),
.Y(n_407)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_391),
.A2(n_392),
.B1(n_395),
.B2(n_406),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_392),
.Y(n_391)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_393),
.B(n_394),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_394),
.C(n_406),
.Y(n_409)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_395),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_402),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_396),
.B(n_403),
.C(n_404),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_404),
.Y(n_402)
);

INVxp67_ASAP7_75t_L g423 ( 
.A(n_405),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_410),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g454 ( 
.A(n_409),
.B(n_410),
.Y(n_454)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_432),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g411 ( 
.A1(n_412),
.A2(n_429),
.B1(n_430),
.B2(n_431),
.Y(n_411)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_412),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_413),
.A2(n_414),
.B1(n_421),
.B2(n_422),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_414),
.Y(n_413)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_414),
.B(n_421),
.Y(n_488)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_417),
.Y(n_416)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_426),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_428),
.Y(n_427)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_429),
.Y(n_431)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_429),
.B(n_430),
.C(n_432),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g432 ( 
.A1(n_433),
.A2(n_434),
.B1(n_440),
.B2(n_453),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_433),
.B(n_441),
.C(n_445),
.Y(n_502)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_434),
.Y(n_433)
);

INVx3_ASAP7_75t_L g436 ( 
.A(n_437),
.Y(n_436)
);

INVx4_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_440),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_441),
.B(n_445),
.Y(n_440)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_442),
.Y(n_490)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_444),
.Y(n_443)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_449),
.Y(n_448)
);

INVx2_ASAP7_75t_L g450 ( 
.A(n_451),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

NAND2xp33_ASAP7_75t_SL g455 ( 
.A(n_456),
.B(n_478),
.Y(n_455)
);

A2O1A1Ixp33_ASAP7_75t_SL g512 ( 
.A1(n_456),
.A2(n_478),
.B(n_513),
.C(n_516),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g456 ( 
.A(n_457),
.B(n_475),
.Y(n_456)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_457),
.B(n_475),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_460),
.C(n_462),
.Y(n_457)
);

XNOR2xp5_ASAP7_75t_L g492 ( 
.A(n_458),
.B(n_460),
.Y(n_492)
);

XOR2xp5_ASAP7_75t_L g491 ( 
.A(n_462),
.B(n_492),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g462 ( 
.A(n_463),
.B(n_468),
.C(n_473),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_463),
.B(n_482),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g463 ( 
.A(n_464),
.B(n_466),
.Y(n_463)
);

XOR2xp5_ASAP7_75t_L g501 ( 
.A(n_464),
.B(n_466),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_SL g482 ( 
.A1(n_468),
.A2(n_469),
.B1(n_473),
.B2(n_483),
.Y(n_482)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_472),
.Y(n_471)
);

INVx1_ASAP7_75t_SL g483 ( 
.A(n_473),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g478 ( 
.A(n_479),
.B(n_491),
.Y(n_478)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_479),
.B(n_491),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_480),
.B(n_484),
.C(n_485),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_SL g504 ( 
.A1(n_480),
.A2(n_481),
.B1(n_484),
.B2(n_505),
.Y(n_504)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_484),
.Y(n_505)
);

XNOR2xp5_ASAP7_75t_L g503 ( 
.A(n_485),
.B(n_504),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_486),
.B(n_488),
.C(n_489),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g498 ( 
.A1(n_486),
.A2(n_487),
.B1(n_489),
.B2(n_499),
.Y(n_498)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_487),
.Y(n_486)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_488),
.B(n_498),
.Y(n_497)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_489),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g493 ( 
.A(n_494),
.B(n_506),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_495),
.Y(n_494)
);

OAI21xp5_ASAP7_75t_L g513 ( 
.A1(n_495),
.A2(n_514),
.B(n_515),
.Y(n_513)
);

NOR2x1_ASAP7_75t_L g495 ( 
.A(n_496),
.B(n_503),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_496),
.B(n_503),
.Y(n_515)
);

MAJIxp5_ASAP7_75t_L g496 ( 
.A(n_497),
.B(n_500),
.C(n_502),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g508 ( 
.A(n_497),
.B(n_509),
.Y(n_508)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_500),
.A2(n_501),
.B1(n_502),
.B2(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_501),
.Y(n_500)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_502),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_507),
.B(n_508),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_L g514 ( 
.A(n_507),
.B(n_508),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g520 ( 
.A(n_521),
.B(n_524),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_521),
.B(n_524),
.Y(n_525)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_523),
.Y(n_522)
);

INVxp67_ASAP7_75t_L g530 ( 
.A(n_531),
.Y(n_530)
);


endmodule