module fake_jpeg_21787_n_338 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_338);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_338;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_8),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx12_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_3),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVxp67_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_10),
.B(n_16),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

BUFx5_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_19),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_36),
.B(n_31),
.Y(n_68)
);

AND2x6_ASAP7_75t_L g37 ( 
.A(n_32),
.B(n_0),
.Y(n_37)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_37),
.B(n_26),
.C(n_22),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_38),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_22),
.B(n_0),
.Y(n_39)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_39),
.B(n_45),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_20),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_40),
.B(n_43),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

CKINVDCx6p67_ASAP7_75t_R g59 ( 
.A(n_41),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_33),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_44),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_22),
.B(n_0),
.Y(n_45)
);

INVx13_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

INVx11_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_46),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_48),
.A2(n_52),
.B1(n_63),
.B2(n_36),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_39),
.B(n_27),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_49),
.B(n_55),
.Y(n_81)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_61),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_46),
.A2(n_19),
.B1(n_24),
.B2(n_26),
.Y(n_52)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_53),
.A2(n_37),
.B(n_34),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_54),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_45),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

INVx3_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_38),
.Y(n_61)
);

BUFx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_62),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g63 ( 
.A1(n_46),
.A2(n_24),
.B1(n_27),
.B2(n_35),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_68),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_37),
.A2(n_35),
.B1(n_31),
.B2(n_25),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g95 ( 
.A1(n_65),
.A2(n_30),
.B1(n_25),
.B2(n_28),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_17),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_66),
.B(n_36),
.Y(n_71)
);

BUFx12f_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

CKINVDCx11_ASAP7_75t_R g82 ( 
.A(n_67),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_69),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_71),
.B(n_47),
.Y(n_108)
);

CKINVDCx12_ASAP7_75t_R g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_73),
.B(n_77),
.Y(n_101)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_66),
.B(n_55),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g116 ( 
.A1(n_74),
.A2(n_91),
.B(n_81),
.Y(n_116)
);

NAND2x1_ASAP7_75t_SL g76 ( 
.A(n_70),
.B(n_41),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_SL g114 ( 
.A(n_76),
.B(n_71),
.C(n_87),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_58),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_78),
.B(n_83),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_40),
.Y(n_79)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_79),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_70),
.B(n_43),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_40),
.Y(n_84)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_84),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_65),
.B(n_43),
.Y(n_85)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_85),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_86),
.A2(n_57),
.B1(n_59),
.B2(n_67),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_70),
.A2(n_37),
.B1(n_21),
.B2(n_29),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_87),
.A2(n_94),
.B1(n_50),
.B2(n_61),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_30),
.Y(n_89)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_89),
.Y(n_110)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_90),
.B(n_93),
.Y(n_123)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_57),
.A2(n_17),
.B1(n_18),
.B2(n_28),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_95),
.A2(n_18),
.B1(n_17),
.B2(n_28),
.Y(n_122)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_98),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_23),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g149 ( 
.A1(n_99),
.A2(n_113),
.B(n_114),
.Y(n_149)
);

NOR3xp33_ASAP7_75t_L g100 ( 
.A(n_91),
.B(n_67),
.C(n_62),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_100),
.B(n_103),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_102),
.A2(n_127),
.B1(n_98),
.B2(n_96),
.Y(n_141)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_80),
.Y(n_103)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_97),
.Y(n_105)
);

INVx6_ASAP7_75t_L g131 ( 
.A(n_105),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_SL g130 ( 
.A(n_108),
.B(n_75),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g109 ( 
.A(n_79),
.B(n_67),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_115),
.Y(n_134)
);

AND2x6_ASAP7_75t_L g111 ( 
.A(n_74),
.B(n_14),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_116),
.Y(n_157)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_80),
.Y(n_112)
);

HB1xp67_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_85),
.A2(n_64),
.B(n_44),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_81),
.B(n_69),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_72),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_117),
.Y(n_128)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_83),
.B(n_69),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_120),
.B(n_126),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_72),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_121),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g148 ( 
.A1(n_122),
.A2(n_94),
.B1(n_88),
.B2(n_92),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_23),
.Y(n_125)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_125),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_78),
.B(n_23),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_91),
.A2(n_42),
.B1(n_44),
.B2(n_17),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_130),
.B(n_140),
.Y(n_161)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_132),
.B(n_133),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

INVx1_ASAP7_75t_SL g136 ( 
.A(n_126),
.Y(n_136)
);

OA22x2_ASAP7_75t_L g159 ( 
.A1(n_136),
.A2(n_121),
.B1(n_82),
.B2(n_80),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_127),
.A2(n_95),
.B1(n_86),
.B2(n_76),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_138),
.A2(n_110),
.B1(n_101),
.B2(n_109),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_115),
.B(n_95),
.Y(n_140)
);

OAI21xp33_ASAP7_75t_SL g174 ( 
.A1(n_141),
.A2(n_148),
.B(n_102),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_116),
.B(n_76),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_143),
.B(n_150),
.Y(n_172)
);

OAI32xp33_ASAP7_75t_L g144 ( 
.A1(n_114),
.A2(n_76),
.A3(n_75),
.B1(n_84),
.B2(n_89),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_144),
.B(n_140),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_124),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_117),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_146),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_104),
.B(n_90),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_120),
.B(n_82),
.C(n_80),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_151),
.B(n_110),
.C(n_122),
.Y(n_176)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_108),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_152),
.B(n_153),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_104),
.B(n_56),
.Y(n_153)
);

AOI21xp33_ASAP7_75t_L g154 ( 
.A1(n_118),
.A2(n_16),
.B(n_10),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g166 ( 
.A(n_154),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_56),
.Y(n_155)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_155),
.Y(n_158)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_124),
.Y(n_156)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_156),
.Y(n_170)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_159),
.A2(n_171),
.B(n_182),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_L g163 ( 
.A1(n_143),
.A2(n_107),
.B(n_113),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_163),
.A2(n_168),
.B(n_169),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_147),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_147),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_165),
.B(n_173),
.Y(n_213)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_157),
.B(n_111),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_176),
.C(n_178),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g168 ( 
.A1(n_149),
.A2(n_107),
.B(n_113),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_149),
.A2(n_111),
.B(n_106),
.Y(n_169)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_142),
.A2(n_101),
.B(n_125),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_153),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_174),
.A2(n_180),
.B1(n_187),
.B2(n_141),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g177 ( 
.A(n_128),
.B(n_106),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_177),
.B(n_155),
.Y(n_208)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_150),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_SL g217 ( 
.A(n_179),
.B(n_181),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_128),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_137),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_142),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_183),
.B(n_186),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_134),
.A2(n_135),
.B(n_136),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g200 ( 
.A1(n_184),
.A2(n_189),
.B(n_130),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_134),
.A2(n_109),
.B1(n_93),
.B2(n_88),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_137),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_188),
.A2(n_97),
.B(n_105),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_135),
.A2(n_73),
.B(n_97),
.Y(n_189)
);

HB1xp67_ASAP7_75t_L g190 ( 
.A(n_164),
.Y(n_190)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_190),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_185),
.A2(n_148),
.B1(n_157),
.B2(n_146),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_191),
.A2(n_196),
.B1(n_210),
.B2(n_159),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_192),
.A2(n_159),
.B1(n_160),
.B2(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_194),
.B(n_195),
.Y(n_224)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_177),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_173),
.A2(n_156),
.B1(n_152),
.B2(n_132),
.Y(n_196)
);

INVx13_ASAP7_75t_L g197 ( 
.A(n_165),
.Y(n_197)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_197),
.Y(n_235)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_198),
.A2(n_203),
.B(n_205),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_200),
.A2(n_214),
.B(n_42),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_172),
.B(n_138),
.C(n_129),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_201),
.B(n_207),
.C(n_209),
.Y(n_219)
);

OR2x2_ASAP7_75t_L g202 ( 
.A(n_162),
.B(n_144),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_202),
.Y(n_227)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_175),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_187),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_184),
.C(n_178),
.Y(n_207)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_208),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_161),
.B(n_129),
.C(n_136),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g210 ( 
.A1(n_169),
.A2(n_112),
.B1(n_119),
.B2(n_103),
.Y(n_210)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_212),
.A2(n_139),
.B1(n_131),
.B2(n_92),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_139),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_215),
.A2(n_218),
.B1(n_179),
.B2(n_158),
.Y(n_223)
);

INVx13_ASAP7_75t_L g216 ( 
.A(n_162),
.Y(n_216)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_216),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g218 ( 
.A(n_180),
.B(n_97),
.Y(n_218)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_193),
.B(n_168),
.C(n_163),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_SL g262 ( 
.A(n_220),
.B(n_202),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_199),
.B(n_176),
.C(n_158),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_221),
.B(n_225),
.C(n_229),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_167),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_222),
.B(n_226),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g255 ( 
.A1(n_223),
.A2(n_230),
.B(n_238),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_207),
.B(n_171),
.C(n_160),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_193),
.B(n_159),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g265 ( 
.A(n_228),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_170),
.C(n_182),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_206),
.B(n_188),
.C(n_181),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_231),
.B(n_233),
.C(n_240),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_200),
.B(n_159),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_236),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_97),
.C(n_166),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_234),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_191),
.B(n_44),
.Y(n_236)
);

AOI322xp5_ASAP7_75t_L g237 ( 
.A1(n_218),
.A2(n_44),
.A3(n_42),
.B1(n_47),
.B2(n_51),
.C1(n_131),
.C2(n_88),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_237),
.B(n_244),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_209),
.B(n_42),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_192),
.A2(n_131),
.B1(n_92),
.B2(n_28),
.Y(n_243)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_51),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_216),
.Y(n_248)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_248),
.Y(n_278)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_251),
.B(n_254),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_221),
.B(n_215),
.C(n_214),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_253),
.C(n_240),
.Y(n_274)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_219),
.B(n_194),
.C(n_213),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

A2O1A1O1Ixp25_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_202),
.B(n_218),
.C(n_211),
.D(n_213),
.Y(n_257)
);

XOR2xp5_ASAP7_75t_L g272 ( 
.A(n_257),
.B(n_260),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_239),
.B(n_216),
.Y(n_258)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_235),
.B(n_217),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_259),
.B(n_263),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_219),
.B(n_210),
.Y(n_260)
);

BUFx12f_ASAP7_75t_SL g261 ( 
.A(n_244),
.Y(n_261)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_261),
.A2(n_242),
.B(n_229),
.Y(n_269)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_262),
.B(n_266),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_232),
.B(n_195),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_217),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_264),
.B(n_18),
.Y(n_283)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_261),
.Y(n_268)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_268),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_273),
.B(n_283),
.Y(n_288)
);

AOI22xp5_ASAP7_75t_L g270 ( 
.A1(n_265),
.A2(n_205),
.B1(n_227),
.B2(n_204),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g290 ( 
.A1(n_270),
.A2(n_263),
.B1(n_257),
.B2(n_255),
.Y(n_290)
);

OAI21xp5_ASAP7_75t_SL g273 ( 
.A1(n_267),
.A2(n_204),
.B(n_212),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_274),
.B(n_275),
.C(n_246),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_253),
.B(n_225),
.C(n_222),
.Y(n_275)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_252),
.A2(n_223),
.B1(n_236),
.B2(n_226),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_280),
.B1(n_281),
.B2(n_246),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_250),
.A2(n_198),
.B1(n_203),
.B2(n_245),
.Y(n_280)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_255),
.A2(n_197),
.B1(n_196),
.B2(n_208),
.Y(n_281)
);

FAx1_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_233),
.CI(n_197),
.CON(n_282),
.SN(n_282)
);

NAND2xp5_ASAP7_75t_SL g292 ( 
.A(n_282),
.B(n_266),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_284),
.B(n_256),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_283),
.B(n_279),
.Y(n_286)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_286),
.A2(n_291),
.B(n_292),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g287 ( 
.A(n_270),
.B(n_247),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g302 ( 
.A(n_287),
.B(n_290),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_295),
.Y(n_312)
);

INVxp67_ASAP7_75t_L g291 ( 
.A(n_277),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_277),
.B(n_260),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_293),
.B(n_294),
.Y(n_308)
);

NOR2x1_ASAP7_75t_SL g294 ( 
.A(n_269),
.B(n_256),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_281),
.B(n_247),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_296),
.B(n_285),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_SL g297 ( 
.A(n_271),
.B(n_249),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_SL g311 ( 
.A(n_297),
.B(n_293),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_249),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g309 ( 
.A1(n_298),
.A2(n_272),
.B(n_284),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g300 ( 
.A(n_299),
.B(n_274),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_300),
.B(n_304),
.Y(n_319)
);

HB1xp67_ASAP7_75t_L g301 ( 
.A(n_285),
.Y(n_301)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_301),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g303 ( 
.A1(n_288),
.A2(n_271),
.B(n_273),
.Y(n_303)
);

CKINVDCx20_ASAP7_75t_R g320 ( 
.A(n_303),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_SL g304 ( 
.A(n_295),
.B(n_272),
.Y(n_304)
);

INVxp67_ASAP7_75t_L g316 ( 
.A(n_305),
.Y(n_316)
);

XNOR2xp5_ASAP7_75t_L g307 ( 
.A(n_289),
.B(n_275),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_307),
.A2(n_309),
.B(n_311),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_291),
.B(n_282),
.Y(n_310)
);

OAI22xp5_ASAP7_75t_L g315 ( 
.A1(n_310),
.A2(n_51),
.B1(n_47),
.B2(n_14),
.Y(n_315)
);

AO21x1_ASAP7_75t_L g313 ( 
.A1(n_301),
.A2(n_276),
.B(n_282),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_313),
.B(n_314),
.Y(n_326)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_315),
.A2(n_318),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.C1(n_3),
.C2(n_4),
.Y(n_325)
);

OAI21xp5_ASAP7_75t_L g317 ( 
.A1(n_302),
.A2(n_18),
.B(n_15),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_317),
.B(n_1),
.C(n_2),
.Y(n_330)
);

FAx1_ASAP7_75t_SL g318 ( 
.A(n_308),
.B(n_15),
.CI(n_14),
.CON(n_318),
.SN(n_318)
);

INVxp33_ASAP7_75t_L g322 ( 
.A(n_308),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g324 ( 
.A1(n_322),
.A2(n_316),
.B(n_321),
.Y(n_324)
);

AOI322xp5_ASAP7_75t_L g323 ( 
.A1(n_320),
.A2(n_306),
.A3(n_312),
.B1(n_13),
.B2(n_12),
.C1(n_11),
.C2(n_5),
.Y(n_323)
);

AOI322xp5_ASAP7_75t_L g333 ( 
.A1(n_323),
.A2(n_325),
.A3(n_327),
.B1(n_328),
.B2(n_318),
.C1(n_5),
.C2(n_6),
.Y(n_333)
);

AOI21xp5_ASAP7_75t_L g331 ( 
.A1(n_324),
.A2(n_326),
.B(n_329),
.Y(n_331)
);

AOI322xp5_ASAP7_75t_L g327 ( 
.A1(n_322),
.A2(n_312),
.A3(n_13),
.B1(n_12),
.B2(n_11),
.C1(n_4),
.C2(n_5),
.Y(n_327)
);

AOI322xp5_ASAP7_75t_L g328 ( 
.A1(n_319),
.A2(n_0),
.A3(n_1),
.B1(n_2),
.B2(n_3),
.C1(n_4),
.C2(n_5),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_313),
.B(n_23),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_330),
.B(n_1),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

AOI321xp33_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_334),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_23),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_323),
.B(n_1),
.C(n_7),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g337 ( 
.A(n_335),
.B(n_331),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_336),
.C(n_8),
.Y(n_338)
);


endmodule