module fake_aes_6757_n_715 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_715);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_715;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_563;
wire n_540;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_648;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_235;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_420;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_195;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_606;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_44), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_49), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_71), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_39), .Y(n_83) );
CKINVDCx5p33_ASAP7_75t_R g84 ( .A(n_3), .Y(n_84) );
BUFx2_ASAP7_75t_L g85 ( .A(n_28), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_57), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_63), .Y(n_87) );
INVx1_ASAP7_75t_SL g88 ( .A(n_56), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_16), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_48), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_21), .Y(n_91) );
CKINVDCx16_ASAP7_75t_R g92 ( .A(n_15), .Y(n_92) );
INVxp33_ASAP7_75t_L g93 ( .A(n_62), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_19), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_64), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_34), .Y(n_96) );
INVxp33_ASAP7_75t_SL g97 ( .A(n_36), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_43), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_37), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_24), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_74), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_26), .Y(n_102) );
INVx1_ASAP7_75t_SL g103 ( .A(n_41), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_66), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_18), .Y(n_105) );
INVxp67_ASAP7_75t_L g106 ( .A(n_42), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_75), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_47), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_70), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_79), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_27), .Y(n_111) );
BUFx2_ASAP7_75t_SL g112 ( .A(n_33), .Y(n_112) );
INVxp67_ASAP7_75t_SL g113 ( .A(n_2), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_1), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_38), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_15), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_29), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_59), .Y(n_118) );
INVxp67_ASAP7_75t_L g119 ( .A(n_5), .Y(n_119) );
INVxp67_ASAP7_75t_SL g120 ( .A(n_51), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_54), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_30), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_18), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_16), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_23), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_46), .Y(n_126) );
INVxp67_ASAP7_75t_SL g127 ( .A(n_67), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_17), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_83), .Y(n_129) );
BUFx2_ASAP7_75t_SL g130 ( .A(n_85), .Y(n_130) );
INVx2_ASAP7_75t_L g131 ( .A(n_83), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
BUFx2_ASAP7_75t_L g133 ( .A(n_85), .Y(n_133) );
CKINVDCx20_ASAP7_75t_R g134 ( .A(n_92), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_86), .Y(n_135) );
BUFx6f_ASAP7_75t_L g136 ( .A(n_87), .Y(n_136) );
INVx1_ASAP7_75t_SL g137 ( .A(n_84), .Y(n_137) );
AND2x2_ASAP7_75t_L g138 ( .A(n_90), .B(n_0), .Y(n_138) );
CKINVDCx5p33_ASAP7_75t_R g139 ( .A(n_91), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_95), .Y(n_141) );
INVx3_ASAP7_75t_L g142 ( .A(n_95), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g143 ( .A(n_89), .B(n_0), .Y(n_143) );
CKINVDCx20_ASAP7_75t_R g144 ( .A(n_84), .Y(n_144) );
NOR2xp33_ASAP7_75t_R g145 ( .A(n_91), .B(n_31), .Y(n_145) );
CKINVDCx5p33_ASAP7_75t_R g146 ( .A(n_115), .Y(n_146) );
CKINVDCx5p33_ASAP7_75t_R g147 ( .A(n_115), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_96), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_97), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_97), .Y(n_150) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_89), .B(n_1), .Y(n_151) );
OAI22xp5_ASAP7_75t_L g152 ( .A1(n_105), .A2(n_2), .B1(n_3), .B2(n_4), .Y(n_152) );
BUFx3_ASAP7_75t_L g153 ( .A(n_96), .Y(n_153) );
AND2x2_ASAP7_75t_L g154 ( .A(n_93), .B(n_4), .Y(n_154) );
INVx3_ASAP7_75t_L g155 ( .A(n_99), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_94), .B(n_5), .Y(n_156) );
HB1xp67_ASAP7_75t_L g157 ( .A(n_105), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_99), .Y(n_158) );
HB1xp67_ASAP7_75t_L g159 ( .A(n_94), .Y(n_159) );
INVx3_ASAP7_75t_L g160 ( .A(n_100), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_112), .Y(n_161) );
NOR2xp33_ASAP7_75t_R g162 ( .A(n_80), .B(n_40), .Y(n_162) );
HB1xp67_ASAP7_75t_L g163 ( .A(n_124), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_100), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g165 ( .A(n_124), .B(n_6), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_108), .Y(n_166) );
BUFx3_ASAP7_75t_L g167 ( .A(n_108), .Y(n_167) );
CKINVDCx5p33_ASAP7_75t_R g168 ( .A(n_112), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_117), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_117), .Y(n_170) );
OR2x2_ASAP7_75t_L g171 ( .A(n_114), .B(n_6), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_88), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_116), .B(n_7), .Y(n_173) );
CKINVDCx5p33_ASAP7_75t_R g174 ( .A(n_98), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_142), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_136), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_136), .Y(n_177) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_157), .Y(n_178) );
NAND2xp5_ASAP7_75t_SL g179 ( .A(n_139), .B(n_104), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_136), .Y(n_180) );
INVx2_ASAP7_75t_L g181 ( .A(n_136), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_136), .Y(n_182) );
INVx1_ASAP7_75t_L g183 ( .A(n_142), .Y(n_183) );
BUFx6f_ASAP7_75t_L g184 ( .A(n_136), .Y(n_184) );
NOR2xp33_ASAP7_75t_L g185 ( .A(n_133), .B(n_106), .Y(n_185) );
INVx1_ASAP7_75t_L g186 ( .A(n_136), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_133), .B(n_128), .Y(n_187) );
AND2x2_ASAP7_75t_L g188 ( .A(n_130), .B(n_119), .Y(n_188) );
BUFx6f_ASAP7_75t_L g189 ( .A(n_170), .Y(n_189) );
INVx1_ASAP7_75t_L g190 ( .A(n_170), .Y(n_190) );
BUFx6f_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
OR2x2_ASAP7_75t_L g192 ( .A(n_130), .B(n_113), .Y(n_192) );
BUFx2_ASAP7_75t_L g193 ( .A(n_157), .Y(n_193) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_149), .B(n_111), .Y(n_194) );
INVx2_ASAP7_75t_L g195 ( .A(n_170), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_159), .B(n_123), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_170), .Y(n_197) );
INVx4_ASAP7_75t_L g198 ( .A(n_142), .Y(n_198) );
INVx8_ASAP7_75t_L g199 ( .A(n_161), .Y(n_199) );
AO22x2_ASAP7_75t_L g200 ( .A1(n_152), .A2(n_125), .B1(n_126), .B2(n_110), .Y(n_200) );
INVx1_ASAP7_75t_L g201 ( .A(n_142), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_138), .B(n_109), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_170), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_148), .Y(n_204) );
BUFx6f_ASAP7_75t_L g205 ( .A(n_170), .Y(n_205) );
NOR2xp33_ASAP7_75t_L g206 ( .A(n_150), .B(n_118), .Y(n_206) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_138), .B(n_107), .Y(n_207) );
BUFx6f_ASAP7_75t_L g208 ( .A(n_153), .Y(n_208) );
INVx2_ASAP7_75t_SL g209 ( .A(n_153), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_148), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_148), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_137), .B(n_125), .Y(n_212) );
INVx4_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
BUFx6f_ASAP7_75t_L g214 ( .A(n_153), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_155), .Y(n_215) );
NOR2xp33_ASAP7_75t_L g216 ( .A(n_168), .B(n_81), .Y(n_216) );
NOR2xp33_ASAP7_75t_L g217 ( .A(n_146), .B(n_82), .Y(n_217) );
INVx4_ASAP7_75t_L g218 ( .A(n_155), .Y(n_218) );
AOI22xp33_ASAP7_75t_L g219 ( .A1(n_159), .A2(n_126), .B1(n_101), .B2(n_122), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_129), .Y(n_220) );
NAND2xp5_ASAP7_75t_SL g221 ( .A(n_147), .B(n_172), .Y(n_221) );
INVx4_ASAP7_75t_L g222 ( .A(n_155), .Y(n_222) );
NAND2xp5_ASAP7_75t_L g223 ( .A(n_138), .B(n_121), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_154), .B(n_102), .Y(n_224) );
AND2x2_ASAP7_75t_L g225 ( .A(n_163), .B(n_127), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_155), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_129), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_160), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_163), .B(n_120), .Y(n_229) );
AND2x4_ASAP7_75t_L g230 ( .A(n_132), .B(n_103), .Y(n_230) );
BUFx6f_ASAP7_75t_L g231 ( .A(n_167), .Y(n_231) );
CKINVDCx5p33_ASAP7_75t_R g232 ( .A(n_144), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_129), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_174), .B(n_45), .Y(n_234) );
HB1xp67_ASAP7_75t_L g235 ( .A(n_193), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_198), .Y(n_236) );
AND2x4_ASAP7_75t_L g237 ( .A(n_230), .B(n_154), .Y(n_237) );
INVx1_ASAP7_75t_SL g238 ( .A(n_193), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_230), .B(n_154), .Y(n_239) );
BUFx6f_ASAP7_75t_L g240 ( .A(n_208), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_230), .B(n_137), .Y(n_241) );
NOR2x1_ASAP7_75t_L g242 ( .A(n_221), .B(n_171), .Y(n_242) );
BUFx8_ASAP7_75t_L g243 ( .A(n_187), .Y(n_243) );
BUFx4f_ASAP7_75t_SL g244 ( .A(n_187), .Y(n_244) );
INVxp67_ASAP7_75t_SL g245 ( .A(n_198), .Y(n_245) );
INVx2_ASAP7_75t_L g246 ( .A(n_198), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_196), .B(n_171), .Y(n_247) );
AND2x2_ASAP7_75t_L g248 ( .A(n_187), .B(n_134), .Y(n_248) );
INVx2_ASAP7_75t_L g249 ( .A(n_213), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_213), .Y(n_250) );
BUFx2_ASAP7_75t_L g251 ( .A(n_178), .Y(n_251) );
CKINVDCx11_ASAP7_75t_R g252 ( .A(n_199), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_213), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_218), .Y(n_254) );
INVxp33_ASAP7_75t_SL g255 ( .A(n_232), .Y(n_255) );
AND2x2_ASAP7_75t_L g256 ( .A(n_225), .B(n_173), .Y(n_256) );
INVx2_ASAP7_75t_L g257 ( .A(n_218), .Y(n_257) );
CKINVDCx5p33_ASAP7_75t_R g258 ( .A(n_232), .Y(n_258) );
AND2x4_ASAP7_75t_L g259 ( .A(n_196), .B(n_173), .Y(n_259) );
AND3x1_ASAP7_75t_SL g260 ( .A(n_200), .B(n_152), .C(n_164), .Y(n_260) );
INVx2_ASAP7_75t_L g261 ( .A(n_218), .Y(n_261) );
INVx3_ASAP7_75t_L g262 ( .A(n_222), .Y(n_262) );
INVx2_ASAP7_75t_L g263 ( .A(n_222), .Y(n_263) );
OAI22xp5_ASAP7_75t_L g264 ( .A1(n_192), .A2(n_156), .B1(n_143), .B2(n_151), .Y(n_264) );
AND2x2_ASAP7_75t_L g265 ( .A(n_225), .B(n_156), .Y(n_265) );
INVx1_ASAP7_75t_L g266 ( .A(n_222), .Y(n_266) );
INVx2_ASAP7_75t_L g267 ( .A(n_210), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_202), .B(n_169), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_208), .Y(n_269) );
INVx5_ASAP7_75t_L g270 ( .A(n_208), .Y(n_270) );
NOR3xp33_ASAP7_75t_SL g271 ( .A(n_179), .B(n_143), .C(n_165), .Y(n_271) );
NOR3xp33_ASAP7_75t_SL g272 ( .A(n_194), .B(n_151), .C(n_165), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_207), .B(n_223), .Y(n_273) );
NOR3xp33_ASAP7_75t_SL g274 ( .A(n_206), .B(n_169), .C(n_164), .Y(n_274) );
NAND2xp33_ASAP7_75t_SL g275 ( .A(n_212), .B(n_145), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_220), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_224), .B(n_141), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_220), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_208), .Y(n_279) );
INVx5_ASAP7_75t_L g280 ( .A(n_208), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_229), .B(n_141), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_192), .Y(n_282) );
BUFx3_ASAP7_75t_L g283 ( .A(n_214), .Y(n_283) );
INVx2_ASAP7_75t_L g284 ( .A(n_210), .Y(n_284) );
NOR2xp33_ASAP7_75t_R g285 ( .A(n_199), .B(n_160), .Y(n_285) );
AOI22xp5_ASAP7_75t_L g286 ( .A1(n_188), .A2(n_158), .B1(n_132), .B2(n_135), .Y(n_286) );
BUFx6f_ASAP7_75t_L g287 ( .A(n_214), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_229), .B(n_158), .Y(n_288) );
OR2x6_ASAP7_75t_L g289 ( .A(n_200), .B(n_140), .Y(n_289) );
BUFx2_ASAP7_75t_L g290 ( .A(n_199), .Y(n_290) );
CKINVDCx5p33_ASAP7_75t_R g291 ( .A(n_199), .Y(n_291) );
BUFx6f_ASAP7_75t_L g292 ( .A(n_214), .Y(n_292) );
INVx1_ASAP7_75t_L g293 ( .A(n_227), .Y(n_293) );
INVx1_ASAP7_75t_L g294 ( .A(n_227), .Y(n_294) );
INVx5_ASAP7_75t_L g295 ( .A(n_214), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_233), .Y(n_296) );
NAND2xp5_ASAP7_75t_L g297 ( .A(n_185), .B(n_140), .Y(n_297) );
AND2x4_ASAP7_75t_L g298 ( .A(n_188), .B(n_135), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_233), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_212), .B(n_167), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_209), .B(n_167), .Y(n_301) );
INVx2_ASAP7_75t_L g302 ( .A(n_267), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_240), .Y(n_303) );
INVx3_ASAP7_75t_L g304 ( .A(n_262), .Y(n_304) );
INVx5_ASAP7_75t_L g305 ( .A(n_262), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_298), .B(n_234), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_282), .A2(n_219), .B1(n_200), .B2(n_209), .Y(n_307) );
OR2x6_ASAP7_75t_L g308 ( .A(n_289), .B(n_200), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_298), .Y(n_309) );
INVx2_ASAP7_75t_SL g310 ( .A(n_243), .Y(n_310) );
BUFx2_ASAP7_75t_L g311 ( .A(n_243), .Y(n_311) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_244), .B(n_217), .Y(n_312) );
INVx1_ASAP7_75t_L g313 ( .A(n_298), .Y(n_313) );
INVx3_ASAP7_75t_L g314 ( .A(n_262), .Y(n_314) );
OR2x6_ASAP7_75t_L g315 ( .A(n_289), .B(n_211), .Y(n_315) );
NAND2xp33_ASAP7_75t_L g316 ( .A(n_285), .B(n_211), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_259), .B(n_216), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g318 ( .A1(n_238), .A2(n_183), .B1(n_228), .B2(n_215), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g319 ( .A(n_259), .B(n_175), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_301), .A2(n_201), .B(n_204), .Y(n_320) );
INVx2_ASAP7_75t_L g321 ( .A(n_267), .Y(n_321) );
BUFx3_ASAP7_75t_L g322 ( .A(n_243), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g323 ( .A(n_259), .B(n_226), .Y(n_323) );
BUFx3_ASAP7_75t_L g324 ( .A(n_290), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_269), .Y(n_325) );
OR2x2_ASAP7_75t_L g326 ( .A(n_251), .B(n_160), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_273), .Y(n_327) );
INVxp67_ASAP7_75t_SL g328 ( .A(n_235), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_265), .B(n_226), .Y(n_329) );
INVxp67_ASAP7_75t_SL g330 ( .A(n_245), .Y(n_330) );
BUFx3_ASAP7_75t_L g331 ( .A(n_269), .Y(n_331) );
NOR2xp33_ASAP7_75t_L g332 ( .A(n_247), .B(n_160), .Y(n_332) );
BUFx6f_ASAP7_75t_L g333 ( .A(n_240), .Y(n_333) );
BUFx6f_ASAP7_75t_L g334 ( .A(n_240), .Y(n_334) );
NAND2xp5_ASAP7_75t_SL g335 ( .A(n_285), .B(n_236), .Y(n_335) );
INVx5_ASAP7_75t_L g336 ( .A(n_240), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_284), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_252), .Y(n_338) );
BUFx8_ASAP7_75t_L g339 ( .A(n_248), .Y(n_339) );
INVx3_ASAP7_75t_SL g340 ( .A(n_291), .Y(n_340) );
NAND2xp5_ASAP7_75t_L g341 ( .A(n_256), .B(n_231), .Y(n_341) );
INVx3_ASAP7_75t_L g342 ( .A(n_236), .Y(n_342) );
INVx2_ASAP7_75t_SL g343 ( .A(n_241), .Y(n_343) );
NAND2x1p5_ASAP7_75t_L g344 ( .A(n_241), .B(n_231), .Y(n_344) );
INVx1_ASAP7_75t_SL g345 ( .A(n_241), .Y(n_345) );
BUFx8_ASAP7_75t_SL g346 ( .A(n_258), .Y(n_346) );
INVx3_ASAP7_75t_L g347 ( .A(n_246), .Y(n_347) );
INVx2_ASAP7_75t_L g348 ( .A(n_284), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_279), .Y(n_349) );
AOI22xp5_ASAP7_75t_L g350 ( .A1(n_237), .A2(n_231), .B1(n_214), .B2(n_131), .Y(n_350) );
AND2x4_ASAP7_75t_L g351 ( .A(n_272), .B(n_166), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_246), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_268), .Y(n_353) );
NAND2xp5_ASAP7_75t_SL g354 ( .A(n_249), .B(n_231), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_289), .Y(n_355) );
OAI21xp5_ASAP7_75t_L g356 ( .A1(n_276), .A2(n_190), .B(n_186), .Y(n_356) );
INVx1_ASAP7_75t_SL g357 ( .A(n_252), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_327), .Y(n_358) );
BUFx2_ASAP7_75t_SL g359 ( .A(n_322), .Y(n_359) );
AOI22xp33_ASAP7_75t_SL g360 ( .A1(n_308), .A2(n_255), .B1(n_289), .B2(n_258), .Y(n_360) );
OAI22xp33_ASAP7_75t_L g361 ( .A1(n_308), .A2(n_255), .B1(n_291), .B2(n_286), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_308), .A2(n_237), .B1(n_247), .B2(n_239), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_353), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_308), .B(n_247), .Y(n_364) );
INVx1_ASAP7_75t_L g365 ( .A(n_302), .Y(n_365) );
NAND2xp5_ASAP7_75t_L g366 ( .A(n_351), .B(n_264), .Y(n_366) );
CKINVDCx5p33_ASAP7_75t_R g367 ( .A(n_346), .Y(n_367) );
AO31x2_ASAP7_75t_L g368 ( .A1(n_307), .A2(n_166), .A3(n_131), .B(n_294), .Y(n_368) );
NOR2xp33_ASAP7_75t_L g369 ( .A(n_317), .B(n_239), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_302), .Y(n_370) );
OR2x6_ASAP7_75t_L g371 ( .A(n_315), .B(n_237), .Y(n_371) );
INVx2_ASAP7_75t_L g372 ( .A(n_321), .Y(n_372) );
INVxp33_ASAP7_75t_L g373 ( .A(n_346), .Y(n_373) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_351), .B(n_277), .Y(n_374) );
AOI22xp33_ASAP7_75t_SL g375 ( .A1(n_355), .A2(n_260), .B1(n_300), .B2(n_297), .Y(n_375) );
AOI22xp33_ASAP7_75t_L g376 ( .A1(n_351), .A2(n_275), .B1(n_242), .B2(n_281), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_329), .B(n_288), .Y(n_377) );
BUFx3_ASAP7_75t_L g378 ( .A(n_315), .Y(n_378) );
INVx2_ASAP7_75t_L g379 ( .A(n_321), .Y(n_379) );
AND2x2_ASAP7_75t_L g380 ( .A(n_315), .B(n_278), .Y(n_380) );
AND2x4_ASAP7_75t_L g381 ( .A(n_322), .B(n_274), .Y(n_381) );
AOI21xp33_ASAP7_75t_L g382 ( .A1(n_343), .A2(n_299), .B(n_296), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g383 ( .A1(n_343), .A2(n_275), .B1(n_266), .B2(n_254), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_337), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_315), .B(n_293), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_323), .B(n_271), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_337), .Y(n_387) );
OAI21xp33_ASAP7_75t_L g388 ( .A1(n_332), .A2(n_131), .B(n_166), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_348), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_348), .Y(n_390) );
AOI221xp5_ASAP7_75t_L g391 ( .A1(n_309), .A2(n_162), .B1(n_250), .B2(n_253), .C(n_231), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_352), .Y(n_392) );
OAI221xp5_ASAP7_75t_SL g393 ( .A1(n_361), .A2(n_357), .B1(n_311), .B2(n_310), .C(n_326), .Y(n_393) );
AOI22xp33_ASAP7_75t_SL g394 ( .A1(n_359), .A2(n_339), .B1(n_338), .B2(n_310), .Y(n_394) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_381), .A2(n_339), .B1(n_306), .B2(n_328), .Y(n_395) );
OAI22xp33_ASAP7_75t_L g396 ( .A1(n_371), .A2(n_338), .B1(n_340), .B2(n_345), .Y(n_396) );
NAND2x1_ASAP7_75t_L g397 ( .A(n_372), .B(n_303), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_377), .B(n_319), .Y(n_398) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_378), .Y(n_399) );
BUFx6f_ASAP7_75t_L g400 ( .A(n_378), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_358), .Y(n_401) );
AOI221xp5_ASAP7_75t_L g402 ( .A1(n_369), .A2(n_313), .B1(n_312), .B2(n_306), .C(n_341), .Y(n_402) );
OAI211xp5_ASAP7_75t_L g403 ( .A1(n_375), .A2(n_318), .B(n_324), .C(n_350), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_377), .B(n_352), .Y(n_404) );
OAI22xp5_ASAP7_75t_L g405 ( .A1(n_360), .A2(n_344), .B1(n_324), .B2(n_340), .Y(n_405) );
OAI211xp5_ASAP7_75t_L g406 ( .A1(n_375), .A2(n_354), .B(n_335), .C(n_330), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_362), .A2(n_344), .B1(n_316), .B2(n_335), .C(n_304), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_358), .B(n_306), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_365), .Y(n_409) );
NOR2x1_ASAP7_75t_SL g410 ( .A(n_371), .B(n_303), .Y(n_410) );
AND2x4_ASAP7_75t_L g411 ( .A(n_363), .B(n_305), .Y(n_411) );
AOI22xp33_ASAP7_75t_L g412 ( .A1(n_381), .A2(n_339), .B1(n_314), .B2(n_304), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_365), .Y(n_413) );
OAI22xp33_ASAP7_75t_L g414 ( .A1(n_371), .A2(n_305), .B1(n_347), .B2(n_342), .Y(n_414) );
INVx3_ASAP7_75t_SL g415 ( .A(n_371), .Y(n_415) );
AOI221xp5_ASAP7_75t_L g416 ( .A1(n_363), .A2(n_320), .B1(n_347), .B2(n_342), .C(n_304), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_364), .B(n_342), .Y(n_417) );
AOI21xp5_ASAP7_75t_SL g418 ( .A1(n_378), .A2(n_303), .B(n_349), .Y(n_418) );
AND2x2_ASAP7_75t_L g419 ( .A(n_374), .B(n_347), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_372), .Y(n_420) );
AOI222xp33_ASAP7_75t_L g421 ( .A1(n_386), .A2(n_316), .B1(n_314), .B2(n_354), .C1(n_356), .C2(n_305), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_393), .A2(n_376), .B1(n_366), .B2(n_374), .C(n_383), .Y(n_422) );
AOI221xp5_ASAP7_75t_L g423 ( .A1(n_402), .A2(n_386), .B1(n_381), .B2(n_366), .C(n_364), .Y(n_423) );
INVx2_ASAP7_75t_SL g424 ( .A(n_404), .Y(n_424) );
BUFx10_ASAP7_75t_L g425 ( .A(n_411), .Y(n_425) );
NAND2xp33_ASAP7_75t_R g426 ( .A(n_411), .B(n_367), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_398), .A2(n_381), .B1(n_371), .B2(n_385), .Y(n_427) );
INVx2_ASAP7_75t_L g428 ( .A(n_420), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_404), .B(n_370), .Y(n_429) );
OAI221xp5_ASAP7_75t_L g430 ( .A1(n_395), .A2(n_359), .B1(n_388), .B2(n_391), .C(n_382), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_420), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g432 ( .A(n_398), .B(n_380), .Y(n_432) );
AO21x2_ASAP7_75t_L g433 ( .A1(n_406), .A2(n_382), .B(n_388), .Y(n_433) );
AOI22xp33_ASAP7_75t_L g434 ( .A1(n_396), .A2(n_380), .B1(n_385), .B2(n_391), .Y(n_434) );
AOI221xp5_ASAP7_75t_L g435 ( .A1(n_401), .A2(n_373), .B1(n_392), .B2(n_370), .C(n_387), .Y(n_435) );
AND2x2_ASAP7_75t_L g436 ( .A(n_409), .B(n_384), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_409), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g438 ( .A1(n_408), .A2(n_390), .B1(n_387), .B2(n_384), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_413), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_413), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_415), .A2(n_392), .B1(n_390), .B2(n_314), .Y(n_441) );
AOI22xp33_ASAP7_75t_L g442 ( .A1(n_415), .A2(n_389), .B1(n_379), .B2(n_372), .Y(n_442) );
NOR2x1_ASAP7_75t_SL g443 ( .A(n_405), .B(n_379), .Y(n_443) );
OAI33xp33_ASAP7_75t_L g444 ( .A1(n_417), .A2(n_186), .A3(n_203), .B1(n_197), .B2(n_177), .B3(n_190), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_410), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_397), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g447 ( .A1(n_408), .A2(n_412), .B1(n_403), .B2(n_394), .C(n_419), .Y(n_447) );
NAND2xp33_ASAP7_75t_R g448 ( .A(n_411), .B(n_379), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_419), .Y(n_449) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_415), .A2(n_389), .B1(n_305), .B2(n_325), .Y(n_450) );
NOR2xp33_ASAP7_75t_R g451 ( .A(n_399), .B(n_7), .Y(n_451) );
OR2x2_ASAP7_75t_L g452 ( .A(n_417), .B(n_368), .Y(n_452) );
AND2x4_ASAP7_75t_L g453 ( .A(n_410), .B(n_389), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_399), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_399), .Y(n_455) );
INVx3_ASAP7_75t_L g456 ( .A(n_399), .Y(n_456) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_429), .B(n_399), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_429), .B(n_368), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_440), .Y(n_459) );
INVx1_ASAP7_75t_SL g460 ( .A(n_451), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g461 ( .A1(n_423), .A2(n_421), .B1(n_416), .B2(n_414), .Y(n_461) );
INVx1_ASAP7_75t_L g462 ( .A(n_440), .Y(n_462) );
OAI221xp5_ASAP7_75t_L g463 ( .A1(n_427), .A2(n_407), .B1(n_400), .B2(n_397), .C(n_418), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_447), .A2(n_400), .B1(n_325), .B2(n_331), .Y(n_464) );
AO21x2_ASAP7_75t_L g465 ( .A1(n_433), .A2(n_418), .B(n_368), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_440), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_437), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_449), .B(n_368), .Y(n_468) );
NAND4xp25_ASAP7_75t_L g469 ( .A(n_435), .B(n_8), .C(n_9), .D(n_10), .Y(n_469) );
INVx2_ASAP7_75t_L g470 ( .A(n_428), .Y(n_470) );
NAND4xp25_ASAP7_75t_L g471 ( .A(n_434), .B(n_177), .C(n_203), .D(n_197), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_437), .Y(n_472) );
OAI221xp5_ASAP7_75t_L g473 ( .A1(n_422), .A2(n_400), .B1(n_280), .B2(n_270), .C(n_295), .Y(n_473) );
INVx5_ASAP7_75t_L g474 ( .A(n_425), .Y(n_474) );
HB1xp67_ASAP7_75t_L g475 ( .A(n_424), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_452), .B(n_368), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_424), .B(n_400), .Y(n_477) );
OAI22xp33_ASAP7_75t_L g478 ( .A1(n_448), .A2(n_400), .B1(n_305), .B2(n_336), .Y(n_478) );
BUFx2_ASAP7_75t_L g479 ( .A(n_445), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_449), .B(n_368), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_436), .B(n_8), .Y(n_481) );
HB1xp67_ASAP7_75t_L g482 ( .A(n_436), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_439), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_428), .Y(n_484) );
BUFx3_ASAP7_75t_L g485 ( .A(n_425), .Y(n_485) );
INVxp67_ASAP7_75t_L g486 ( .A(n_426), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_432), .B(n_9), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_439), .B(n_10), .Y(n_488) );
AOI211x1_ASAP7_75t_L g489 ( .A1(n_430), .A2(n_11), .B(n_12), .C(n_13), .Y(n_489) );
INVx4_ASAP7_75t_L g490 ( .A(n_425), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
INVx3_ASAP7_75t_L g492 ( .A(n_453), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_431), .B(n_11), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_452), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_431), .B(n_12), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_438), .B(n_13), .Y(n_496) );
INVx2_ASAP7_75t_L g497 ( .A(n_446), .Y(n_497) );
INVx1_ASAP7_75t_SL g498 ( .A(n_425), .Y(n_498) );
AOI22xp5_ASAP7_75t_L g499 ( .A1(n_438), .A2(n_331), .B1(n_336), .B2(n_334), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_453), .B(n_14), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_453), .B(n_14), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_453), .B(n_17), .Y(n_502) );
INVx1_ASAP7_75t_L g503 ( .A(n_446), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_454), .B(n_19), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_441), .B(n_20), .Y(n_505) );
OR2x2_ASAP7_75t_L g506 ( .A(n_482), .B(n_455), .Y(n_506) );
NAND2xp33_ASAP7_75t_R g507 ( .A(n_479), .B(n_455), .Y(n_507) );
OR2x2_ASAP7_75t_L g508 ( .A(n_494), .B(n_454), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_458), .B(n_456), .Y(n_509) );
INVx2_ASAP7_75t_SL g510 ( .A(n_479), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_467), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_458), .B(n_456), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_467), .Y(n_513) );
INVxp67_ASAP7_75t_L g514 ( .A(n_475), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_481), .B(n_456), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_492), .B(n_446), .Y(n_516) );
OAI321xp33_ASAP7_75t_L g517 ( .A1(n_469), .A2(n_442), .A3(n_450), .B1(n_443), .B2(n_176), .C(n_189), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_481), .B(n_456), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_472), .Y(n_519) );
NOR2xp33_ASAP7_75t_R g520 ( .A(n_474), .B(n_20), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_494), .B(n_433), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_472), .Y(n_522) );
AND2x2_ASAP7_75t_SL g523 ( .A(n_490), .B(n_443), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_468), .B(n_433), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_483), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_470), .Y(n_526) );
OR2x2_ASAP7_75t_L g527 ( .A(n_457), .B(n_22), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_460), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_488), .B(n_483), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_500), .B(n_25), .Y(n_530) );
AND2x2_ASAP7_75t_L g531 ( .A(n_500), .B(n_32), .Y(n_531) );
INVx1_ASAP7_75t_L g532 ( .A(n_459), .Y(n_532) );
INVx2_ASAP7_75t_L g533 ( .A(n_470), .Y(n_533) );
NAND4xp25_ASAP7_75t_L g534 ( .A(n_469), .B(n_176), .C(n_180), .D(n_181), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_459), .Y(n_535) );
INVx2_ASAP7_75t_L g536 ( .A(n_470), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_488), .B(n_336), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_462), .Y(n_538) );
INVx1_ASAP7_75t_SL g539 ( .A(n_498), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_468), .B(n_35), .Y(n_540) );
OR2x2_ASAP7_75t_L g541 ( .A(n_476), .B(n_50), .Y(n_541) );
HB1xp67_ASAP7_75t_L g542 ( .A(n_484), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g543 ( .A(n_501), .B(n_336), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_480), .B(n_52), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g545 ( .A(n_489), .B(n_205), .C(n_191), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_501), .B(n_336), .Y(n_546) );
AND2x4_ASAP7_75t_SL g547 ( .A(n_490), .B(n_303), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_462), .Y(n_548) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_480), .B(n_280), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_476), .B(n_53), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_504), .B(n_280), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_504), .B(n_280), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_466), .Y(n_553) );
INVx1_ASAP7_75t_L g554 ( .A(n_466), .Y(n_554) );
NAND4xp25_ASAP7_75t_L g555 ( .A(n_464), .B(n_180), .C(n_181), .D(n_182), .Y(n_555) );
NOR2xp33_ASAP7_75t_L g556 ( .A(n_486), .B(n_487), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_485), .B(n_55), .Y(n_557) );
INVxp67_ASAP7_75t_L g558 ( .A(n_485), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_492), .B(n_58), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_493), .B(n_295), .Y(n_560) );
INVx1_ASAP7_75t_L g561 ( .A(n_493), .Y(n_561) );
HB1xp67_ASAP7_75t_L g562 ( .A(n_484), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_478), .B(n_349), .Y(n_563) );
OAI22xp33_ASAP7_75t_SL g564 ( .A1(n_510), .A2(n_490), .B1(n_485), .B2(n_474), .Y(n_564) );
INVx2_ASAP7_75t_L g565 ( .A(n_542), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_529), .B(n_495), .Y(n_566) );
NOR2xp67_ASAP7_75t_L g567 ( .A(n_510), .B(n_474), .Y(n_567) );
AOI21xp5_ASAP7_75t_L g568 ( .A1(n_563), .A2(n_473), .B(n_463), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_561), .B(n_495), .Y(n_570) );
AOI221xp5_ASAP7_75t_L g571 ( .A1(n_556), .A2(n_489), .B1(n_496), .B2(n_502), .C(n_505), .Y(n_571) );
AOI32xp33_ASAP7_75t_L g572 ( .A1(n_528), .A2(n_490), .A3(n_492), .B1(n_503), .B2(n_477), .Y(n_572) );
AND2x2_ASAP7_75t_L g573 ( .A(n_509), .B(n_492), .Y(n_573) );
OAI31xp33_ASAP7_75t_L g574 ( .A1(n_534), .A2(n_471), .A3(n_503), .B(n_497), .Y(n_574) );
AOI221xp5_ASAP7_75t_L g575 ( .A1(n_556), .A2(n_461), .B1(n_497), .B2(n_444), .C(n_465), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_509), .B(n_491), .Y(n_576) );
OAI32xp33_ASAP7_75t_L g577 ( .A1(n_507), .A2(n_497), .A3(n_491), .B1(n_484), .B2(n_474), .Y(n_577) );
OAI22xp5_ASAP7_75t_SL g578 ( .A1(n_523), .A2(n_474), .B1(n_461), .B2(n_499), .Y(n_578) );
OAI221xp5_ASAP7_75t_SL g579 ( .A1(n_541), .A2(n_499), .B1(n_491), .B2(n_474), .C(n_465), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_513), .Y(n_580) );
AOI31xp33_ASAP7_75t_L g581 ( .A1(n_507), .A2(n_465), .A3(n_61), .B(n_65), .Y(n_581) );
INVx1_ASAP7_75t_SL g582 ( .A(n_539), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_519), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_522), .Y(n_584) );
A2O1A1Ixp33_ASAP7_75t_L g585 ( .A1(n_517), .A2(n_349), .B(n_334), .C(n_333), .Y(n_585) );
INVx1_ASAP7_75t_SL g586 ( .A(n_520), .Y(n_586) );
OAI22xp33_ASAP7_75t_L g587 ( .A1(n_545), .A2(n_349), .B1(n_334), .B2(n_333), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_542), .Y(n_588) );
AOI221xp5_ASAP7_75t_L g589 ( .A1(n_514), .A2(n_205), .B1(n_191), .B2(n_189), .C(n_184), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_525), .B(n_524), .Y(n_590) );
INVxp67_ASAP7_75t_L g591 ( .A(n_521), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_512), .B(n_60), .Y(n_592) );
INVx2_ASAP7_75t_L g593 ( .A(n_562), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_532), .Y(n_594) );
NAND2xp33_ASAP7_75t_L g595 ( .A(n_520), .B(n_334), .Y(n_595) );
NOR4xp25_ASAP7_75t_SL g596 ( .A(n_563), .B(n_68), .C(n_69), .D(n_72), .Y(n_596) );
AND2x2_ASAP7_75t_SL g597 ( .A(n_523), .B(n_333), .Y(n_597) );
AOI22xp33_ASAP7_75t_L g598 ( .A1(n_550), .A2(n_292), .B1(n_287), .B2(n_279), .Y(n_598) );
OAI221xp5_ASAP7_75t_L g599 ( .A1(n_558), .A2(n_195), .B1(n_182), .B2(n_270), .C(n_295), .Y(n_599) );
AOI221xp5_ASAP7_75t_L g600 ( .A1(n_524), .A2(n_205), .B1(n_191), .B2(n_189), .C(n_184), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_535), .Y(n_601) );
OR2x2_ASAP7_75t_L g602 ( .A(n_506), .B(n_73), .Y(n_602) );
AND4x1_ASAP7_75t_L g603 ( .A(n_530), .B(n_76), .C(n_77), .D(n_78), .Y(n_603) );
NAND3xp33_ASAP7_75t_L g604 ( .A(n_550), .B(n_184), .C(n_189), .Y(n_604) );
OAI21xp33_ASAP7_75t_L g605 ( .A1(n_512), .A2(n_195), .B(n_189), .Y(n_605) );
INVx1_ASAP7_75t_SL g606 ( .A(n_547), .Y(n_606) );
OAI31xp33_ASAP7_75t_L g607 ( .A1(n_531), .A2(n_283), .A3(n_249), .B(n_257), .Y(n_607) );
NOR2xp33_ASAP7_75t_L g608 ( .A(n_515), .B(n_184), .Y(n_608) );
AOI22xp5_ASAP7_75t_L g609 ( .A1(n_518), .A2(n_270), .B1(n_295), .B2(n_292), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_538), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_548), .Y(n_611) );
AOI21xp33_ASAP7_75t_SL g612 ( .A1(n_557), .A2(n_263), .B(n_257), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_540), .B(n_295), .Y(n_613) );
CKINVDCx16_ASAP7_75t_R g614 ( .A(n_540), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_553), .Y(n_615) );
OAI21xp5_ASAP7_75t_L g616 ( .A1(n_544), .A2(n_270), .B(n_283), .Y(n_616) );
INVx1_ASAP7_75t_L g617 ( .A(n_554), .Y(n_617) );
NOR2xp67_ASAP7_75t_SL g618 ( .A(n_614), .B(n_544), .Y(n_618) );
XNOR2xp5_ASAP7_75t_L g619 ( .A(n_582), .B(n_543), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_590), .B(n_508), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_569), .Y(n_621) );
XNOR2xp5_ASAP7_75t_L g622 ( .A(n_586), .B(n_597), .Y(n_622) );
BUFx2_ASAP7_75t_L g623 ( .A(n_597), .Y(n_623) );
AND2x2_ASAP7_75t_L g624 ( .A(n_576), .B(n_516), .Y(n_624) );
INVx1_ASAP7_75t_L g625 ( .A(n_580), .Y(n_625) );
NOR3xp33_ASAP7_75t_SL g626 ( .A(n_578), .B(n_549), .C(n_537), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_583), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_591), .B(n_562), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_591), .B(n_526), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_588), .B(n_565), .Y(n_630) );
INVxp67_ASAP7_75t_L g631 ( .A(n_565), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_584), .Y(n_632) );
XOR2xp5_ASAP7_75t_L g633 ( .A(n_566), .B(n_546), .Y(n_633) );
INVx1_ASAP7_75t_SL g634 ( .A(n_606), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_594), .B(n_536), .Y(n_635) );
OAI21xp5_ASAP7_75t_SL g636 ( .A1(n_581), .A2(n_547), .B(n_559), .Y(n_636) );
INVxp67_ASAP7_75t_L g637 ( .A(n_593), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_601), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_610), .Y(n_639) );
OR2x2_ASAP7_75t_L g640 ( .A(n_593), .B(n_536), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_611), .B(n_526), .Y(n_641) );
OAI21xp5_ASAP7_75t_L g642 ( .A1(n_574), .A2(n_559), .B(n_551), .Y(n_642) );
NOR2xp67_ASAP7_75t_SL g643 ( .A(n_604), .B(n_527), .Y(n_643) );
AND2x2_ASAP7_75t_L g644 ( .A(n_573), .B(n_516), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_615), .B(n_516), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_617), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_570), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g648 ( .A(n_575), .B(n_533), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_564), .Y(n_649) );
OR2x2_ASAP7_75t_L g650 ( .A(n_567), .B(n_533), .Y(n_650) );
NOR2xp33_ASAP7_75t_L g651 ( .A(n_612), .B(n_602), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_608), .Y(n_652) );
NOR2x1_ASAP7_75t_L g653 ( .A(n_595), .B(n_555), .Y(n_653) );
NOR4xp25_ASAP7_75t_SL g654 ( .A(n_579), .B(n_552), .C(n_560), .D(n_270), .Y(n_654) );
NOR4xp25_ASAP7_75t_SL g655 ( .A(n_579), .B(n_184), .C(n_191), .D(n_205), .Y(n_655) );
AND2x2_ASAP7_75t_L g656 ( .A(n_608), .B(n_191), .Y(n_656) );
INVx1_ASAP7_75t_SL g657 ( .A(n_634), .Y(n_657) );
AOI21xp33_ASAP7_75t_L g658 ( .A1(n_649), .A2(n_571), .B(n_592), .Y(n_658) );
AOI222xp33_ASAP7_75t_L g659 ( .A1(n_648), .A2(n_577), .B1(n_616), .B2(n_613), .C1(n_585), .C2(n_605), .Y(n_659) );
INVx1_ASAP7_75t_L g660 ( .A(n_621), .Y(n_660) );
OAI22xp5_ASAP7_75t_L g661 ( .A1(n_636), .A2(n_572), .B1(n_598), .B2(n_568), .Y(n_661) );
INVx2_ASAP7_75t_L g662 ( .A(n_630), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g663 ( .A(n_647), .B(n_645), .Y(n_663) );
NAND3xp33_ASAP7_75t_L g664 ( .A(n_626), .B(n_585), .C(n_603), .Y(n_664) );
AOI22xp5_ASAP7_75t_L g665 ( .A1(n_618), .A2(n_609), .B1(n_587), .B2(n_598), .Y(n_665) );
XOR2xp5_ASAP7_75t_L g666 ( .A(n_622), .B(n_587), .Y(n_666) );
INVx2_ASAP7_75t_SL g667 ( .A(n_624), .Y(n_667) );
INVx1_ASAP7_75t_L g668 ( .A(n_625), .Y(n_668) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_647), .B(n_600), .Y(n_669) );
XNOR2xp5_ASAP7_75t_L g670 ( .A(n_633), .B(n_599), .Y(n_670) );
NAND2xp5_ASAP7_75t_L g671 ( .A(n_627), .B(n_589), .Y(n_671) );
INVx1_ASAP7_75t_L g672 ( .A(n_632), .Y(n_672) );
CKINVDCx20_ASAP7_75t_R g673 ( .A(n_619), .Y(n_673) );
NAND3x2_ASAP7_75t_L g674 ( .A(n_623), .B(n_607), .C(n_596), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_638), .Y(n_675) );
XNOR2xp5_ASAP7_75t_L g676 ( .A(n_626), .B(n_261), .Y(n_676) );
NAND3xp33_ASAP7_75t_L g677 ( .A(n_642), .B(n_205), .C(n_279), .Y(n_677) );
AND2x2_ASAP7_75t_L g678 ( .A(n_644), .B(n_279), .Y(n_678) );
INVx2_ASAP7_75t_SL g679 ( .A(n_624), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_639), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_660), .Y(n_681) );
AOI321xp33_ASAP7_75t_L g682 ( .A1(n_661), .A2(n_652), .A3(n_651), .B1(n_653), .B2(n_645), .C(n_620), .Y(n_682) );
HB1xp67_ASAP7_75t_L g683 ( .A(n_657), .Y(n_683) );
AO22x2_ASAP7_75t_L g684 ( .A1(n_661), .A2(n_646), .B1(n_637), .B2(n_631), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_668), .Y(n_685) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_667), .A2(n_651), .B(n_650), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_672), .Y(n_687) );
NAND2xp5_ASAP7_75t_SL g688 ( .A(n_659), .B(n_637), .Y(n_688) );
INVx1_ASAP7_75t_SL g689 ( .A(n_673), .Y(n_689) );
OAI211xp5_ASAP7_75t_SL g690 ( .A1(n_658), .A2(n_628), .B(n_631), .C(n_629), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_671), .B(n_641), .Y(n_691) );
OAI21xp33_ASAP7_75t_SL g692 ( .A1(n_679), .A2(n_644), .B(n_635), .Y(n_692) );
INVx2_ASAP7_75t_SL g693 ( .A(n_662), .Y(n_693) );
NAND2xp5_ASAP7_75t_L g694 ( .A(n_675), .B(n_640), .Y(n_694) );
AOI21xp33_ASAP7_75t_L g695 ( .A1(n_674), .A2(n_671), .B(n_664), .Y(n_695) );
NOR3xp33_ASAP7_75t_L g696 ( .A(n_658), .B(n_656), .C(n_654), .Y(n_696) );
NAND5xp2_ASAP7_75t_L g697 ( .A(n_665), .B(n_656), .C(n_655), .D(n_643), .E(n_292), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_669), .A2(n_261), .B(n_263), .C(n_287), .Y(n_698) );
AOI221xp5_ASAP7_75t_L g699 ( .A1(n_680), .A2(n_287), .B1(n_666), .B2(n_670), .C(n_663), .Y(n_699) );
O2A1O1Ixp5_ASAP7_75t_L g700 ( .A1(n_677), .A2(n_658), .B(n_649), .C(n_661), .Y(n_700) );
NAND2x1p5_ASAP7_75t_L g701 ( .A(n_678), .B(n_676), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_695), .B(n_691), .Y(n_702) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_689), .Y(n_703) );
NAND3xp33_ASAP7_75t_SL g704 ( .A(n_700), .B(n_682), .C(n_699), .Y(n_704) );
OAI21x1_ASAP7_75t_L g705 ( .A1(n_688), .A2(n_683), .B(n_701), .Y(n_705) );
INVx1_ASAP7_75t_SL g706 ( .A(n_693), .Y(n_706) );
NAND2xp5_ASAP7_75t_L g707 ( .A(n_702), .B(n_696), .Y(n_707) );
NOR3xp33_ASAP7_75t_SL g708 ( .A(n_704), .B(n_690), .C(n_697), .Y(n_708) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_703), .B(n_698), .Y(n_709) );
INVxp67_ASAP7_75t_SL g710 ( .A(n_709), .Y(n_710) );
AND2x4_ASAP7_75t_L g711 ( .A(n_708), .B(n_706), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_711), .Y(n_712) );
OAI21xp5_ASAP7_75t_L g713 ( .A1(n_710), .A2(n_707), .B(n_705), .Y(n_713) );
AOI322xp5_ASAP7_75t_L g714 ( .A1(n_712), .A2(n_711), .A3(n_686), .B1(n_692), .B2(n_684), .C1(n_681), .C2(n_685), .Y(n_714) );
AOI221xp5_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_713), .B1(n_684), .B2(n_687), .C(n_694), .Y(n_715) );
endmodule