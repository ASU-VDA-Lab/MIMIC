module fake_jpeg_26596_n_341 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_341);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_341;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx11_ASAP7_75t_R g18 ( 
.A(n_4),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

INVx11_ASAP7_75t_SL g20 ( 
.A(n_5),
.Y(n_20)
);

INVx8_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_16),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_2),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_6),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx5_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_14),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVxp67_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

INVx3_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx6_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_32),
.B(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_38),
.B(n_39),
.Y(n_49)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_32),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

CKINVDCx16_ASAP7_75t_R g41 ( 
.A(n_20),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_41),
.B(n_48),
.Y(n_66)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_17),
.Y(n_42)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_42),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_7),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_43),
.B(n_29),
.Y(n_54)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

INVx6_ASAP7_75t_L g61 ( 
.A(n_44),
.Y(n_61)
);

BUFx12_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_45),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

BUFx2_ASAP7_75t_SL g59 ( 
.A(n_46),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

INVx6_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_53),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_56),
.Y(n_73)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_47),
.Y(n_55)
);

INVx1_ASAP7_75t_SL g78 ( 
.A(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_24),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_48),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_67),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_60),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_42),
.B(n_47),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_63),
.B(n_26),
.Y(n_88)
);

CKINVDCx14_ASAP7_75t_R g64 ( 
.A(n_38),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_64),
.B(n_28),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_70),
.B(n_41),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_63),
.A2(n_22),
.B1(n_42),
.B2(n_21),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_L g106 ( 
.A1(n_71),
.A2(n_98),
.B1(n_40),
.B2(n_44),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_72),
.Y(n_108)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_76),
.B(n_82),
.Y(n_112)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_79),
.Y(n_105)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_49),
.Y(n_82)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_83),
.Y(n_126)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2x1_ASAP7_75t_L g86 ( 
.A(n_55),
.B(n_46),
.Y(n_86)
);

AND2x2_ASAP7_75t_L g104 ( 
.A(n_86),
.B(n_88),
.Y(n_104)
);

CKINVDCx12_ASAP7_75t_R g87 ( 
.A(n_69),
.Y(n_87)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_87),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_89),
.Y(n_125)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_90),
.B(n_91),
.Y(n_115)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_92),
.B(n_96),
.Y(n_119)
);

INVx11_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_93),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_50),
.A2(n_22),
.B1(n_40),
.B2(n_18),
.Y(n_94)
);

OAI21xp33_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_30),
.B(n_70),
.Y(n_107)
);

INVx6_ASAP7_75t_SL g95 ( 
.A(n_53),
.Y(n_95)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_95),
.Y(n_124)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_56),
.Y(n_97)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_97),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g98 ( 
.A1(n_57),
.A2(n_22),
.B1(n_21),
.B2(n_37),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_99),
.B(n_31),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_54),
.C(n_39),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_101),
.B(n_116),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_85),
.A2(n_44),
.B1(n_37),
.B2(n_61),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_102),
.A2(n_118),
.B1(n_74),
.B2(n_77),
.Y(n_147)
);

OAI32xp33_ASAP7_75t_L g103 ( 
.A1(n_97),
.A2(n_30),
.A3(n_39),
.B1(n_61),
.B2(n_18),
.Y(n_103)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_103),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_106),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g153 ( 
.A1(n_107),
.A2(n_34),
.B1(n_95),
.B2(n_77),
.Y(n_153)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_75),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g142 ( 
.A(n_109),
.Y(n_142)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_75),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_113),
.B(n_93),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_114),
.B(n_33),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_73),
.B(n_46),
.Y(n_116)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_87),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_117),
.A2(n_90),
.B1(n_84),
.B2(n_74),
.Y(n_135)
);

AO22x1_ASAP7_75t_SL g118 ( 
.A1(n_86),
.A2(n_46),
.B1(n_40),
.B2(n_26),
.Y(n_118)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_120),
.Y(n_143)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_84),
.Y(n_122)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_122),
.Y(n_148)
);

AND2x2_ASAP7_75t_SL g123 ( 
.A(n_86),
.B(n_26),
.Y(n_123)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_123),
.A2(n_78),
.B(n_91),
.Y(n_144)
);

MAJx2_ASAP7_75t_L g127 ( 
.A(n_76),
.B(n_28),
.C(n_31),
.Y(n_127)
);

AND2x6_ASAP7_75t_L g137 ( 
.A(n_127),
.B(n_10),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_100),
.B(n_73),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_129),
.B(n_139),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_123),
.A2(n_81),
.B1(n_96),
.B2(n_83),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_130),
.A2(n_131),
.B1(n_147),
.B2(n_113),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g131 ( 
.A1(n_123),
.A2(n_81),
.B1(n_79),
.B2(n_92),
.Y(n_131)
);

INVx2_ASAP7_75t_SL g132 ( 
.A(n_110),
.Y(n_132)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_132),
.Y(n_172)
);

AND2x2_ASAP7_75t_SL g133 ( 
.A(n_104),
.B(n_26),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_SL g181 ( 
.A1(n_133),
.A2(n_137),
.B(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_116),
.B(n_78),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_134),
.B(n_150),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g164 ( 
.A(n_135),
.Y(n_164)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_136),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_122),
.Y(n_139)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_117),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_141),
.B(n_145),
.Y(n_165)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_105),
.Y(n_145)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_146),
.Y(n_184)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_119),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_149),
.B(n_157),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_100),
.B(n_121),
.Y(n_150)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_126),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_151),
.B(n_126),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_104),
.B(n_24),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_152),
.B(n_154),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g190 ( 
.A1(n_153),
.A2(n_65),
.B(n_60),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_104),
.B(n_24),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_121),
.B(n_19),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_155),
.B(n_156),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_101),
.B(n_23),
.Y(n_156)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_SL g195 ( 
.A(n_158),
.B(n_166),
.C(n_141),
.Y(n_195)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_142),
.Y(n_159)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_159),
.Y(n_192)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_128),
.A2(n_102),
.B1(n_112),
.B2(n_118),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_162),
.A2(n_163),
.B1(n_167),
.B2(n_177),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_128),
.A2(n_118),
.B1(n_103),
.B2(n_109),
.Y(n_163)
);

OAI21xp5_ASAP7_75t_L g166 ( 
.A1(n_152),
.A2(n_127),
.B(n_125),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_105),
.B1(n_124),
.B2(n_108),
.Y(n_167)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_168),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_156),
.C(n_133),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_170),
.B(n_175),
.C(n_23),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_124),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_148),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g174 ( 
.A1(n_133),
.A2(n_111),
.B(n_1),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_174),
.A2(n_190),
.B(n_148),
.Y(n_191)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_133),
.B(n_134),
.C(n_154),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g176 ( 
.A(n_130),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g201 ( 
.A(n_176),
.B(n_180),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_138),
.A2(n_110),
.B1(n_34),
.B2(n_30),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_111),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_27),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_182),
.B(n_146),
.Y(n_196)
);

INVxp67_ASAP7_75t_L g183 ( 
.A(n_131),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_183),
.B(n_142),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_144),
.A2(n_153),
.B1(n_137),
.B2(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_185),
.A2(n_186),
.B1(n_189),
.B2(n_28),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_157),
.A2(n_34),
.B1(n_25),
.B2(n_29),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_33),
.B1(n_23),
.B2(n_27),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g204 ( 
.A(n_187),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_155),
.B(n_25),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g219 ( 
.A(n_188),
.B(n_8),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_143),
.A2(n_23),
.B1(n_36),
.B2(n_31),
.Y(n_189)
);

NAND2xp33_ASAP7_75t_SL g234 ( 
.A(n_191),
.B(n_195),
.Y(n_234)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_193),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_196),
.B(n_202),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g246 ( 
.A(n_197),
.B(n_214),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_184),
.B(n_141),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_SL g222 ( 
.A(n_198),
.B(n_200),
.Y(n_222)
);

AOI22x1_ASAP7_75t_L g199 ( 
.A1(n_176),
.A2(n_142),
.B1(n_151),
.B2(n_132),
.Y(n_199)
);

AOI22xp5_ASAP7_75t_L g231 ( 
.A1(n_199),
.A2(n_164),
.B1(n_172),
.B2(n_177),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_179),
.B(n_178),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_145),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_208),
.C(n_216),
.Y(n_224)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_165),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_206),
.Y(n_232)
);

INVxp67_ASAP7_75t_SL g206 ( 
.A(n_182),
.Y(n_206)
);

OR2x4_ASAP7_75t_L g207 ( 
.A(n_163),
.B(n_132),
.Y(n_207)
);

AO22x1_ASAP7_75t_L g227 ( 
.A1(n_207),
.A2(n_183),
.B1(n_167),
.B2(n_190),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g208 ( 
.A(n_170),
.B(n_171),
.C(n_175),
.Y(n_208)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_164),
.A2(n_0),
.B(n_2),
.Y(n_209)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_209),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_179),
.B(n_36),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_210),
.B(n_217),
.Y(n_228)
);

CKINVDCx14_ASAP7_75t_R g211 ( 
.A(n_161),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_211),
.B(n_215),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_185),
.B(n_162),
.Y(n_212)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_212),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_181),
.A2(n_174),
.B(n_166),
.Y(n_214)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_52),
.C(n_69),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_178),
.B(n_36),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_159),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_219),
.Y(n_241)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_172),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_220),
.B(n_0),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_173),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g248 ( 
.A(n_223),
.B(n_214),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_160),
.C(n_173),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_225),
.B(n_226),
.C(n_237),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_169),
.C(n_158),
.Y(n_226)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_231),
.Y(n_254)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_202),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_233),
.B(n_236),
.Y(n_263)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_196),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_216),
.B(n_189),
.C(n_188),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_201),
.Y(n_238)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_238),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_199),
.Y(n_240)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_240),
.Y(n_262)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_199),
.Y(n_242)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_220),
.B(n_186),
.Y(n_243)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_243),
.Y(n_269)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_212),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_244),
.B(n_207),
.Y(n_255)
);

AND2x2_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_0),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_194),
.B(n_0),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_219),
.Y(n_261)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_248),
.B(n_258),
.C(n_259),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_223),
.B(n_215),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_249),
.B(n_253),
.Y(n_275)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_250),
.Y(n_278)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_224),
.B(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_255),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g256 ( 
.A(n_246),
.B(n_195),
.Y(n_256)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_257),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_246),
.B(n_213),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_224),
.B(n_212),
.C(n_213),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_226),
.B(n_209),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_261),
.B(n_266),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_235),
.A2(n_221),
.B1(n_230),
.B2(n_229),
.Y(n_264)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_221),
.B1(n_231),
.B2(n_243),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g265 ( 
.A(n_225),
.B(n_204),
.Y(n_265)
);

AOI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_265),
.A2(n_268),
.B1(n_234),
.B2(n_227),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g266 ( 
.A(n_222),
.B(n_192),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_SL g268 ( 
.A(n_234),
.B(n_192),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_261),
.B(n_232),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_270),
.B(n_274),
.Y(n_296)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_263),
.Y(n_271)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_271),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_252),
.B(n_239),
.C(n_237),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_250),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g291 ( 
.A(n_276),
.B(n_281),
.Y(n_291)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_258),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_279),
.B(n_280),
.Y(n_289)
);

INVx1_ASAP7_75t_SL g280 ( 
.A(n_251),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_252),
.B(n_239),
.C(n_230),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_260),
.Y(n_282)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_282),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_269),
.B(n_247),
.Y(n_284)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_284),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_285),
.A2(n_262),
.B1(n_254),
.B2(n_280),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_286),
.B(n_268),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g287 ( 
.A(n_272),
.B(n_256),
.Y(n_287)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_287),
.B(n_297),
.Y(n_302)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_288),
.Y(n_309)
);

AOI221xp5_ASAP7_75t_L g292 ( 
.A1(n_283),
.A2(n_265),
.B1(n_259),
.B2(n_241),
.C(n_257),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_292),
.B(n_9),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_228),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_295),
.B(n_299),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_SL g298 ( 
.A1(n_286),
.A2(n_267),
.B1(n_240),
.B2(n_227),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g303 ( 
.A1(n_298),
.A2(n_300),
.B1(n_279),
.B2(n_277),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_L g299 ( 
.A(n_273),
.B(n_278),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_282),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_274),
.B(n_248),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_301),
.B(n_272),
.C(n_275),
.Y(n_304)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_303),
.B(n_307),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_304),
.B(n_312),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_305),
.B(n_311),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_9),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_291),
.A2(n_9),
.B(n_13),
.Y(n_308)
);

OAI21xp5_ASAP7_75t_L g316 ( 
.A1(n_308),
.A2(n_293),
.B(n_7),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_289),
.B(n_296),
.C(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_310),
.B(n_314),
.C(n_11),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_8),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_289),
.B(n_10),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_294),
.A2(n_10),
.B1(n_13),
.B2(n_12),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_313),
.B(n_11),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_7),
.C(n_12),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_306),
.B(n_290),
.Y(n_315)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_315),
.Y(n_325)
);

AOI31xp67_ASAP7_75t_L g328 ( 
.A1(n_316),
.A2(n_311),
.A3(n_16),
.B(n_5),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g317 ( 
.A1(n_309),
.A2(n_300),
.B(n_6),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_3),
.B(n_4),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_310),
.B(n_6),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_322),
.B(n_3),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_314),
.B(n_11),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_302),
.C(n_4),
.Y(n_331)
);

INVx11_ASAP7_75t_L g326 ( 
.A(n_324),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_320),
.B(n_307),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_327),
.B(n_329),
.Y(n_332)
);

NAND3xp33_ASAP7_75t_L g334 ( 
.A(n_328),
.B(n_331),
.C(n_3),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_330),
.A2(n_319),
.B1(n_323),
.B2(n_5),
.Y(n_333)
);

AOI21x1_ASAP7_75t_L g335 ( 
.A1(n_333),
.A2(n_334),
.B(n_326),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_336),
.B(n_320),
.Y(n_337)
);

AOI322xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_325),
.A3(n_327),
.B1(n_332),
.B2(n_321),
.C1(n_302),
.C2(n_326),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_338),
.Y(n_339)
);

OAI21xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_5),
.B(n_3),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g341 ( 
.A(n_340),
.B(n_4),
.Y(n_341)
);


endmodule