module fake_jpeg_2449_n_97 (n_13, n_21, n_1, n_10, n_23, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_24, n_26, n_9, n_5, n_11, n_17, n_25, n_2, n_12, n_8, n_15, n_7, n_97);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_24;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_97;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_57;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_22),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_11),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_3),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_26),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_13),
.B(n_19),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_4),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_23),
.Y(n_37)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_34),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_39)
);

OAI22xp33_ASAP7_75t_SL g47 ( 
.A1(n_39),
.A2(n_41),
.B1(n_29),
.B2(n_35),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_40),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_34),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

INVx5_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2x1_ASAP7_75t_L g48 ( 
.A(n_44),
.B(n_33),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_47),
.A2(n_28),
.B(n_44),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g54 ( 
.A(n_48),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_43),
.B(n_27),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_50),
.B(n_51),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_38),
.B(n_36),
.Y(n_51)
);

NOR4xp25_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_30),
.C(n_36),
.D(n_7),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_53),
.B(n_56),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_55),
.A2(n_49),
.B1(n_46),
.B2(n_28),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_51),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_45),
.A2(n_42),
.B1(n_40),
.B2(n_35),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_57),
.A2(n_49),
.B1(n_32),
.B2(n_17),
.Y(n_66)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_52),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_58),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_37),
.B(n_29),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_59),
.B(n_5),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_61),
.Y(n_72)
);

NAND2x1_ASAP7_75t_SL g62 ( 
.A(n_45),
.B(n_28),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_62),
.B(n_6),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_63),
.A2(n_65),
.B1(n_69),
.B2(n_16),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_64),
.B(n_70),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g65 ( 
.A1(n_57),
.A2(n_49),
.B1(n_46),
.B2(n_28),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_66),
.A2(n_54),
.B1(n_59),
.B2(n_61),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_54),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_8),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_71),
.B(n_15),
.Y(n_77)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_72),
.Y(n_73)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_73),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_77),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_63),
.A2(n_62),
.B1(n_58),
.B2(n_9),
.Y(n_75)
);

INVxp67_ASAP7_75t_L g84 ( 
.A(n_75),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_65),
.A2(n_18),
.B1(n_24),
.B2(n_14),
.Y(n_76)
);

XNOR2xp5_ASAP7_75t_L g86 ( 
.A(n_76),
.B(n_79),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_78),
.B(n_81),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_67),
.B(n_9),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_64),
.A2(n_10),
.B(n_20),
.Y(n_82)
);

NOR4xp25_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_21),
.C(n_25),
.D(n_10),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_89),
.B(n_90),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_88),
.B(n_80),
.C(n_82),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_91),
.A2(n_83),
.B(n_80),
.Y(n_92)
);

OAI31xp33_ASAP7_75t_L g93 ( 
.A1(n_92),
.A2(n_87),
.A3(n_82),
.B(n_74),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_93),
.A2(n_86),
.B(n_84),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_84),
.C(n_76),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_66),
.B(n_68),
.Y(n_96)
);

BUFx24_ASAP7_75t_SL g97 ( 
.A(n_96),
.Y(n_97)
);


endmodule