module fake_netlist_5_462_n_3322 (n_54, n_29, n_16, n_43, n_0, n_12, n_9, n_47, n_58, n_36, n_25, n_53, n_18, n_27, n_42, n_64, n_22, n_1, n_8, n_45, n_10, n_24, n_28, n_46, n_21, n_44, n_40, n_34, n_62, n_38, n_61, n_4, n_32, n_35, n_41, n_65, n_56, n_51, n_63, n_11, n_17, n_19, n_57, n_7, n_37, n_59, n_15, n_26, n_30, n_20, n_5, n_33, n_55, n_14, n_48, n_2, n_31, n_23, n_13, n_50, n_66, n_3, n_49, n_52, n_60, n_6, n_39, n_3322);

input n_54;
input n_29;
input n_16;
input n_43;
input n_0;
input n_12;
input n_9;
input n_47;
input n_58;
input n_36;
input n_25;
input n_53;
input n_18;
input n_27;
input n_42;
input n_64;
input n_22;
input n_1;
input n_8;
input n_45;
input n_10;
input n_24;
input n_28;
input n_46;
input n_21;
input n_44;
input n_40;
input n_34;
input n_62;
input n_38;
input n_61;
input n_4;
input n_32;
input n_35;
input n_41;
input n_65;
input n_56;
input n_51;
input n_63;
input n_11;
input n_17;
input n_19;
input n_57;
input n_7;
input n_37;
input n_59;
input n_15;
input n_26;
input n_30;
input n_20;
input n_5;
input n_33;
input n_55;
input n_14;
input n_48;
input n_2;
input n_31;
input n_23;
input n_13;
input n_50;
input n_66;
input n_3;
input n_49;
input n_52;
input n_60;
input n_6;
input n_39;

output n_3322;

wire n_924;
wire n_1263;
wire n_3304;
wire n_977;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_611;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_469;
wire n_1508;
wire n_82;
wire n_2771;
wire n_785;
wire n_3241;
wire n_549;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_532;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_226;
wire n_1780;
wire n_3256;
wire n_1488;
wire n_667;
wire n_2899;
wire n_2955;
wire n_790;
wire n_1055;
wire n_2386;
wire n_1501;
wire n_111;
wire n_2395;
wire n_880;
wire n_3086;
wire n_3297;
wire n_544;
wire n_1007;
wire n_2369;
wire n_155;
wire n_2927;
wire n_552;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2347;
wire n_2520;
wire n_2821;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_956;
wire n_564;
wire n_423;
wire n_1738;
wire n_2021;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_105;
wire n_3088;
wire n_1021;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_551;
wire n_2143;
wire n_2853;
wire n_2059;
wire n_1323;
wire n_1466;
wire n_688;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_800;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_2389;
wire n_671;
wire n_819;
wire n_1451;
wire n_1022;
wire n_2302;
wire n_915;
wire n_1545;
wire n_2374;
wire n_864;
wire n_173;
wire n_859;
wire n_951;
wire n_1947;
wire n_1264;
wire n_2114;
wire n_447;
wire n_247;
wire n_2001;
wire n_1494;
wire n_292;
wire n_625;
wire n_854;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_1580;
wire n_674;
wire n_417;
wire n_1939;
wire n_2486;
wire n_1806;
wire n_516;
wire n_933;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_497;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_606;
wire n_3019;
wire n_275;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_877;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_755;
wire n_1118;
wire n_1686;
wire n_947;
wire n_1285;
wire n_373;
wire n_307;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_530;
wire n_87;
wire n_150;
wire n_1107;
wire n_1728;
wire n_556;
wire n_2076;
wire n_3036;
wire n_2482;
wire n_2031;
wire n_2677;
wire n_1230;
wire n_668;
wire n_375;
wire n_301;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_929;
wire n_3010;
wire n_3180;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_902;
wire n_1576;
wire n_191;
wire n_1705;
wire n_1294;
wire n_659;
wire n_1104;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_171;
wire n_1182;
wire n_3188;
wire n_3107;
wire n_579;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_938;
wire n_1098;
wire n_2963;
wire n_2142;
wire n_3186;
wire n_3082;
wire n_320;
wire n_1154;
wire n_2189;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_406;
wire n_519;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1016;
wire n_1243;
wire n_546;
wire n_2959;
wire n_101;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_1845;
wire n_281;
wire n_240;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_291;
wire n_231;
wire n_257;
wire n_2761;
wire n_731;
wire n_371;
wire n_1483;
wire n_2888;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_709;
wire n_1490;
wire n_317;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_569;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_227;
wire n_2306;
wire n_920;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2635;
wire n_2652;
wire n_94;
wire n_335;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_1669;
wire n_2566;
wire n_370;
wire n_976;
wire n_1949;
wire n_343;
wire n_1449;
wire n_308;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_297;
wire n_2587;
wire n_156;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_775;
wire n_219;
wire n_3060;
wire n_157;
wire n_2651;
wire n_600;
wire n_1484;
wire n_2071;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_223;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_2099;
wire n_2408;
wire n_264;
wire n_1877;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_955;
wire n_1850;
wire n_163;
wire n_3028;
wire n_339;
wire n_1146;
wire n_882;
wire n_183;
wire n_243;
wire n_2384;
wire n_1036;
wire n_1097;
wire n_1749;
wire n_347;
wire n_3156;
wire n_550;
wire n_696;
wire n_3101;
wire n_897;
wire n_215;
wire n_350;
wire n_196;
wire n_798;
wire n_646;
wire n_1428;
wire n_2663;
wire n_436;
wire n_1394;
wire n_2659;
wire n_1414;
wire n_1216;
wire n_290;
wire n_580;
wire n_2693;
wire n_1040;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_1852;
wire n_2159;
wire n_578;
wire n_2976;
wire n_926;
wire n_2249;
wire n_2180;
wire n_344;
wire n_2353;
wire n_1218;
wire n_2439;
wire n_1931;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_422;
wire n_475;
wire n_777;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_1030;
wire n_72;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_415;
wire n_1071;
wire n_485;
wire n_1561;
wire n_1267;
wire n_1165;
wire n_496;
wire n_1801;
wire n_1391;
wire n_958;
wire n_1034;
wire n_670;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_1600;
wire n_521;
wire n_663;
wire n_845;
wire n_2235;
wire n_1862;
wire n_673;
wire n_837;
wire n_1239;
wire n_2915;
wire n_528;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_680;
wire n_1473;
wire n_1587;
wire n_2682;
wire n_395;
wire n_164;
wire n_553;
wire n_901;
wire n_2432;
wire n_813;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_214;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_675;
wire n_2699;
wire n_888;
wire n_1880;
wire n_2769;
wire n_2337;
wire n_1167;
wire n_1626;
wire n_637;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_184;
wire n_446;
wire n_1863;
wire n_1064;
wire n_144;
wire n_858;
wire n_2079;
wire n_2238;
wire n_114;
wire n_96;
wire n_923;
wire n_2118;
wire n_691;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_881;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_468;
wire n_213;
wire n_129;
wire n_342;
wire n_2932;
wire n_2753;
wire n_464;
wire n_2980;
wire n_363;
wire n_1582;
wire n_197;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_1459;
wire n_460;
wire n_889;
wire n_2358;
wire n_973;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_477;
wire n_3191;
wire n_571;
wire n_1585;
wire n_461;
wire n_2684;
wire n_2712;
wire n_3193;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3273;
wire n_2713;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_907;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_190;
wire n_989;
wire n_2544;
wire n_1039;
wire n_2214;
wire n_2055;
wire n_228;
wire n_283;
wire n_3025;
wire n_1403;
wire n_2248;
wire n_2356;
wire n_488;
wire n_736;
wire n_892;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1000;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_1002;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_310;
wire n_3310;
wire n_593;
wire n_2258;
wire n_748;
wire n_586;
wire n_1058;
wire n_1667;
wire n_838;
wire n_2784;
wire n_2919;
wire n_332;
wire n_3092;
wire n_1053;
wire n_1224;
wire n_2865;
wire n_349;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_230;
wire n_1331;
wire n_953;
wire n_279;
wire n_1014;
wire n_1241;
wire n_70;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_289;
wire n_963;
wire n_1052;
wire n_954;
wire n_627;
wire n_1385;
wire n_440;
wire n_793;
wire n_478;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_476;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_534;
wire n_3106;
wire n_1882;
wire n_884;
wire n_345;
wire n_944;
wire n_1754;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_91;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_2828;
wire n_1809;
wire n_1856;
wire n_182;
wire n_143;
wire n_647;
wire n_237;
wire n_407;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_857;
wire n_832;
wire n_2305;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_207;
wire n_561;
wire n_1319;
wire n_2379;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_1027;
wire n_971;
wire n_1156;
wire n_117;
wire n_326;
wire n_794;
wire n_404;
wire n_2798;
wire n_2331;
wire n_2945;
wire n_2293;
wire n_686;
wire n_2837;
wire n_847;
wire n_1393;
wire n_2319;
wire n_596;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_2762;
wire n_558;
wire n_2808;
wire n_702;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_822;
wire n_1412;
wire n_2679;
wire n_1709;
wire n_2676;
wire n_2108;
wire n_728;
wire n_266;
wire n_1162;
wire n_272;
wire n_1538;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3116;
wire n_352;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_1038;
wire n_2967;
wire n_520;
wire n_1369;
wire n_409;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_887;
wire n_1905;
wire n_2553;
wire n_154;
wire n_3207;
wire n_2581;
wire n_71;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_300;
wire n_2698;
wire n_809;
wire n_870;
wire n_931;
wire n_599;
wire n_1711;
wire n_1662;
wire n_1891;
wire n_1481;
wire n_2626;
wire n_3042;
wire n_1942;
wire n_434;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_868;
wire n_2454;
wire n_639;
wire n_2804;
wire n_914;
wire n_2120;
wire n_411;
wire n_414;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_965;
wire n_1876;
wire n_1743;
wire n_935;
wire n_817;
wire n_121;
wire n_1175;
wire n_2763;
wire n_360;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_2009;
wire n_1888;
wire n_759;
wire n_2222;
wire n_1892;
wire n_806;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_1477;
wire n_3142;
wire n_324;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_187;
wire n_1189;
wire n_2690;
wire n_103;
wire n_97;
wire n_2215;
wire n_1259;
wire n_1690;
wire n_706;
wire n_746;
wire n_1649;
wire n_3150;
wire n_747;
wire n_2064;
wire n_784;
wire n_110;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_2413;
wire n_431;
wire n_1194;
wire n_1925;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_615;
wire n_851;
wire n_1759;
wire n_843;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_523;
wire n_913;
wire n_1537;
wire n_705;
wire n_865;
wire n_2227;
wire n_678;
wire n_2671;
wire n_697;
wire n_127;
wire n_1222;
wire n_75;
wire n_1679;
wire n_2190;
wire n_776;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_367;
wire n_2629;
wire n_2592;
wire n_452;
wire n_525;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_649;
wire n_547;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_1833;
wire n_116;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_284;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_139;
wire n_1734;
wire n_3038;
wire n_744;
wire n_590;
wire n_629;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_254;
wire n_1680;
wire n_1233;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_526;
wire n_1916;
wire n_3317;
wire n_293;
wire n_372;
wire n_677;
wire n_244;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_314;
wire n_368;
wire n_433;
wire n_604;
wire n_2007;
wire n_3220;
wire n_949;
wire n_2539;
wire n_3263;
wire n_100;
wire n_2582;
wire n_1443;
wire n_1008;
wire n_946;
wire n_1539;
wire n_2736;
wire n_1001;
wire n_1503;
wire n_2054;
wire n_498;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_1866;
wire n_689;
wire n_3158;
wire n_738;
wire n_1624;
wire n_3000;
wire n_640;
wire n_1510;
wire n_252;
wire n_624;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_295;
wire n_133;
wire n_1010;
wire n_3113;
wire n_1231;
wire n_739;
wire n_1406;
wire n_1279;
wire n_3108;
wire n_1994;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_610;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_936;
wire n_568;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_757;
wire n_3280;
wire n_2342;
wire n_633;
wire n_2856;
wire n_439;
wire n_106;
wire n_1832;
wire n_259;
wire n_448;
wire n_1851;
wire n_758;
wire n_999;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3003;
wire n_1933;
wire n_2290;
wire n_93;
wire n_1656;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_563;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_1145;
wire n_878;
wire n_524;
wire n_204;
wire n_394;
wire n_1678;
wire n_1049;
wire n_1153;
wire n_2145;
wire n_741;
wire n_1639;
wire n_1306;
wire n_1068;
wire n_3030;
wire n_1871;
wire n_2580;
wire n_2545;
wire n_2787;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_122;
wire n_331;
wire n_906;
wire n_1163;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_919;
wire n_908;
wire n_2412;
wire n_2406;
wire n_90;
wire n_2846;
wire n_724;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_2035;
wire n_658;
wire n_2061;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_456;
wire n_959;
wire n_2459;
wire n_3031;
wire n_535;
wire n_152;
wire n_940;
wire n_1445;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_592;
wire n_3243;
wire n_1169;
wire n_1692;
wire n_1596;
wire n_2666;
wire n_2982;
wire n_1017;
wire n_2481;
wire n_2947;
wire n_2171;
wire n_123;
wire n_978;
wire n_2768;
wire n_2314;
wire n_2116;
wire n_1434;
wire n_1054;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_267;
wire n_514;
wire n_457;
wire n_1079;
wire n_1045;
wire n_1208;
wire n_2093;
wire n_2038;
wire n_2320;
wire n_2473;
wire n_3287;
wire n_2137;
wire n_603;
wire n_1431;
wire n_2583;
wire n_484;
wire n_1593;
wire n_1033;
wire n_442;
wire n_2299;
wire n_131;
wire n_2540;
wire n_2873;
wire n_636;
wire n_660;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_1009;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_109;
wire n_742;
wire n_750;
wire n_2029;
wire n_995;
wire n_454;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_374;
wire n_3021;
wire n_1989;
wire n_185;
wire n_2359;
wire n_2941;
wire n_396;
wire n_1887;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_255;
wire n_2346;
wire n_2457;
wire n_662;
wire n_459;
wire n_2312;
wire n_218;
wire n_962;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_723;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_2339;
wire n_1336;
wire n_2882;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_473;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_1043;
wire n_2585;
wire n_355;
wire n_486;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_614;
wire n_337;
wire n_1421;
wire n_88;
wire n_2571;
wire n_1286;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_168;
wire n_974;
wire n_2565;
wire n_727;
wire n_1159;
wire n_957;
wire n_773;
wire n_208;
wire n_142;
wire n_2124;
wire n_743;
wire n_3001;
wire n_2081;
wire n_299;
wire n_303;
wire n_3149;
wire n_296;
wire n_613;
wire n_1119;
wire n_2156;
wire n_1240;
wire n_2729;
wire n_1820;
wire n_2261;
wire n_3268;
wire n_2418;
wire n_829;
wire n_2519;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_2897;
wire n_2077;
wire n_1416;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_361;
wire n_700;
wire n_1237;
wire n_573;
wire n_69;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_388;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_761;
wire n_2477;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_1006;
wire n_2110;
wire n_329;
wire n_274;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_582;
wire n_1332;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_73;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_309;
wire n_512;
wire n_2367;
wire n_2033;
wire n_1591;
wire n_84;
wire n_130;
wire n_322;
wire n_1682;
wire n_2628;
wire n_2390;
wire n_1980;
wire n_1249;
wire n_2896;
wire n_652;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_288;
wire n_2400;
wire n_1031;
wire n_263;
wire n_609;
wire n_1041;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_224;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_383;
wire n_3103;
wire n_834;
wire n_112;
wire n_765;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_893;
wire n_1015;
wire n_1140;
wire n_891;
wire n_1651;
wire n_1965;
wire n_239;
wire n_630;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_504;
wire n_1823;
wire n_511;
wire n_874;
wire n_2464;
wire n_358;
wire n_1101;
wire n_2831;
wire n_77;
wire n_102;
wire n_1106;
wire n_1456;
wire n_2230;
wire n_2015;
wire n_2365;
wire n_1982;
wire n_1875;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_987;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_261;
wire n_174;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_767;
wire n_993;
wire n_2490;
wire n_1903;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_545;
wire n_441;
wire n_860;
wire n_3229;
wire n_450;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_429;
wire n_948;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_628;
wire n_365;
wire n_1849;
wire n_2410;
wire n_729;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_970;
wire n_1935;
wire n_911;
wire n_2922;
wire n_1430;
wire n_83;
wire n_3275;
wire n_2645;
wire n_2467;
wire n_513;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_560;
wire n_1534;
wire n_340;
wire n_2288;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_1044;
wire n_2436;
wire n_346;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_495;
wire n_602;
wire n_574;
wire n_2593;
wire n_1435;
wire n_879;
wire n_2416;
wire n_2405;
wire n_623;
wire n_3286;
wire n_2088;
wire n_405;
wire n_2953;
wire n_824;
wire n_359;
wire n_1645;
wire n_2461;
wire n_490;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_996;
wire n_921;
wire n_1684;
wire n_233;
wire n_2658;
wire n_1717;
wire n_572;
wire n_366;
wire n_2895;
wire n_815;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_128;
wire n_1821;
wire n_120;
wire n_2929;
wire n_327;
wire n_135;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_1037;
wire n_2368;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_2890;
wire n_3059;
wire n_2554;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_426;
wire n_1438;
wire n_1082;
wire n_1840;
wire n_589;
wire n_716;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_562;
wire n_1436;
wire n_1691;
wire n_952;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_391;
wire n_701;
wire n_1437;
wire n_1023;
wire n_2075;
wire n_645;
wire n_539;
wire n_803;
wire n_1092;
wire n_2694;
wire n_238;
wire n_1776;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2789;
wire n_2131;
wire n_3026;
wire n_2216;
wire n_531;
wire n_3020;
wire n_1757;
wire n_890;
wire n_1897;
wire n_764;
wire n_1919;
wire n_1056;
wire n_1424;
wire n_162;
wire n_960;
wire n_2933;
wire n_2308;
wire n_1893;
wire n_2910;
wire n_222;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_1047;
wire n_2053;
wire n_2163;
wire n_634;
wire n_2328;
wire n_199;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_348;
wire n_1382;
wire n_1029;
wire n_925;
wire n_1206;
wire n_424;
wire n_2647;
wire n_3160;
wire n_1311;
wire n_2969;
wire n_2864;
wire n_2191;
wire n_3195;
wire n_1519;
wire n_256;
wire n_950;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_380;
wire n_419;
wire n_1346;
wire n_3053;
wire n_444;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_316;
wire n_2266;
wire n_389;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_418;
wire n_248;
wire n_136;
wire n_146;
wire n_86;
wire n_912;
wire n_315;
wire n_968;
wire n_451;
wire n_619;
wire n_408;
wire n_2440;
wire n_1386;
wire n_1699;
wire n_376;
wire n_967;
wire n_1442;
wire n_2923;
wire n_2541;
wire n_74;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_515;
wire n_2333;
wire n_351;
wire n_885;
wire n_2916;
wire n_3166;
wire n_397;
wire n_1432;
wire n_1357;
wire n_483;
wire n_2125;
wire n_683;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1057;
wire n_1051;
wire n_1085;
wire n_1066;
wire n_721;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_1050;
wire n_841;
wire n_802;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_983;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_2870;
wire n_280;
wire n_1305;
wire n_3178;
wire n_873;
wire n_1826;
wire n_378;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_762;
wire n_1283;
wire n_1644;
wire n_2637;
wire n_2334;
wire n_690;
wire n_1974;
wire n_2463;
wire n_583;
wire n_2086;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_302;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_2881;
wire n_1203;
wire n_1631;
wire n_3282;
wire n_2472;
wire n_821;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_1768;
wire n_321;
wire n_2294;
wire n_1179;
wire n_621;
wire n_753;
wire n_2475;
wire n_2733;
wire n_455;
wire n_1048;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_212;
wire n_385;
wire n_2785;
wire n_2556;
wire n_507;
wire n_2269;
wire n_2732;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3274;
wire n_3041;
wire n_3299;
wire n_2646;
wire n_1560;
wire n_1605;
wire n_2236;
wire n_330;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_972;
wire n_692;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_820;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_2460;
wire n_2589;
wire n_3203;
wire n_1301;
wire n_1363;
wire n_1668;
wire n_1185;
wire n_991;
wire n_2903;
wire n_828;
wire n_1967;
wire n_779;
wire n_576;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_804;
wire n_537;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_945;
wire n_2997;
wire n_492;
wire n_153;
wire n_1504;
wire n_943;
wire n_341;
wire n_250;
wire n_992;
wire n_3067;
wire n_1932;
wire n_2755;
wire n_543;
wire n_260;
wire n_842;
wire n_650;
wire n_984;
wire n_694;
wire n_3237;
wire n_2082;
wire n_286;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_883;
wire n_1983;
wire n_3167;
wire n_470;
wire n_325;
wire n_449;
wire n_1594;
wire n_132;
wire n_1214;
wire n_1342;
wire n_1400;
wire n_900;
wire n_2362;
wire n_856;
wire n_2609;
wire n_1793;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_918;
wire n_942;
wire n_2169;
wire n_1804;
wire n_189;
wire n_1147;
wire n_1557;
wire n_1977;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1422;
wire n_1077;
wire n_3196;
wire n_3078;
wire n_2533;
wire n_2364;
wire n_540;
wire n_618;
wire n_3094;
wire n_896;
wire n_2310;
wire n_2780;
wire n_323;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_195;
wire n_356;
wire n_2291;
wire n_3099;
wire n_2596;
wire n_894;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_831;
wire n_2280;
wire n_2192;
wire n_964;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_234;
wire n_1575;
wire n_1735;
wire n_1697;
wire n_833;
wire n_2318;
wire n_2393;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_225;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_988;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_814;
wire n_2751;
wire n_2793;
wire n_2707;
wire n_192;
wire n_2971;
wire n_1549;
wire n_2311;
wire n_1934;
wire n_1201;
wire n_1114;
wire n_655;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_669;
wire n_472;
wire n_1458;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_2471;
wire n_1807;
wire n_387;
wire n_1149;
wire n_2618;
wire n_398;
wire n_1671;
wire n_635;
wire n_2559;
wire n_763;
wire n_3230;
wire n_1020;
wire n_1062;
wire n_211;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_1204;
wire n_2840;
wire n_2810;
wire n_2325;
wire n_178;
wire n_2747;
wire n_2446;
wire n_1814;
wire n_1035;
wire n_2822;
wire n_287;
wire n_555;
wire n_783;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_661;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_849;
wire n_2795;
wire n_336;
wire n_584;
wire n_681;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_430;
wire n_2002;
wire n_2282;
wire n_510;
wire n_2800;
wire n_216;
wire n_2371;
wire n_2935;
wire n_311;
wire n_3233;
wire n_3177;
wire n_830;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_2352;
wire n_1413;
wire n_801;
wire n_2207;
wire n_2080;
wire n_2619;
wire n_2377;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_241;
wire n_875;
wire n_357;
wire n_1110;
wire n_1655;
wire n_445;
wire n_2641;
wire n_3198;
wire n_749;
wire n_1895;
wire n_3123;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_717;
wire n_165;
wire n_939;
wire n_482;
wire n_2361;
wire n_1088;
wire n_588;
wire n_1173;
wire n_789;
wire n_1232;
wire n_1603;
wire n_734;
wire n_638;
wire n_2638;
wire n_866;
wire n_107;
wire n_969;
wire n_1401;
wire n_2492;
wire n_1019;
wire n_1105;
wire n_249;
wire n_1998;
wire n_304;
wire n_1338;
wire n_577;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_338;
wire n_149;
wire n_1653;
wire n_693;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_836;
wire n_990;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_975;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_567;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_778;
wire n_1122;
wire n_151;
wire n_3192;
wire n_2608;
wire n_306;
wire n_2657;
wire n_770;
wire n_458;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_2649;
wire n_1102;
wire n_2852;
wire n_2392;
wire n_3093;
wire n_1843;
wire n_711;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_85;
wire n_1187;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1392;
wire n_1597;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1834;
wire n_1659;
wire n_2097;
wire n_2313;
wire n_2542;
wire n_489;
wire n_1174;
wire n_2431;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_617;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_876;
wire n_1516;
wire n_1190;
wire n_1736;
wire n_1685;
wire n_118;
wire n_2409;
wire n_601;
wire n_917;
wire n_1714;
wire n_966;
wire n_253;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_206;
wire n_172;
wire n_217;
wire n_726;
wire n_3174;
wire n_982;
wire n_2575;
wire n_2988;
wire n_1573;
wire n_1453;
wire n_1731;
wire n_2217;
wire n_818;
wire n_2373;
wire n_1970;
wire n_861;
wire n_1713;
wire n_1183;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_899;
wire n_1253;
wire n_210;
wire n_1737;
wire n_2201;
wire n_2722;
wire n_2117;
wire n_2745;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_774;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_1335;
wire n_1777;
wire n_1514;
wire n_1957;
wire n_1345;
wire n_1059;
wire n_176;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_1899;
wire n_3226;
wire n_557;
wire n_1410;
wire n_1005;
wire n_607;
wire n_1003;
wire n_679;
wire n_710;
wire n_3090;
wire n_2067;
wire n_527;
wire n_1168;
wire n_707;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_2877;
wire n_3318;
wire n_2148;
wire n_937;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_393;
wire n_108;
wire n_487;
wire n_1726;
wire n_665;
wire n_1835;
wire n_1584;
wire n_3035;
wire n_1440;
wire n_177;
wire n_2164;
wire n_421;
wire n_1988;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_910;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_768;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_205;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_754;
wire n_2811;
wire n_1496;
wire n_179;
wire n_1125;
wire n_125;
wire n_410;
wire n_2547;
wire n_3014;
wire n_708;
wire n_529;
wire n_1812;
wire n_735;
wire n_2501;
wire n_3079;
wire n_232;
wire n_1915;
wire n_1109;
wire n_126;
wire n_895;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_2121;
wire n_1803;
wire n_202;
wire n_3308;
wire n_2665;
wire n_427;
wire n_1399;
wire n_1991;
wire n_1543;
wire n_1979;
wire n_791;
wire n_732;
wire n_1533;
wire n_2224;
wire n_193;
wire n_2924;
wire n_808;
wire n_2484;
wire n_797;
wire n_1025;
wire n_1930;
wire n_1955;
wire n_2765;
wire n_500;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_148;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_435;
wire n_2003;
wire n_159;
wire n_766;
wire n_1457;
wire n_541;
wire n_2692;
wire n_3148;
wire n_538;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_799;
wire n_2264;
wire n_2754;
wire n_687;
wire n_715;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_536;
wire n_872;
wire n_2012;
wire n_594;
wire n_200;
wire n_1291;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_1155;
wire n_1418;
wire n_89;
wire n_1972;
wire n_1524;
wire n_1689;
wire n_1485;
wire n_2806;
wire n_115;
wire n_1011;
wire n_1184;
wire n_2184;
wire n_985;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_869;
wire n_810;
wire n_2965;
wire n_416;
wire n_827;
wire n_3217;
wire n_401;
wire n_1703;
wire n_3312;
wire n_1352;
wire n_2926;
wire n_626;
wire n_2197;
wire n_2199;
wire n_1650;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_305;
wire n_2023;
wire n_2213;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_137;
wire n_676;
wire n_294;
wire n_318;
wire n_2103;
wire n_653;
wire n_2160;
wire n_642;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_194;
wire n_855;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_850;
wire n_684;
wire n_3074;
wire n_124;
wire n_3204;
wire n_268;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_664;
wire n_1999;
wire n_503;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_2480;
wire n_235;
wire n_1372;
wire n_2861;
wire n_605;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_353;
wire n_620;
wire n_643;
wire n_2430;
wire n_2363;
wire n_916;
wire n_1081;
wire n_2549;
wire n_493;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_703;
wire n_698;
wire n_980;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_780;
wire n_2977;
wire n_2601;
wire n_3043;
wire n_998;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_467;
wire n_1227;
wire n_1531;
wire n_840;
wire n_1334;
wire n_1907;
wire n_501;
wire n_823;
wire n_245;
wire n_2686;
wire n_2528;
wire n_725;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_672;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3315;
wire n_581;
wire n_2906;
wire n_382;
wire n_554;
wire n_1625;
wire n_2130;
wire n_2187;
wire n_2284;
wire n_898;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_1762;
wire n_1013;
wire n_1452;
wire n_718;
wire n_2687;
wire n_265;
wire n_3023;
wire n_1120;
wire n_719;
wire n_443;
wire n_1791;
wire n_198;
wire n_1890;
wire n_1747;
wire n_714;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_909;
wire n_1944;
wire n_1497;
wire n_1530;
wire n_2654;
wire n_997;
wire n_3104;
wire n_932;
wire n_3169;
wire n_3151;
wire n_612;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_788;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_119;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_559;
wire n_825;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_508;
wire n_2186;
wire n_506;
wire n_1320;
wire n_1663;
wire n_737;
wire n_1718;
wire n_986;
wire n_2315;
wire n_509;
wire n_3228;
wire n_1317;
wire n_147;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_2562;
wire n_1281;
wire n_67;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_1024;
wire n_1063;
wire n_1889;
wire n_209;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_733;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_941;
wire n_2326;
wire n_981;
wire n_2560;
wire n_1569;
wire n_2188;
wire n_68;
wire n_867;
wire n_186;
wire n_2348;
wire n_2422;
wire n_134;
wire n_2239;
wire n_587;
wire n_2950;
wire n_792;
wire n_756;
wire n_1429;
wire n_399;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_548;
wire n_3170;
wire n_812;
wire n_298;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_518;
wire n_505;
wire n_2057;
wire n_3272;
wire n_3011;
wire n_1772;
wire n_282;
wire n_752;
wire n_905;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_782;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_862;
wire n_1425;
wire n_760;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_381;
wire n_2889;
wire n_220;
wire n_390;
wire n_1330;
wire n_1867;
wire n_1945;
wire n_2772;
wire n_481;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_769;
wire n_2497;
wire n_2006;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1046;
wire n_271;
wire n_934;
wire n_1618;
wire n_2260;
wire n_826;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_886;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_654;
wire n_1172;
wire n_167;
wire n_2535;
wire n_379;
wire n_428;
wire n_1341;
wire n_2774;
wire n_570;
wire n_2726;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_853;
wire n_3062;
wire n_3161;
wire n_377;
wire n_2317;
wire n_751;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_786;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_392;
wire n_2579;
wire n_3017;
wire n_158;
wire n_2476;
wire n_704;
wire n_787;
wire n_1770;
wire n_138;
wire n_2781;
wire n_2456;
wire n_961;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_771;
wire n_2778;
wire n_276;
wire n_95;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_169;
wire n_2887;
wire n_522;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_400;
wire n_930;
wire n_181;
wire n_1873;
wire n_1411;
wire n_3201;
wire n_3054;
wire n_221;
wire n_622;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_1087;
wire n_2526;
wire n_2854;
wire n_386;
wire n_994;
wire n_1701;
wire n_2194;
wire n_848;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_104;
wire n_682;
wire n_1567;
wire n_141;
wire n_2567;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_922;
wire n_3122;
wire n_816;
wire n_1648;
wire n_591;
wire n_145;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_313;
wire n_631;
wire n_479;
wire n_1246;
wire n_1339;
wire n_1478;
wire n_1797;
wire n_432;
wire n_1769;
wire n_2957;
wire n_839;
wire n_1210;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_328;
wire n_140;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_369;
wire n_1842;
wire n_871;
wire n_2442;
wire n_3309;
wire n_598;
wire n_685;
wire n_608;
wire n_928;
wire n_1367;
wire n_78;
wire n_1943;
wire n_1460;
wire n_772;
wire n_2018;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_499;
wire n_2531;
wire n_1589;
wire n_517;
wire n_98;
wire n_2961;
wire n_402;
wire n_413;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_796;
wire n_1858;
wire n_1619;
wire n_2815;
wire n_236;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1012;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_903;
wire n_2453;
wire n_1525;
wire n_1752;
wire n_2397;
wire n_740;
wire n_2883;
wire n_3115;
wire n_203;
wire n_384;
wire n_3076;
wire n_2208;
wire n_1404;
wire n_80;
wire n_3063;
wire n_2912;
wire n_1794;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_277;
wire n_1061;
wire n_3251;
wire n_92;
wire n_1910;
wire n_333;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_462;
wire n_2050;
wire n_2809;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_258;
wire n_1113;
wire n_3118;
wire n_79;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_1226;
wire n_722;
wire n_1277;
wire n_2591;
wire n_188;
wire n_2146;
wire n_844;
wire n_201;
wire n_471;
wire n_852;
wire n_1487;
wire n_1864;
wire n_1028;
wire n_1601;
wire n_781;
wire n_474;
wire n_2940;
wire n_542;
wire n_463;
wire n_1546;
wire n_595;
wire n_502;
wire n_466;
wire n_2612;
wire n_420;
wire n_1337;
wire n_1495;
wire n_632;
wire n_699;
wire n_979;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_1245;
wire n_846;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_465;
wire n_2832;
wire n_76;
wire n_362;
wire n_1321;
wire n_170;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_161;
wire n_273;
wire n_1937;
wire n_585;
wire n_2112;
wire n_3250;
wire n_1739;
wire n_3181;
wire n_270;
wire n_2958;
wire n_616;
wire n_2278;
wire n_81;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_745;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_648;
wire n_1379;
wire n_2734;
wire n_312;
wire n_2196;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_494;
wire n_1761;
wire n_641;
wire n_3238;
wire n_3210;
wire n_730;
wire n_3175;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_354;
wire n_575;
wire n_480;
wire n_425;
wire n_795;
wire n_2404;
wire n_2083;
wire n_695;
wire n_180;
wire n_3281;
wire n_656;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3266;
wire n_2485;
wire n_229;
wire n_1956;
wire n_1936;
wire n_437;
wire n_1642;
wire n_2279;
wire n_2655;
wire n_2027;
wire n_403;
wire n_453;
wire n_2642;
wire n_1130;
wire n_720;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_863;
wire n_2210;
wire n_805;
wire n_3247;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_2892;
wire n_3057;
wire n_3194;
wire n_3066;
wire n_113;
wire n_712;
wire n_2414;
wire n_2907;
wire n_246;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_1042;
wire n_1402;
wire n_2820;
wire n_269;
wire n_2049;
wire n_2273;
wire n_285;
wire n_412;
wire n_2719;
wire n_1493;
wire n_657;
wire n_644;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_491;
wire n_1258;
wire n_1074;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_251;
wire n_160;
wire n_566;
wire n_565;
wire n_2586;
wire n_1448;
wire n_2225;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_597;
wire n_1996;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_651;
wire n_1340;
wire n_2972;
wire n_2274;
wire n_334;
wire n_811;
wire n_1558;
wire n_3225;
wire n_807;
wire n_3321;
wire n_2166;
wire n_2938;
wire n_3212;
wire n_835;
wire n_175;
wire n_666;
wire n_3319;
wire n_262;
wire n_1433;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_99;
wire n_1254;
wire n_1026;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_319;
wire n_364;
wire n_1138;
wire n_927;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2044;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_1004;
wire n_1186;
wire n_242;
wire n_1032;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2991;
wire n_2010;
wire n_1018;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_2975;
wire n_438;
wire n_2599;
wire n_713;
wire n_2704;
wire n_904;
wire n_2839;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_166;
wire n_1180;
wire n_1827;
wire n_2524;
wire n_1271;
wire n_2802;
wire n_533;
wire n_1542;
wire n_1251;
wire n_3159;
wire n_278;
wire n_2728;
wire n_2268;

CKINVDCx5p33_ASAP7_75t_R g67 ( 
.A(n_58),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx5p33_ASAP7_75t_R g69 ( 
.A(n_47),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_50),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_48),
.Y(n_71)
);

CKINVDCx5p33_ASAP7_75t_R g72 ( 
.A(n_61),
.Y(n_72)
);

CKINVDCx5p33_ASAP7_75t_R g73 ( 
.A(n_27),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_66),
.Y(n_74)
);

CKINVDCx5p33_ASAP7_75t_R g75 ( 
.A(n_26),
.Y(n_75)
);

CKINVDCx5p33_ASAP7_75t_R g76 ( 
.A(n_23),
.Y(n_76)
);

CKINVDCx5p33_ASAP7_75t_R g77 ( 
.A(n_49),
.Y(n_77)
);

CKINVDCx5p33_ASAP7_75t_R g78 ( 
.A(n_7),
.Y(n_78)
);

CKINVDCx5p33_ASAP7_75t_R g79 ( 
.A(n_48),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_60),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_9),
.Y(n_81)
);

CKINVDCx5p33_ASAP7_75t_R g82 ( 
.A(n_56),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_49),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_41),
.Y(n_84)
);

CKINVDCx5p33_ASAP7_75t_R g85 ( 
.A(n_62),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_5),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_6),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_55),
.Y(n_88)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_1),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_12),
.Y(n_90)
);

CKINVDCx5p33_ASAP7_75t_R g91 ( 
.A(n_17),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_27),
.Y(n_92)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_20),
.Y(n_93)
);

BUFx3_ASAP7_75t_L g94 ( 
.A(n_11),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g95 ( 
.A(n_21),
.Y(n_95)
);

CKINVDCx5p33_ASAP7_75t_R g96 ( 
.A(n_52),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_30),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_30),
.Y(n_98)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_35),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_43),
.Y(n_100)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_44),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_24),
.Y(n_103)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_16),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_33),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g106 ( 
.A(n_13),
.Y(n_106)
);

CKINVDCx5p33_ASAP7_75t_R g107 ( 
.A(n_45),
.Y(n_107)
);

CKINVDCx5p33_ASAP7_75t_R g108 ( 
.A(n_15),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_33),
.Y(n_109)
);

CKINVDCx5p33_ASAP7_75t_R g110 ( 
.A(n_4),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_57),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_4),
.Y(n_112)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_21),
.Y(n_113)
);

CKINVDCx5p33_ASAP7_75t_R g114 ( 
.A(n_44),
.Y(n_114)
);

CKINVDCx5p33_ASAP7_75t_R g115 ( 
.A(n_32),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_16),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_39),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_23),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_1),
.Y(n_119)
);

CKINVDCx5p33_ASAP7_75t_R g120 ( 
.A(n_32),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_64),
.Y(n_121)
);

BUFx2_ASAP7_75t_L g122 ( 
.A(n_18),
.Y(n_122)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_29),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_3),
.Y(n_124)
);

CKINVDCx5p33_ASAP7_75t_R g125 ( 
.A(n_20),
.Y(n_125)
);

CKINVDCx5p33_ASAP7_75t_R g126 ( 
.A(n_45),
.Y(n_126)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_36),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_28),
.Y(n_128)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_50),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_41),
.Y(n_130)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_31),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_6),
.Y(n_132)
);

CKINVDCx5p33_ASAP7_75t_R g133 ( 
.A(n_37),
.Y(n_133)
);

INVxp33_ASAP7_75t_L g134 ( 
.A(n_122),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_99),
.Y(n_135)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_99),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_99),
.Y(n_137)
);

INVxp67_ASAP7_75t_SL g138 ( 
.A(n_93),
.Y(n_138)
);

CKINVDCx5p33_ASAP7_75t_R g139 ( 
.A(n_73),
.Y(n_139)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_74),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_99),
.Y(n_141)
);

INVxp33_ASAP7_75t_L g142 ( 
.A(n_122),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_122),
.Y(n_143)
);

CKINVDCx5p33_ASAP7_75t_R g144 ( 
.A(n_75),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_74),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_99),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_129),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_101),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_129),
.Y(n_150)
);

INVxp33_ASAP7_75t_L g151 ( 
.A(n_68),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_129),
.Y(n_152)
);

CKINVDCx5p33_ASAP7_75t_R g153 ( 
.A(n_76),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_129),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_135),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_135),
.Y(n_156)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_135),
.Y(n_157)
);

AND2x4_ASAP7_75t_L g158 ( 
.A(n_135),
.B(n_101),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_136),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_138),
.B(n_94),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_140),
.Y(n_161)
);

HB1xp67_ASAP7_75t_L g162 ( 
.A(n_143),
.Y(n_162)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_136),
.Y(n_164)
);

NAND2xp33_ASAP7_75t_L g165 ( 
.A(n_134),
.B(n_93),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_140),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_134),
.A2(n_117),
.B1(n_131),
.B2(n_130),
.Y(n_167)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_136),
.Y(n_168)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_140),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_140),
.B(n_121),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_137),
.Y(n_171)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_137),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_137),
.Y(n_173)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_137),
.Y(n_174)
);

HB1xp67_ASAP7_75t_L g175 ( 
.A(n_143),
.Y(n_175)
);

HB1xp67_ASAP7_75t_L g176 ( 
.A(n_143),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_121),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_145),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_141),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_145),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_141),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_145),
.B(n_94),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_141),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g184 ( 
.A(n_145),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g185 ( 
.A(n_141),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_145),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_146),
.Y(n_187)
);

AND2x2_ASAP7_75t_SL g188 ( 
.A(n_149),
.B(n_93),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_162),
.Y(n_190)
);

BUFx6f_ASAP7_75t_L g191 ( 
.A(n_185),
.Y(n_191)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_162),
.Y(n_192)
);

CKINVDCx6p67_ASAP7_75t_R g193 ( 
.A(n_162),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_185),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_167),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_167),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_167),
.Y(n_197)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_157),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_175),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_175),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_176),
.Y(n_203)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_157),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_176),
.Y(n_205)
);

BUFx10_ASAP7_75t_L g206 ( 
.A(n_160),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_176),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g208 ( 
.A(n_185),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_160),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g211 ( 
.A(n_160),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_185),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_188),
.Y(n_213)
);

HB1xp67_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_188),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_188),
.B(n_146),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_188),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_R g218 ( 
.A(n_165),
.B(n_139),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_188),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_188),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_157),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_182),
.Y(n_222)
);

AOI21x1_ASAP7_75t_L g223 ( 
.A1(n_170),
.A2(n_154),
.B(n_152),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_158),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_158),
.Y(n_225)
);

NAND2xp33_ASAP7_75t_R g226 ( 
.A(n_158),
.B(n_139),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g227 ( 
.A(n_158),
.B(n_144),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_158),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_158),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_158),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_182),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_170),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_158),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_170),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_177),
.B(n_144),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_177),
.Y(n_236)
);

BUFx16f_ASAP7_75t_R g237 ( 
.A(n_165),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_155),
.B(n_134),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_155),
.Y(n_239)
);

NAND2xp33_ASAP7_75t_R g240 ( 
.A(n_177),
.B(n_153),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_157),
.Y(n_241)
);

BUFx2_ASAP7_75t_L g242 ( 
.A(n_155),
.Y(n_242)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_157),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_155),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_156),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_R g246 ( 
.A(n_156),
.B(n_153),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_157),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_156),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_156),
.Y(n_249)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_159),
.A2(n_154),
.B(n_152),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_159),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_159),
.B(n_72),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g253 ( 
.A(n_159),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_164),
.Y(n_254)
);

BUFx2_ASAP7_75t_L g255 ( 
.A(n_164),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_164),
.B(n_111),
.Y(n_256)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_163),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_164),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_171),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_171),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_171),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_171),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_173),
.Y(n_263)
);

AND2x4_ASAP7_75t_L g264 ( 
.A(n_173),
.B(n_149),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_R g265 ( 
.A(n_173),
.B(n_80),
.Y(n_265)
);

INVx1_ASAP7_75t_SL g266 ( 
.A(n_173),
.Y(n_266)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_163),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_187),
.Y(n_268)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_187),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_187),
.Y(n_270)
);

INVxp33_ASAP7_75t_SL g271 ( 
.A(n_187),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_194),
.Y(n_272)
);

OR2x6_ASAP7_75t_L g273 ( 
.A(n_227),
.B(n_94),
.Y(n_273)
);

INVx2_ASAP7_75t_SL g274 ( 
.A(n_214),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_214),
.B(n_266),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_194),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_230),
.B(n_138),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_210),
.B(n_142),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_240),
.Y(n_279)
);

NAND2xp33_ASAP7_75t_SL g280 ( 
.A(n_218),
.B(n_80),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_191),
.Y(n_281)
);

INVx4_ASAP7_75t_SL g282 ( 
.A(n_191),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_200),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_163),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_213),
.A2(n_142),
.B1(n_67),
.B2(n_82),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_239),
.Y(n_286)
);

INVx4_ASAP7_75t_L g287 ( 
.A(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_200),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_209),
.Y(n_289)
);

NAND2x1p5_ASAP7_75t_L g290 ( 
.A(n_230),
.B(n_222),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_209),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_211),
.B(n_163),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_211),
.B(n_151),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_218),
.B(n_265),
.Y(n_294)
);

BUFx3_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

AND2x6_ASAP7_75t_L g296 ( 
.A(n_222),
.B(n_94),
.Y(n_296)
);

BUFx10_ASAP7_75t_L g297 ( 
.A(n_238),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_212),
.Y(n_298)
);

INVx2_ASAP7_75t_SL g299 ( 
.A(n_206),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_212),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_217),
.B(n_219),
.Y(n_301)
);

OR2x6_ASAP7_75t_L g302 ( 
.A(n_227),
.B(n_106),
.Y(n_302)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_191),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g304 ( 
.A(n_191),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_235),
.B(n_232),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_220),
.B(n_163),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_242),
.Y(n_307)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_255),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_239),
.Y(n_309)
);

INVx1_ASAP7_75t_SL g310 ( 
.A(n_203),
.Y(n_310)
);

BUFx2_ASAP7_75t_L g311 ( 
.A(n_236),
.Y(n_311)
);

INVx2_ASAP7_75t_L g312 ( 
.A(n_245),
.Y(n_312)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_245),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_249),
.Y(n_314)
);

INVx3_ASAP7_75t_L g315 ( 
.A(n_191),
.Y(n_315)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_249),
.Y(n_316)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_224),
.B(n_138),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_251),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_235),
.B(n_151),
.Y(n_319)
);

AND2x6_ASAP7_75t_L g320 ( 
.A(n_231),
.B(n_106),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_234),
.B(n_67),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_251),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_231),
.B(n_163),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_254),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_254),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_265),
.B(n_82),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_240),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_238),
.B(n_146),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_206),
.B(n_168),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g330 ( 
.A(n_190),
.B(n_146),
.Y(n_330)
);

INVx4_ASAP7_75t_L g331 ( 
.A(n_191),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_246),
.B(n_85),
.Y(n_332)
);

INVx1_ASAP7_75t_SL g333 ( 
.A(n_205),
.Y(n_333)
);

INVx4_ASAP7_75t_L g334 ( 
.A(n_191),
.Y(n_334)
);

CKINVDCx5p33_ASAP7_75t_R g335 ( 
.A(n_246),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_260),
.Y(n_336)
);

INVx3_ASAP7_75t_L g337 ( 
.A(n_208),
.Y(n_337)
);

BUFx3_ASAP7_75t_L g338 ( 
.A(n_255),
.Y(n_338)
);

INVx8_ASAP7_75t_L g339 ( 
.A(n_225),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_260),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_226),
.Y(n_341)
);

INVx2_ASAP7_75t_L g342 ( 
.A(n_263),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_SL g343 ( 
.A(n_236),
.B(n_85),
.Y(n_343)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_263),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g345 ( 
.A(n_208),
.Y(n_345)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_269),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_269),
.Y(n_347)
);

AO21x2_ASAP7_75t_L g348 ( 
.A1(n_216),
.A2(n_149),
.B(n_148),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_206),
.B(n_168),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g350 ( 
.A(n_190),
.B(n_147),
.Y(n_350)
);

NAND2xp33_ASAP7_75t_L g351 ( 
.A(n_228),
.B(n_149),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_253),
.A2(n_117),
.B1(n_84),
.B2(n_116),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_226),
.Y(n_353)
);

AND2x4_ASAP7_75t_L g354 ( 
.A(n_229),
.B(n_147),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_253),
.A2(n_84),
.B1(n_116),
.B2(n_87),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_244),
.B(n_147),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_264),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_271),
.B(n_95),
.Y(n_358)
);

INVx1_ASAP7_75t_SL g359 ( 
.A(n_202),
.Y(n_359)
);

BUFx3_ASAP7_75t_L g360 ( 
.A(n_233),
.Y(n_360)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_208),
.Y(n_361)
);

INVx5_ASAP7_75t_L g362 ( 
.A(n_208),
.Y(n_362)
);

AND2x4_ASAP7_75t_L g363 ( 
.A(n_216),
.B(n_147),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_264),
.Y(n_364)
);

INVxp33_ASAP7_75t_L g365 ( 
.A(n_192),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_264),
.Y(n_366)
);

INVx2_ASAP7_75t_L g367 ( 
.A(n_250),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_264),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_250),
.Y(n_369)
);

AND2x6_ASAP7_75t_L g370 ( 
.A(n_237),
.B(n_106),
.Y(n_370)
);

HB1xp67_ASAP7_75t_L g371 ( 
.A(n_192),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_206),
.B(n_168),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g373 ( 
.A(n_248),
.B(n_148),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_264),
.Y(n_374)
);

AND2x4_ASAP7_75t_L g375 ( 
.A(n_261),
.B(n_148),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_206),
.B(n_168),
.Y(n_376)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_268),
.B(n_168),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_223),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_270),
.B(n_77),
.Y(n_379)
);

INVx1_ASAP7_75t_SL g380 ( 
.A(n_202),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_193),
.B(n_148),
.Y(n_381)
);

AND2x2_ASAP7_75t_L g382 ( 
.A(n_193),
.B(n_150),
.Y(n_382)
);

BUFx2_ASAP7_75t_L g383 ( 
.A(n_193),
.Y(n_383)
);

HAxp5_ASAP7_75t_SL g384 ( 
.A(n_195),
.B(n_68),
.CON(n_384),
.SN(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_208),
.B(n_168),
.Y(n_385)
);

INVx5_ASAP7_75t_L g386 ( 
.A(n_208),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_223),
.Y(n_387)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_199),
.Y(n_388)
);

AND2x6_ASAP7_75t_L g389 ( 
.A(n_237),
.B(n_106),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_198),
.Y(n_390)
);

INVx2_ASAP7_75t_SL g391 ( 
.A(n_259),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_208),
.B(n_172),
.Y(n_392)
);

AND2x4_ASAP7_75t_L g393 ( 
.A(n_252),
.B(n_150),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_198),
.Y(n_394)
);

OR2x2_ASAP7_75t_L g395 ( 
.A(n_201),
.B(n_95),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_198),
.Y(n_396)
);

AND2x2_ASAP7_75t_L g397 ( 
.A(n_207),
.B(n_150),
.Y(n_397)
);

BUFx2_ASAP7_75t_L g398 ( 
.A(n_258),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_258),
.B(n_150),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_204),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_252),
.B(n_172),
.Y(n_401)
);

INVx4_ASAP7_75t_L g402 ( 
.A(n_204),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_256),
.B(n_172),
.Y(n_403)
);

BUFx6f_ASAP7_75t_L g404 ( 
.A(n_204),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_256),
.B(n_172),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_221),
.Y(n_406)
);

AND2x6_ASAP7_75t_L g407 ( 
.A(n_221),
.B(n_70),
.Y(n_407)
);

BUFx10_ASAP7_75t_L g408 ( 
.A(n_196),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_221),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_241),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g411 ( 
.A(n_241),
.B(n_70),
.Y(n_411)
);

AND2x2_ASAP7_75t_L g412 ( 
.A(n_262),
.B(n_152),
.Y(n_412)
);

INVx4_ASAP7_75t_L g413 ( 
.A(n_241),
.Y(n_413)
);

AND2x4_ASAP7_75t_L g414 ( 
.A(n_243),
.B(n_152),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g415 ( 
.A(n_197),
.B(n_123),
.Y(n_415)
);

BUFx3_ASAP7_75t_L g416 ( 
.A(n_243),
.Y(n_416)
);

OR2x2_ASAP7_75t_L g417 ( 
.A(n_243),
.B(n_123),
.Y(n_417)
);

BUFx2_ASAP7_75t_L g418 ( 
.A(n_247),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_247),
.Y(n_419)
);

AND2x4_ASAP7_75t_L g420 ( 
.A(n_267),
.B(n_154),
.Y(n_420)
);

BUFx3_ASAP7_75t_L g421 ( 
.A(n_247),
.Y(n_421)
);

BUFx6f_ASAP7_75t_L g422 ( 
.A(n_257),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_257),
.Y(n_423)
);

INVx2_ASAP7_75t_SL g424 ( 
.A(n_277),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_357),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_357),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_287),
.B(n_83),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g428 ( 
.A(n_278),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_356),
.B(n_154),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_364),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_335),
.Y(n_431)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_286),
.Y(n_432)
);

AO22x2_ASAP7_75t_L g433 ( 
.A1(n_384),
.A2(n_97),
.B1(n_92),
.B2(n_100),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_364),
.Y(n_434)
);

INVx2_ASAP7_75t_L g435 ( 
.A(n_286),
.Y(n_435)
);

INVx2_ASAP7_75t_SL g436 ( 
.A(n_277),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_279),
.B(n_327),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_286),
.Y(n_438)
);

NAND2x1p5_ASAP7_75t_L g439 ( 
.A(n_331),
.B(n_257),
.Y(n_439)
);

INVxp67_ASAP7_75t_SL g440 ( 
.A(n_303),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_312),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_328),
.B(n_267),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_366),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_312),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g445 ( 
.A(n_328),
.B(n_267),
.Y(n_445)
);

AOI22xp33_ASAP7_75t_L g446 ( 
.A1(n_363),
.A2(n_87),
.B1(n_130),
.B2(n_131),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g447 ( 
.A(n_277),
.B(n_172),
.Y(n_447)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_303),
.Y(n_448)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_301),
.A2(n_71),
.B1(n_181),
.B2(n_183),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_366),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_277),
.B(n_275),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_274),
.B(n_172),
.Y(n_452)
);

NAND2xp5_ASAP7_75t_SL g453 ( 
.A(n_341),
.B(n_71),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g454 ( 
.A(n_274),
.B(n_174),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_312),
.Y(n_455)
);

INVx4_ASAP7_75t_L g456 ( 
.A(n_303),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_313),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_313),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_313),
.Y(n_459)
);

CKINVDCx5p33_ASAP7_75t_R g460 ( 
.A(n_383),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_314),
.Y(n_461)
);

INVx3_ASAP7_75t_L g462 ( 
.A(n_303),
.Y(n_462)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_314),
.Y(n_463)
);

INVx1_ASAP7_75t_L g464 ( 
.A(n_314),
.Y(n_464)
);

INVxp67_ASAP7_75t_L g465 ( 
.A(n_371),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g466 ( 
.A(n_356),
.B(n_174),
.Y(n_466)
);

HB1xp67_ASAP7_75t_L g467 ( 
.A(n_412),
.Y(n_467)
);

AO22x2_ASAP7_75t_L g468 ( 
.A1(n_384),
.A2(n_83),
.B1(n_132),
.B2(n_86),
.Y(n_468)
);

INVxp67_ASAP7_75t_L g469 ( 
.A(n_321),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_316),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_316),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_316),
.Y(n_472)
);

INVxp67_ASAP7_75t_SL g473 ( 
.A(n_303),
.Y(n_473)
);

AO22x2_ASAP7_75t_L g474 ( 
.A1(n_287),
.A2(n_105),
.B1(n_103),
.B2(n_102),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_336),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_336),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_SL g477 ( 
.A(n_353),
.B(n_78),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_336),
.Y(n_478)
);

NAND2x1p5_ASAP7_75t_L g479 ( 
.A(n_331),
.B(n_174),
.Y(n_479)
);

BUFx4f_ASAP7_75t_L g480 ( 
.A(n_339),
.Y(n_480)
);

AND2x4_ASAP7_75t_L g481 ( 
.A(n_360),
.B(n_59),
.Y(n_481)
);

NOR2xp33_ASAP7_75t_L g482 ( 
.A(n_358),
.B(n_128),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_342),
.Y(n_483)
);

AO22x2_ASAP7_75t_L g484 ( 
.A1(n_287),
.A2(n_86),
.B1(n_132),
.B2(n_89),
.Y(n_484)
);

NAND3x1_ASAP7_75t_L g485 ( 
.A(n_352),
.B(n_103),
.C(n_89),
.Y(n_485)
);

INVx2_ASAP7_75t_L g486 ( 
.A(n_342),
.Y(n_486)
);

INVx2_ASAP7_75t_L g487 ( 
.A(n_342),
.Y(n_487)
);

AO22x2_ASAP7_75t_L g488 ( 
.A1(n_287),
.A2(n_118),
.B1(n_113),
.B2(n_109),
.Y(n_488)
);

BUFx3_ASAP7_75t_L g489 ( 
.A(n_295),
.Y(n_489)
);

AND2x2_ASAP7_75t_L g490 ( 
.A(n_373),
.B(n_174),
.Y(n_490)
);

AND2x4_ASAP7_75t_L g491 ( 
.A(n_360),
.B(n_368),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_293),
.B(n_174),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_368),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g494 ( 
.A(n_319),
.B(n_174),
.Y(n_494)
);

OR2x6_ASAP7_75t_L g495 ( 
.A(n_339),
.B(n_90),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_317),
.B(n_179),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_317),
.B(n_179),
.Y(n_497)
);

INVx3_ASAP7_75t_L g498 ( 
.A(n_303),
.Y(n_498)
);

BUFx2_ASAP7_75t_L g499 ( 
.A(n_391),
.Y(n_499)
);

INVxp67_ASAP7_75t_L g500 ( 
.A(n_305),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_346),
.Y(n_501)
);

NAND2x1p5_ASAP7_75t_L g502 ( 
.A(n_331),
.B(n_179),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_374),
.Y(n_503)
);

AO22x2_ASAP7_75t_L g504 ( 
.A1(n_299),
.A2(n_295),
.B1(n_308),
.B2(n_307),
.Y(n_504)
);

INVx5_ASAP7_75t_L g505 ( 
.A(n_304),
.Y(n_505)
);

INVx2_ASAP7_75t_L g506 ( 
.A(n_346),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_304),
.Y(n_507)
);

AOI22xp33_ASAP7_75t_L g508 ( 
.A1(n_363),
.A2(n_128),
.B1(n_179),
.B2(n_181),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_374),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_309),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g511 ( 
.A(n_317),
.B(n_179),
.Y(n_511)
);

INVxp67_ASAP7_75t_L g512 ( 
.A(n_397),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_SL g513 ( 
.A(n_297),
.B(n_79),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_309),
.Y(n_514)
);

INVx1_ASAP7_75t_L g515 ( 
.A(n_318),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_318),
.Y(n_516)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_322),
.Y(n_517)
);

NOR2x1p5_ASAP7_75t_L g518 ( 
.A(n_395),
.B(n_69),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_322),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_325),
.Y(n_520)
);

AND2x4_ASAP7_75t_L g521 ( 
.A(n_360),
.B(n_65),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_325),
.Y(n_522)
);

AND2x2_ASAP7_75t_L g523 ( 
.A(n_373),
.B(n_179),
.Y(n_523)
);

AO22x2_ASAP7_75t_L g524 ( 
.A1(n_299),
.A2(n_105),
.B1(n_102),
.B2(n_100),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_304),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_317),
.B(n_363),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_340),
.Y(n_527)
);

INVx5_ASAP7_75t_L g528 ( 
.A(n_304),
.Y(n_528)
);

AND2x4_ASAP7_75t_L g529 ( 
.A(n_354),
.B(n_90),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_340),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_344),
.Y(n_531)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_344),
.Y(n_532)
);

AND2x4_ASAP7_75t_L g533 ( 
.A(n_354),
.B(n_92),
.Y(n_533)
);

INVx1_ASAP7_75t_L g534 ( 
.A(n_347),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_347),
.Y(n_535)
);

BUFx3_ASAP7_75t_L g536 ( 
.A(n_295),
.Y(n_536)
);

BUFx6f_ASAP7_75t_L g537 ( 
.A(n_304),
.Y(n_537)
);

OAI221xp5_ASAP7_75t_L g538 ( 
.A1(n_415),
.A2(n_118),
.B1(n_113),
.B2(n_97),
.C(n_127),
.Y(n_538)
);

AOI22xp5_ASAP7_75t_L g539 ( 
.A1(n_297),
.A2(n_181),
.B1(n_183),
.B2(n_169),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_346),
.Y(n_540)
);

NAND2x1p5_ASAP7_75t_L g541 ( 
.A(n_331),
.B(n_334),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_363),
.B(n_181),
.Y(n_542)
);

NAND2xp5_ASAP7_75t_L g543 ( 
.A(n_375),
.B(n_181),
.Y(n_543)
);

NOR2xp33_ASAP7_75t_L g544 ( 
.A(n_365),
.B(n_96),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_324),
.Y(n_545)
);

AOI22xp33_ASAP7_75t_L g546 ( 
.A1(n_393),
.A2(n_181),
.B1(n_183),
.B2(n_109),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_324),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_418),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_330),
.B(n_183),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_418),
.Y(n_550)
);

NOR2xp67_ASAP7_75t_L g551 ( 
.A(n_388),
.B(n_69),
.Y(n_551)
);

AOI22xp33_ASAP7_75t_L g552 ( 
.A1(n_393),
.A2(n_183),
.B1(n_127),
.B2(n_104),
.Y(n_552)
);

BUFx3_ASAP7_75t_L g553 ( 
.A(n_307),
.Y(n_553)
);

AO22x2_ASAP7_75t_L g554 ( 
.A1(n_307),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_554)
);

AND2x2_ASAP7_75t_L g555 ( 
.A(n_330),
.B(n_183),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_350),
.B(n_81),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g557 ( 
.A(n_375),
.B(n_169),
.Y(n_557)
);

INVx2_ASAP7_75t_L g558 ( 
.A(n_414),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_272),
.Y(n_559)
);

INVx1_ASAP7_75t_SL g560 ( 
.A(n_310),
.Y(n_560)
);

AND2x4_ASAP7_75t_L g561 ( 
.A(n_354),
.B(n_169),
.Y(n_561)
);

INVx1_ASAP7_75t_L g562 ( 
.A(n_272),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_276),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_414),
.Y(n_564)
);

AND2x2_ASAP7_75t_SL g565 ( 
.A(n_393),
.B(n_186),
.Y(n_565)
);

NAND2x1p5_ASAP7_75t_L g566 ( 
.A(n_334),
.B(n_169),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_283),
.Y(n_567)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_375),
.B(n_169),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_414),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_352),
.A2(n_133),
.B1(n_126),
.B2(n_125),
.Y(n_570)
);

OAI221xp5_ASAP7_75t_L g571 ( 
.A1(n_285),
.A2(n_120),
.B1(n_98),
.B2(n_107),
.C(n_108),
.Y(n_571)
);

INVx1_ASAP7_75t_L g572 ( 
.A(n_283),
.Y(n_572)
);

AOI22xp33_ASAP7_75t_L g573 ( 
.A1(n_393),
.A2(n_110),
.B1(n_112),
.B2(n_114),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_414),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_375),
.B(n_169),
.Y(n_575)
);

OAI22xp33_ASAP7_75t_L g576 ( 
.A1(n_273),
.A2(n_133),
.B1(n_88),
.B2(n_91),
.Y(n_576)
);

NAND2x1p5_ASAP7_75t_L g577 ( 
.A(n_334),
.B(n_361),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_420),
.Y(n_578)
);

INVx1_ASAP7_75t_L g579 ( 
.A(n_420),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_308),
.A2(n_338),
.B1(n_381),
.B2(n_382),
.Y(n_580)
);

INVx1_ASAP7_75t_L g581 ( 
.A(n_420),
.Y(n_581)
);

INVx2_ASAP7_75t_L g582 ( 
.A(n_420),
.Y(n_582)
);

BUFx2_ASAP7_75t_L g583 ( 
.A(n_391),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g584 ( 
.A(n_308),
.B(n_115),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_377),
.B(n_169),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_354),
.B(n_338),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_288),
.Y(n_587)
);

NAND2x1p5_ASAP7_75t_L g588 ( 
.A(n_334),
.B(n_169),
.Y(n_588)
);

NOR2xp33_ASAP7_75t_L g589 ( 
.A(n_338),
.B(n_124),
.Y(n_589)
);

NAND2xp33_ASAP7_75t_L g590 ( 
.A(n_304),
.B(n_161),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_L g591 ( 
.A(n_297),
.B(n_119),
.Y(n_591)
);

AOI22xp33_ASAP7_75t_L g592 ( 
.A1(n_273),
.A2(n_81),
.B1(n_88),
.B2(n_91),
.Y(n_592)
);

A2O1A1Ixp33_ASAP7_75t_L g593 ( 
.A1(n_381),
.A2(n_125),
.B(n_126),
.C(n_184),
.Y(n_593)
);

INVx2_ASAP7_75t_SL g594 ( 
.A(n_417),
.Y(n_594)
);

AND2x4_ASAP7_75t_L g595 ( 
.A(n_382),
.B(n_0),
.Y(n_595)
);

NOR2xp33_ASAP7_75t_L g596 ( 
.A(n_395),
.B(n_2),
.Y(n_596)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_288),
.Y(n_597)
);

INVx2_ASAP7_75t_L g598 ( 
.A(n_289),
.Y(n_598)
);

O2A1O1Ixp33_ASAP7_75t_L g599 ( 
.A1(n_482),
.A2(n_294),
.B(n_379),
.C(n_326),
.Y(n_599)
);

AND2x2_ASAP7_75t_SL g600 ( 
.A(n_480),
.B(n_383),
.Y(n_600)
);

NAND2xp5_ASAP7_75t_L g601 ( 
.A(n_451),
.B(n_297),
.Y(n_601)
);

INVx2_ASAP7_75t_L g602 ( 
.A(n_432),
.Y(n_602)
);

HB1xp67_ASAP7_75t_L g603 ( 
.A(n_467),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_594),
.B(n_350),
.Y(n_604)
);

BUFx2_ASAP7_75t_L g605 ( 
.A(n_499),
.Y(n_605)
);

AOI21x1_ASAP7_75t_L g606 ( 
.A1(n_494),
.A2(n_376),
.B(n_372),
.Y(n_606)
);

BUFx6f_ASAP7_75t_L g607 ( 
.A(n_525),
.Y(n_607)
);

OAI21xp5_ASAP7_75t_L g608 ( 
.A1(n_526),
.A2(n_306),
.B(n_329),
.Y(n_608)
);

OAI22xp5_ASAP7_75t_L g609 ( 
.A1(n_424),
.A2(n_290),
.B1(n_339),
.B2(n_349),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_550),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_550),
.Y(n_611)
);

OAI22xp5_ASAP7_75t_L g612 ( 
.A1(n_424),
.A2(n_290),
.B1(n_339),
.B2(n_284),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_594),
.B(n_397),
.Y(n_613)
);

AOI21xp5_ASAP7_75t_L g614 ( 
.A1(n_505),
.A2(n_351),
.B(n_386),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_432),
.Y(n_615)
);

AOI21xp5_ASAP7_75t_L g616 ( 
.A1(n_505),
.A2(n_386),
.B(n_362),
.Y(n_616)
);

NOR2xp33_ASAP7_75t_L g617 ( 
.A(n_500),
.B(n_311),
.Y(n_617)
);

NOR2xp67_ASAP7_75t_L g618 ( 
.A(n_431),
.B(n_417),
.Y(n_618)
);

HB1xp67_ASAP7_75t_L g619 ( 
.A(n_489),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_429),
.B(n_399),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_429),
.B(n_399),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_433),
.A2(n_370),
.B1(n_389),
.B2(n_273),
.Y(n_622)
);

INVx1_ASAP7_75t_SL g623 ( 
.A(n_560),
.Y(n_623)
);

AOI22xp33_ASAP7_75t_L g624 ( 
.A1(n_433),
.A2(n_370),
.B1(n_389),
.B2(n_273),
.Y(n_624)
);

AOI21xp5_ASAP7_75t_L g625 ( 
.A1(n_505),
.A2(n_362),
.B(n_386),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_436),
.B(n_412),
.Y(n_626)
);

AND2x2_ASAP7_75t_L g627 ( 
.A(n_512),
.B(n_408),
.Y(n_627)
);

NAND2xp5_ASAP7_75t_L g628 ( 
.A(n_436),
.B(n_290),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_466),
.B(n_370),
.Y(n_629)
);

INVx2_ASAP7_75t_L g630 ( 
.A(n_435),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_L g631 ( 
.A(n_466),
.B(n_490),
.Y(n_631)
);

AND2x2_ASAP7_75t_L g632 ( 
.A(n_556),
.B(n_408),
.Y(n_632)
);

AOI21xp5_ASAP7_75t_L g633 ( 
.A1(n_505),
.A2(n_386),
.B(n_362),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_SL g634 ( 
.A(n_565),
.B(n_345),
.Y(n_634)
);

OAI21xp5_ASAP7_75t_L g635 ( 
.A1(n_447),
.A2(n_403),
.B(n_405),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_505),
.A2(n_362),
.B(n_386),
.Y(n_636)
);

AOI22xp5_ASAP7_75t_L g637 ( 
.A1(n_586),
.A2(n_280),
.B1(n_339),
.B2(n_370),
.Y(n_637)
);

HB1xp67_ASAP7_75t_L g638 ( 
.A(n_489),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_490),
.B(n_523),
.Y(n_639)
);

O2A1O1Ixp33_ASAP7_75t_L g640 ( 
.A1(n_596),
.A2(n_428),
.B(n_571),
.C(n_538),
.Y(n_640)
);

NOR2xp33_ASAP7_75t_L g641 ( 
.A(n_469),
.B(n_311),
.Y(n_641)
);

AOI21xp5_ASAP7_75t_L g642 ( 
.A1(n_528),
.A2(n_541),
.B(n_577),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_525),
.Y(n_643)
);

NAND2xp5_ASAP7_75t_L g644 ( 
.A(n_523),
.B(n_370),
.Y(n_644)
);

AOI21xp5_ASAP7_75t_L g645 ( 
.A1(n_528),
.A2(n_386),
.B(n_362),
.Y(n_645)
);

AOI21xp5_ASAP7_75t_L g646 ( 
.A1(n_528),
.A2(n_362),
.B(n_361),
.Y(n_646)
);

A2O1A1Ixp33_ASAP7_75t_L g647 ( 
.A1(n_449),
.A2(n_292),
.B(n_289),
.C(n_300),
.Y(n_647)
);

OAI22xp5_ASAP7_75t_L g648 ( 
.A1(n_565),
.A2(n_273),
.B1(n_302),
.B2(n_291),
.Y(n_648)
);

AOI21xp5_ASAP7_75t_L g649 ( 
.A1(n_528),
.A2(n_361),
.B(n_345),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_435),
.Y(n_650)
);

AOI21xp5_ASAP7_75t_L g651 ( 
.A1(n_528),
.A2(n_345),
.B(n_367),
.Y(n_651)
);

AOI21x1_ASAP7_75t_L g652 ( 
.A1(n_438),
.A2(n_291),
.B(n_300),
.Y(n_652)
);

AND2x4_ASAP7_75t_L g653 ( 
.A(n_586),
.B(n_298),
.Y(n_653)
);

A2O1A1Ixp33_ASAP7_75t_L g654 ( 
.A1(n_510),
.A2(n_298),
.B(n_323),
.C(n_355),
.Y(n_654)
);

INVx1_ASAP7_75t_L g655 ( 
.A(n_598),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_548),
.B(n_370),
.Y(n_656)
);

AND2x2_ASAP7_75t_L g657 ( 
.A(n_556),
.B(n_408),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_L g658 ( 
.A(n_437),
.B(n_408),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_598),
.Y(n_659)
);

AOI21xp5_ASAP7_75t_L g660 ( 
.A1(n_541),
.A2(n_345),
.B(n_369),
.Y(n_660)
);

BUFx6f_ASAP7_75t_L g661 ( 
.A(n_525),
.Y(n_661)
);

BUFx6f_ASAP7_75t_L g662 ( 
.A(n_525),
.Y(n_662)
);

AND2x2_ASAP7_75t_SL g663 ( 
.A(n_480),
.B(n_398),
.Y(n_663)
);

CKINVDCx5p33_ASAP7_75t_R g664 ( 
.A(n_431),
.Y(n_664)
);

AOI22xp5_ASAP7_75t_L g665 ( 
.A1(n_586),
.A2(n_389),
.B1(n_370),
.B2(n_332),
.Y(n_665)
);

AOI21xp5_ASAP7_75t_L g666 ( 
.A1(n_541),
.A2(n_345),
.B(n_367),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_465),
.B(n_343),
.Y(n_667)
);

NAND2xp5_ASAP7_75t_SL g668 ( 
.A(n_427),
.B(n_402),
.Y(n_668)
);

BUFx6f_ASAP7_75t_L g669 ( 
.A(n_525),
.Y(n_669)
);

NAND2xp5_ASAP7_75t_L g670 ( 
.A(n_549),
.B(n_389),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_461),
.Y(n_671)
);

AOI21xp5_ASAP7_75t_L g672 ( 
.A1(n_577),
.A2(n_387),
.B(n_378),
.Y(n_672)
);

INVx2_ASAP7_75t_L g673 ( 
.A(n_461),
.Y(n_673)
);

BUFx6f_ASAP7_75t_L g674 ( 
.A(n_537),
.Y(n_674)
);

NAND2xp5_ASAP7_75t_L g675 ( 
.A(n_549),
.B(n_389),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_555),
.B(n_389),
.Y(n_676)
);

AOI22xp5_ASAP7_75t_L g677 ( 
.A1(n_427),
.A2(n_389),
.B1(n_302),
.B2(n_333),
.Y(n_677)
);

NOR2xp33_ASAP7_75t_L g678 ( 
.A(n_453),
.B(n_398),
.Y(n_678)
);

NAND3xp33_ASAP7_75t_L g679 ( 
.A(n_584),
.B(n_355),
.C(n_302),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_491),
.B(n_402),
.Y(n_680)
);

AOI21xp5_ASAP7_75t_L g681 ( 
.A1(n_442),
.A2(n_445),
.B(n_456),
.Y(n_681)
);

AOI21xp5_ASAP7_75t_L g682 ( 
.A1(n_456),
.A2(n_387),
.B(n_378),
.Y(n_682)
);

INVx3_ASAP7_75t_SL g683 ( 
.A(n_460),
.Y(n_683)
);

OAI21xp33_ASAP7_75t_L g684 ( 
.A1(n_446),
.A2(n_359),
.B(n_380),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_L g685 ( 
.A(n_555),
.B(n_296),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_559),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_529),
.B(n_296),
.Y(n_687)
);

AND2x2_ASAP7_75t_L g688 ( 
.A(n_589),
.B(n_302),
.Y(n_688)
);

AOI21xp5_ASAP7_75t_L g689 ( 
.A1(n_456),
.A2(n_387),
.B(n_402),
.Y(n_689)
);

NOR2xp33_ASAP7_75t_L g690 ( 
.A(n_595),
.B(n_302),
.Y(n_690)
);

AND2x6_ASAP7_75t_L g691 ( 
.A(n_481),
.B(n_281),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_L g692 ( 
.A(n_529),
.B(n_296),
.Y(n_692)
);

NOR2xp33_ASAP7_75t_L g693 ( 
.A(n_595),
.B(n_402),
.Y(n_693)
);

AOI21xp5_ASAP7_75t_L g694 ( 
.A1(n_590),
.A2(n_413),
.B(n_337),
.Y(n_694)
);

OAI21x1_ASAP7_75t_L g695 ( 
.A1(n_439),
.A2(n_281),
.B(n_315),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_529),
.B(n_533),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_590),
.A2(n_413),
.B(n_337),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_533),
.B(n_296),
.Y(n_698)
);

NOR2xp33_ASAP7_75t_L g699 ( 
.A(n_595),
.B(n_413),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_533),
.B(n_296),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_L g701 ( 
.A(n_492),
.B(n_514),
.Y(n_701)
);

OAI22xp5_ASAP7_75t_L g702 ( 
.A1(n_580),
.A2(n_597),
.B1(n_562),
.B2(n_587),
.Y(n_702)
);

AOI21xp5_ASAP7_75t_L g703 ( 
.A1(n_440),
.A2(n_281),
.B(n_337),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_470),
.Y(n_704)
);

HB1xp67_ASAP7_75t_L g705 ( 
.A(n_536),
.Y(n_705)
);

AOI21x1_ASAP7_75t_L g706 ( 
.A1(n_438),
.A2(n_401),
.B(n_385),
.Y(n_706)
);

AOI21x1_ASAP7_75t_L g707 ( 
.A1(n_441),
.A2(n_392),
.B(n_390),
.Y(n_707)
);

OAI22xp5_ASAP7_75t_L g708 ( 
.A1(n_580),
.A2(n_337),
.B1(n_315),
.B2(n_421),
.Y(n_708)
);

NAND2xp5_ASAP7_75t_SL g709 ( 
.A(n_491),
.B(n_404),
.Y(n_709)
);

NOR2xp33_ASAP7_75t_L g710 ( 
.A(n_591),
.B(n_421),
.Y(n_710)
);

AOI21xp5_ASAP7_75t_L g711 ( 
.A1(n_473),
.A2(n_315),
.B(n_421),
.Y(n_711)
);

O2A1O1Ixp5_ASAP7_75t_L g712 ( 
.A1(n_513),
.A2(n_593),
.B(n_585),
.C(n_543),
.Y(n_712)
);

NAND3xp33_ASAP7_75t_L g713 ( 
.A(n_544),
.B(n_422),
.C(n_404),
.Y(n_713)
);

INVx1_ASAP7_75t_L g714 ( 
.A(n_563),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_515),
.B(n_296),
.Y(n_715)
);

CKINVDCx11_ASAP7_75t_R g716 ( 
.A(n_499),
.Y(n_716)
);

AOI21xp5_ASAP7_75t_L g717 ( 
.A1(n_507),
.A2(n_416),
.B(n_348),
.Y(n_717)
);

NOR2xp33_ASAP7_75t_L g718 ( 
.A(n_477),
.B(n_416),
.Y(n_718)
);

A2O1A1Ixp33_ASAP7_75t_L g719 ( 
.A1(n_516),
.A2(n_406),
.B(n_390),
.C(n_394),
.Y(n_719)
);

O2A1O1Ixp33_ASAP7_75t_L g720 ( 
.A1(n_576),
.A2(n_406),
.B(n_394),
.C(n_409),
.Y(n_720)
);

INVx4_ASAP7_75t_L g721 ( 
.A(n_536),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_518),
.B(n_348),
.Y(n_722)
);

AOI21xp5_ASAP7_75t_L g723 ( 
.A1(n_496),
.A2(n_416),
.B(n_348),
.Y(n_723)
);

OAI21xp5_ASAP7_75t_L g724 ( 
.A1(n_542),
.A2(n_409),
.B(n_410),
.Y(n_724)
);

AOI21xp5_ASAP7_75t_L g725 ( 
.A1(n_497),
.A2(n_396),
.B(n_419),
.Y(n_725)
);

OAI22xp5_ASAP7_75t_L g726 ( 
.A1(n_580),
.A2(n_422),
.B1(n_404),
.B2(n_419),
.Y(n_726)
);

O2A1O1Ixp33_ASAP7_75t_L g727 ( 
.A1(n_517),
.A2(n_410),
.B(n_423),
.C(n_400),
.Y(n_727)
);

AOI22xp33_ASAP7_75t_L g728 ( 
.A1(n_433),
.A2(n_296),
.B1(n_320),
.B2(n_407),
.Y(n_728)
);

AOI22xp5_ASAP7_75t_L g729 ( 
.A1(n_491),
.A2(n_320),
.B1(n_422),
.B2(n_404),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_519),
.B(n_320),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_553),
.B(n_320),
.Y(n_731)
);

CKINVDCx20_ASAP7_75t_R g732 ( 
.A(n_460),
.Y(n_732)
);

INVx3_ASAP7_75t_L g733 ( 
.A(n_558),
.Y(n_733)
);

AOI21xp5_ASAP7_75t_L g734 ( 
.A1(n_511),
.A2(n_396),
.B(n_419),
.Y(n_734)
);

NAND2xp5_ASAP7_75t_L g735 ( 
.A(n_520),
.B(n_522),
.Y(n_735)
);

OAI22xp5_ASAP7_75t_L g736 ( 
.A1(n_580),
.A2(n_422),
.B1(n_404),
.B2(n_419),
.Y(n_736)
);

NAND3xp33_ASAP7_75t_L g737 ( 
.A(n_573),
.B(n_422),
.C(n_404),
.Y(n_737)
);

OAI21xp5_ASAP7_75t_L g738 ( 
.A1(n_557),
.A2(n_320),
.B(n_423),
.Y(n_738)
);

AOI21xp5_ASAP7_75t_L g739 ( 
.A1(n_537),
.A2(n_396),
.B(n_422),
.Y(n_739)
);

NAND2xp5_ASAP7_75t_L g740 ( 
.A(n_527),
.B(n_320),
.Y(n_740)
);

NOR2xp33_ASAP7_75t_L g741 ( 
.A(n_583),
.B(n_553),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_530),
.A2(n_423),
.B(n_400),
.C(n_396),
.Y(n_742)
);

HB1xp67_ASAP7_75t_L g743 ( 
.A(n_583),
.Y(n_743)
);

NOR2xp33_ASAP7_75t_L g744 ( 
.A(n_531),
.B(n_400),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_532),
.B(n_320),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_567),
.Y(n_746)
);

AND2x2_ASAP7_75t_L g747 ( 
.A(n_551),
.B(n_411),
.Y(n_747)
);

AOI21xp5_ASAP7_75t_L g748 ( 
.A1(n_537),
.A2(n_282),
.B(n_189),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_R g749 ( 
.A(n_574),
.B(n_411),
.Y(n_749)
);

INVx2_ASAP7_75t_L g750 ( 
.A(n_470),
.Y(n_750)
);

NAND2xp5_ASAP7_75t_L g751 ( 
.A(n_534),
.B(n_411),
.Y(n_751)
);

O2A1O1Ixp5_ASAP7_75t_L g752 ( 
.A1(n_545),
.A2(n_547),
.B(n_535),
.C(n_572),
.Y(n_752)
);

AND2x2_ASAP7_75t_L g753 ( 
.A(n_592),
.B(n_411),
.Y(n_753)
);

INVx4_ASAP7_75t_L g754 ( 
.A(n_537),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_481),
.B(n_282),
.Y(n_755)
);

NAND2xp5_ASAP7_75t_L g756 ( 
.A(n_425),
.B(n_411),
.Y(n_756)
);

AND2x2_ASAP7_75t_L g757 ( 
.A(n_433),
.B(n_411),
.Y(n_757)
);

AOI21xp5_ASAP7_75t_L g758 ( 
.A1(n_537),
.A2(n_282),
.B(n_189),
.Y(n_758)
);

AOI21xp5_ASAP7_75t_L g759 ( 
.A1(n_566),
.A2(n_282),
.B(n_189),
.Y(n_759)
);

INVx2_ASAP7_75t_L g760 ( 
.A(n_483),
.Y(n_760)
);

NOR3xp33_ASAP7_75t_L g761 ( 
.A(n_570),
.B(n_411),
.C(n_407),
.Y(n_761)
);

HB1xp67_ASAP7_75t_L g762 ( 
.A(n_481),
.Y(n_762)
);

BUFx6f_ASAP7_75t_L g763 ( 
.A(n_448),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_426),
.B(n_407),
.Y(n_764)
);

AOI21xp5_ASAP7_75t_L g765 ( 
.A1(n_566),
.A2(n_282),
.B(n_189),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_430),
.B(n_407),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_566),
.A2(n_189),
.B(n_180),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_588),
.A2(n_189),
.B(n_180),
.Y(n_768)
);

INVx2_ASAP7_75t_SL g769 ( 
.A(n_521),
.Y(n_769)
);

AOI21xp5_ASAP7_75t_L g770 ( 
.A1(n_588),
.A2(n_439),
.B(n_479),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_588),
.A2(n_189),
.B(n_180),
.Y(n_771)
);

NAND3xp33_ASAP7_75t_L g772 ( 
.A(n_552),
.B(n_180),
.C(n_166),
.Y(n_772)
);

OR2x2_ASAP7_75t_L g773 ( 
.A(n_452),
.B(n_5),
.Y(n_773)
);

BUFx6f_ASAP7_75t_L g774 ( 
.A(n_448),
.Y(n_774)
);

AOI21xp33_ASAP7_75t_L g775 ( 
.A1(n_568),
.A2(n_7),
.B(n_8),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_434),
.B(n_443),
.Y(n_776)
);

AOI21xp5_ASAP7_75t_L g777 ( 
.A1(n_439),
.A2(n_189),
.B(n_180),
.Y(n_777)
);

AOI21xp5_ASAP7_75t_L g778 ( 
.A1(n_479),
.A2(n_189),
.B(n_180),
.Y(n_778)
);

INVx1_ASAP7_75t_L g779 ( 
.A(n_441),
.Y(n_779)
);

AOI21xp5_ASAP7_75t_L g780 ( 
.A1(n_479),
.A2(n_189),
.B(n_180),
.Y(n_780)
);

AOI21xp5_ASAP7_75t_L g781 ( 
.A1(n_502),
.A2(n_189),
.B(n_180),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_558),
.B(n_407),
.Y(n_782)
);

INVx2_ASAP7_75t_SL g783 ( 
.A(n_521),
.Y(n_783)
);

AOI21xp5_ASAP7_75t_L g784 ( 
.A1(n_502),
.A2(n_575),
.B(n_582),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_SL g785 ( 
.A(n_521),
.B(n_180),
.Y(n_785)
);

AOI21xp5_ASAP7_75t_L g786 ( 
.A1(n_502),
.A2(n_582),
.B(n_564),
.Y(n_786)
);

AOI21xp5_ASAP7_75t_L g787 ( 
.A1(n_564),
.A2(n_189),
.B(n_180),
.Y(n_787)
);

A2O1A1Ixp33_ASAP7_75t_L g788 ( 
.A1(n_450),
.A2(n_407),
.B(n_186),
.C(n_184),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_454),
.A2(n_407),
.B(n_9),
.C(n_10),
.Y(n_789)
);

INVx1_ASAP7_75t_L g790 ( 
.A(n_444),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_493),
.B(n_8),
.Y(n_791)
);

AOI21xp5_ASAP7_75t_L g792 ( 
.A1(n_569),
.A2(n_189),
.B(n_186),
.Y(n_792)
);

AOI21xp5_ASAP7_75t_L g793 ( 
.A1(n_569),
.A2(n_186),
.B(n_184),
.Y(n_793)
);

INVx2_ASAP7_75t_L g794 ( 
.A(n_483),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_503),
.B(n_10),
.Y(n_795)
);

O2A1O1Ixp33_ASAP7_75t_L g796 ( 
.A1(n_509),
.A2(n_495),
.B(n_540),
.C(n_444),
.Y(n_796)
);

INVx1_ASAP7_75t_L g797 ( 
.A(n_455),
.Y(n_797)
);

INVx1_ASAP7_75t_L g798 ( 
.A(n_455),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_561),
.B(n_186),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_448),
.A2(n_186),
.B(n_184),
.Y(n_800)
);

NOR2xp33_ASAP7_75t_L g801 ( 
.A(n_574),
.B(n_11),
.Y(n_801)
);

BUFx2_ASAP7_75t_L g802 ( 
.A(n_605),
.Y(n_802)
);

INVx1_ASAP7_75t_L g803 ( 
.A(n_686),
.Y(n_803)
);

INVx3_ASAP7_75t_L g804 ( 
.A(n_653),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_602),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_620),
.B(n_578),
.Y(n_806)
);

INVx2_ASAP7_75t_L g807 ( 
.A(n_602),
.Y(n_807)
);

NOR2xp33_ASAP7_75t_L g808 ( 
.A(n_617),
.B(n_578),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_601),
.B(n_457),
.Y(n_809)
);

INVx4_ASAP7_75t_L g810 ( 
.A(n_607),
.Y(n_810)
);

AOI21xp5_ASAP7_75t_L g811 ( 
.A1(n_770),
.A2(n_457),
.B(n_458),
.Y(n_811)
);

INVx1_ASAP7_75t_L g812 ( 
.A(n_714),
.Y(n_812)
);

NOR2xp33_ASAP7_75t_L g813 ( 
.A(n_617),
.B(n_579),
.Y(n_813)
);

O2A1O1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_640),
.A2(n_495),
.B(n_581),
.C(n_579),
.Y(n_814)
);

AO21x1_ASAP7_75t_L g815 ( 
.A1(n_668),
.A2(n_796),
.B(n_702),
.Y(n_815)
);

INVx2_ASAP7_75t_L g816 ( 
.A(n_615),
.Y(n_816)
);

AOI21xp5_ASAP7_75t_L g817 ( 
.A1(n_642),
.A2(n_458),
.B(n_459),
.Y(n_817)
);

AOI21xp5_ASAP7_75t_L g818 ( 
.A1(n_689),
.A2(n_459),
.B(n_478),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_SL g819 ( 
.A(n_688),
.B(n_475),
.Y(n_819)
);

NOR2xp33_ASAP7_75t_L g820 ( 
.A(n_679),
.B(n_581),
.Y(n_820)
);

CKINVDCx5p33_ASAP7_75t_R g821 ( 
.A(n_664),
.Y(n_821)
);

A2O1A1Ixp33_ASAP7_75t_L g822 ( 
.A1(n_599),
.A2(n_561),
.B(n_463),
.C(n_464),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_621),
.B(n_468),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_746),
.Y(n_824)
);

OAI22xp5_ASAP7_75t_L g825 ( 
.A1(n_693),
.A2(n_504),
.B1(n_463),
.B2(n_476),
.Y(n_825)
);

INVx2_ASAP7_75t_L g826 ( 
.A(n_615),
.Y(n_826)
);

AOI21xp5_ASAP7_75t_L g827 ( 
.A1(n_694),
.A2(n_475),
.B(n_464),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_604),
.B(n_468),
.Y(n_828)
);

AND2x4_ASAP7_75t_L g829 ( 
.A(n_721),
.B(n_561),
.Y(n_829)
);

OAI22x1_ASAP7_75t_L g830 ( 
.A1(n_677),
.A2(n_468),
.B1(n_554),
.B2(n_485),
.Y(n_830)
);

OR2x2_ASAP7_75t_L g831 ( 
.A(n_613),
.B(n_495),
.Y(n_831)
);

AOI21xp5_ASAP7_75t_L g832 ( 
.A1(n_697),
.A2(n_476),
.B(n_478),
.Y(n_832)
);

NAND3xp33_ASAP7_75t_SL g833 ( 
.A(n_658),
.B(n_508),
.C(n_539),
.Y(n_833)
);

NAND3xp33_ASAP7_75t_SL g834 ( 
.A(n_658),
.B(n_471),
.C(n_472),
.Y(n_834)
);

NAND2xp5_ASAP7_75t_L g835 ( 
.A(n_632),
.B(n_468),
.Y(n_835)
);

NAND2xp5_ASAP7_75t_L g836 ( 
.A(n_657),
.B(n_693),
.Y(n_836)
);

OAI22xp5_ASAP7_75t_L g837 ( 
.A1(n_699),
.A2(n_504),
.B1(n_472),
.B2(n_471),
.Y(n_837)
);

INVx3_ASAP7_75t_L g838 ( 
.A(n_653),
.Y(n_838)
);

CKINVDCx20_ASAP7_75t_R g839 ( 
.A(n_732),
.Y(n_839)
);

NAND2x1p5_ASAP7_75t_L g840 ( 
.A(n_754),
.B(n_462),
.Y(n_840)
);

AOI21xp5_ASAP7_75t_L g841 ( 
.A1(n_660),
.A2(n_462),
.B(n_498),
.Y(n_841)
);

INVx3_ASAP7_75t_L g842 ( 
.A(n_653),
.Y(n_842)
);

OAI21x1_ASAP7_75t_L g843 ( 
.A1(n_695),
.A2(n_486),
.B(n_487),
.Y(n_843)
);

NOR2xp33_ASAP7_75t_L g844 ( 
.A(n_641),
.B(n_506),
.Y(n_844)
);

OR2x2_ASAP7_75t_L g845 ( 
.A(n_603),
.B(n_495),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_716),
.Y(n_846)
);

OAI22xp5_ASAP7_75t_L g847 ( 
.A1(n_699),
.A2(n_504),
.B1(n_546),
.B2(n_487),
.Y(n_847)
);

OAI22xp5_ASAP7_75t_L g848 ( 
.A1(n_769),
.A2(n_504),
.B1(n_486),
.B2(n_506),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_610),
.B(n_501),
.Y(n_849)
);

BUFx6f_ASAP7_75t_L g850 ( 
.A(n_607),
.Y(n_850)
);

AOI22xp33_ASAP7_75t_L g851 ( 
.A1(n_775),
.A2(n_554),
.B1(n_474),
.B2(n_488),
.Y(n_851)
);

NOR2xp33_ASAP7_75t_L g852 ( 
.A(n_641),
.B(n_501),
.Y(n_852)
);

OAI21x1_ASAP7_75t_L g853 ( 
.A1(n_666),
.A2(n_462),
.B(n_498),
.Y(n_853)
);

AOI22xp33_ASAP7_75t_L g854 ( 
.A1(n_622),
.A2(n_554),
.B1(n_474),
.B2(n_488),
.Y(n_854)
);

NAND2xp5_ASAP7_75t_L g855 ( 
.A(n_611),
.B(n_488),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_655),
.Y(n_856)
);

OAI21xp33_ASAP7_75t_SL g857 ( 
.A1(n_668),
.A2(n_634),
.B(n_624),
.Y(n_857)
);

NAND2xp5_ASAP7_75t_L g858 ( 
.A(n_626),
.B(n_488),
.Y(n_858)
);

O2A1O1Ixp33_ASAP7_75t_SL g859 ( 
.A1(n_647),
.A2(n_554),
.B(n_498),
.C(n_484),
.Y(n_859)
);

BUFx6f_ASAP7_75t_L g860 ( 
.A(n_607),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_672),
.A2(n_524),
.B(n_474),
.Y(n_861)
);

NAND2xp5_ASAP7_75t_SL g862 ( 
.A(n_710),
.B(n_474),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_659),
.Y(n_863)
);

AOI21xp5_ASAP7_75t_L g864 ( 
.A1(n_681),
.A2(n_524),
.B(n_484),
.Y(n_864)
);

OR2x2_ASAP7_75t_L g865 ( 
.A(n_623),
.B(n_485),
.Y(n_865)
);

AND2x4_ASAP7_75t_L g866 ( 
.A(n_721),
.B(n_12),
.Y(n_866)
);

AO21x1_ASAP7_75t_L g867 ( 
.A1(n_710),
.A2(n_524),
.B(n_484),
.Y(n_867)
);

NAND2x1_ASAP7_75t_L g868 ( 
.A(n_691),
.B(n_754),
.Y(n_868)
);

AOI21xp5_ASAP7_75t_L g869 ( 
.A1(n_608),
.A2(n_524),
.B(n_484),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_SL g870 ( 
.A(n_631),
.B(n_186),
.Y(n_870)
);

INVx1_ASAP7_75t_L g871 ( 
.A(n_735),
.Y(n_871)
);

INVx2_ASAP7_75t_L g872 ( 
.A(n_630),
.Y(n_872)
);

NOR2xp33_ASAP7_75t_L g873 ( 
.A(n_678),
.B(n_13),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_630),
.Y(n_874)
);

AOI21xp5_ASAP7_75t_L g875 ( 
.A1(n_635),
.A2(n_186),
.B(n_184),
.Y(n_875)
);

O2A1O1Ixp5_ASAP7_75t_L g876 ( 
.A1(n_606),
.A2(n_14),
.B(n_15),
.C(n_17),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_716),
.Y(n_877)
);

BUFx8_ASAP7_75t_L g878 ( 
.A(n_627),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_779),
.Y(n_879)
);

AOI21xp5_ASAP7_75t_L g880 ( 
.A1(n_651),
.A2(n_186),
.B(n_184),
.Y(n_880)
);

AOI21xp5_ASAP7_75t_L g881 ( 
.A1(n_682),
.A2(n_186),
.B(n_184),
.Y(n_881)
);

CKINVDCx11_ASAP7_75t_R g882 ( 
.A(n_732),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_650),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_701),
.A2(n_186),
.B(n_184),
.Y(n_884)
);

NOR2xp33_ASAP7_75t_L g885 ( 
.A(n_678),
.B(n_14),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_650),
.Y(n_886)
);

AOI22xp5_ASAP7_75t_L g887 ( 
.A1(n_618),
.A2(n_186),
.B1(n_184),
.B2(n_180),
.Y(n_887)
);

INVx3_ASAP7_75t_L g888 ( 
.A(n_754),
.Y(n_888)
);

O2A1O1Ixp33_ASAP7_75t_L g889 ( 
.A1(n_654),
.A2(n_18),
.B(n_19),
.C(n_22),
.Y(n_889)
);

O2A1O1Ixp33_ASAP7_75t_L g890 ( 
.A1(n_654),
.A2(n_19),
.B(n_22),
.C(n_24),
.Y(n_890)
);

NAND2x1_ASAP7_75t_L g891 ( 
.A(n_691),
.B(n_184),
.Y(n_891)
);

INVx1_ASAP7_75t_SL g892 ( 
.A(n_743),
.Y(n_892)
);

AOI21xp5_ASAP7_75t_L g893 ( 
.A1(n_639),
.A2(n_178),
.B(n_166),
.Y(n_893)
);

BUFx3_ASAP7_75t_L g894 ( 
.A(n_683),
.Y(n_894)
);

NAND2xp5_ASAP7_75t_SL g895 ( 
.A(n_718),
.B(n_184),
.Y(n_895)
);

NOR3xp33_ASAP7_75t_SL g896 ( 
.A(n_684),
.B(n_667),
.C(n_690),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_691),
.B(n_25),
.Y(n_897)
);

OA22x2_ASAP7_75t_L g898 ( 
.A1(n_665),
.A2(n_25),
.B1(n_26),
.B2(n_28),
.Y(n_898)
);

INVx2_ASAP7_75t_SL g899 ( 
.A(n_683),
.Y(n_899)
);

NOR2xp33_ASAP7_75t_L g900 ( 
.A(n_696),
.B(n_29),
.Y(n_900)
);

NAND2xp5_ASAP7_75t_L g901 ( 
.A(n_691),
.B(n_31),
.Y(n_901)
);

AND2x2_ASAP7_75t_L g902 ( 
.A(n_722),
.B(n_34),
.Y(n_902)
);

BUFx6f_ASAP7_75t_L g903 ( 
.A(n_607),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_718),
.B(n_178),
.Y(n_904)
);

NAND2x1p5_ASAP7_75t_L g905 ( 
.A(n_680),
.B(n_178),
.Y(n_905)
);

BUFx6f_ASAP7_75t_L g906 ( 
.A(n_643),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_SL g907 ( 
.A(n_600),
.B(n_663),
.Y(n_907)
);

INVx2_ASAP7_75t_L g908 ( 
.A(n_671),
.Y(n_908)
);

O2A1O1Ixp33_ASAP7_75t_L g909 ( 
.A1(n_647),
.A2(n_667),
.B(n_795),
.C(n_791),
.Y(n_909)
);

BUFx6f_ASAP7_75t_L g910 ( 
.A(n_643),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_680),
.A2(n_166),
.B(n_161),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_649),
.A2(n_166),
.B(n_161),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_656),
.A2(n_34),
.B(n_35),
.C(n_36),
.Y(n_913)
);

AOI21xp5_ASAP7_75t_L g914 ( 
.A1(n_614),
.A2(n_178),
.B(n_166),
.Y(n_914)
);

NOR2xp67_ASAP7_75t_L g915 ( 
.A(n_619),
.B(n_37),
.Y(n_915)
);

NOR2xp33_ASAP7_75t_L g916 ( 
.A(n_629),
.B(n_38),
.Y(n_916)
);

AOI21xp5_ASAP7_75t_L g917 ( 
.A1(n_784),
.A2(n_166),
.B(n_161),
.Y(n_917)
);

INVx6_ASAP7_75t_L g918 ( 
.A(n_643),
.Y(n_918)
);

BUFx4f_ASAP7_75t_L g919 ( 
.A(n_663),
.Y(n_919)
);

NAND2xp5_ASAP7_75t_L g920 ( 
.A(n_691),
.B(n_38),
.Y(n_920)
);

INVx8_ASAP7_75t_L g921 ( 
.A(n_643),
.Y(n_921)
);

AOI22xp5_ASAP7_75t_L g922 ( 
.A1(n_783),
.A2(n_178),
.B1(n_166),
.B2(n_161),
.Y(n_922)
);

O2A1O1Ixp33_ASAP7_75t_L g923 ( 
.A1(n_789),
.A2(n_39),
.B(n_40),
.C(n_42),
.Y(n_923)
);

OAI22x1_ASAP7_75t_L g924 ( 
.A1(n_757),
.A2(n_40),
.B1(n_42),
.B2(n_43),
.Y(n_924)
);

OAI22xp5_ASAP7_75t_L g925 ( 
.A1(n_762),
.A2(n_178),
.B1(n_166),
.B2(n_161),
.Y(n_925)
);

CKINVDCx14_ASAP7_75t_R g926 ( 
.A(n_741),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_671),
.Y(n_927)
);

CKINVDCx8_ASAP7_75t_R g928 ( 
.A(n_741),
.Y(n_928)
);

AOI221x1_ASAP7_75t_L g929 ( 
.A1(n_648),
.A2(n_708),
.B1(n_737),
.B2(n_761),
.C(n_612),
.Y(n_929)
);

BUFx6f_ASAP7_75t_L g930 ( 
.A(n_661),
.Y(n_930)
);

AO32x1_ASAP7_75t_L g931 ( 
.A1(n_609),
.A2(n_46),
.A3(n_47),
.B1(n_51),
.B2(n_52),
.Y(n_931)
);

AOI21xp5_ASAP7_75t_L g932 ( 
.A1(n_724),
.A2(n_738),
.B(n_685),
.Y(n_932)
);

BUFx6f_ASAP7_75t_L g933 ( 
.A(n_661),
.Y(n_933)
);

INVx3_ASAP7_75t_L g934 ( 
.A(n_763),
.Y(n_934)
);

BUFx6f_ASAP7_75t_L g935 ( 
.A(n_661),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_L g936 ( 
.A(n_690),
.B(n_46),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_SL g937 ( 
.A(n_600),
.B(n_161),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_SL g938 ( 
.A(n_628),
.B(n_161),
.Y(n_938)
);

O2A1O1Ixp33_ASAP7_75t_L g939 ( 
.A1(n_801),
.A2(n_53),
.B(n_54),
.C(n_55),
.Y(n_939)
);

O2A1O1Ixp5_ASAP7_75t_SL g940 ( 
.A1(n_726),
.A2(n_53),
.B(n_54),
.C(n_161),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_723),
.A2(n_161),
.B(n_166),
.Y(n_941)
);

OR2x2_ASAP7_75t_L g942 ( 
.A(n_638),
.B(n_161),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_790),
.Y(n_943)
);

O2A1O1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_801),
.A2(n_166),
.B(n_178),
.C(n_773),
.Y(n_944)
);

A2O1A1Ixp33_ASAP7_75t_L g945 ( 
.A1(n_712),
.A2(n_166),
.B(n_178),
.C(n_752),
.Y(n_945)
);

OAI21x1_ASAP7_75t_L g946 ( 
.A1(n_652),
.A2(n_706),
.B(n_707),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_776),
.B(n_733),
.Y(n_947)
);

BUFx3_ASAP7_75t_L g948 ( 
.A(n_705),
.Y(n_948)
);

AND2x2_ASAP7_75t_L g949 ( 
.A(n_733),
.B(n_178),
.Y(n_949)
);

A2O1A1Ixp33_ASAP7_75t_L g950 ( 
.A1(n_786),
.A2(n_178),
.B(n_687),
.C(n_692),
.Y(n_950)
);

BUFx6f_ASAP7_75t_L g951 ( 
.A(n_661),
.Y(n_951)
);

INVxp67_ASAP7_75t_L g952 ( 
.A(n_670),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_797),
.Y(n_953)
);

INVx4_ASAP7_75t_L g954 ( 
.A(n_662),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_L g955 ( 
.A(n_644),
.B(n_178),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_717),
.A2(n_178),
.B(n_755),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_675),
.B(n_676),
.Y(n_957)
);

INVx2_ASAP7_75t_L g958 ( 
.A(n_673),
.Y(n_958)
);

INVx2_ASAP7_75t_L g959 ( 
.A(n_673),
.Y(n_959)
);

NAND2xp5_ASAP7_75t_SL g960 ( 
.A(n_637),
.B(n_728),
.Y(n_960)
);

AOI22xp5_ASAP7_75t_L g961 ( 
.A1(n_755),
.A2(n_698),
.B1(n_700),
.B2(n_747),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_728),
.B(n_713),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_R g963 ( 
.A(n_731),
.B(n_782),
.Y(n_963)
);

OAI22x1_ASAP7_75t_L g964 ( 
.A1(n_634),
.A2(n_753),
.B1(n_798),
.B2(n_624),
.Y(n_964)
);

A2O1A1Ixp33_ASAP7_75t_L g965 ( 
.A1(n_622),
.A2(n_720),
.B(n_730),
.C(n_740),
.Y(n_965)
);

BUFx6f_ASAP7_75t_L g966 ( 
.A(n_662),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_704),
.Y(n_967)
);

CKINVDCx14_ASAP7_75t_R g968 ( 
.A(n_749),
.Y(n_968)
);

OAI22xp5_ASAP7_75t_L g969 ( 
.A1(n_729),
.A2(n_709),
.B1(n_745),
.B2(n_715),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_763),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_799),
.B(n_760),
.Y(n_971)
);

NOR2x1_ASAP7_75t_L g972 ( 
.A(n_709),
.B(n_760),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_744),
.A2(n_736),
.B1(n_785),
.B2(n_719),
.Y(n_973)
);

BUFx6f_ASAP7_75t_L g974 ( 
.A(n_662),
.Y(n_974)
);

A2O1A1Ixp33_ASAP7_75t_L g975 ( 
.A1(n_744),
.A2(n_727),
.B(n_782),
.C(n_756),
.Y(n_975)
);

NOR2xp67_ASAP7_75t_SL g976 ( 
.A(n_662),
.B(n_674),
.Y(n_976)
);

BUFx2_ASAP7_75t_L g977 ( 
.A(n_763),
.Y(n_977)
);

INVxp67_ASAP7_75t_L g978 ( 
.A(n_799),
.Y(n_978)
);

O2A1O1Ixp33_ASAP7_75t_SL g979 ( 
.A1(n_742),
.A2(n_788),
.B(n_719),
.C(n_751),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_704),
.Y(n_980)
);

NAND2xp5_ASAP7_75t_SL g981 ( 
.A(n_764),
.B(n_766),
.Y(n_981)
);

OR2x2_ASAP7_75t_L g982 ( 
.A(n_750),
.B(n_794),
.Y(n_982)
);

OAI21xp5_ASAP7_75t_L g983 ( 
.A1(n_725),
.A2(n_734),
.B(n_772),
.Y(n_983)
);

INVx4_ASAP7_75t_L g984 ( 
.A(n_669),
.Y(n_984)
);

BUFx2_ASAP7_75t_L g985 ( 
.A(n_763),
.Y(n_985)
);

OAI22xp5_ASAP7_75t_L g986 ( 
.A1(n_785),
.A2(n_674),
.B1(n_669),
.B2(n_794),
.Y(n_986)
);

BUFx3_ASAP7_75t_L g987 ( 
.A(n_774),
.Y(n_987)
);

INVx1_ASAP7_75t_L g988 ( 
.A(n_750),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_774),
.B(n_711),
.Y(n_989)
);

HB1xp67_ASAP7_75t_L g990 ( 
.A(n_669),
.Y(n_990)
);

NOR2xp33_ASAP7_75t_L g991 ( 
.A(n_774),
.B(n_674),
.Y(n_991)
);

HB1xp67_ASAP7_75t_L g992 ( 
.A(n_669),
.Y(n_992)
);

OAI21x1_ASAP7_75t_L g993 ( 
.A1(n_703),
.A2(n_739),
.B(n_646),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_616),
.A2(n_625),
.B(n_633),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_788),
.A2(n_742),
.B(n_792),
.C(n_787),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_774),
.Y(n_996)
);

AND2x4_ASAP7_75t_L g997 ( 
.A(n_674),
.B(n_748),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_L g998 ( 
.A(n_749),
.B(n_793),
.Y(n_998)
);

NAND2xp5_ASAP7_75t_L g999 ( 
.A(n_758),
.B(n_800),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_636),
.A2(n_645),
.B(n_759),
.Y(n_1000)
);

INVx1_ASAP7_75t_L g1001 ( 
.A(n_777),
.Y(n_1001)
);

NAND2xp5_ASAP7_75t_SL g1002 ( 
.A(n_765),
.B(n_778),
.Y(n_1002)
);

NAND3xp33_ASAP7_75t_L g1003 ( 
.A(n_780),
.B(n_781),
.C(n_768),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_767),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_771),
.A2(n_482),
.B(n_640),
.C(n_428),
.Y(n_1005)
);

NOR2xp33_ASAP7_75t_R g1006 ( 
.A(n_664),
.B(n_341),
.Y(n_1006)
);

INVx1_ASAP7_75t_L g1007 ( 
.A(n_686),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_640),
.A2(n_599),
.B(n_482),
.C(n_679),
.Y(n_1008)
);

INVx1_ASAP7_75t_L g1009 ( 
.A(n_686),
.Y(n_1009)
);

OAI21xp33_ASAP7_75t_L g1010 ( 
.A1(n_684),
.A2(n_482),
.B(n_415),
.Y(n_1010)
);

NOR2xp33_ASAP7_75t_L g1011 ( 
.A(n_617),
.B(n_500),
.Y(n_1011)
);

A2O1A1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_640),
.A2(n_599),
.B(n_482),
.C(n_679),
.Y(n_1012)
);

INVx1_ASAP7_75t_L g1013 ( 
.A(n_686),
.Y(n_1013)
);

AOI21xp5_ASAP7_75t_L g1014 ( 
.A1(n_770),
.A2(n_541),
.B(n_528),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_601),
.B(n_427),
.Y(n_1015)
);

NAND2xp33_ASAP7_75t_L g1016 ( 
.A(n_691),
.B(n_341),
.Y(n_1016)
);

AOI21xp5_ASAP7_75t_L g1017 ( 
.A1(n_770),
.A2(n_541),
.B(n_528),
.Y(n_1017)
);

NOR2xp33_ASAP7_75t_L g1018 ( 
.A(n_617),
.B(n_500),
.Y(n_1018)
);

OAI22xp5_ASAP7_75t_L g1019 ( 
.A1(n_693),
.A2(n_301),
.B1(n_353),
.B2(n_341),
.Y(n_1019)
);

AOI21xp5_ASAP7_75t_L g1020 ( 
.A1(n_770),
.A2(n_541),
.B(n_528),
.Y(n_1020)
);

AOI22xp5_ASAP7_75t_L g1021 ( 
.A1(n_632),
.A2(n_482),
.B1(n_341),
.B2(n_353),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_664),
.Y(n_1022)
);

INVx1_ASAP7_75t_L g1023 ( 
.A(n_686),
.Y(n_1023)
);

INVx2_ASAP7_75t_L g1024 ( 
.A(n_602),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_SL g1025 ( 
.A(n_601),
.B(n_427),
.Y(n_1025)
);

BUFx2_ASAP7_75t_L g1026 ( 
.A(n_605),
.Y(n_1026)
);

AO32x2_ASAP7_75t_L g1027 ( 
.A1(n_702),
.A2(n_708),
.A3(n_612),
.B1(n_609),
.B2(n_648),
.Y(n_1027)
);

INVx3_ASAP7_75t_L g1028 ( 
.A(n_653),
.Y(n_1028)
);

AOI21xp5_ASAP7_75t_L g1029 ( 
.A1(n_770),
.A2(n_541),
.B(n_528),
.Y(n_1029)
);

NAND3x1_ASAP7_75t_L g1030 ( 
.A(n_658),
.B(n_355),
.C(n_352),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_L g1031 ( 
.A(n_620),
.B(n_210),
.Y(n_1031)
);

AOI22xp5_ASAP7_75t_L g1032 ( 
.A1(n_632),
.A2(n_482),
.B1(n_341),
.B2(n_353),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_686),
.Y(n_1033)
);

BUFx6f_ASAP7_75t_L g1034 ( 
.A(n_607),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_686),
.Y(n_1035)
);

A2O1A1Ixp33_ASAP7_75t_L g1036 ( 
.A1(n_640),
.A2(n_599),
.B(n_482),
.C(n_679),
.Y(n_1036)
);

O2A1O1Ixp5_ASAP7_75t_SL g1037 ( 
.A1(n_775),
.A2(n_702),
.B(n_513),
.C(n_612),
.Y(n_1037)
);

NOR2xp33_ASAP7_75t_SL g1038 ( 
.A(n_664),
.B(n_431),
.Y(n_1038)
);

AND2x2_ASAP7_75t_L g1039 ( 
.A(n_632),
.B(n_467),
.Y(n_1039)
);

A2O1A1Ixp33_ASAP7_75t_L g1040 ( 
.A1(n_640),
.A2(n_599),
.B(n_482),
.C(n_679),
.Y(n_1040)
);

INVx2_ASAP7_75t_L g1041 ( 
.A(n_805),
.Y(n_1041)
);

AND2x2_ASAP7_75t_L g1042 ( 
.A(n_971),
.B(n_823),
.Y(n_1042)
);

BUFx3_ASAP7_75t_L g1043 ( 
.A(n_802),
.Y(n_1043)
);

INVx2_ASAP7_75t_SL g1044 ( 
.A(n_921),
.Y(n_1044)
);

BUFx6f_ASAP7_75t_L g1045 ( 
.A(n_850),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_1031),
.B(n_871),
.Y(n_1046)
);

AO21x2_ASAP7_75t_L g1047 ( 
.A1(n_864),
.A2(n_869),
.B(n_861),
.Y(n_1047)
);

INVx1_ASAP7_75t_SL g1048 ( 
.A(n_1026),
.Y(n_1048)
);

AND2x4_ASAP7_75t_L g1049 ( 
.A(n_804),
.B(n_838),
.Y(n_1049)
);

NOR2xp33_ASAP7_75t_L g1050 ( 
.A(n_1021),
.B(n_1032),
.Y(n_1050)
);

NAND2x1p5_ASAP7_75t_L g1051 ( 
.A(n_868),
.B(n_819),
.Y(n_1051)
);

AND2x4_ASAP7_75t_L g1052 ( 
.A(n_804),
.B(n_838),
.Y(n_1052)
);

NAND2xp5_ASAP7_75t_L g1053 ( 
.A(n_1010),
.B(n_1011),
.Y(n_1053)
);

BUFx8_ASAP7_75t_SL g1054 ( 
.A(n_839),
.Y(n_1054)
);

INVx3_ASAP7_75t_L g1055 ( 
.A(n_840),
.Y(n_1055)
);

INVx3_ASAP7_75t_L g1056 ( 
.A(n_840),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_902),
.B(n_896),
.Y(n_1057)
);

AND2x4_ASAP7_75t_L g1058 ( 
.A(n_842),
.B(n_1028),
.Y(n_1058)
);

BUFx6f_ASAP7_75t_L g1059 ( 
.A(n_850),
.Y(n_1059)
);

CKINVDCx6p67_ASAP7_75t_R g1060 ( 
.A(n_882),
.Y(n_1060)
);

INVx5_ASAP7_75t_SL g1061 ( 
.A(n_829),
.Y(n_1061)
);

INVx6_ASAP7_75t_L g1062 ( 
.A(n_878),
.Y(n_1062)
);

INVx5_ASAP7_75t_L g1063 ( 
.A(n_850),
.Y(n_1063)
);

INVx2_ASAP7_75t_L g1064 ( 
.A(n_807),
.Y(n_1064)
);

AOI22xp5_ASAP7_75t_L g1065 ( 
.A1(n_873),
.A2(n_885),
.B1(n_1030),
.B2(n_900),
.Y(n_1065)
);

NAND2x1p5_ASAP7_75t_L g1066 ( 
.A(n_819),
.B(n_962),
.Y(n_1066)
);

INVx3_ASAP7_75t_L g1067 ( 
.A(n_888),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_988),
.Y(n_1068)
);

INVx5_ASAP7_75t_SL g1069 ( 
.A(n_829),
.Y(n_1069)
);

BUFx3_ASAP7_75t_L g1070 ( 
.A(n_894),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_879),
.Y(n_1071)
);

BUFx3_ASAP7_75t_L g1072 ( 
.A(n_878),
.Y(n_1072)
);

BUFx6f_ASAP7_75t_L g1073 ( 
.A(n_850),
.Y(n_1073)
);

BUFx12f_ASAP7_75t_L g1074 ( 
.A(n_821),
.Y(n_1074)
);

BUFx6f_ASAP7_75t_L g1075 ( 
.A(n_860),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_943),
.Y(n_1076)
);

BUFx12f_ASAP7_75t_L g1077 ( 
.A(n_1022),
.Y(n_1077)
);

INVxp67_ASAP7_75t_SL g1078 ( 
.A(n_976),
.Y(n_1078)
);

BUFx2_ASAP7_75t_L g1079 ( 
.A(n_952),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_953),
.Y(n_1080)
);

NAND2xp5_ASAP7_75t_L g1081 ( 
.A(n_1011),
.B(n_1018),
.Y(n_1081)
);

CKINVDCx16_ASAP7_75t_R g1082 ( 
.A(n_1038),
.Y(n_1082)
);

INVx1_ASAP7_75t_L g1083 ( 
.A(n_856),
.Y(n_1083)
);

BUFx6f_ASAP7_75t_L g1084 ( 
.A(n_860),
.Y(n_1084)
);

BUFx3_ASAP7_75t_L g1085 ( 
.A(n_899),
.Y(n_1085)
);

INVx2_ASAP7_75t_SL g1086 ( 
.A(n_921),
.Y(n_1086)
);

NAND2xp5_ASAP7_75t_L g1087 ( 
.A(n_1018),
.B(n_1039),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_896),
.B(n_978),
.Y(n_1088)
);

BUFx2_ASAP7_75t_L g1089 ( 
.A(n_952),
.Y(n_1089)
);

INVxp67_ASAP7_75t_SL g1090 ( 
.A(n_947),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_857),
.Y(n_1091)
);

INVx6_ASAP7_75t_SL g1092 ( 
.A(n_997),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_863),
.Y(n_1093)
);

INVx1_ASAP7_75t_SL g1094 ( 
.A(n_892),
.Y(n_1094)
);

BUFx6f_ASAP7_75t_L g1095 ( 
.A(n_860),
.Y(n_1095)
);

INVx3_ASAP7_75t_SL g1096 ( 
.A(n_921),
.Y(n_1096)
);

OR2x6_ASAP7_75t_L g1097 ( 
.A(n_814),
.B(n_815),
.Y(n_1097)
);

NOR2xp33_ASAP7_75t_SL g1098 ( 
.A(n_919),
.B(n_928),
.Y(n_1098)
);

INVx5_ASAP7_75t_L g1099 ( 
.A(n_860),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_816),
.Y(n_1100)
);

BUFx3_ASAP7_75t_L g1101 ( 
.A(n_948),
.Y(n_1101)
);

BUFx2_ASAP7_75t_SL g1102 ( 
.A(n_903),
.Y(n_1102)
);

NOR2xp33_ASAP7_75t_L g1103 ( 
.A(n_1019),
.B(n_926),
.Y(n_1103)
);

BUFx6f_ASAP7_75t_L g1104 ( 
.A(n_903),
.Y(n_1104)
);

BUFx5_ASAP7_75t_L g1105 ( 
.A(n_1001),
.Y(n_1105)
);

INVx2_ASAP7_75t_SL g1106 ( 
.A(n_918),
.Y(n_1106)
);

NAND2x1p5_ASAP7_75t_L g1107 ( 
.A(n_962),
.B(n_907),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_826),
.Y(n_1108)
);

CKINVDCx8_ASAP7_75t_R g1109 ( 
.A(n_977),
.Y(n_1109)
);

NOR2xp33_ASAP7_75t_L g1110 ( 
.A(n_836),
.B(n_835),
.Y(n_1110)
);

NAND2xp5_ASAP7_75t_L g1111 ( 
.A(n_808),
.B(n_813),
.Y(n_1111)
);

BUFx2_ASAP7_75t_SL g1112 ( 
.A(n_903),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_1006),
.Y(n_1113)
);

INVxp67_ASAP7_75t_SL g1114 ( 
.A(n_808),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_872),
.Y(n_1115)
);

INVx8_ASAP7_75t_L g1116 ( 
.A(n_903),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_1006),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_842),
.Y(n_1118)
);

INVx4_ASAP7_75t_L g1119 ( 
.A(n_906),
.Y(n_1119)
);

BUFx4_ASAP7_75t_SL g1120 ( 
.A(n_846),
.Y(n_1120)
);

BUFx12f_ASAP7_75t_L g1121 ( 
.A(n_865),
.Y(n_1121)
);

BUFx2_ASAP7_75t_SL g1122 ( 
.A(n_906),
.Y(n_1122)
);

INVx3_ASAP7_75t_L g1123 ( 
.A(n_888),
.Y(n_1123)
);

BUFx12f_ASAP7_75t_L g1124 ( 
.A(n_866),
.Y(n_1124)
);

INVx1_ASAP7_75t_L g1125 ( 
.A(n_874),
.Y(n_1125)
);

BUFx5_ASAP7_75t_L g1126 ( 
.A(n_1004),
.Y(n_1126)
);

BUFx3_ASAP7_75t_L g1127 ( 
.A(n_1028),
.Y(n_1127)
);

INVx3_ASAP7_75t_SL g1128 ( 
.A(n_918),
.Y(n_1128)
);

INVxp67_ASAP7_75t_SL g1129 ( 
.A(n_813),
.Y(n_1129)
);

INVx5_ASAP7_75t_L g1130 ( 
.A(n_906),
.Y(n_1130)
);

HB1xp67_ASAP7_75t_L g1131 ( 
.A(n_845),
.Y(n_1131)
);

BUFx6f_ASAP7_75t_L g1132 ( 
.A(n_906),
.Y(n_1132)
);

INVx3_ASAP7_75t_L g1133 ( 
.A(n_910),
.Y(n_1133)
);

NAND2xp5_ASAP7_75t_L g1134 ( 
.A(n_844),
.B(n_852),
.Y(n_1134)
);

INVx3_ASAP7_75t_SL g1135 ( 
.A(n_918),
.Y(n_1135)
);

INVx3_ASAP7_75t_L g1136 ( 
.A(n_910),
.Y(n_1136)
);

CKINVDCx14_ASAP7_75t_R g1137 ( 
.A(n_877),
.Y(n_1137)
);

INVx3_ASAP7_75t_L g1138 ( 
.A(n_910),
.Y(n_1138)
);

AND2x2_ASAP7_75t_L g1139 ( 
.A(n_978),
.B(n_916),
.Y(n_1139)
);

BUFx2_ASAP7_75t_SL g1140 ( 
.A(n_910),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_985),
.Y(n_1141)
);

OAI22xp5_ASAP7_75t_L g1142 ( 
.A1(n_919),
.A2(n_1008),
.B1(n_1036),
.B2(n_1012),
.Y(n_1142)
);

INVx3_ASAP7_75t_SL g1143 ( 
.A(n_831),
.Y(n_1143)
);

INVx2_ASAP7_75t_SL g1144 ( 
.A(n_987),
.Y(n_1144)
);

BUFx3_ASAP7_75t_L g1145 ( 
.A(n_930),
.Y(n_1145)
);

AND2x2_ASAP7_75t_L g1146 ( 
.A(n_916),
.B(n_828),
.Y(n_1146)
);

NAND2xp5_ASAP7_75t_L g1147 ( 
.A(n_844),
.B(n_852),
.Y(n_1147)
);

BUFx6f_ASAP7_75t_SL g1148 ( 
.A(n_866),
.Y(n_1148)
);

INVx2_ASAP7_75t_SL g1149 ( 
.A(n_930),
.Y(n_1149)
);

INVx6_ASAP7_75t_L g1150 ( 
.A(n_810),
.Y(n_1150)
);

BUFx3_ASAP7_75t_L g1151 ( 
.A(n_930),
.Y(n_1151)
);

BUFx4_ASAP7_75t_SL g1152 ( 
.A(n_996),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_883),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_930),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_886),
.Y(n_1155)
);

BUFx6f_ASAP7_75t_L g1156 ( 
.A(n_933),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_908),
.Y(n_1157)
);

BUFx4_ASAP7_75t_SL g1158 ( 
.A(n_803),
.Y(n_1158)
);

BUFx3_ASAP7_75t_L g1159 ( 
.A(n_933),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_927),
.Y(n_1160)
);

AOI22xp33_ASAP7_75t_L g1161 ( 
.A1(n_873),
.A2(n_885),
.B1(n_833),
.B2(n_830),
.Y(n_1161)
);

INVx3_ASAP7_75t_L g1162 ( 
.A(n_933),
.Y(n_1162)
);

BUFx8_ASAP7_75t_L g1163 ( 
.A(n_997),
.Y(n_1163)
);

INVx1_ASAP7_75t_L g1164 ( 
.A(n_958),
.Y(n_1164)
);

BUFx3_ASAP7_75t_L g1165 ( 
.A(n_933),
.Y(n_1165)
);

INVx2_ASAP7_75t_SL g1166 ( 
.A(n_935),
.Y(n_1166)
);

INVx2_ASAP7_75t_L g1167 ( 
.A(n_959),
.Y(n_1167)
);

INVx2_ASAP7_75t_SL g1168 ( 
.A(n_935),
.Y(n_1168)
);

INVx2_ASAP7_75t_L g1169 ( 
.A(n_967),
.Y(n_1169)
);

BUFx3_ASAP7_75t_L g1170 ( 
.A(n_935),
.Y(n_1170)
);

BUFx12f_ASAP7_75t_L g1171 ( 
.A(n_935),
.Y(n_1171)
);

CKINVDCx20_ASAP7_75t_R g1172 ( 
.A(n_968),
.Y(n_1172)
);

BUFx3_ASAP7_75t_L g1173 ( 
.A(n_951),
.Y(n_1173)
);

CKINVDCx6p67_ASAP7_75t_R g1174 ( 
.A(n_924),
.Y(n_1174)
);

AOI22xp33_ASAP7_75t_L g1175 ( 
.A1(n_833),
.A2(n_820),
.B1(n_1025),
.B2(n_1015),
.Y(n_1175)
);

INVx1_ASAP7_75t_SL g1176 ( 
.A(n_942),
.Y(n_1176)
);

BUFx2_ASAP7_75t_L g1177 ( 
.A(n_990),
.Y(n_1177)
);

BUFx3_ASAP7_75t_L g1178 ( 
.A(n_951),
.Y(n_1178)
);

HB1xp67_ASAP7_75t_L g1179 ( 
.A(n_990),
.Y(n_1179)
);

NOR2xp67_ASAP7_75t_L g1180 ( 
.A(n_834),
.B(n_961),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_980),
.Y(n_1181)
);

INVx1_ASAP7_75t_SL g1182 ( 
.A(n_992),
.Y(n_1182)
);

BUFx2_ASAP7_75t_L g1183 ( 
.A(n_992),
.Y(n_1183)
);

BUFx12f_ASAP7_75t_L g1184 ( 
.A(n_966),
.Y(n_1184)
);

INVx3_ASAP7_75t_L g1185 ( 
.A(n_966),
.Y(n_1185)
);

CKINVDCx5p33_ASAP7_75t_R g1186 ( 
.A(n_934),
.Y(n_1186)
);

INVx2_ASAP7_75t_L g1187 ( 
.A(n_1024),
.Y(n_1187)
);

BUFx6f_ASAP7_75t_L g1188 ( 
.A(n_966),
.Y(n_1188)
);

INVx1_ASAP7_75t_L g1189 ( 
.A(n_982),
.Y(n_1189)
);

BUFx3_ASAP7_75t_L g1190 ( 
.A(n_966),
.Y(n_1190)
);

BUFx4_ASAP7_75t_SL g1191 ( 
.A(n_812),
.Y(n_1191)
);

CKINVDCx16_ASAP7_75t_R g1192 ( 
.A(n_963),
.Y(n_1192)
);

BUFx5_ASAP7_75t_L g1193 ( 
.A(n_949),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_946),
.Y(n_1194)
);

BUFx2_ASAP7_75t_L g1195 ( 
.A(n_964),
.Y(n_1195)
);

INVx6_ASAP7_75t_L g1196 ( 
.A(n_810),
.Y(n_1196)
);

BUFx3_ASAP7_75t_L g1197 ( 
.A(n_974),
.Y(n_1197)
);

BUFx3_ASAP7_75t_L g1198 ( 
.A(n_974),
.Y(n_1198)
);

CKINVDCx20_ASAP7_75t_R g1199 ( 
.A(n_936),
.Y(n_1199)
);

BUFx3_ASAP7_75t_L g1200 ( 
.A(n_974),
.Y(n_1200)
);

BUFx2_ASAP7_75t_L g1201 ( 
.A(n_855),
.Y(n_1201)
);

BUFx2_ASAP7_75t_L g1202 ( 
.A(n_963),
.Y(n_1202)
);

INVx5_ASAP7_75t_L g1203 ( 
.A(n_974),
.Y(n_1203)
);

BUFx8_ASAP7_75t_L g1204 ( 
.A(n_1034),
.Y(n_1204)
);

BUFx2_ASAP7_75t_L g1205 ( 
.A(n_972),
.Y(n_1205)
);

CKINVDCx11_ASAP7_75t_R g1206 ( 
.A(n_1034),
.Y(n_1206)
);

AOI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_820),
.A2(n_1025),
.B1(n_1015),
.B2(n_900),
.Y(n_1207)
);

NAND2x1p5_ASAP7_75t_L g1208 ( 
.A(n_907),
.B(n_960),
.Y(n_1208)
);

INVxp67_ASAP7_75t_SL g1209 ( 
.A(n_806),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_897),
.Y(n_1210)
);

AND2x6_ASAP7_75t_L g1211 ( 
.A(n_957),
.B(n_901),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1040),
.B(n_1005),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_898),
.B(n_858),
.Y(n_1213)
);

BUFx2_ASAP7_75t_SL g1214 ( 
.A(n_1034),
.Y(n_1214)
);

INVx2_ASAP7_75t_L g1215 ( 
.A(n_824),
.Y(n_1215)
);

INVx1_ASAP7_75t_L g1216 ( 
.A(n_848),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_1034),
.Y(n_1217)
);

BUFx2_ASAP7_75t_L g1218 ( 
.A(n_1027),
.Y(n_1218)
);

BUFx2_ASAP7_75t_SL g1219 ( 
.A(n_954),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_849),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1007),
.Y(n_1221)
);

BUFx2_ASAP7_75t_SL g1222 ( 
.A(n_954),
.Y(n_1222)
);

BUFx2_ASAP7_75t_L g1223 ( 
.A(n_1027),
.Y(n_1223)
);

INVx1_ASAP7_75t_SL g1224 ( 
.A(n_1009),
.Y(n_1224)
);

BUFx3_ASAP7_75t_L g1225 ( 
.A(n_934),
.Y(n_1225)
);

INVx2_ASAP7_75t_L g1226 ( 
.A(n_1013),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_891),
.Y(n_1227)
);

INVx2_ASAP7_75t_L g1228 ( 
.A(n_1023),
.Y(n_1228)
);

NAND2xp5_ASAP7_75t_L g1229 ( 
.A(n_909),
.B(n_1033),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1035),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_970),
.Y(n_1231)
);

INVx4_ASAP7_75t_L g1232 ( 
.A(n_984),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_984),
.Y(n_1233)
);

BUFx4_ASAP7_75t_SL g1234 ( 
.A(n_1003),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_809),
.Y(n_1235)
);

INVx6_ASAP7_75t_L g1236 ( 
.A(n_1016),
.Y(n_1236)
);

INVx5_ASAP7_75t_L g1237 ( 
.A(n_970),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_979),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_920),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_809),
.Y(n_1240)
);

INVx3_ASAP7_75t_L g1241 ( 
.A(n_853),
.Y(n_1241)
);

BUFx3_ASAP7_75t_L g1242 ( 
.A(n_991),
.Y(n_1242)
);

INVx2_ASAP7_75t_SL g1243 ( 
.A(n_991),
.Y(n_1243)
);

CKINVDCx20_ASAP7_75t_R g1244 ( 
.A(n_937),
.Y(n_1244)
);

INVx2_ASAP7_75t_L g1245 ( 
.A(n_843),
.Y(n_1245)
);

INVx1_ASAP7_75t_SL g1246 ( 
.A(n_937),
.Y(n_1246)
);

INVx2_ASAP7_75t_L g1247 ( 
.A(n_989),
.Y(n_1247)
);

INVx3_ASAP7_75t_L g1248 ( 
.A(n_905),
.Y(n_1248)
);

INVx1_ASAP7_75t_L g1249 ( 
.A(n_1027),
.Y(n_1249)
);

BUFx3_ASAP7_75t_L g1250 ( 
.A(n_998),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_898),
.Y(n_1251)
);

NAND2xp5_ASAP7_75t_L g1252 ( 
.A(n_851),
.B(n_862),
.Y(n_1252)
);

INVx6_ASAP7_75t_L g1253 ( 
.A(n_986),
.Y(n_1253)
);

AND2x4_ASAP7_75t_L g1254 ( 
.A(n_981),
.B(n_822),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_905),
.Y(n_1255)
);

INVx1_ASAP7_75t_SL g1256 ( 
.A(n_895),
.Y(n_1256)
);

BUFx3_ASAP7_75t_L g1257 ( 
.A(n_999),
.Y(n_1257)
);

INVx2_ASAP7_75t_L g1258 ( 
.A(n_955),
.Y(n_1258)
);

NAND2x1p5_ASAP7_75t_L g1259 ( 
.A(n_960),
.B(n_1002),
.Y(n_1259)
);

AOI22xp5_ASAP7_75t_L g1260 ( 
.A1(n_915),
.A2(n_862),
.B1(n_854),
.B2(n_851),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1027),
.Y(n_1261)
);

NAND2xp5_ASAP7_75t_L g1262 ( 
.A(n_854),
.B(n_939),
.Y(n_1262)
);

INVx2_ASAP7_75t_R g1263 ( 
.A(n_929),
.Y(n_1263)
);

BUFx3_ASAP7_75t_L g1264 ( 
.A(n_867),
.Y(n_1264)
);

AO21x2_ASAP7_75t_L g1265 ( 
.A1(n_1194),
.A2(n_834),
.B(n_983),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1235),
.Y(n_1266)
);

OAI21x1_ASAP7_75t_L g1267 ( 
.A1(n_1241),
.A2(n_993),
.B(n_994),
.Y(n_1267)
);

OAI22xp5_ASAP7_75t_L g1268 ( 
.A1(n_1065),
.A2(n_973),
.B1(n_975),
.B2(n_890),
.Y(n_1268)
);

AOI21xp5_ASAP7_75t_L g1269 ( 
.A1(n_1142),
.A2(n_1014),
.B(n_1020),
.Y(n_1269)
);

OAI22xp5_ASAP7_75t_L g1270 ( 
.A1(n_1065),
.A2(n_889),
.B1(n_965),
.B2(n_923),
.Y(n_1270)
);

NOR2x1_ASAP7_75t_R g1271 ( 
.A(n_1062),
.B(n_981),
.Y(n_1271)
);

INVx2_ASAP7_75t_L g1272 ( 
.A(n_1247),
.Y(n_1272)
);

BUFx8_ASAP7_75t_L g1273 ( 
.A(n_1148),
.Y(n_1273)
);

AOI22xp33_ASAP7_75t_L g1274 ( 
.A1(n_1161),
.A2(n_1050),
.B1(n_1174),
.B2(n_1057),
.Y(n_1274)
);

CKINVDCx20_ASAP7_75t_R g1275 ( 
.A(n_1054),
.Y(n_1275)
);

CKINVDCx9p33_ASAP7_75t_R g1276 ( 
.A(n_1202),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1042),
.B(n_825),
.Y(n_1277)
);

AOI22xp33_ASAP7_75t_SL g1278 ( 
.A1(n_1251),
.A2(n_1091),
.B1(n_1192),
.B2(n_1262),
.Y(n_1278)
);

AO21x2_ASAP7_75t_L g1279 ( 
.A1(n_1194),
.A2(n_945),
.B(n_932),
.Y(n_1279)
);

OAI21x1_ASAP7_75t_L g1280 ( 
.A1(n_1241),
.A2(n_1000),
.B(n_1017),
.Y(n_1280)
);

AO31x2_ASAP7_75t_L g1281 ( 
.A1(n_1245),
.A2(n_837),
.A3(n_950),
.B(n_969),
.Y(n_1281)
);

CKINVDCx20_ASAP7_75t_R g1282 ( 
.A(n_1113),
.Y(n_1282)
);

OR2x2_ASAP7_75t_L g1283 ( 
.A(n_1201),
.B(n_904),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1201),
.B(n_904),
.Y(n_1284)
);

OAI21xp5_ASAP7_75t_L g1285 ( 
.A1(n_1212),
.A2(n_1037),
.B(n_944),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1235),
.Y(n_1286)
);

OAI21x1_ASAP7_75t_L g1287 ( 
.A1(n_1241),
.A2(n_1029),
.B(n_941),
.Y(n_1287)
);

O2A1O1Ixp33_ASAP7_75t_SL g1288 ( 
.A1(n_1111),
.A2(n_913),
.B(n_938),
.C(n_895),
.Y(n_1288)
);

OAI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1251),
.A2(n_847),
.B1(n_887),
.B2(n_859),
.Y(n_1289)
);

BUFx2_ASAP7_75t_SL g1290 ( 
.A(n_1148),
.Y(n_1290)
);

INVx1_ASAP7_75t_L g1291 ( 
.A(n_1240),
.Y(n_1291)
);

AOI21xp5_ASAP7_75t_L g1292 ( 
.A1(n_1229),
.A2(n_859),
.B(n_1002),
.Y(n_1292)
);

NAND2x1_ASAP7_75t_L g1293 ( 
.A(n_1236),
.B(n_811),
.Y(n_1293)
);

INVx1_ASAP7_75t_L g1294 ( 
.A(n_1240),
.Y(n_1294)
);

AND2x4_ASAP7_75t_L g1295 ( 
.A(n_1257),
.B(n_938),
.Y(n_1295)
);

O2A1O1Ixp33_ASAP7_75t_L g1296 ( 
.A1(n_1053),
.A2(n_876),
.B(n_979),
.C(n_995),
.Y(n_1296)
);

INVx1_ASAP7_75t_SL g1297 ( 
.A(n_1079),
.Y(n_1297)
);

INVx2_ASAP7_75t_SL g1298 ( 
.A(n_1242),
.Y(n_1298)
);

INVx1_ASAP7_75t_L g1299 ( 
.A(n_1249),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_1215),
.Y(n_1300)
);

INVx1_ASAP7_75t_L g1301 ( 
.A(n_1249),
.Y(n_1301)
);

AOI22xp33_ASAP7_75t_L g1302 ( 
.A1(n_1174),
.A2(n_870),
.B1(n_956),
.B2(n_925),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_SL g1303 ( 
.A1(n_1091),
.A2(n_931),
.B1(n_940),
.B2(n_876),
.Y(n_1303)
);

INVx2_ASAP7_75t_L g1304 ( 
.A(n_1215),
.Y(n_1304)
);

AO21x2_ASAP7_75t_L g1305 ( 
.A1(n_1180),
.A2(n_817),
.B(n_827),
.Y(n_1305)
);

AO21x2_ASAP7_75t_L g1306 ( 
.A1(n_1180),
.A2(n_832),
.B(n_841),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1057),
.A2(n_870),
.B1(n_893),
.B2(n_818),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1226),
.Y(n_1308)
);

AND2x2_ASAP7_75t_L g1309 ( 
.A(n_1042),
.B(n_922),
.Y(n_1309)
);

OAI22x1_ASAP7_75t_L g1310 ( 
.A1(n_1260),
.A2(n_931),
.B1(n_875),
.B2(n_917),
.Y(n_1310)
);

INVx3_ASAP7_75t_L g1311 ( 
.A(n_1257),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_1074),
.Y(n_1312)
);

INVx1_ASAP7_75t_L g1313 ( 
.A(n_1261),
.Y(n_1313)
);

OR2x2_ASAP7_75t_L g1314 ( 
.A(n_1146),
.B(n_884),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_1261),
.Y(n_1315)
);

INVx2_ASAP7_75t_L g1316 ( 
.A(n_1226),
.Y(n_1316)
);

AOI22xp33_ASAP7_75t_L g1317 ( 
.A1(n_1207),
.A2(n_911),
.B1(n_912),
.B2(n_880),
.Y(n_1317)
);

INVxp67_ASAP7_75t_L g1318 ( 
.A(n_1131),
.Y(n_1318)
);

NAND2xp5_ASAP7_75t_L g1319 ( 
.A(n_1046),
.B(n_881),
.Y(n_1319)
);

INVx1_ASAP7_75t_L g1320 ( 
.A(n_1083),
.Y(n_1320)
);

AOI22xp33_ASAP7_75t_L g1321 ( 
.A1(n_1146),
.A2(n_914),
.B1(n_931),
.B2(n_1143),
.Y(n_1321)
);

NOR2x1_ASAP7_75t_SL g1322 ( 
.A(n_1097),
.B(n_1238),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1114),
.B(n_1129),
.Y(n_1323)
);

OAI21xp5_ASAP7_75t_L g1324 ( 
.A1(n_1175),
.A2(n_1209),
.B(n_1259),
.Y(n_1324)
);

OR2x6_ASAP7_75t_L g1325 ( 
.A(n_1097),
.B(n_1259),
.Y(n_1325)
);

OR2x2_ASAP7_75t_L g1326 ( 
.A(n_1218),
.B(n_1223),
.Y(n_1326)
);

AOI21xp5_ASAP7_75t_L g1327 ( 
.A1(n_1257),
.A2(n_1097),
.B(n_1238),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_L g1328 ( 
.A(n_1134),
.B(n_1147),
.Y(n_1328)
);

AOI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1143),
.A2(n_1199),
.B1(n_1121),
.B2(n_1239),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_1228),
.Y(n_1330)
);

OAI21xp5_ASAP7_75t_L g1331 ( 
.A1(n_1259),
.A2(n_1254),
.B(n_1088),
.Y(n_1331)
);

NAND3xp33_ASAP7_75t_SL g1332 ( 
.A(n_1098),
.B(n_1210),
.C(n_1081),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1110),
.B(n_1090),
.Y(n_1333)
);

AND2x6_ASAP7_75t_L g1334 ( 
.A(n_1254),
.B(n_1258),
.Y(n_1334)
);

AOI22x1_ASAP7_75t_L g1335 ( 
.A1(n_1192),
.A2(n_1202),
.B1(n_1220),
.B2(n_1088),
.Y(n_1335)
);

AND2x2_ASAP7_75t_L g1336 ( 
.A(n_1213),
.B(n_1195),
.Y(n_1336)
);

A2O1A1Ixp33_ASAP7_75t_L g1337 ( 
.A1(n_1260),
.A2(n_1238),
.B(n_1103),
.C(n_1254),
.Y(n_1337)
);

AOI22xp33_ASAP7_75t_SL g1338 ( 
.A1(n_1082),
.A2(n_1238),
.B1(n_1148),
.B2(n_1121),
.Y(n_1338)
);

INVx2_ASAP7_75t_L g1339 ( 
.A(n_1228),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1163),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1083),
.Y(n_1341)
);

BUFx2_ASAP7_75t_L g1342 ( 
.A(n_1195),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_L g1343 ( 
.A1(n_1254),
.A2(n_1097),
.B(n_1066),
.Y(n_1343)
);

OAI222xp33_ASAP7_75t_L g1344 ( 
.A1(n_1208),
.A2(n_1097),
.B1(n_1107),
.B2(n_1252),
.C1(n_1066),
.C2(n_1139),
.Y(n_1344)
);

OAI21x1_ASAP7_75t_L g1345 ( 
.A1(n_1051),
.A2(n_1227),
.B(n_1258),
.Y(n_1345)
);

AND2x2_ASAP7_75t_L g1346 ( 
.A(n_1213),
.B(n_1218),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1230),
.Y(n_1347)
);

NAND2xp5_ASAP7_75t_L g1348 ( 
.A(n_1139),
.B(n_1087),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1230),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1093),
.Y(n_1350)
);

OR2x2_ASAP7_75t_L g1351 ( 
.A(n_1223),
.B(n_1047),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1051),
.A2(n_1227),
.B(n_1248),
.Y(n_1352)
);

INVx1_ASAP7_75t_L g1353 ( 
.A(n_1093),
.Y(n_1353)
);

AO21x2_ASAP7_75t_L g1354 ( 
.A1(n_1047),
.A2(n_1216),
.B(n_1076),
.Y(n_1354)
);

AOI22x1_ASAP7_75t_L g1355 ( 
.A1(n_1066),
.A2(n_1208),
.B1(n_1205),
.B2(n_1107),
.Y(n_1355)
);

OA21x2_ASAP7_75t_L g1356 ( 
.A1(n_1216),
.A2(n_1076),
.B(n_1071),
.Y(n_1356)
);

INVxp67_ASAP7_75t_L g1357 ( 
.A(n_1094),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1071),
.Y(n_1358)
);

BUFx2_ASAP7_75t_R g1359 ( 
.A(n_1072),
.Y(n_1359)
);

INVx2_ASAP7_75t_L g1360 ( 
.A(n_1080),
.Y(n_1360)
);

NAND2x1p5_ASAP7_75t_L g1361 ( 
.A(n_1238),
.B(n_1250),
.Y(n_1361)
);

INVx2_ASAP7_75t_SL g1362 ( 
.A(n_1242),
.Y(n_1362)
);

AOI22xp5_ASAP7_75t_L g1363 ( 
.A1(n_1250),
.A2(n_1082),
.B1(n_1079),
.B2(n_1089),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1089),
.B(n_1250),
.Y(n_1364)
);

OAI21x1_ASAP7_75t_SL g1365 ( 
.A1(n_1243),
.A2(n_1068),
.B(n_1080),
.Y(n_1365)
);

OAI21x1_ASAP7_75t_L g1366 ( 
.A1(n_1051),
.A2(n_1227),
.B(n_1248),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_L g1367 ( 
.A1(n_1143),
.A2(n_1211),
.B1(n_1208),
.B2(n_1263),
.Y(n_1367)
);

OAI222xp33_ASAP7_75t_L g1368 ( 
.A1(n_1107),
.A2(n_1246),
.B1(n_1244),
.B2(n_1256),
.C1(n_1048),
.C2(n_1224),
.Y(n_1368)
);

OA21x2_ASAP7_75t_L g1369 ( 
.A1(n_1221),
.A2(n_1205),
.B(n_1263),
.Y(n_1369)
);

INVx1_ASAP7_75t_SL g1370 ( 
.A(n_1182),
.Y(n_1370)
);

INVx3_ASAP7_75t_L g1371 ( 
.A(n_1163),
.Y(n_1371)
);

OAI21x1_ASAP7_75t_L g1372 ( 
.A1(n_1248),
.A2(n_1056),
.B(n_1055),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1221),
.Y(n_1373)
);

OAI21x1_ASAP7_75t_L g1374 ( 
.A1(n_1055),
.A2(n_1056),
.B(n_1067),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1117),
.B(n_1043),
.Y(n_1375)
);

INVx2_ASAP7_75t_L g1376 ( 
.A(n_1105),
.Y(n_1376)
);

OAI21xp5_ASAP7_75t_L g1377 ( 
.A1(n_1211),
.A2(n_1176),
.B(n_1189),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1105),
.Y(n_1378)
);

AOI22xp33_ASAP7_75t_L g1379 ( 
.A1(n_1211),
.A2(n_1263),
.B1(n_1253),
.B2(n_1264),
.Y(n_1379)
);

NOR2xp33_ASAP7_75t_L g1380 ( 
.A(n_1043),
.B(n_1172),
.Y(n_1380)
);

OAI21x1_ASAP7_75t_SL g1381 ( 
.A1(n_1243),
.A2(n_1041),
.B(n_1167),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1189),
.B(n_1141),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1105),
.Y(n_1383)
);

AOI22xp33_ASAP7_75t_SL g1384 ( 
.A1(n_1238),
.A2(n_1253),
.B1(n_1236),
.B2(n_1062),
.Y(n_1384)
);

AOI21xp5_ASAP7_75t_L g1385 ( 
.A1(n_1047),
.A2(n_1234),
.B(n_1130),
.Y(n_1385)
);

AND2x2_ASAP7_75t_L g1386 ( 
.A(n_1264),
.B(n_1242),
.Y(n_1386)
);

OAI21x1_ASAP7_75t_SL g1387 ( 
.A1(n_1041),
.A2(n_1064),
.B(n_1167),
.Y(n_1387)
);

OAI222xp33_ASAP7_75t_L g1388 ( 
.A1(n_1109),
.A2(n_1264),
.B1(n_1164),
.B2(n_1160),
.C1(n_1108),
.C2(n_1115),
.Y(n_1388)
);

AO31x2_ASAP7_75t_L g1389 ( 
.A1(n_1100),
.A2(n_1181),
.A3(n_1153),
.B(n_1164),
.Y(n_1389)
);

BUFx3_ASAP7_75t_L g1390 ( 
.A(n_1163),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1105),
.Y(n_1391)
);

NAND2xp5_ASAP7_75t_L g1392 ( 
.A(n_1211),
.B(n_1049),
.Y(n_1392)
);

INVxp33_ASAP7_75t_L g1393 ( 
.A(n_1101),
.Y(n_1393)
);

OA21x2_ASAP7_75t_L g1394 ( 
.A1(n_1100),
.A2(n_1108),
.B(n_1160),
.Y(n_1394)
);

CKINVDCx11_ASAP7_75t_R g1395 ( 
.A(n_1060),
.Y(n_1395)
);

OAI21x1_ASAP7_75t_L g1396 ( 
.A1(n_1067),
.A2(n_1123),
.B(n_1169),
.Y(n_1396)
);

OAI21x1_ASAP7_75t_SL g1397 ( 
.A1(n_1064),
.A2(n_1169),
.B(n_1187),
.Y(n_1397)
);

OAI21x1_ASAP7_75t_L g1398 ( 
.A1(n_1123),
.A2(n_1187),
.B(n_1115),
.Y(n_1398)
);

AOI21xp5_ASAP7_75t_L g1399 ( 
.A1(n_1063),
.A2(n_1130),
.B(n_1203),
.Y(n_1399)
);

A2O1A1Ixp33_ASAP7_75t_L g1400 ( 
.A1(n_1085),
.A2(n_1078),
.B(n_1118),
.C(n_1127),
.Y(n_1400)
);

AOI21x1_ASAP7_75t_L g1401 ( 
.A1(n_1177),
.A2(n_1183),
.B(n_1125),
.Y(n_1401)
);

AOI21xp5_ASAP7_75t_L g1402 ( 
.A1(n_1063),
.A2(n_1203),
.B(n_1099),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1211),
.A2(n_1153),
.B(n_1181),
.Y(n_1403)
);

NAND3xp33_ASAP7_75t_SL g1404 ( 
.A(n_1109),
.B(n_1186),
.C(n_1191),
.Y(n_1404)
);

INVx4_ASAP7_75t_L g1405 ( 
.A(n_1063),
.Y(n_1405)
);

AOI21x1_ASAP7_75t_L g1406 ( 
.A1(n_1177),
.A2(n_1183),
.B(n_1155),
.Y(n_1406)
);

OAI21x1_ASAP7_75t_L g1407 ( 
.A1(n_1123),
.A2(n_1157),
.B(n_1155),
.Y(n_1407)
);

OAI22xp5_ASAP7_75t_L g1408 ( 
.A1(n_1253),
.A2(n_1085),
.B1(n_1101),
.B2(n_1062),
.Y(n_1408)
);

OAI21x1_ASAP7_75t_L g1409 ( 
.A1(n_1125),
.A2(n_1157),
.B(n_1136),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1133),
.A2(n_1138),
.B(n_1162),
.Y(n_1410)
);

O2A1O1Ixp33_ASAP7_75t_L g1411 ( 
.A1(n_1085),
.A2(n_1101),
.B(n_1070),
.C(n_1072),
.Y(n_1411)
);

AOI21x1_ASAP7_75t_L g1412 ( 
.A1(n_1179),
.A2(n_1049),
.B(n_1052),
.Y(n_1412)
);

OAI21x1_ASAP7_75t_L g1413 ( 
.A1(n_1133),
.A2(n_1162),
.B(n_1185),
.Y(n_1413)
);

OAI21x1_ASAP7_75t_L g1414 ( 
.A1(n_1133),
.A2(n_1162),
.B(n_1185),
.Y(n_1414)
);

AOI21xp5_ASAP7_75t_L g1415 ( 
.A1(n_1063),
.A2(n_1130),
.B(n_1203),
.Y(n_1415)
);

OAI21x1_ASAP7_75t_L g1416 ( 
.A1(n_1136),
.A2(n_1185),
.B(n_1138),
.Y(n_1416)
);

INVx2_ASAP7_75t_L g1417 ( 
.A(n_1105),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1136),
.A2(n_1138),
.B(n_1126),
.Y(n_1418)
);

AOI22xp33_ASAP7_75t_L g1419 ( 
.A1(n_1211),
.A2(n_1253),
.B1(n_1124),
.B2(n_1236),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1105),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1105),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1105),
.A2(n_1126),
.A3(n_1119),
.B(n_1211),
.Y(n_1422)
);

OAI21x1_ASAP7_75t_L g1423 ( 
.A1(n_1105),
.A2(n_1126),
.B(n_1092),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1126),
.Y(n_1424)
);

AND2x4_ASAP7_75t_L g1425 ( 
.A(n_1049),
.B(n_1052),
.Y(n_1425)
);

AO21x2_ASAP7_75t_L g1426 ( 
.A1(n_1126),
.A2(n_1058),
.B(n_1052),
.Y(n_1426)
);

OAI22xp33_ASAP7_75t_L g1427 ( 
.A1(n_1060),
.A2(n_1062),
.B1(n_1124),
.B2(n_1236),
.Y(n_1427)
);

BUFx12f_ASAP7_75t_L g1428 ( 
.A(n_1074),
.Y(n_1428)
);

AOI22x1_ASAP7_75t_L g1429 ( 
.A1(n_1186),
.A2(n_1255),
.B1(n_1233),
.B2(n_1232),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1126),
.A2(n_1092),
.B(n_1163),
.Y(n_1430)
);

INVx4_ASAP7_75t_SL g1431 ( 
.A(n_1045),
.Y(n_1431)
);

OA21x2_ASAP7_75t_L g1432 ( 
.A1(n_1126),
.A2(n_1058),
.B(n_1052),
.Y(n_1432)
);

BUFx2_ASAP7_75t_L g1433 ( 
.A(n_1126),
.Y(n_1433)
);

OAI21x1_ASAP7_75t_L g1434 ( 
.A1(n_1126),
.A2(n_1092),
.B(n_1193),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_1193),
.Y(n_1435)
);

OAI21x1_ASAP7_75t_L g1436 ( 
.A1(n_1092),
.A2(n_1193),
.B(n_1130),
.Y(n_1436)
);

OAI22xp33_ASAP7_75t_SL g1437 ( 
.A1(n_1118),
.A2(n_1127),
.B1(n_1150),
.B2(n_1196),
.Y(n_1437)
);

OR2x6_ASAP7_75t_L g1438 ( 
.A(n_1219),
.B(n_1222),
.Y(n_1438)
);

HB1xp67_ASAP7_75t_L g1439 ( 
.A(n_1225),
.Y(n_1439)
);

OAI21x1_ASAP7_75t_L g1440 ( 
.A1(n_1193),
.A2(n_1203),
.B(n_1130),
.Y(n_1440)
);

CKINVDCx8_ASAP7_75t_R g1441 ( 
.A(n_1102),
.Y(n_1441)
);

BUFx3_ASAP7_75t_L g1442 ( 
.A(n_1204),
.Y(n_1442)
);

NAND2xp5_ASAP7_75t_L g1443 ( 
.A(n_1049),
.B(n_1058),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1193),
.A2(n_1130),
.B(n_1203),
.Y(n_1444)
);

OA21x2_ASAP7_75t_L g1445 ( 
.A1(n_1058),
.A2(n_1149),
.B(n_1168),
.Y(n_1445)
);

OAI21x1_ASAP7_75t_L g1446 ( 
.A1(n_1193),
.A2(n_1099),
.B(n_1203),
.Y(n_1446)
);

OAI21x1_ASAP7_75t_L g1447 ( 
.A1(n_1193),
.A2(n_1099),
.B(n_1063),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1118),
.B(n_1127),
.Y(n_1448)
);

HB1xp67_ASAP7_75t_L g1449 ( 
.A(n_1225),
.Y(n_1449)
);

AO21x2_ASAP7_75t_L g1450 ( 
.A1(n_1255),
.A2(n_1193),
.B(n_1237),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1237),
.Y(n_1451)
);

OR2x2_ASAP7_75t_L g1452 ( 
.A(n_1351),
.B(n_1070),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1320),
.Y(n_1453)
);

INVx1_ASAP7_75t_L g1454 ( 
.A(n_1320),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1341),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1341),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1350),
.Y(n_1457)
);

INVx1_ASAP7_75t_L g1458 ( 
.A(n_1350),
.Y(n_1458)
);

NAND2xp5_ASAP7_75t_L g1459 ( 
.A(n_1333),
.B(n_1193),
.Y(n_1459)
);

INVx6_ASAP7_75t_SL g1460 ( 
.A(n_1438),
.Y(n_1460)
);

OAI22xp5_ASAP7_75t_L g1461 ( 
.A1(n_1337),
.A2(n_1072),
.B1(n_1137),
.B2(n_1061),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1346),
.B(n_1225),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1445),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1353),
.Y(n_1464)
);

OAI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1280),
.A2(n_1099),
.B(n_1237),
.Y(n_1465)
);

OAI21xp5_ASAP7_75t_L g1466 ( 
.A1(n_1270),
.A2(n_1144),
.B(n_1166),
.Y(n_1466)
);

INVx3_ASAP7_75t_L g1467 ( 
.A(n_1432),
.Y(n_1467)
);

INVx1_ASAP7_75t_SL g1468 ( 
.A(n_1297),
.Y(n_1468)
);

BUFx3_ASAP7_75t_L g1469 ( 
.A(n_1445),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1353),
.Y(n_1470)
);

HB1xp67_ASAP7_75t_L g1471 ( 
.A(n_1401),
.Y(n_1471)
);

INVx1_ASAP7_75t_L g1472 ( 
.A(n_1373),
.Y(n_1472)
);

INVx3_ASAP7_75t_L g1473 ( 
.A(n_1432),
.Y(n_1473)
);

OAI22xp5_ASAP7_75t_L g1474 ( 
.A1(n_1274),
.A2(n_1069),
.B1(n_1061),
.B2(n_1099),
.Y(n_1474)
);

INVxp67_ASAP7_75t_SL g1475 ( 
.A(n_1401),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1373),
.Y(n_1476)
);

INVx2_ASAP7_75t_L g1477 ( 
.A(n_1358),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1356),
.Y(n_1478)
);

BUFx3_ASAP7_75t_L g1479 ( 
.A(n_1445),
.Y(n_1479)
);

BUFx6f_ASAP7_75t_L g1480 ( 
.A(n_1423),
.Y(n_1480)
);

INVx2_ASAP7_75t_L g1481 ( 
.A(n_1358),
.Y(n_1481)
);

HB1xp67_ASAP7_75t_SL g1482 ( 
.A(n_1359),
.Y(n_1482)
);

HB1xp67_ASAP7_75t_L g1483 ( 
.A(n_1406),
.Y(n_1483)
);

AO21x1_ASAP7_75t_SL g1484 ( 
.A1(n_1344),
.A2(n_1158),
.B(n_1204),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1360),
.Y(n_1485)
);

INVx6_ASAP7_75t_L g1486 ( 
.A(n_1273),
.Y(n_1486)
);

BUFx3_ASAP7_75t_L g1487 ( 
.A(n_1445),
.Y(n_1487)
);

OAI21x1_ASAP7_75t_L g1488 ( 
.A1(n_1267),
.A2(n_1237),
.B(n_1204),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1406),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1356),
.Y(n_1490)
);

OAI21x1_ASAP7_75t_L g1491 ( 
.A1(n_1267),
.A2(n_1237),
.B(n_1204),
.Y(n_1491)
);

OAI22xp5_ASAP7_75t_L g1492 ( 
.A1(n_1278),
.A2(n_1061),
.B1(n_1069),
.B2(n_1144),
.Y(n_1492)
);

INVx1_ASAP7_75t_L g1493 ( 
.A(n_1356),
.Y(n_1493)
);

HB1xp67_ASAP7_75t_L g1494 ( 
.A(n_1354),
.Y(n_1494)
);

BUFx12f_ASAP7_75t_L g1495 ( 
.A(n_1395),
.Y(n_1495)
);

AOI221xp5_ASAP7_75t_L g1496 ( 
.A1(n_1268),
.A2(n_1106),
.B1(n_1231),
.B2(n_1044),
.C(n_1086),
.Y(n_1496)
);

CKINVDCx20_ASAP7_75t_R g1497 ( 
.A(n_1275),
.Y(n_1497)
);

AND2x2_ASAP7_75t_L g1498 ( 
.A(n_1346),
.B(n_1231),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1356),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1432),
.Y(n_1500)
);

OAI21x1_ASAP7_75t_L g1501 ( 
.A1(n_1287),
.A2(n_1237),
.B(n_1214),
.Y(n_1501)
);

INVx2_ASAP7_75t_L g1502 ( 
.A(n_1398),
.Y(n_1502)
);

BUFx2_ASAP7_75t_L g1503 ( 
.A(n_1432),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1266),
.B(n_1231),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1266),
.Y(n_1505)
);

AO21x2_ASAP7_75t_L g1506 ( 
.A1(n_1269),
.A2(n_1214),
.B(n_1112),
.Y(n_1506)
);

INVx2_ASAP7_75t_L g1507 ( 
.A(n_1398),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_1286),
.Y(n_1508)
);

OAI22xp5_ASAP7_75t_L g1509 ( 
.A1(n_1289),
.A2(n_1069),
.B1(n_1061),
.B2(n_1128),
.Y(n_1509)
);

INVx2_ASAP7_75t_SL g1510 ( 
.A(n_1369),
.Y(n_1510)
);

OAI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1423),
.A2(n_1140),
.B(n_1122),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1286),
.B(n_1188),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1291),
.Y(n_1513)
);

INVx2_ASAP7_75t_L g1514 ( 
.A(n_1291),
.Y(n_1514)
);

AO21x2_ASAP7_75t_L g1515 ( 
.A1(n_1327),
.A2(n_1112),
.B(n_1122),
.Y(n_1515)
);

AND2x4_ASAP7_75t_L g1516 ( 
.A(n_1422),
.B(n_1119),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1294),
.Y(n_1517)
);

OAI21x1_ASAP7_75t_L g1518 ( 
.A1(n_1292),
.A2(n_1140),
.B(n_1102),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1336),
.B(n_1170),
.Y(n_1519)
);

BUFx3_ASAP7_75t_L g1520 ( 
.A(n_1340),
.Y(n_1520)
);

HB1xp67_ASAP7_75t_L g1521 ( 
.A(n_1354),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1336),
.B(n_1170),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1282),
.Y(n_1523)
);

INVx1_ASAP7_75t_L g1524 ( 
.A(n_1294),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1332),
.A2(n_1077),
.B1(n_1069),
.B2(n_1206),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1299),
.Y(n_1526)
);

AOI22xp33_ASAP7_75t_L g1527 ( 
.A1(n_1335),
.A2(n_1077),
.B1(n_1196),
.B2(n_1150),
.Y(n_1527)
);

OAI21x1_ASAP7_75t_L g1528 ( 
.A1(n_1352),
.A2(n_1119),
.B(n_1219),
.Y(n_1528)
);

CKINVDCx20_ASAP7_75t_R g1529 ( 
.A(n_1312),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1323),
.B(n_1364),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1394),
.Y(n_1531)
);

INVx1_ASAP7_75t_L g1532 ( 
.A(n_1299),
.Y(n_1532)
);

INVx2_ASAP7_75t_L g1533 ( 
.A(n_1394),
.Y(n_1533)
);

OAI22xp5_ASAP7_75t_L g1534 ( 
.A1(n_1289),
.A2(n_1135),
.B1(n_1128),
.B2(n_1150),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1301),
.Y(n_1535)
);

BUFx2_ASAP7_75t_L g1536 ( 
.A(n_1361),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1394),
.Y(n_1537)
);

INVx2_ASAP7_75t_SL g1538 ( 
.A(n_1369),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1422),
.B(n_1190),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1394),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1301),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1396),
.Y(n_1542)
);

INVx2_ASAP7_75t_L g1543 ( 
.A(n_1396),
.Y(n_1543)
);

AND2x2_ASAP7_75t_L g1544 ( 
.A(n_1422),
.B(n_1190),
.Y(n_1544)
);

INVx2_ASAP7_75t_SL g1545 ( 
.A(n_1369),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1272),
.B(n_1156),
.Y(n_1546)
);

INVx1_ASAP7_75t_L g1547 ( 
.A(n_1313),
.Y(n_1547)
);

HB1xp67_ASAP7_75t_L g1548 ( 
.A(n_1354),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_1313),
.Y(n_1549)
);

AOI22xp33_ASAP7_75t_L g1550 ( 
.A1(n_1335),
.A2(n_1150),
.B1(n_1196),
.B2(n_1106),
.Y(n_1550)
);

HB1xp67_ASAP7_75t_L g1551 ( 
.A(n_1369),
.Y(n_1551)
);

AOI22xp33_ASAP7_75t_L g1552 ( 
.A1(n_1324),
.A2(n_1196),
.B1(n_1232),
.B2(n_1233),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1315),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1315),
.Y(n_1554)
);

OA21x2_ASAP7_75t_L g1555 ( 
.A1(n_1285),
.A2(n_1149),
.B(n_1044),
.Y(n_1555)
);

INVx1_ASAP7_75t_L g1556 ( 
.A(n_1365),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1365),
.Y(n_1557)
);

OAI21x1_ASAP7_75t_L g1558 ( 
.A1(n_1352),
.A2(n_1366),
.B(n_1345),
.Y(n_1558)
);

INVx1_ASAP7_75t_L g1559 ( 
.A(n_1300),
.Y(n_1559)
);

INVx1_ASAP7_75t_L g1560 ( 
.A(n_1300),
.Y(n_1560)
);

HB1xp67_ASAP7_75t_L g1561 ( 
.A(n_1412),
.Y(n_1561)
);

AOI21x1_ASAP7_75t_L g1562 ( 
.A1(n_1293),
.A2(n_1086),
.B(n_1222),
.Y(n_1562)
);

AOI22xp33_ASAP7_75t_L g1563 ( 
.A1(n_1324),
.A2(n_1342),
.B1(n_1329),
.B2(n_1425),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1304),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1422),
.B(n_1200),
.Y(n_1565)
);

BUFx2_ASAP7_75t_L g1566 ( 
.A(n_1361),
.Y(n_1566)
);

NAND2x1p5_ASAP7_75t_L g1567 ( 
.A(n_1433),
.B(n_1119),
.Y(n_1567)
);

HB1xp67_ASAP7_75t_L g1568 ( 
.A(n_1412),
.Y(n_1568)
);

AOI22xp33_ASAP7_75t_L g1569 ( 
.A1(n_1328),
.A2(n_1233),
.B1(n_1232),
.B2(n_1200),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1422),
.B(n_1200),
.Y(n_1570)
);

OAI22xp5_ASAP7_75t_L g1571 ( 
.A1(n_1321),
.A2(n_1135),
.B1(n_1128),
.B2(n_1096),
.Y(n_1571)
);

AOI22xp33_ASAP7_75t_L g1572 ( 
.A1(n_1285),
.A2(n_1348),
.B1(n_1318),
.B2(n_1303),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1331),
.B(n_1198),
.Y(n_1573)
);

BUFx2_ASAP7_75t_L g1574 ( 
.A(n_1361),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1308),
.Y(n_1575)
);

BUFx3_ASAP7_75t_L g1576 ( 
.A(n_1340),
.Y(n_1576)
);

INVx1_ASAP7_75t_L g1577 ( 
.A(n_1308),
.Y(n_1577)
);

AOI22xp33_ASAP7_75t_L g1578 ( 
.A1(n_1310),
.A2(n_1233),
.B1(n_1232),
.B2(n_1198),
.Y(n_1578)
);

INVx1_ASAP7_75t_L g1579 ( 
.A(n_1316),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1331),
.B(n_1351),
.Y(n_1580)
);

BUFx2_ASAP7_75t_SL g1581 ( 
.A(n_1441),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1316),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1330),
.Y(n_1583)
);

INVx1_ASAP7_75t_L g1584 ( 
.A(n_1330),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1343),
.B(n_1198),
.Y(n_1585)
);

OAI21x1_ASAP7_75t_L g1586 ( 
.A1(n_1366),
.A2(n_1116),
.B(n_1059),
.Y(n_1586)
);

INVx3_ASAP7_75t_L g1587 ( 
.A(n_1426),
.Y(n_1587)
);

INVx1_ASAP7_75t_L g1588 ( 
.A(n_1339),
.Y(n_1588)
);

INVx1_ASAP7_75t_L g1589 ( 
.A(n_1347),
.Y(n_1589)
);

OR2x2_ASAP7_75t_L g1590 ( 
.A(n_1326),
.B(n_1197),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1347),
.Y(n_1591)
);

BUFx2_ASAP7_75t_L g1592 ( 
.A(n_1426),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1349),
.Y(n_1593)
);

AND2x4_ASAP7_75t_L g1594 ( 
.A(n_1426),
.B(n_1197),
.Y(n_1594)
);

OAI21x1_ASAP7_75t_L g1595 ( 
.A1(n_1345),
.A2(n_1116),
.B(n_1059),
.Y(n_1595)
);

INVx1_ASAP7_75t_L g1596 ( 
.A(n_1349),
.Y(n_1596)
);

CKINVDCx6p67_ASAP7_75t_R g1597 ( 
.A(n_1276),
.Y(n_1597)
);

AND2x4_ASAP7_75t_L g1598 ( 
.A(n_1434),
.B(n_1197),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1389),
.Y(n_1599)
);

INVx1_ASAP7_75t_L g1600 ( 
.A(n_1389),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1389),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1389),
.Y(n_1602)
);

AO21x1_ASAP7_75t_SL g1603 ( 
.A1(n_1343),
.A2(n_1152),
.B(n_1120),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1272),
.B(n_1217),
.Y(n_1604)
);

INVx2_ASAP7_75t_L g1605 ( 
.A(n_1389),
.Y(n_1605)
);

INVx1_ASAP7_75t_L g1606 ( 
.A(n_1407),
.Y(n_1606)
);

INVx2_ASAP7_75t_L g1607 ( 
.A(n_1407),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1293),
.A2(n_1184),
.B(n_1171),
.Y(n_1608)
);

OR2x2_ASAP7_75t_L g1609 ( 
.A(n_1326),
.B(n_1190),
.Y(n_1609)
);

AND2x2_ASAP7_75t_L g1610 ( 
.A(n_1325),
.B(n_1178),
.Y(n_1610)
);

BUFx6f_ASAP7_75t_L g1611 ( 
.A(n_1434),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1418),
.Y(n_1612)
);

INVx3_ASAP7_75t_L g1613 ( 
.A(n_1418),
.Y(n_1613)
);

INVx3_ASAP7_75t_L g1614 ( 
.A(n_1372),
.Y(n_1614)
);

AOI22xp33_ASAP7_75t_L g1615 ( 
.A1(n_1342),
.A2(n_1145),
.B1(n_1178),
.B2(n_1159),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1325),
.B(n_1178),
.Y(n_1616)
);

HB1xp67_ASAP7_75t_L g1617 ( 
.A(n_1311),
.Y(n_1617)
);

INVx2_ASAP7_75t_L g1618 ( 
.A(n_1409),
.Y(n_1618)
);

AOI22xp33_ASAP7_75t_SL g1619 ( 
.A1(n_1355),
.A2(n_1184),
.B1(n_1171),
.B2(n_1116),
.Y(n_1619)
);

HB1xp67_ASAP7_75t_L g1620 ( 
.A(n_1311),
.Y(n_1620)
);

INVx2_ASAP7_75t_L g1621 ( 
.A(n_1409),
.Y(n_1621)
);

BUFx12f_ASAP7_75t_L g1622 ( 
.A(n_1312),
.Y(n_1622)
);

CKINVDCx6p67_ASAP7_75t_R g1623 ( 
.A(n_1428),
.Y(n_1623)
);

AOI22xp33_ASAP7_75t_L g1624 ( 
.A1(n_1425),
.A2(n_1145),
.B1(n_1151),
.B2(n_1170),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1383),
.Y(n_1625)
);

AOI21xp5_ASAP7_75t_L g1626 ( 
.A1(n_1506),
.A2(n_1385),
.B(n_1296),
.Y(n_1626)
);

OAI222xp33_ASAP7_75t_L g1627 ( 
.A1(n_1572),
.A2(n_1363),
.B1(n_1338),
.B2(n_1384),
.C1(n_1379),
.C2(n_1408),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1462),
.B(n_1386),
.Y(n_1628)
);

BUFx3_ASAP7_75t_L g1629 ( 
.A(n_1495),
.Y(n_1629)
);

HB1xp67_ASAP7_75t_L g1630 ( 
.A(n_1617),
.Y(n_1630)
);

A2O1A1Ixp33_ASAP7_75t_L g1631 ( 
.A1(n_1534),
.A2(n_1363),
.B(n_1403),
.C(n_1400),
.Y(n_1631)
);

AND3x1_ASAP7_75t_L g1632 ( 
.A(n_1525),
.B(n_1380),
.C(n_1375),
.Y(n_1632)
);

AOI22xp33_ASAP7_75t_L g1633 ( 
.A1(n_1572),
.A2(n_1534),
.B1(n_1509),
.B2(n_1461),
.Y(n_1633)
);

AOI22xp33_ASAP7_75t_L g1634 ( 
.A1(n_1509),
.A2(n_1310),
.B1(n_1309),
.B2(n_1325),
.Y(n_1634)
);

AOI21xp33_ASAP7_75t_L g1635 ( 
.A1(n_1563),
.A2(n_1271),
.B(n_1355),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1526),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_R g1637 ( 
.A(n_1503),
.B(n_1438),
.Y(n_1637)
);

CKINVDCx5p33_ASAP7_75t_R g1638 ( 
.A(n_1497),
.Y(n_1638)
);

NAND2xp33_ASAP7_75t_R g1639 ( 
.A(n_1503),
.B(n_1555),
.Y(n_1639)
);

INVx3_ASAP7_75t_L g1640 ( 
.A(n_1463),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_R g1641 ( 
.A(n_1482),
.B(n_1404),
.Y(n_1641)
);

OAI22xp5_ASAP7_75t_SL g1642 ( 
.A1(n_1495),
.A2(n_1428),
.B1(n_1290),
.B2(n_1419),
.Y(n_1642)
);

NAND2xp5_ASAP7_75t_L g1643 ( 
.A(n_1530),
.B(n_1297),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1452),
.B(n_1392),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1462),
.B(n_1386),
.Y(n_1645)
);

HB1xp67_ASAP7_75t_L g1646 ( 
.A(n_1617),
.Y(n_1646)
);

OAI21xp33_ASAP7_75t_L g1647 ( 
.A1(n_1578),
.A2(n_1377),
.B(n_1367),
.Y(n_1647)
);

OR2x2_ASAP7_75t_L g1648 ( 
.A(n_1452),
.B(n_1377),
.Y(n_1648)
);

INVx4_ASAP7_75t_L g1649 ( 
.A(n_1486),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1462),
.B(n_1425),
.Y(n_1650)
);

HB1xp67_ASAP7_75t_L g1651 ( 
.A(n_1620),
.Y(n_1651)
);

BUFx6f_ASAP7_75t_L g1652 ( 
.A(n_1603),
.Y(n_1652)
);

CKINVDCx5p33_ASAP7_75t_R g1653 ( 
.A(n_1523),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_L g1654 ( 
.A(n_1530),
.B(n_1370),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1580),
.B(n_1311),
.Y(n_1655)
);

NAND2xp33_ASAP7_75t_R g1656 ( 
.A(n_1555),
.B(n_1438),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1459),
.B(n_1370),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1498),
.B(n_1425),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_SL g1659 ( 
.A(n_1461),
.B(n_1427),
.C(n_1368),
.Y(n_1659)
);

INVxp33_ASAP7_75t_SL g1660 ( 
.A(n_1581),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_R g1661 ( 
.A(n_1482),
.B(n_1441),
.Y(n_1661)
);

OR2x2_ASAP7_75t_L g1662 ( 
.A(n_1580),
.B(n_1325),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1498),
.B(n_1325),
.Y(n_1663)
);

NOR3xp33_ASAP7_75t_SL g1664 ( 
.A(n_1466),
.B(n_1411),
.C(n_1388),
.Y(n_1664)
);

NAND2xp33_ASAP7_75t_R g1665 ( 
.A(n_1555),
.B(n_1438),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1580),
.B(n_1314),
.Y(n_1666)
);

AOI21xp5_ASAP7_75t_SL g1667 ( 
.A1(n_1492),
.A2(n_1271),
.B(n_1438),
.Y(n_1667)
);

CKINVDCx5p33_ASAP7_75t_R g1668 ( 
.A(n_1495),
.Y(n_1668)
);

HB1xp67_ASAP7_75t_L g1669 ( 
.A(n_1620),
.Y(n_1669)
);

OAI21x1_ASAP7_75t_L g1670 ( 
.A1(n_1488),
.A2(n_1430),
.B(n_1446),
.Y(n_1670)
);

BUFx10_ASAP7_75t_L g1671 ( 
.A(n_1486),
.Y(n_1671)
);

AO31x2_ASAP7_75t_L g1672 ( 
.A1(n_1601),
.A2(n_1322),
.A3(n_1605),
.B(n_1602),
.Y(n_1672)
);

AND2x2_ASAP7_75t_L g1673 ( 
.A(n_1498),
.B(n_1519),
.Y(n_1673)
);

AND2x2_ASAP7_75t_L g1674 ( 
.A(n_1519),
.B(n_1298),
.Y(n_1674)
);

BUFx12f_ASAP7_75t_L g1675 ( 
.A(n_1622),
.Y(n_1675)
);

INVx2_ASAP7_75t_L g1676 ( 
.A(n_1531),
.Y(n_1676)
);

AOI22xp33_ASAP7_75t_SL g1677 ( 
.A1(n_1492),
.A2(n_1322),
.B1(n_1290),
.B2(n_1273),
.Y(n_1677)
);

AO32x2_ASAP7_75t_L g1678 ( 
.A1(n_1510),
.A2(n_1298),
.A3(n_1362),
.B1(n_1405),
.B2(n_1403),
.Y(n_1678)
);

AND2x4_ASAP7_75t_SL g1679 ( 
.A(n_1597),
.B(n_1371),
.Y(n_1679)
);

OR2x2_ASAP7_75t_L g1680 ( 
.A(n_1459),
.B(n_1314),
.Y(n_1680)
);

INVx2_ASAP7_75t_L g1681 ( 
.A(n_1531),
.Y(n_1681)
);

NAND2xp33_ASAP7_75t_R g1682 ( 
.A(n_1555),
.B(n_1592),
.Y(n_1682)
);

INVx1_ASAP7_75t_L g1683 ( 
.A(n_1526),
.Y(n_1683)
);

AND2x2_ASAP7_75t_L g1684 ( 
.A(n_1519),
.B(n_1362),
.Y(n_1684)
);

NAND2x1p5_ASAP7_75t_L g1685 ( 
.A(n_1518),
.B(n_1430),
.Y(n_1685)
);

OR2x6_ASAP7_75t_L g1686 ( 
.A(n_1581),
.B(n_1486),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1532),
.Y(n_1687)
);

NOR2xp33_ASAP7_75t_R g1688 ( 
.A(n_1529),
.B(n_1597),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_R g1689 ( 
.A(n_1597),
.B(n_1371),
.Y(n_1689)
);

BUFx10_ASAP7_75t_L g1690 ( 
.A(n_1486),
.Y(n_1690)
);

NOR2xp33_ASAP7_75t_R g1691 ( 
.A(n_1622),
.B(n_1371),
.Y(n_1691)
);

NAND2xp33_ASAP7_75t_R g1692 ( 
.A(n_1555),
.B(n_1433),
.Y(n_1692)
);

CKINVDCx5p33_ASAP7_75t_R g1693 ( 
.A(n_1622),
.Y(n_1693)
);

AND2x2_ASAP7_75t_L g1694 ( 
.A(n_1522),
.B(n_1573),
.Y(n_1694)
);

NAND2xp5_ASAP7_75t_L g1695 ( 
.A(n_1468),
.B(n_1382),
.Y(n_1695)
);

INVx2_ASAP7_75t_L g1696 ( 
.A(n_1531),
.Y(n_1696)
);

NOR2xp33_ASAP7_75t_R g1697 ( 
.A(n_1623),
.B(n_1273),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1468),
.B(n_1283),
.Y(n_1698)
);

OR2x6_ASAP7_75t_L g1699 ( 
.A(n_1486),
.B(n_1436),
.Y(n_1699)
);

INVx2_ASAP7_75t_L g1700 ( 
.A(n_1533),
.Y(n_1700)
);

AND2x2_ASAP7_75t_L g1701 ( 
.A(n_1522),
.B(n_1393),
.Y(n_1701)
);

NOR3xp33_ASAP7_75t_SL g1702 ( 
.A(n_1466),
.B(n_1448),
.C(n_1319),
.Y(n_1702)
);

CKINVDCx16_ASAP7_75t_R g1703 ( 
.A(n_1522),
.Y(n_1703)
);

NAND2xp5_ASAP7_75t_L g1704 ( 
.A(n_1504),
.B(n_1573),
.Y(n_1704)
);

CKINVDCx16_ASAP7_75t_R g1705 ( 
.A(n_1520),
.Y(n_1705)
);

CKINVDCx20_ASAP7_75t_R g1706 ( 
.A(n_1623),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1504),
.B(n_1573),
.Y(n_1707)
);

HB1xp67_ASAP7_75t_L g1708 ( 
.A(n_1590),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1590),
.B(n_1283),
.Y(n_1709)
);

BUFx3_ASAP7_75t_L g1710 ( 
.A(n_1623),
.Y(n_1710)
);

BUFx3_ASAP7_75t_L g1711 ( 
.A(n_1520),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1533),
.Y(n_1712)
);

OAI21xp5_ASAP7_75t_L g1713 ( 
.A1(n_1527),
.A2(n_1288),
.B(n_1357),
.Y(n_1713)
);

AND2x2_ASAP7_75t_L g1714 ( 
.A(n_1585),
.B(n_1435),
.Y(n_1714)
);

INVx2_ASAP7_75t_L g1715 ( 
.A(n_1533),
.Y(n_1715)
);

NAND2xp5_ASAP7_75t_L g1716 ( 
.A(n_1609),
.B(n_1284),
.Y(n_1716)
);

AND2x4_ASAP7_75t_SL g1717 ( 
.A(n_1594),
.B(n_1439),
.Y(n_1717)
);

BUFx2_ASAP7_75t_L g1718 ( 
.A(n_1460),
.Y(n_1718)
);

INVx1_ASAP7_75t_L g1719 ( 
.A(n_1532),
.Y(n_1719)
);

BUFx3_ASAP7_75t_L g1720 ( 
.A(n_1520),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1535),
.Y(n_1721)
);

CKINVDCx16_ASAP7_75t_R g1722 ( 
.A(n_1576),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1460),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1609),
.B(n_1284),
.Y(n_1724)
);

NOR2xp33_ASAP7_75t_R g1725 ( 
.A(n_1608),
.B(n_1273),
.Y(n_1725)
);

OA21x2_ASAP7_75t_L g1726 ( 
.A1(n_1478),
.A2(n_1383),
.B(n_1391),
.Y(n_1726)
);

INVx2_ASAP7_75t_L g1727 ( 
.A(n_1537),
.Y(n_1727)
);

AO31x2_ASAP7_75t_L g1728 ( 
.A1(n_1601),
.A2(n_1421),
.A3(n_1391),
.B(n_1378),
.Y(n_1728)
);

OAI22xp5_ASAP7_75t_L g1729 ( 
.A1(n_1552),
.A2(n_1550),
.B1(n_1569),
.B2(n_1619),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1594),
.B(n_1435),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1594),
.B(n_1421),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1546),
.B(n_1295),
.Y(n_1732)
);

INVx2_ASAP7_75t_L g1733 ( 
.A(n_1537),
.Y(n_1733)
);

AO31x2_ASAP7_75t_L g1734 ( 
.A1(n_1601),
.A2(n_1376),
.A3(n_1378),
.B(n_1417),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1585),
.B(n_1443),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_R g1736 ( 
.A(n_1608),
.B(n_1340),
.Y(n_1736)
);

BUFx3_ASAP7_75t_L g1737 ( 
.A(n_1576),
.Y(n_1737)
);

AND2x2_ASAP7_75t_L g1738 ( 
.A(n_1585),
.B(n_1277),
.Y(n_1738)
);

NOR2xp33_ASAP7_75t_R g1739 ( 
.A(n_1576),
.B(n_1390),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1546),
.B(n_1295),
.Y(n_1740)
);

INVx2_ASAP7_75t_L g1741 ( 
.A(n_1537),
.Y(n_1741)
);

BUFx6f_ASAP7_75t_SL g1742 ( 
.A(n_1598),
.Y(n_1742)
);

AND2x4_ASAP7_75t_L g1743 ( 
.A(n_1594),
.B(n_1376),
.Y(n_1743)
);

HB1xp67_ASAP7_75t_L g1744 ( 
.A(n_1539),
.Y(n_1744)
);

INVx2_ASAP7_75t_L g1745 ( 
.A(n_1540),
.Y(n_1745)
);

NAND2xp33_ASAP7_75t_R g1746 ( 
.A(n_1592),
.B(n_1399),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1604),
.B(n_1512),
.Y(n_1747)
);

NOR3xp33_ASAP7_75t_SL g1748 ( 
.A(n_1496),
.B(n_1451),
.C(n_1415),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1540),
.Y(n_1749)
);

INVx2_ASAP7_75t_L g1750 ( 
.A(n_1540),
.Y(n_1750)
);

CKINVDCx16_ASAP7_75t_R g1751 ( 
.A(n_1610),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1604),
.B(n_1512),
.Y(n_1752)
);

INVx1_ASAP7_75t_L g1753 ( 
.A(n_1535),
.Y(n_1753)
);

BUFx12f_ASAP7_75t_L g1754 ( 
.A(n_1598),
.Y(n_1754)
);

AND2x2_ASAP7_75t_L g1755 ( 
.A(n_1610),
.B(n_1277),
.Y(n_1755)
);

NAND2xp5_ASAP7_75t_L g1756 ( 
.A(n_1559),
.B(n_1295),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1541),
.Y(n_1757)
);

CKINVDCx16_ASAP7_75t_R g1758 ( 
.A(n_1610),
.Y(n_1758)
);

INVx1_ASAP7_75t_L g1759 ( 
.A(n_1541),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_R g1760 ( 
.A(n_1536),
.B(n_1566),
.Y(n_1760)
);

OR2x2_ASAP7_75t_L g1761 ( 
.A(n_1625),
.B(n_1265),
.Y(n_1761)
);

NOR2xp33_ASAP7_75t_R g1762 ( 
.A(n_1562),
.B(n_1390),
.Y(n_1762)
);

HB1xp67_ASAP7_75t_L g1763 ( 
.A(n_1539),
.Y(n_1763)
);

INVx2_ASAP7_75t_L g1764 ( 
.A(n_1625),
.Y(n_1764)
);

AND2x4_ASAP7_75t_L g1765 ( 
.A(n_1594),
.B(n_1390),
.Y(n_1765)
);

NOR2xp33_ASAP7_75t_R g1766 ( 
.A(n_1562),
.B(n_1442),
.Y(n_1766)
);

OAI22xp33_ASAP7_75t_L g1767 ( 
.A1(n_1571),
.A2(n_1442),
.B1(n_1309),
.B2(n_1429),
.Y(n_1767)
);

HB1xp67_ASAP7_75t_L g1768 ( 
.A(n_1539),
.Y(n_1768)
);

NAND3xp33_ASAP7_75t_SL g1769 ( 
.A(n_1496),
.B(n_1302),
.C(n_1307),
.Y(n_1769)
);

INVx1_ASAP7_75t_L g1770 ( 
.A(n_1547),
.Y(n_1770)
);

CKINVDCx20_ASAP7_75t_R g1771 ( 
.A(n_1603),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1559),
.B(n_1295),
.Y(n_1772)
);

NAND2xp5_ASAP7_75t_L g1773 ( 
.A(n_1560),
.B(n_1334),
.Y(n_1773)
);

INVx3_ASAP7_75t_L g1774 ( 
.A(n_1463),
.Y(n_1774)
);

NAND2xp33_ASAP7_75t_R g1775 ( 
.A(n_1536),
.B(n_1402),
.Y(n_1775)
);

NAND2xp33_ASAP7_75t_SL g1776 ( 
.A(n_1569),
.B(n_1096),
.Y(n_1776)
);

BUFx3_ASAP7_75t_L g1777 ( 
.A(n_1567),
.Y(n_1777)
);

NOR2xp33_ASAP7_75t_R g1778 ( 
.A(n_1552),
.B(n_1442),
.Y(n_1778)
);

INVx1_ASAP7_75t_SL g1779 ( 
.A(n_1616),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1547),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1549),
.Y(n_1781)
);

NAND3xp33_ASAP7_75t_L g1782 ( 
.A(n_1578),
.B(n_1317),
.C(n_1449),
.Y(n_1782)
);

INVx1_ASAP7_75t_L g1783 ( 
.A(n_1549),
.Y(n_1783)
);

INVx5_ASAP7_75t_SL g1784 ( 
.A(n_1515),
.Y(n_1784)
);

INVx2_ASAP7_75t_L g1785 ( 
.A(n_1625),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_L g1786 ( 
.A(n_1560),
.B(n_1334),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1553),
.Y(n_1787)
);

INVx2_ASAP7_75t_L g1788 ( 
.A(n_1467),
.Y(n_1788)
);

INVx1_ASAP7_75t_L g1789 ( 
.A(n_1553),
.Y(n_1789)
);

AOI22xp33_ASAP7_75t_SL g1790 ( 
.A1(n_1474),
.A2(n_1334),
.B1(n_1437),
.B2(n_1429),
.Y(n_1790)
);

BUFx3_ASAP7_75t_L g1791 ( 
.A(n_1567),
.Y(n_1791)
);

AND2x4_ASAP7_75t_SL g1792 ( 
.A(n_1598),
.B(n_1405),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1554),
.Y(n_1793)
);

OAI22xp5_ASAP7_75t_L g1794 ( 
.A1(n_1619),
.A2(n_1405),
.B1(n_1451),
.B2(n_1135),
.Y(n_1794)
);

BUFx10_ASAP7_75t_L g1795 ( 
.A(n_1598),
.Y(n_1795)
);

AND2x2_ASAP7_75t_L g1796 ( 
.A(n_1616),
.B(n_1372),
.Y(n_1796)
);

AND2x2_ASAP7_75t_L g1797 ( 
.A(n_1616),
.B(n_1436),
.Y(n_1797)
);

NOR2xp33_ASAP7_75t_R g1798 ( 
.A(n_1624),
.B(n_1096),
.Y(n_1798)
);

CKINVDCx5p33_ASAP7_75t_R g1799 ( 
.A(n_1598),
.Y(n_1799)
);

NAND2xp33_ASAP7_75t_R g1800 ( 
.A(n_1566),
.B(n_1447),
.Y(n_1800)
);

HB1xp67_ASAP7_75t_L g1801 ( 
.A(n_1544),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_L g1802 ( 
.A(n_1564),
.B(n_1334),
.Y(n_1802)
);

OR2x6_ASAP7_75t_L g1803 ( 
.A(n_1574),
.B(n_1447),
.Y(n_1803)
);

AND2x2_ASAP7_75t_L g1804 ( 
.A(n_1544),
.B(n_1450),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1564),
.B(n_1334),
.Y(n_1805)
);

HB1xp67_ASAP7_75t_L g1806 ( 
.A(n_1544),
.Y(n_1806)
);

NOR2xp33_ASAP7_75t_R g1807 ( 
.A(n_1574),
.B(n_1116),
.Y(n_1807)
);

O2A1O1Ixp5_ASAP7_75t_L g1808 ( 
.A1(n_1571),
.A2(n_1420),
.B(n_1424),
.C(n_1405),
.Y(n_1808)
);

NAND2xp33_ASAP7_75t_R g1809 ( 
.A(n_1467),
.B(n_1446),
.Y(n_1809)
);

INVx2_ASAP7_75t_L g1810 ( 
.A(n_1467),
.Y(n_1810)
);

AOI22xp33_ASAP7_75t_L g1811 ( 
.A1(n_1474),
.A2(n_1334),
.B1(n_1305),
.B2(n_1265),
.Y(n_1811)
);

NAND2xp33_ASAP7_75t_R g1812 ( 
.A(n_1467),
.B(n_1473),
.Y(n_1812)
);

INVx5_ASAP7_75t_L g1813 ( 
.A(n_1473),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1554),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1565),
.Y(n_1815)
);

NAND2xp33_ASAP7_75t_R g1816 ( 
.A(n_1473),
.B(n_1444),
.Y(n_1816)
);

BUFx12f_ASAP7_75t_L g1817 ( 
.A(n_1567),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1453),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1565),
.Y(n_1819)
);

INVx2_ASAP7_75t_L g1820 ( 
.A(n_1473),
.Y(n_1820)
);

AND2x2_ASAP7_75t_L g1821 ( 
.A(n_1565),
.B(n_1450),
.Y(n_1821)
);

AND2x2_ASAP7_75t_L g1822 ( 
.A(n_1570),
.B(n_1450),
.Y(n_1822)
);

AOI22xp33_ASAP7_75t_L g1823 ( 
.A1(n_1484),
.A2(n_1334),
.B1(n_1305),
.B2(n_1306),
.Y(n_1823)
);

AND2x2_ASAP7_75t_L g1824 ( 
.A(n_1570),
.B(n_1374),
.Y(n_1824)
);

NAND2xp5_ASAP7_75t_SL g1825 ( 
.A(n_1556),
.B(n_1437),
.Y(n_1825)
);

INVx2_ASAP7_75t_SL g1826 ( 
.A(n_1570),
.Y(n_1826)
);

OR2x6_ASAP7_75t_L g1827 ( 
.A(n_1488),
.B(n_1444),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1575),
.B(n_1281),
.Y(n_1828)
);

INVx2_ASAP7_75t_L g1829 ( 
.A(n_1500),
.Y(n_1829)
);

INVx2_ASAP7_75t_L g1830 ( 
.A(n_1500),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1453),
.Y(n_1831)
);

NAND2xp5_ASAP7_75t_L g1832 ( 
.A(n_1575),
.B(n_1281),
.Y(n_1832)
);

CKINVDCx20_ASAP7_75t_R g1833 ( 
.A(n_1484),
.Y(n_1833)
);

INVx2_ASAP7_75t_L g1834 ( 
.A(n_1500),
.Y(n_1834)
);

AND2x2_ASAP7_75t_L g1835 ( 
.A(n_1477),
.B(n_1374),
.Y(n_1835)
);

CKINVDCx5p33_ASAP7_75t_R g1836 ( 
.A(n_1460),
.Y(n_1836)
);

OR2x6_ASAP7_75t_L g1837 ( 
.A(n_1488),
.B(n_1440),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1454),
.Y(n_1838)
);

AOI22xp33_ASAP7_75t_L g1839 ( 
.A1(n_1506),
.A2(n_1306),
.B1(n_1279),
.B2(n_1381),
.Y(n_1839)
);

AND2x4_ASAP7_75t_SL g1840 ( 
.A(n_1516),
.B(n_1615),
.Y(n_1840)
);

AOI22xp33_ASAP7_75t_SL g1841 ( 
.A1(n_1506),
.A2(n_1440),
.B1(n_1381),
.B2(n_1279),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1500),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1454),
.Y(n_1843)
);

INVx3_ASAP7_75t_L g1844 ( 
.A(n_1754),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1795),
.Y(n_1845)
);

HB1xp67_ASAP7_75t_L g1846 ( 
.A(n_1630),
.Y(n_1846)
);

AND2x2_ASAP7_75t_L g1847 ( 
.A(n_1703),
.B(n_1516),
.Y(n_1847)
);

HB1xp67_ASAP7_75t_L g1848 ( 
.A(n_1646),
.Y(n_1848)
);

AND2x2_ASAP7_75t_L g1849 ( 
.A(n_1744),
.B(n_1516),
.Y(n_1849)
);

AO31x2_ASAP7_75t_L g1850 ( 
.A1(n_1626),
.A2(n_1490),
.A3(n_1493),
.B(n_1478),
.Y(n_1850)
);

AO21x2_ASAP7_75t_L g1851 ( 
.A1(n_1762),
.A2(n_1548),
.B(n_1494),
.Y(n_1851)
);

INVx2_ASAP7_75t_L g1852 ( 
.A(n_1726),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1726),
.Y(n_1853)
);

AND2x2_ASAP7_75t_L g1854 ( 
.A(n_1763),
.B(n_1768),
.Y(n_1854)
);

OR2x2_ASAP7_75t_L g1855 ( 
.A(n_1815),
.B(n_1471),
.Y(n_1855)
);

HB1xp67_ASAP7_75t_L g1856 ( 
.A(n_1651),
.Y(n_1856)
);

INVx1_ASAP7_75t_L g1857 ( 
.A(n_1764),
.Y(n_1857)
);

OR2x2_ASAP7_75t_L g1858 ( 
.A(n_1819),
.B(n_1471),
.Y(n_1858)
);

OR2x2_ASAP7_75t_L g1859 ( 
.A(n_1801),
.B(n_1483),
.Y(n_1859)
);

INVx1_ASAP7_75t_SL g1860 ( 
.A(n_1717),
.Y(n_1860)
);

INVx2_ASAP7_75t_L g1861 ( 
.A(n_1726),
.Y(n_1861)
);

HB1xp67_ASAP7_75t_L g1862 ( 
.A(n_1669),
.Y(n_1862)
);

INVx2_ASAP7_75t_SL g1863 ( 
.A(n_1795),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1764),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1806),
.B(n_1516),
.Y(n_1865)
);

HB1xp67_ASAP7_75t_L g1866 ( 
.A(n_1708),
.Y(n_1866)
);

AOI222xp33_ASAP7_75t_L g1867 ( 
.A1(n_1627),
.A2(n_1475),
.B1(n_1524),
.B2(n_1505),
.C1(n_1508),
.C2(n_1513),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1826),
.B(n_1516),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1785),
.Y(n_1869)
);

AND2x4_ASAP7_75t_L g1870 ( 
.A(n_1803),
.B(n_1463),
.Y(n_1870)
);

BUFx6f_ASAP7_75t_L g1871 ( 
.A(n_1652),
.Y(n_1871)
);

AND2x2_ASAP7_75t_L g1872 ( 
.A(n_1751),
.B(n_1469),
.Y(n_1872)
);

AND2x2_ASAP7_75t_L g1873 ( 
.A(n_1758),
.B(n_1469),
.Y(n_1873)
);

INVx2_ASAP7_75t_L g1874 ( 
.A(n_1676),
.Y(n_1874)
);

NAND2xp5_ASAP7_75t_L g1875 ( 
.A(n_1704),
.B(n_1483),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1785),
.Y(n_1876)
);

OR2x2_ASAP7_75t_L g1877 ( 
.A(n_1707),
.B(n_1666),
.Y(n_1877)
);

AND2x2_ASAP7_75t_L g1878 ( 
.A(n_1694),
.B(n_1469),
.Y(n_1878)
);

INVx1_ASAP7_75t_L g1879 ( 
.A(n_1636),
.Y(n_1879)
);

NAND2xp5_ASAP7_75t_L g1880 ( 
.A(n_1747),
.B(n_1489),
.Y(n_1880)
);

INVx2_ASAP7_75t_L g1881 ( 
.A(n_1676),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1681),
.Y(n_1882)
);

INVx2_ASAP7_75t_L g1883 ( 
.A(n_1681),
.Y(n_1883)
);

BUFx2_ASAP7_75t_L g1884 ( 
.A(n_1762),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1683),
.Y(n_1885)
);

BUFx3_ASAP7_75t_L g1886 ( 
.A(n_1629),
.Y(n_1886)
);

BUFx6f_ASAP7_75t_L g1887 ( 
.A(n_1652),
.Y(n_1887)
);

OR2x2_ASAP7_75t_L g1888 ( 
.A(n_1655),
.B(n_1489),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1804),
.B(n_1479),
.Y(n_1889)
);

OR2x2_ASAP7_75t_L g1890 ( 
.A(n_1657),
.B(n_1680),
.Y(n_1890)
);

INVx2_ASAP7_75t_L g1891 ( 
.A(n_1696),
.Y(n_1891)
);

INVx2_ASAP7_75t_L g1892 ( 
.A(n_1696),
.Y(n_1892)
);

INVx2_ASAP7_75t_SL g1893 ( 
.A(n_1717),
.Y(n_1893)
);

INVx2_ASAP7_75t_SL g1894 ( 
.A(n_1754),
.Y(n_1894)
);

AOI33xp33_ASAP7_75t_L g1895 ( 
.A1(n_1633),
.A2(n_1556),
.A3(n_1557),
.B1(n_1510),
.B2(n_1545),
.B3(n_1538),
.Y(n_1895)
);

INVx2_ASAP7_75t_L g1896 ( 
.A(n_1700),
.Y(n_1896)
);

INVx4_ASAP7_75t_L g1897 ( 
.A(n_1652),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1687),
.Y(n_1898)
);

AND2x2_ASAP7_75t_L g1899 ( 
.A(n_1821),
.B(n_1822),
.Y(n_1899)
);

INVx3_ASAP7_75t_L g1900 ( 
.A(n_1813),
.Y(n_1900)
);

NAND2xp5_ASAP7_75t_L g1901 ( 
.A(n_1752),
.B(n_1475),
.Y(n_1901)
);

AOI22xp33_ASAP7_75t_L g1902 ( 
.A1(n_1769),
.A2(n_1557),
.B1(n_1460),
.B2(n_1506),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1700),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1719),
.Y(n_1904)
);

AND2x2_ASAP7_75t_L g1905 ( 
.A(n_1796),
.B(n_1479),
.Y(n_1905)
);

AND2x2_ASAP7_75t_L g1906 ( 
.A(n_1797),
.B(n_1479),
.Y(n_1906)
);

NOR2x1_ASAP7_75t_L g1907 ( 
.A(n_1667),
.B(n_1487),
.Y(n_1907)
);

INVx2_ASAP7_75t_L g1908 ( 
.A(n_1712),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1824),
.B(n_1487),
.Y(n_1909)
);

INVxp67_ASAP7_75t_SL g1910 ( 
.A(n_1639),
.Y(n_1910)
);

AND2x2_ASAP7_75t_L g1911 ( 
.A(n_1779),
.B(n_1487),
.Y(n_1911)
);

AND2x2_ASAP7_75t_L g1912 ( 
.A(n_1673),
.B(n_1731),
.Y(n_1912)
);

AND2x2_ASAP7_75t_L g1913 ( 
.A(n_1731),
.B(n_1587),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1721),
.Y(n_1914)
);

BUFx3_ASAP7_75t_L g1915 ( 
.A(n_1629),
.Y(n_1915)
);

INVx2_ASAP7_75t_L g1916 ( 
.A(n_1712),
.Y(n_1916)
);

AND2x4_ASAP7_75t_L g1917 ( 
.A(n_1803),
.B(n_1611),
.Y(n_1917)
);

AND2x2_ASAP7_75t_L g1918 ( 
.A(n_1731),
.B(n_1587),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1753),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1757),
.Y(n_1920)
);

OR2x2_ASAP7_75t_L g1921 ( 
.A(n_1698),
.B(n_1587),
.Y(n_1921)
);

AND2x2_ASAP7_75t_L g1922 ( 
.A(n_1714),
.B(n_1587),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_L g1923 ( 
.A(n_1643),
.B(n_1599),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1803),
.B(n_1611),
.Y(n_1924)
);

BUFx2_ASAP7_75t_L g1925 ( 
.A(n_1766),
.Y(n_1925)
);

INVx1_ASAP7_75t_L g1926 ( 
.A(n_1759),
.Y(n_1926)
);

INVx2_ASAP7_75t_L g1927 ( 
.A(n_1715),
.Y(n_1927)
);

INVx2_ASAP7_75t_L g1928 ( 
.A(n_1715),
.Y(n_1928)
);

BUFx2_ASAP7_75t_L g1929 ( 
.A(n_1766),
.Y(n_1929)
);

AOI221xp5_ASAP7_75t_L g1930 ( 
.A1(n_1713),
.A2(n_1568),
.B1(n_1561),
.B2(n_1551),
.C(n_1510),
.Y(n_1930)
);

INVx2_ASAP7_75t_L g1931 ( 
.A(n_1727),
.Y(n_1931)
);

OA21x2_ASAP7_75t_L g1932 ( 
.A1(n_1808),
.A2(n_1490),
.B(n_1493),
.Y(n_1932)
);

OR2x2_ASAP7_75t_L g1933 ( 
.A(n_1709),
.B(n_1561),
.Y(n_1933)
);

INVx2_ASAP7_75t_L g1934 ( 
.A(n_1727),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1770),
.Y(n_1935)
);

INVx5_ASAP7_75t_L g1936 ( 
.A(n_1784),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1780),
.Y(n_1937)
);

INVx2_ASAP7_75t_L g1938 ( 
.A(n_1733),
.Y(n_1938)
);

BUFx2_ASAP7_75t_L g1939 ( 
.A(n_1736),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1781),
.Y(n_1940)
);

INVx1_ASAP7_75t_L g1941 ( 
.A(n_1783),
.Y(n_1941)
);

AND2x2_ASAP7_75t_L g1942 ( 
.A(n_1730),
.B(n_1612),
.Y(n_1942)
);

OR2x2_ASAP7_75t_L g1943 ( 
.A(n_1716),
.B(n_1568),
.Y(n_1943)
);

AND2x4_ASAP7_75t_L g1944 ( 
.A(n_1699),
.B(n_1611),
.Y(n_1944)
);

INVx3_ASAP7_75t_L g1945 ( 
.A(n_1813),
.Y(n_1945)
);

INVx1_ASAP7_75t_L g1946 ( 
.A(n_1787),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1789),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1730),
.B(n_1612),
.Y(n_1948)
);

INVx2_ASAP7_75t_L g1949 ( 
.A(n_1733),
.Y(n_1949)
);

NOR2xp33_ASAP7_75t_L g1950 ( 
.A(n_1710),
.B(n_1638),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1743),
.B(n_1612),
.Y(n_1951)
);

INVx1_ASAP7_75t_L g1952 ( 
.A(n_1793),
.Y(n_1952)
);

AOI22xp5_ASAP7_75t_L g1953 ( 
.A1(n_1633),
.A2(n_1515),
.B1(n_1518),
.B2(n_1524),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1729),
.A2(n_1515),
.B1(n_1518),
.B2(n_1513),
.Y(n_1954)
);

AND2x2_ASAP7_75t_L g1955 ( 
.A(n_1743),
.B(n_1612),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1814),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1699),
.B(n_1611),
.Y(n_1957)
);

AND2x2_ASAP7_75t_L g1958 ( 
.A(n_1743),
.B(n_1613),
.Y(n_1958)
);

AND2x2_ASAP7_75t_L g1959 ( 
.A(n_1735),
.B(n_1613),
.Y(n_1959)
);

OR2x2_ASAP7_75t_L g1960 ( 
.A(n_1724),
.B(n_1551),
.Y(n_1960)
);

INVx1_ASAP7_75t_L g1961 ( 
.A(n_1818),
.Y(n_1961)
);

INVx1_ASAP7_75t_L g1962 ( 
.A(n_1831),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1838),
.Y(n_1963)
);

AND2x2_ASAP7_75t_L g1964 ( 
.A(n_1738),
.B(n_1613),
.Y(n_1964)
);

OAI21x1_ASAP7_75t_L g1965 ( 
.A1(n_1670),
.A2(n_1558),
.B(n_1685),
.Y(n_1965)
);

INVx2_ASAP7_75t_L g1966 ( 
.A(n_1741),
.Y(n_1966)
);

INVx2_ASAP7_75t_L g1967 ( 
.A(n_1741),
.Y(n_1967)
);

INVx2_ASAP7_75t_L g1968 ( 
.A(n_1745),
.Y(n_1968)
);

INVx5_ASAP7_75t_L g1969 ( 
.A(n_1784),
.Y(n_1969)
);

OR2x2_ASAP7_75t_L g1970 ( 
.A(n_1761),
.B(n_1605),
.Y(n_1970)
);

INVx1_ASAP7_75t_L g1971 ( 
.A(n_1843),
.Y(n_1971)
);

INVx2_ASAP7_75t_L g1972 ( 
.A(n_1745),
.Y(n_1972)
);

INVx3_ASAP7_75t_L g1973 ( 
.A(n_1813),
.Y(n_1973)
);

BUFx4f_ASAP7_75t_SL g1974 ( 
.A(n_1706),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1755),
.B(n_1613),
.Y(n_1975)
);

INVx2_ASAP7_75t_L g1976 ( 
.A(n_1749),
.Y(n_1976)
);

INVx1_ASAP7_75t_SL g1977 ( 
.A(n_1835),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1749),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1813),
.Y(n_1979)
);

INVx2_ASAP7_75t_L g1980 ( 
.A(n_1750),
.Y(n_1980)
);

BUFx2_ASAP7_75t_L g1981 ( 
.A(n_1736),
.Y(n_1981)
);

OAI21xp5_ASAP7_75t_L g1982 ( 
.A1(n_1664),
.A2(n_1528),
.B(n_1511),
.Y(n_1982)
);

HB1xp67_ASAP7_75t_L g1983 ( 
.A(n_1644),
.Y(n_1983)
);

INVx1_ASAP7_75t_L g1984 ( 
.A(n_1750),
.Y(n_1984)
);

AND2x4_ASAP7_75t_SL g1985 ( 
.A(n_1652),
.B(n_1611),
.Y(n_1985)
);

OAI31xp33_ASAP7_75t_L g1986 ( 
.A1(n_1631),
.A2(n_1635),
.A3(n_1647),
.B(n_1776),
.Y(n_1986)
);

HB1xp67_ASAP7_75t_L g1987 ( 
.A(n_1760),
.Y(n_1987)
);

AND2x2_ASAP7_75t_L g1988 ( 
.A(n_1799),
.B(n_1614),
.Y(n_1988)
);

OR2x2_ASAP7_75t_L g1989 ( 
.A(n_1756),
.B(n_1605),
.Y(n_1989)
);

NAND2x1p5_ASAP7_75t_L g1990 ( 
.A(n_1825),
.B(n_1528),
.Y(n_1990)
);

NAND2xp33_ASAP7_75t_R g1991 ( 
.A(n_1688),
.B(n_1577),
.Y(n_1991)
);

AOI22xp33_ASAP7_75t_SL g1992 ( 
.A1(n_1778),
.A2(n_1515),
.B1(n_1611),
.B2(n_1480),
.Y(n_1992)
);

AND2x2_ASAP7_75t_L g1993 ( 
.A(n_1650),
.B(n_1614),
.Y(n_1993)
);

INVx2_ASAP7_75t_L g1994 ( 
.A(n_1788),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1654),
.B(n_1599),
.Y(n_1995)
);

AND2x2_ASAP7_75t_L g1996 ( 
.A(n_1658),
.B(n_1614),
.Y(n_1996)
);

INVx2_ASAP7_75t_L g1997 ( 
.A(n_1788),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1728),
.Y(n_1998)
);

BUFx6f_ASAP7_75t_L g1999 ( 
.A(n_1710),
.Y(n_1999)
);

AND2x2_ASAP7_75t_L g2000 ( 
.A(n_1628),
.B(n_1614),
.Y(n_2000)
);

INVx2_ASAP7_75t_L g2001 ( 
.A(n_1810),
.Y(n_2001)
);

AND2x2_ASAP7_75t_L g2002 ( 
.A(n_1645),
.B(n_1538),
.Y(n_2002)
);

INVx2_ASAP7_75t_L g2003 ( 
.A(n_1810),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1840),
.B(n_1538),
.Y(n_2004)
);

AND2x2_ASAP7_75t_L g2005 ( 
.A(n_1840),
.B(n_1545),
.Y(n_2005)
);

OR2x2_ASAP7_75t_L g2006 ( 
.A(n_1772),
.B(n_1600),
.Y(n_2006)
);

AND2x4_ASAP7_75t_SL g2007 ( 
.A(n_1686),
.B(n_1611),
.Y(n_2007)
);

INVx1_ASAP7_75t_L g2008 ( 
.A(n_1728),
.Y(n_2008)
);

BUFx2_ASAP7_75t_L g2009 ( 
.A(n_1739),
.Y(n_2009)
);

INVx2_ASAP7_75t_L g2010 ( 
.A(n_1820),
.Y(n_2010)
);

INVx1_ASAP7_75t_L g2011 ( 
.A(n_1728),
.Y(n_2011)
);

INVx8_ASAP7_75t_L g2012 ( 
.A(n_1675),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1728),
.Y(n_2013)
);

INVx3_ASAP7_75t_L g2014 ( 
.A(n_1820),
.Y(n_2014)
);

INVx1_ASAP7_75t_L g2015 ( 
.A(n_1828),
.Y(n_2015)
);

AOI22xp33_ASAP7_75t_L g2016 ( 
.A1(n_1776),
.A2(n_1460),
.B1(n_1279),
.B2(n_1480),
.Y(n_2016)
);

AND2x2_ASAP7_75t_L g2017 ( 
.A(n_1765),
.B(n_1545),
.Y(n_2017)
);

INVx2_ASAP7_75t_L g2018 ( 
.A(n_1829),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1765),
.B(n_1480),
.Y(n_2019)
);

AND2x2_ASAP7_75t_L g2020 ( 
.A(n_1663),
.B(n_1480),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_L g2021 ( 
.A(n_1695),
.B(n_1600),
.Y(n_2021)
);

AND2x4_ASAP7_75t_L g2022 ( 
.A(n_1699),
.B(n_1480),
.Y(n_2022)
);

HB1xp67_ASAP7_75t_L g2023 ( 
.A(n_1760),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1829),
.Y(n_2024)
);

NAND2xp33_ASAP7_75t_R g2025 ( 
.A(n_1688),
.B(n_1577),
.Y(n_2025)
);

AND2x2_ASAP7_75t_L g2026 ( 
.A(n_1674),
.B(n_1480),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1832),
.Y(n_2027)
);

HB1xp67_ASAP7_75t_L g2028 ( 
.A(n_1732),
.Y(n_2028)
);

INVx1_ASAP7_75t_L g2029 ( 
.A(n_1830),
.Y(n_2029)
);

HB1xp67_ASAP7_75t_L g2030 ( 
.A(n_1740),
.Y(n_2030)
);

AND2x2_ASAP7_75t_L g2031 ( 
.A(n_1684),
.B(n_1480),
.Y(n_2031)
);

INVx1_ASAP7_75t_L g2032 ( 
.A(n_1830),
.Y(n_2032)
);

OAI222xp33_ASAP7_75t_L g2033 ( 
.A1(n_1677),
.A2(n_1567),
.B1(n_1508),
.B2(n_1505),
.C1(n_1470),
.C2(n_1455),
.Y(n_2033)
);

INVx3_ASAP7_75t_L g2034 ( 
.A(n_1834),
.Y(n_2034)
);

INVx2_ASAP7_75t_L g2035 ( 
.A(n_1834),
.Y(n_2035)
);

OA21x2_ASAP7_75t_L g2036 ( 
.A1(n_1842),
.A2(n_1499),
.B(n_1558),
.Y(n_2036)
);

NOR2xp33_ASAP7_75t_L g2037 ( 
.A(n_1675),
.B(n_1579),
.Y(n_2037)
);

BUFx2_ASAP7_75t_L g2038 ( 
.A(n_1739),
.Y(n_2038)
);

AND2x4_ASAP7_75t_L g2039 ( 
.A(n_1792),
.B(n_1558),
.Y(n_2039)
);

NOR3xp33_ASAP7_75t_L g2040 ( 
.A(n_1642),
.B(n_1528),
.C(n_1606),
.Y(n_2040)
);

INVx2_ASAP7_75t_L g2041 ( 
.A(n_1842),
.Y(n_2041)
);

BUFx3_ASAP7_75t_L g2042 ( 
.A(n_1668),
.Y(n_2042)
);

INVxp67_ASAP7_75t_SL g2043 ( 
.A(n_1639),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1792),
.B(n_1491),
.Y(n_2044)
);

INVx2_ASAP7_75t_L g2045 ( 
.A(n_1672),
.Y(n_2045)
);

INVx4_ASAP7_75t_L g2046 ( 
.A(n_1686),
.Y(n_2046)
);

INVx1_ASAP7_75t_L g2047 ( 
.A(n_1734),
.Y(n_2047)
);

BUFx2_ASAP7_75t_L g2048 ( 
.A(n_1817),
.Y(n_2048)
);

INVx1_ASAP7_75t_L g2049 ( 
.A(n_1734),
.Y(n_2049)
);

INVx2_ASAP7_75t_L g2050 ( 
.A(n_1672),
.Y(n_2050)
);

AND2x2_ASAP7_75t_L g2051 ( 
.A(n_1640),
.B(n_1477),
.Y(n_2051)
);

BUFx2_ASAP7_75t_L g2052 ( 
.A(n_1817),
.Y(n_2052)
);

AND2x4_ASAP7_75t_L g2053 ( 
.A(n_1827),
.B(n_1491),
.Y(n_2053)
);

BUFx2_ASAP7_75t_L g2054 ( 
.A(n_1718),
.Y(n_2054)
);

AND2x2_ASAP7_75t_L g2055 ( 
.A(n_1640),
.B(n_1477),
.Y(n_2055)
);

HB1xp67_ASAP7_75t_L g2056 ( 
.A(n_1773),
.Y(n_2056)
);

INVx1_ASAP7_75t_L g2057 ( 
.A(n_1734),
.Y(n_2057)
);

AND2x2_ASAP7_75t_L g2058 ( 
.A(n_1774),
.B(n_1481),
.Y(n_2058)
);

INVx2_ASAP7_75t_L g2059 ( 
.A(n_1852),
.Y(n_2059)
);

AO21x2_ASAP7_75t_L g2060 ( 
.A1(n_1910),
.A2(n_1825),
.B(n_1499),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_L g2061 ( 
.A(n_2028),
.B(n_1701),
.Y(n_2061)
);

OR2x2_ASAP7_75t_L g2062 ( 
.A(n_1877),
.B(n_1648),
.Y(n_2062)
);

OAI21x1_ASAP7_75t_L g2063 ( 
.A1(n_1965),
.A2(n_1685),
.B(n_1774),
.Y(n_2063)
);

INVx2_ASAP7_75t_L g2064 ( 
.A(n_1852),
.Y(n_2064)
);

AND2x2_ASAP7_75t_L g2065 ( 
.A(n_1847),
.B(n_1705),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_2042),
.Y(n_2066)
);

OAI22xp33_ASAP7_75t_L g2067 ( 
.A1(n_1991),
.A2(n_1686),
.B1(n_1794),
.B2(n_1767),
.Y(n_2067)
);

AOI21xp5_ASAP7_75t_L g2068 ( 
.A1(n_1986),
.A2(n_1631),
.B(n_1767),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_L g2069 ( 
.A(n_2030),
.B(n_1901),
.Y(n_2069)
);

A2O1A1Ixp33_ASAP7_75t_L g2070 ( 
.A1(n_1986),
.A2(n_1659),
.B(n_1702),
.C(n_1748),
.Y(n_2070)
);

AOI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1867),
.A2(n_1790),
.B(n_1782),
.Y(n_2071)
);

AOI222xp33_ASAP7_75t_L g2072 ( 
.A1(n_1930),
.A2(n_1634),
.B1(n_1811),
.B2(n_1660),
.C1(n_1679),
.C2(n_1823),
.Y(n_2072)
);

INVx1_ASAP7_75t_L g2073 ( 
.A(n_1879),
.Y(n_2073)
);

INVx2_ASAP7_75t_SL g2074 ( 
.A(n_1886),
.Y(n_2074)
);

INVx2_ASAP7_75t_L g2075 ( 
.A(n_1852),
.Y(n_2075)
);

OAI21xp33_ASAP7_75t_L g2076 ( 
.A1(n_1867),
.A2(n_1634),
.B(n_1811),
.Y(n_2076)
);

AOI21xp5_ASAP7_75t_L g2077 ( 
.A1(n_2012),
.A2(n_1907),
.B(n_1982),
.Y(n_2077)
);

INVx2_ASAP7_75t_L g2078 ( 
.A(n_1853),
.Y(n_2078)
);

INVx1_ASAP7_75t_L g2079 ( 
.A(n_1879),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1901),
.B(n_1786),
.Y(n_2080)
);

INVx1_ASAP7_75t_L g2081 ( 
.A(n_1885),
.Y(n_2081)
);

BUFx2_ASAP7_75t_L g2082 ( 
.A(n_2009),
.Y(n_2082)
);

BUFx3_ASAP7_75t_L g2083 ( 
.A(n_2042),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1846),
.Y(n_2084)
);

AND2x2_ASAP7_75t_L g2085 ( 
.A(n_1987),
.B(n_1722),
.Y(n_2085)
);

INVx2_ASAP7_75t_L g2086 ( 
.A(n_1853),
.Y(n_2086)
);

INVxp67_ASAP7_75t_SL g2087 ( 
.A(n_2023),
.Y(n_2087)
);

INVx1_ASAP7_75t_L g2088 ( 
.A(n_1885),
.Y(n_2088)
);

INVx2_ASAP7_75t_L g2089 ( 
.A(n_1853),
.Y(n_2089)
);

A2O1A1Ixp33_ASAP7_75t_L g2090 ( 
.A1(n_1895),
.A2(n_1823),
.B(n_1771),
.C(n_1679),
.Y(n_2090)
);

INVx1_ASAP7_75t_L g2091 ( 
.A(n_1898),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_L g2092 ( 
.A(n_1875),
.B(n_1802),
.Y(n_2092)
);

AND2x2_ASAP7_75t_L g2093 ( 
.A(n_1884),
.B(n_1723),
.Y(n_2093)
);

OA21x2_ASAP7_75t_L g2094 ( 
.A1(n_1982),
.A2(n_1521),
.B(n_1548),
.Y(n_2094)
);

OAI21xp5_ASAP7_75t_L g2095 ( 
.A1(n_1954),
.A2(n_1632),
.B(n_1841),
.Y(n_2095)
);

AOI21xp5_ASAP7_75t_L g2096 ( 
.A1(n_2012),
.A2(n_1839),
.B(n_1805),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1886),
.B(n_1693),
.Y(n_2097)
);

AO21x2_ASAP7_75t_L g2098 ( 
.A1(n_2043),
.A2(n_1494),
.B(n_1521),
.Y(n_2098)
);

INVx1_ASAP7_75t_SL g2099 ( 
.A(n_1974),
.Y(n_2099)
);

INVx2_ASAP7_75t_L g2100 ( 
.A(n_1861),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_L g2101 ( 
.A(n_1875),
.B(n_1662),
.Y(n_2101)
);

INVx1_ASAP7_75t_L g2102 ( 
.A(n_1898),
.Y(n_2102)
);

OAI211xp5_ASAP7_75t_L g2103 ( 
.A1(n_1954),
.A2(n_1953),
.B(n_1992),
.C(n_1902),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1884),
.B(n_1777),
.Y(n_2104)
);

BUFx2_ASAP7_75t_L g2105 ( 
.A(n_2009),
.Y(n_2105)
);

OAI22xp5_ASAP7_75t_L g2106 ( 
.A1(n_1953),
.A2(n_2038),
.B1(n_1833),
.B2(n_2016),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1904),
.Y(n_2107)
);

INVx1_ASAP7_75t_L g2108 ( 
.A(n_1904),
.Y(n_2108)
);

BUFx3_ASAP7_75t_L g2109 ( 
.A(n_2042),
.Y(n_2109)
);

AOI21xp5_ASAP7_75t_L g2110 ( 
.A1(n_2012),
.A2(n_1839),
.B(n_1837),
.Y(n_2110)
);

INVx1_ASAP7_75t_L g2111 ( 
.A(n_1914),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1861),
.Y(n_2112)
);

INVx2_ASAP7_75t_L g2113 ( 
.A(n_1861),
.Y(n_2113)
);

A2O1A1Ixp33_ASAP7_75t_L g2114 ( 
.A1(n_1907),
.A2(n_1929),
.B(n_1925),
.C(n_1939),
.Y(n_2114)
);

INVx1_ASAP7_75t_L g2115 ( 
.A(n_1914),
.Y(n_2115)
);

AO31x2_ASAP7_75t_L g2116 ( 
.A1(n_1925),
.A2(n_1649),
.A3(n_1621),
.B(n_1618),
.Y(n_2116)
);

INVxp67_ASAP7_75t_L g2117 ( 
.A(n_2025),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_L g2118 ( 
.A(n_2056),
.B(n_1777),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1919),
.Y(n_2119)
);

INVx4_ASAP7_75t_SL g2120 ( 
.A(n_1871),
.Y(n_2120)
);

INVx1_ASAP7_75t_L g2121 ( 
.A(n_1919),
.Y(n_2121)
);

BUFx3_ASAP7_75t_L g2122 ( 
.A(n_2012),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_SL g2123 ( 
.A(n_1929),
.B(n_1689),
.Y(n_2123)
);

BUFx2_ASAP7_75t_L g2124 ( 
.A(n_2038),
.Y(n_2124)
);

OAI21x1_ASAP7_75t_L g2125 ( 
.A1(n_1965),
.A2(n_1618),
.B(n_1621),
.Y(n_2125)
);

A2O1A1Ixp33_ASAP7_75t_L g2126 ( 
.A1(n_1939),
.A2(n_1791),
.B(n_1665),
.C(n_1656),
.Y(n_2126)
);

A2O1A1Ixp33_ASAP7_75t_L g2127 ( 
.A1(n_1981),
.A2(n_1791),
.B(n_1665),
.C(n_1656),
.Y(n_2127)
);

INVxp67_ASAP7_75t_SL g2128 ( 
.A(n_1990),
.Y(n_2128)
);

HB1xp67_ASAP7_75t_L g2129 ( 
.A(n_1848),
.Y(n_2129)
);

AO31x2_ASAP7_75t_L g2130 ( 
.A1(n_1981),
.A2(n_1649),
.A3(n_1621),
.B(n_1618),
.Y(n_2130)
);

INVx2_ASAP7_75t_L g2131 ( 
.A(n_2047),
.Y(n_2131)
);

HB1xp67_ASAP7_75t_L g2132 ( 
.A(n_1856),
.Y(n_2132)
);

NAND2x1_ASAP7_75t_L g2133 ( 
.A(n_2046),
.B(n_1827),
.Y(n_2133)
);

OR2x2_ASAP7_75t_L g2134 ( 
.A(n_1877),
.B(n_1784),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1983),
.B(n_1455),
.Y(n_2135)
);

BUFx6f_ASAP7_75t_L g2136 ( 
.A(n_2012),
.Y(n_2136)
);

INVx1_ASAP7_75t_L g2137 ( 
.A(n_1920),
.Y(n_2137)
);

OAI21xp33_ASAP7_75t_L g2138 ( 
.A1(n_1880),
.A2(n_1778),
.B(n_1641),
.Y(n_2138)
);

AOI22xp33_ASAP7_75t_L g2139 ( 
.A1(n_1886),
.A2(n_1641),
.B1(n_1798),
.B2(n_1697),
.Y(n_2139)
);

INVx2_ASAP7_75t_L g2140 ( 
.A(n_2047),
.Y(n_2140)
);

INVx1_ASAP7_75t_SL g2141 ( 
.A(n_1915),
.Y(n_2141)
);

INVx1_ASAP7_75t_L g2142 ( 
.A(n_1920),
.Y(n_2142)
);

INVx1_ASAP7_75t_L g2143 ( 
.A(n_1926),
.Y(n_2143)
);

INVx2_ASAP7_75t_L g2144 ( 
.A(n_2049),
.Y(n_2144)
);

NAND4xp25_ASAP7_75t_L g2145 ( 
.A(n_2040),
.B(n_1682),
.C(n_1746),
.D(n_1692),
.Y(n_2145)
);

OAI21x1_ASAP7_75t_L g2146 ( 
.A1(n_1990),
.A2(n_1945),
.B(n_1900),
.Y(n_2146)
);

INVx1_ASAP7_75t_L g2147 ( 
.A(n_1926),
.Y(n_2147)
);

INVxp67_ASAP7_75t_L g2148 ( 
.A(n_1866),
.Y(n_2148)
);

AOI22xp33_ASAP7_75t_L g2149 ( 
.A1(n_1915),
.A2(n_1798),
.B1(n_1697),
.B2(n_1661),
.Y(n_2149)
);

INVx4_ASAP7_75t_L g2150 ( 
.A(n_1871),
.Y(n_2150)
);

AND2x2_ASAP7_75t_L g2151 ( 
.A(n_2019),
.B(n_1827),
.Y(n_2151)
);

HB1xp67_ASAP7_75t_L g2152 ( 
.A(n_1862),
.Y(n_2152)
);

OR2x2_ASAP7_75t_L g2153 ( 
.A(n_1890),
.B(n_1481),
.Y(n_2153)
);

INVxp67_ASAP7_75t_L g2154 ( 
.A(n_2037),
.Y(n_2154)
);

AOI22xp33_ASAP7_75t_L g2155 ( 
.A1(n_1915),
.A2(n_1661),
.B1(n_1689),
.B2(n_1691),
.Y(n_2155)
);

AND2x4_ASAP7_75t_L g2156 ( 
.A(n_2046),
.B(n_1837),
.Y(n_2156)
);

AOI21x1_ASAP7_75t_L g2157 ( 
.A1(n_2054),
.A2(n_1837),
.B(n_1606),
.Y(n_2157)
);

OAI22xp33_ASAP7_75t_L g2158 ( 
.A1(n_1871),
.A2(n_1692),
.B1(n_1637),
.B2(n_1682),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_2049),
.Y(n_2159)
);

OAI22xp33_ASAP7_75t_L g2160 ( 
.A1(n_1871),
.A2(n_1637),
.B1(n_1775),
.B2(n_1800),
.Y(n_2160)
);

INVx2_ASAP7_75t_L g2161 ( 
.A(n_2057),
.Y(n_2161)
);

INVx4_ASAP7_75t_L g2162 ( 
.A(n_1871),
.Y(n_2162)
);

A2O1A1Ixp33_ASAP7_75t_L g2163 ( 
.A1(n_1950),
.A2(n_1711),
.B(n_1720),
.C(n_1737),
.Y(n_2163)
);

AOI21xp5_ASAP7_75t_L g2164 ( 
.A1(n_2033),
.A2(n_1836),
.B(n_1491),
.Y(n_2164)
);

OAI21xp33_ASAP7_75t_L g2165 ( 
.A1(n_1880),
.A2(n_1691),
.B(n_1725),
.Y(n_2165)
);

NAND2xp5_ASAP7_75t_L g2166 ( 
.A(n_1890),
.B(n_1456),
.Y(n_2166)
);

INVx1_ASAP7_75t_L g2167 ( 
.A(n_1935),
.Y(n_2167)
);

AO21x2_ASAP7_75t_L g2168 ( 
.A1(n_1851),
.A2(n_1607),
.B(n_1725),
.Y(n_2168)
);

OAI21x1_ASAP7_75t_L g2169 ( 
.A1(n_1990),
.A2(n_1607),
.B(n_1543),
.Y(n_2169)
);

AOI221xp5_ASAP7_75t_L g2170 ( 
.A1(n_2015),
.A2(n_1742),
.B1(n_1476),
.B2(n_1472),
.C(n_1470),
.Y(n_2170)
);

A2O1A1Ixp33_ASAP7_75t_L g2171 ( 
.A1(n_2007),
.A2(n_1720),
.B(n_1737),
.C(n_1711),
.Y(n_2171)
);

BUFx3_ASAP7_75t_L g2172 ( 
.A(n_1999),
.Y(n_2172)
);

AOI21xp33_ASAP7_75t_L g2173 ( 
.A1(n_1933),
.A2(n_1746),
.B(n_1775),
.Y(n_2173)
);

INVxp67_ASAP7_75t_L g2174 ( 
.A(n_1995),
.Y(n_2174)
);

AOI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1995),
.A2(n_1586),
.B(n_1653),
.Y(n_2175)
);

BUFx6f_ASAP7_75t_L g2176 ( 
.A(n_1871),
.Y(n_2176)
);

OAI31xp33_ASAP7_75t_L g2177 ( 
.A1(n_2048),
.A2(n_1456),
.A3(n_1472),
.B(n_1464),
.Y(n_2177)
);

OAI211xp5_ASAP7_75t_L g2178 ( 
.A1(n_2046),
.A2(n_1807),
.B(n_1458),
.C(n_1464),
.Y(n_2178)
);

OAI21x1_ASAP7_75t_L g2179 ( 
.A1(n_1900),
.A2(n_1607),
.B(n_1543),
.Y(n_2179)
);

NAND2x1_ASAP7_75t_L g2180 ( 
.A(n_2046),
.B(n_1514),
.Y(n_2180)
);

AND2x2_ASAP7_75t_L g2181 ( 
.A(n_2019),
.B(n_1678),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1935),
.Y(n_2182)
);

BUFx2_ASAP7_75t_L g2183 ( 
.A(n_1887),
.Y(n_2183)
);

OR2x2_ASAP7_75t_L g2184 ( 
.A(n_1933),
.B(n_1481),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_SL g2185 ( 
.A(n_1999),
.B(n_1807),
.Y(n_2185)
);

AND2x2_ASAP7_75t_L g2186 ( 
.A(n_1872),
.B(n_1678),
.Y(n_2186)
);

AOI22xp33_ASAP7_75t_L g2187 ( 
.A1(n_1887),
.A2(n_1742),
.B1(n_1671),
.B2(n_1690),
.Y(n_2187)
);

NOR2xp33_ASAP7_75t_L g2188 ( 
.A(n_1999),
.B(n_1457),
.Y(n_2188)
);

INVx1_ASAP7_75t_L g2189 ( 
.A(n_1937),
.Y(n_2189)
);

AO21x2_ASAP7_75t_L g2190 ( 
.A1(n_1851),
.A2(n_2008),
.B(n_1998),
.Y(n_2190)
);

OA21x2_ASAP7_75t_L g2191 ( 
.A1(n_1998),
.A2(n_1543),
.B(n_1542),
.Y(n_2191)
);

INVx1_ASAP7_75t_L g2192 ( 
.A(n_1937),
.Y(n_2192)
);

INVx1_ASAP7_75t_L g2193 ( 
.A(n_1940),
.Y(n_2193)
);

INVx1_ASAP7_75t_L g2194 ( 
.A(n_1940),
.Y(n_2194)
);

OAI22xp33_ASAP7_75t_L g2195 ( 
.A1(n_1887),
.A2(n_1800),
.B1(n_1812),
.B2(n_1809),
.Y(n_2195)
);

INVx1_ASAP7_75t_L g2196 ( 
.A(n_1941),
.Y(n_2196)
);

INVx1_ASAP7_75t_L g2197 ( 
.A(n_1941),
.Y(n_2197)
);

INVx1_ASAP7_75t_L g2198 ( 
.A(n_1946),
.Y(n_2198)
);

INVxp67_ASAP7_75t_L g2199 ( 
.A(n_2021),
.Y(n_2199)
);

OAI22xp33_ASAP7_75t_L g2200 ( 
.A1(n_1887),
.A2(n_1812),
.B1(n_1816),
.B2(n_1809),
.Y(n_2200)
);

INVx1_ASAP7_75t_L g2201 ( 
.A(n_1946),
.Y(n_2201)
);

OAI21x1_ASAP7_75t_L g2202 ( 
.A1(n_1900),
.A2(n_1542),
.B(n_1502),
.Y(n_2202)
);

OAI21xp33_ASAP7_75t_L g2203 ( 
.A1(n_1943),
.A2(n_1457),
.B(n_1458),
.Y(n_2203)
);

O2A1O1Ixp5_ASAP7_75t_L g2204 ( 
.A1(n_1870),
.A2(n_1923),
.B(n_1924),
.C(n_1917),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_1947),
.Y(n_2205)
);

OAI221xp5_ASAP7_75t_L g2206 ( 
.A1(n_1943),
.A2(n_1816),
.B1(n_1476),
.B2(n_1593),
.C(n_1591),
.Y(n_2206)
);

OR2x2_ASAP7_75t_L g2207 ( 
.A(n_1960),
.B(n_1485),
.Y(n_2207)
);

INVx2_ASAP7_75t_L g2208 ( 
.A(n_2057),
.Y(n_2208)
);

AOI22xp33_ASAP7_75t_L g2209 ( 
.A1(n_1887),
.A2(n_1690),
.B1(n_1671),
.B2(n_1502),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1947),
.Y(n_2210)
);

INVx1_ASAP7_75t_SL g2211 ( 
.A(n_1999),
.Y(n_2211)
);

INVx2_ASAP7_75t_L g2212 ( 
.A(n_2008),
.Y(n_2212)
);

NOR2xp33_ASAP7_75t_L g2213 ( 
.A(n_1999),
.B(n_1894),
.Y(n_2213)
);

BUFx2_ASAP7_75t_L g2214 ( 
.A(n_1887),
.Y(n_2214)
);

AOI22xp33_ASAP7_75t_L g2215 ( 
.A1(n_1844),
.A2(n_1502),
.B1(n_1507),
.B2(n_1542),
.Y(n_2215)
);

AOI221xp5_ASAP7_75t_L g2216 ( 
.A1(n_2015),
.A2(n_1583),
.B1(n_1584),
.B2(n_1582),
.C(n_1579),
.Y(n_2216)
);

AOI21xp5_ASAP7_75t_L g2217 ( 
.A1(n_1923),
.A2(n_1586),
.B(n_1595),
.Y(n_2217)
);

INVx2_ASAP7_75t_L g2218 ( 
.A(n_2011),
.Y(n_2218)
);

OR2x2_ASAP7_75t_L g2219 ( 
.A(n_1960),
.B(n_1888),
.Y(n_2219)
);

AO21x2_ASAP7_75t_L g2220 ( 
.A1(n_1851),
.A2(n_1507),
.B(n_1501),
.Y(n_2220)
);

INVx1_ASAP7_75t_L g2221 ( 
.A(n_1952),
.Y(n_2221)
);

AOI22xp33_ASAP7_75t_L g2222 ( 
.A1(n_1844),
.A2(n_1507),
.B1(n_1387),
.B2(n_1397),
.Y(n_2222)
);

OR2x2_ASAP7_75t_L g2223 ( 
.A(n_1888),
.B(n_1485),
.Y(n_2223)
);

INVx2_ASAP7_75t_L g2224 ( 
.A(n_2011),
.Y(n_2224)
);

OAI21xp5_ASAP7_75t_L g2225 ( 
.A1(n_2021),
.A2(n_1586),
.B(n_1511),
.Y(n_2225)
);

INVx3_ASAP7_75t_L g2226 ( 
.A(n_1900),
.Y(n_2226)
);

AOI22xp5_ASAP7_75t_L g2227 ( 
.A1(n_1894),
.A2(n_1517),
.B1(n_1514),
.B2(n_1591),
.Y(n_2227)
);

AOI22xp33_ASAP7_75t_L g2228 ( 
.A1(n_1844),
.A2(n_1387),
.B1(n_1397),
.B2(n_1514),
.Y(n_2228)
);

AOI211xp5_ASAP7_75t_L g2229 ( 
.A1(n_1917),
.A2(n_1588),
.B(n_1582),
.C(n_1584),
.Y(n_2229)
);

INVx2_ASAP7_75t_SL g2230 ( 
.A(n_1999),
.Y(n_2230)
);

BUFx6f_ASAP7_75t_L g2231 ( 
.A(n_1897),
.Y(n_2231)
);

AO21x2_ASAP7_75t_L g2232 ( 
.A1(n_1851),
.A2(n_1501),
.B(n_1465),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2027),
.B(n_1596),
.Y(n_2233)
);

BUFx2_ASAP7_75t_L g2234 ( 
.A(n_1897),
.Y(n_2234)
);

INVx1_ASAP7_75t_L g2235 ( 
.A(n_1952),
.Y(n_2235)
);

INVx2_ASAP7_75t_L g2236 ( 
.A(n_2013),
.Y(n_2236)
);

INVx1_ASAP7_75t_L g2237 ( 
.A(n_1956),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_1945),
.Y(n_2238)
);

NOR2xp33_ASAP7_75t_L g2239 ( 
.A(n_2048),
.B(n_1593),
.Y(n_2239)
);

AND2x2_ASAP7_75t_L g2240 ( 
.A(n_1872),
.B(n_1678),
.Y(n_2240)
);

INVx1_ASAP7_75t_L g2241 ( 
.A(n_1956),
.Y(n_2241)
);

INVx1_ASAP7_75t_L g2242 ( 
.A(n_1961),
.Y(n_2242)
);

AND2x2_ASAP7_75t_L g2243 ( 
.A(n_1873),
.B(n_1678),
.Y(n_2243)
);

INVx1_ASAP7_75t_L g2244 ( 
.A(n_2073),
.Y(n_2244)
);

NAND3xp33_ASAP7_75t_L g2245 ( 
.A(n_2068),
.B(n_1969),
.C(n_1936),
.Y(n_2245)
);

AND2x2_ASAP7_75t_L g2246 ( 
.A(n_2093),
.B(n_1913),
.Y(n_2246)
);

NAND3xp33_ASAP7_75t_L g2247 ( 
.A(n_2070),
.B(n_1969),
.C(n_1936),
.Y(n_2247)
);

AOI22xp33_ASAP7_75t_L g2248 ( 
.A1(n_2095),
.A2(n_1844),
.B1(n_2052),
.B2(n_1897),
.Y(n_2248)
);

HB1xp67_ASAP7_75t_L g2249 ( 
.A(n_2082),
.Y(n_2249)
);

AND2x2_ASAP7_75t_L g2250 ( 
.A(n_2093),
.B(n_1913),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_2146),
.Y(n_2251)
);

OAI33xp33_ASAP7_75t_L g2252 ( 
.A1(n_2106),
.A2(n_2027),
.A3(n_1859),
.B1(n_2006),
.B2(n_1858),
.B3(n_1855),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_2148),
.B(n_1899),
.Y(n_2253)
);

BUFx2_ASAP7_75t_L g2254 ( 
.A(n_2120),
.Y(n_2254)
);

AND2x2_ASAP7_75t_L g2255 ( 
.A(n_2105),
.B(n_1918),
.Y(n_2255)
);

AOI33xp33_ASAP7_75t_L g2256 ( 
.A1(n_2158),
.A2(n_1870),
.A3(n_2053),
.B1(n_1917),
.B2(n_1924),
.B3(n_1977),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_2124),
.B(n_1918),
.Y(n_2257)
);

INVx5_ASAP7_75t_L g2258 ( 
.A(n_2176),
.Y(n_2258)
);

INVxp33_ASAP7_75t_SL g2259 ( 
.A(n_2097),
.Y(n_2259)
);

NAND2xp5_ASAP7_75t_L g2260 ( 
.A(n_2071),
.B(n_1899),
.Y(n_2260)
);

INVx2_ASAP7_75t_L g2261 ( 
.A(n_2190),
.Y(n_2261)
);

INVx4_ASAP7_75t_L g2262 ( 
.A(n_2066),
.Y(n_2262)
);

NAND3xp33_ASAP7_75t_SL g2263 ( 
.A(n_2070),
.B(n_2052),
.C(n_2054),
.Y(n_2263)
);

AOI221xp5_ASAP7_75t_L g2264 ( 
.A1(n_2103),
.A2(n_1870),
.B1(n_2053),
.B2(n_1917),
.C(n_1924),
.Y(n_2264)
);

INVx2_ASAP7_75t_L g2265 ( 
.A(n_2190),
.Y(n_2265)
);

INVx1_ASAP7_75t_L g2266 ( 
.A(n_2079),
.Y(n_2266)
);

AND2x2_ASAP7_75t_L g2267 ( 
.A(n_2104),
.B(n_2020),
.Y(n_2267)
);

INVx2_ASAP7_75t_SL g2268 ( 
.A(n_2066),
.Y(n_2268)
);

NAND2xp5_ASAP7_75t_L g2269 ( 
.A(n_2084),
.B(n_1959),
.Y(n_2269)
);

INVx2_ASAP7_75t_SL g2270 ( 
.A(n_2066),
.Y(n_2270)
);

INVxp67_ASAP7_75t_L g2271 ( 
.A(n_2087),
.Y(n_2271)
);

AOI22xp33_ASAP7_75t_SL g2272 ( 
.A1(n_2117),
.A2(n_1897),
.B1(n_1873),
.B2(n_2007),
.Y(n_2272)
);

NAND2xp5_ASAP7_75t_L g2273 ( 
.A(n_2129),
.B(n_1959),
.Y(n_2273)
);

INVx2_ASAP7_75t_L g2274 ( 
.A(n_2059),
.Y(n_2274)
);

AND2x2_ASAP7_75t_L g2275 ( 
.A(n_2104),
.B(n_2020),
.Y(n_2275)
);

BUFx3_ASAP7_75t_L g2276 ( 
.A(n_2083),
.Y(n_2276)
);

INVx5_ASAP7_75t_SL g2277 ( 
.A(n_2136),
.Y(n_2277)
);

OR2x2_ASAP7_75t_L g2278 ( 
.A(n_2219),
.B(n_1859),
.Y(n_2278)
);

NAND3xp33_ASAP7_75t_L g2279 ( 
.A(n_2072),
.B(n_1969),
.C(n_1936),
.Y(n_2279)
);

NAND3xp33_ASAP7_75t_L g2280 ( 
.A(n_2090),
.B(n_1969),
.C(n_1936),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2081),
.Y(n_2281)
);

AND2x2_ASAP7_75t_L g2282 ( 
.A(n_2151),
.B(n_1951),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2088),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2059),
.Y(n_2284)
);

NAND3xp33_ASAP7_75t_L g2285 ( 
.A(n_2090),
.B(n_1969),
.C(n_1936),
.Y(n_2285)
);

AOI22xp33_ASAP7_75t_L g2286 ( 
.A1(n_2076),
.A2(n_1870),
.B1(n_1924),
.B2(n_1957),
.Y(n_2286)
);

BUFx2_ASAP7_75t_L g2287 ( 
.A(n_2120),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_2139),
.A2(n_2149),
.B1(n_2155),
.B2(n_2114),
.Y(n_2288)
);

AND2x4_ASAP7_75t_L g2289 ( 
.A(n_2120),
.B(n_1944),
.Y(n_2289)
);

OR2x2_ASAP7_75t_L g2290 ( 
.A(n_2062),
.B(n_2006),
.Y(n_2290)
);

AND2x2_ASAP7_75t_L g2291 ( 
.A(n_2151),
.B(n_1951),
.Y(n_2291)
);

INVx1_ASAP7_75t_L g2292 ( 
.A(n_2091),
.Y(n_2292)
);

NOR3xp33_ASAP7_75t_L g2293 ( 
.A(n_2114),
.B(n_1973),
.C(n_1945),
.Y(n_2293)
);

AOI221xp5_ASAP7_75t_L g2294 ( 
.A1(n_2145),
.A2(n_2053),
.B1(n_1977),
.B2(n_1961),
.C(n_1971),
.Y(n_2294)
);

OAI33xp33_ASAP7_75t_L g2295 ( 
.A1(n_2195),
.A2(n_1855),
.A3(n_1858),
.B1(n_1921),
.B2(n_1963),
.B3(n_1971),
.Y(n_2295)
);

NAND2xp5_ASAP7_75t_L g2296 ( 
.A(n_2132),
.B(n_2002),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2156),
.B(n_1955),
.Y(n_2297)
);

NOR2x1_ASAP7_75t_L g2298 ( 
.A(n_2083),
.B(n_2109),
.Y(n_2298)
);

NAND2xp5_ASAP7_75t_L g2299 ( 
.A(n_2152),
.B(n_2002),
.Y(n_2299)
);

NAND2xp5_ASAP7_75t_L g2300 ( 
.A(n_2141),
.B(n_2239),
.Y(n_2300)
);

INVx1_ASAP7_75t_L g2301 ( 
.A(n_2102),
.Y(n_2301)
);

AND2x2_ASAP7_75t_L g2302 ( 
.A(n_2156),
.B(n_1955),
.Y(n_2302)
);

AND2x2_ASAP7_75t_L g2303 ( 
.A(n_2156),
.B(n_1958),
.Y(n_2303)
);

AND2x2_ASAP7_75t_L g2304 ( 
.A(n_2085),
.B(n_1958),
.Y(n_2304)
);

OR2x2_ASAP7_75t_L g2305 ( 
.A(n_2174),
.B(n_1921),
.Y(n_2305)
);

BUFx2_ASAP7_75t_L g2306 ( 
.A(n_2150),
.Y(n_2306)
);

AOI31xp33_ASAP7_75t_SL g2307 ( 
.A1(n_2077),
.A2(n_1989),
.A3(n_1970),
.B(n_2050),
.Y(n_2307)
);

AOI21xp5_ASAP7_75t_L g2308 ( 
.A1(n_2123),
.A2(n_2007),
.B(n_1985),
.Y(n_2308)
);

OR2x2_ASAP7_75t_L g2309 ( 
.A(n_2199),
.B(n_1989),
.Y(n_2309)
);

BUFx6f_ASAP7_75t_L g2310 ( 
.A(n_2066),
.Y(n_2310)
);

NOR2x1_ASAP7_75t_SL g2311 ( 
.A(n_2060),
.B(n_1893),
.Y(n_2311)
);

HB1xp67_ASAP7_75t_L g2312 ( 
.A(n_2085),
.Y(n_2312)
);

NAND4xp25_ASAP7_75t_L g2313 ( 
.A(n_2139),
.B(n_2053),
.C(n_1944),
.D(n_1957),
.Y(n_2313)
);

BUFx2_ASAP7_75t_L g2314 ( 
.A(n_2150),
.Y(n_2314)
);

AND2x2_ASAP7_75t_L g2315 ( 
.A(n_2123),
.B(n_1847),
.Y(n_2315)
);

INVx1_ASAP7_75t_L g2316 ( 
.A(n_2107),
.Y(n_2316)
);

HB1xp67_ASAP7_75t_L g2317 ( 
.A(n_2060),
.Y(n_2317)
);

OAI22xp5_ASAP7_75t_L g2318 ( 
.A1(n_2149),
.A2(n_1860),
.B1(n_1893),
.B2(n_1863),
.Y(n_2318)
);

AOI221xp5_ASAP7_75t_L g2319 ( 
.A1(n_2175),
.A2(n_1963),
.B1(n_1962),
.B2(n_1957),
.C(n_1944),
.Y(n_2319)
);

OR2x2_ASAP7_75t_L g2320 ( 
.A(n_2069),
.B(n_1970),
.Y(n_2320)
);

BUFx2_ASAP7_75t_L g2321 ( 
.A(n_2150),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2067),
.A2(n_2127),
.B(n_2126),
.Y(n_2322)
);

NAND2xp5_ASAP7_75t_L g2323 ( 
.A(n_2239),
.B(n_1964),
.Y(n_2323)
);

AND2x2_ASAP7_75t_L g2324 ( 
.A(n_2183),
.B(n_1942),
.Y(n_2324)
);

INVx1_ASAP7_75t_L g2325 ( 
.A(n_2108),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_2162),
.Y(n_2326)
);

INVxp67_ASAP7_75t_SL g2327 ( 
.A(n_2200),
.Y(n_2327)
);

AND2x2_ASAP7_75t_L g2328 ( 
.A(n_2214),
.B(n_1942),
.Y(n_2328)
);

CKINVDCx5p33_ASAP7_75t_R g2329 ( 
.A(n_2109),
.Y(n_2329)
);

AOI221xp5_ASAP7_75t_L g2330 ( 
.A1(n_2173),
.A2(n_2160),
.B1(n_2225),
.B2(n_2206),
.C(n_2126),
.Y(n_2330)
);

OAI221xp5_ASAP7_75t_L g2331 ( 
.A1(n_2127),
.A2(n_1863),
.B1(n_1845),
.B2(n_1860),
.C(n_1945),
.Y(n_2331)
);

AND2x2_ASAP7_75t_L g2332 ( 
.A(n_2186),
.B(n_1948),
.Y(n_2332)
);

BUFx3_ASAP7_75t_L g2333 ( 
.A(n_2136),
.Y(n_2333)
);

INVx2_ASAP7_75t_L g2334 ( 
.A(n_2064),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2111),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_2115),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2064),
.Y(n_2337)
);

AND2x2_ASAP7_75t_L g2338 ( 
.A(n_2186),
.B(n_1948),
.Y(n_2338)
);

INVx2_ASAP7_75t_L g2339 ( 
.A(n_2075),
.Y(n_2339)
);

AND2x2_ASAP7_75t_L g2340 ( 
.A(n_2240),
.B(n_1889),
.Y(n_2340)
);

INVx2_ASAP7_75t_L g2341 ( 
.A(n_2075),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2078),
.Y(n_2342)
);

BUFx2_ASAP7_75t_L g2343 ( 
.A(n_2162),
.Y(n_2343)
);

BUFx3_ASAP7_75t_L g2344 ( 
.A(n_2136),
.Y(n_2344)
);

AND2x2_ASAP7_75t_L g2345 ( 
.A(n_2240),
.B(n_1889),
.Y(n_2345)
);

INVx1_ASAP7_75t_L g2346 ( 
.A(n_2119),
.Y(n_2346)
);

INVx1_ASAP7_75t_L g2347 ( 
.A(n_2121),
.Y(n_2347)
);

AND2x2_ASAP7_75t_L g2348 ( 
.A(n_2243),
.B(n_2017),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_L g2349 ( 
.A(n_2080),
.B(n_1964),
.Y(n_2349)
);

AND2x2_ASAP7_75t_L g2350 ( 
.A(n_2243),
.B(n_2181),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_2137),
.Y(n_2351)
);

NAND2xp5_ASAP7_75t_L g2352 ( 
.A(n_2213),
.B(n_1878),
.Y(n_2352)
);

NAND2xp5_ASAP7_75t_L g2353 ( 
.A(n_2213),
.B(n_1878),
.Y(n_2353)
);

INVx2_ASAP7_75t_L g2354 ( 
.A(n_2078),
.Y(n_2354)
);

INVx2_ASAP7_75t_L g2355 ( 
.A(n_2086),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_2181),
.B(n_2017),
.Y(n_2356)
);

HB1xp67_ASAP7_75t_L g2357 ( 
.A(n_2234),
.Y(n_2357)
);

AND2x2_ASAP7_75t_L g2358 ( 
.A(n_2172),
.B(n_1909),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_2142),
.Y(n_2359)
);

BUFx3_ASAP7_75t_L g2360 ( 
.A(n_2136),
.Y(n_2360)
);

AND2x4_ASAP7_75t_L g2361 ( 
.A(n_2162),
.B(n_1944),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2143),
.Y(n_2362)
);

OAI21x1_ASAP7_75t_L g2363 ( 
.A1(n_2146),
.A2(n_1979),
.B(n_1973),
.Y(n_2363)
);

INVx2_ASAP7_75t_L g2364 ( 
.A(n_2086),
.Y(n_2364)
);

INVx1_ASAP7_75t_L g2365 ( 
.A(n_2147),
.Y(n_2365)
);

BUFx3_ASAP7_75t_L g2366 ( 
.A(n_2122),
.Y(n_2366)
);

INVx2_ASAP7_75t_L g2367 ( 
.A(n_2089),
.Y(n_2367)
);

INVx2_ASAP7_75t_L g2368 ( 
.A(n_2089),
.Y(n_2368)
);

INVx1_ASAP7_75t_L g2369 ( 
.A(n_2167),
.Y(n_2369)
);

INVx3_ASAP7_75t_L g2370 ( 
.A(n_2176),
.Y(n_2370)
);

OR2x2_ASAP7_75t_L g2371 ( 
.A(n_2092),
.B(n_1850),
.Y(n_2371)
);

OR2x2_ASAP7_75t_L g2372 ( 
.A(n_2101),
.B(n_1850),
.Y(n_2372)
);

BUFx3_ASAP7_75t_L g2373 ( 
.A(n_2122),
.Y(n_2373)
);

OAI211xp5_ASAP7_75t_SL g2374 ( 
.A1(n_2154),
.A2(n_1962),
.B(n_2013),
.C(n_1979),
.Y(n_2374)
);

INVx1_ASAP7_75t_L g2375 ( 
.A(n_2182),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2189),
.Y(n_2376)
);

INVx2_ASAP7_75t_L g2377 ( 
.A(n_2100),
.Y(n_2377)
);

BUFx3_ASAP7_75t_L g2378 ( 
.A(n_2097),
.Y(n_2378)
);

AOI21xp5_ASAP7_75t_L g2379 ( 
.A1(n_2163),
.A2(n_1985),
.B(n_2044),
.Y(n_2379)
);

AOI22xp33_ASAP7_75t_SL g2380 ( 
.A1(n_2178),
.A2(n_2005),
.B1(n_2004),
.B2(n_1969),
.Y(n_2380)
);

BUFx6f_ASAP7_75t_L g2381 ( 
.A(n_2176),
.Y(n_2381)
);

AND2x4_ASAP7_75t_L g2382 ( 
.A(n_2171),
.B(n_1957),
.Y(n_2382)
);

INVxp67_ASAP7_75t_L g2383 ( 
.A(n_2188),
.Y(n_2383)
);

INVx3_ASAP7_75t_SL g2384 ( 
.A(n_2231),
.Y(n_2384)
);

AND4x1_ASAP7_75t_L g2385 ( 
.A(n_2155),
.B(n_2005),
.C(n_2004),
.D(n_1988),
.Y(n_2385)
);

NOR2xp67_ASAP7_75t_L g2386 ( 
.A(n_2226),
.B(n_1973),
.Y(n_2386)
);

AND2x2_ASAP7_75t_L g2387 ( 
.A(n_2172),
.B(n_1909),
.Y(n_2387)
);

OAI21xp33_ASAP7_75t_L g2388 ( 
.A1(n_2138),
.A2(n_1911),
.B(n_2022),
.Y(n_2388)
);

BUFx2_ASAP7_75t_L g2389 ( 
.A(n_2231),
.Y(n_2389)
);

NAND2xp5_ASAP7_75t_L g2390 ( 
.A(n_2188),
.B(n_1912),
.Y(n_2390)
);

INVxp67_ASAP7_75t_SL g2391 ( 
.A(n_2074),
.Y(n_2391)
);

AOI221xp5_ASAP7_75t_L g2392 ( 
.A1(n_2204),
.A2(n_2022),
.B1(n_1911),
.B2(n_1854),
.C(n_1922),
.Y(n_2392)
);

AOI22xp33_ASAP7_75t_L g2393 ( 
.A1(n_2165),
.A2(n_2022),
.B1(n_2044),
.B2(n_1988),
.Y(n_2393)
);

AND2x2_ASAP7_75t_L g2394 ( 
.A(n_2230),
.B(n_1906),
.Y(n_2394)
);

AND2x2_ASAP7_75t_L g2395 ( 
.A(n_2230),
.B(n_1906),
.Y(n_2395)
);

AO21x2_ASAP7_75t_L g2396 ( 
.A1(n_2098),
.A2(n_2218),
.B(n_2212),
.Y(n_2396)
);

BUFx2_ASAP7_75t_L g2397 ( 
.A(n_2231),
.Y(n_2397)
);

AND2x2_ASAP7_75t_L g2398 ( 
.A(n_2211),
.B(n_1905),
.Y(n_2398)
);

AND2x2_ASAP7_75t_L g2399 ( 
.A(n_2065),
.B(n_1905),
.Y(n_2399)
);

AND2x4_ASAP7_75t_L g2400 ( 
.A(n_2171),
.B(n_2022),
.Y(n_2400)
);

AND2x2_ASAP7_75t_L g2401 ( 
.A(n_2315),
.B(n_2176),
.Y(n_2401)
);

AND2x2_ASAP7_75t_L g2402 ( 
.A(n_2315),
.B(n_2231),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_2312),
.B(n_2074),
.Y(n_2403)
);

AND2x2_ASAP7_75t_L g2404 ( 
.A(n_2289),
.B(n_2226),
.Y(n_2404)
);

INVx1_ASAP7_75t_L g2405 ( 
.A(n_2244),
.Y(n_2405)
);

INVx1_ASAP7_75t_L g2406 ( 
.A(n_2244),
.Y(n_2406)
);

AND2x2_ASAP7_75t_L g2407 ( 
.A(n_2289),
.B(n_2226),
.Y(n_2407)
);

AND2x2_ASAP7_75t_L g2408 ( 
.A(n_2289),
.B(n_2238),
.Y(n_2408)
);

AND2x2_ASAP7_75t_L g2409 ( 
.A(n_2267),
.B(n_2238),
.Y(n_2409)
);

AND2x2_ASAP7_75t_L g2410 ( 
.A(n_2267),
.B(n_2238),
.Y(n_2410)
);

OR2x2_ASAP7_75t_L g2411 ( 
.A(n_2271),
.B(n_2166),
.Y(n_2411)
);

INVx1_ASAP7_75t_L g2412 ( 
.A(n_2266),
.Y(n_2412)
);

AND2x2_ASAP7_75t_L g2413 ( 
.A(n_2275),
.B(n_2128),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2249),
.Y(n_2414)
);

AND2x2_ASAP7_75t_L g2415 ( 
.A(n_2275),
.B(n_2133),
.Y(n_2415)
);

AND2x2_ASAP7_75t_L g2416 ( 
.A(n_2304),
.B(n_2163),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_2396),
.Y(n_2417)
);

INVx2_ASAP7_75t_L g2418 ( 
.A(n_2396),
.Y(n_2418)
);

INVx1_ASAP7_75t_L g2419 ( 
.A(n_2266),
.Y(n_2419)
);

NAND2xp5_ASAP7_75t_L g2420 ( 
.A(n_2260),
.B(n_2203),
.Y(n_2420)
);

INVx1_ASAP7_75t_SL g2421 ( 
.A(n_2329),
.Y(n_2421)
);

NAND2x1_ASAP7_75t_SL g2422 ( 
.A(n_2298),
.B(n_2157),
.Y(n_2422)
);

INVxp67_ASAP7_75t_L g2423 ( 
.A(n_2357),
.Y(n_2423)
);

INVx2_ASAP7_75t_L g2424 ( 
.A(n_2396),
.Y(n_2424)
);

NAND2xp5_ASAP7_75t_L g2425 ( 
.A(n_2383),
.B(n_2177),
.Y(n_2425)
);

OR2x2_ASAP7_75t_L g2426 ( 
.A(n_2290),
.B(n_2135),
.Y(n_2426)
);

AND2x2_ASAP7_75t_L g2427 ( 
.A(n_2304),
.B(n_1912),
.Y(n_2427)
);

AND2x2_ASAP7_75t_L g2428 ( 
.A(n_2380),
.B(n_2094),
.Y(n_2428)
);

AND2x2_ASAP7_75t_L g2429 ( 
.A(n_2246),
.B(n_2094),
.Y(n_2429)
);

INVx2_ASAP7_75t_L g2430 ( 
.A(n_2381),
.Y(n_2430)
);

INVx1_ASAP7_75t_L g2431 ( 
.A(n_2281),
.Y(n_2431)
);

NAND2xp5_ASAP7_75t_L g2432 ( 
.A(n_2276),
.B(n_2170),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2276),
.B(n_2229),
.Y(n_2433)
);

NAND2xp5_ASAP7_75t_L g2434 ( 
.A(n_2327),
.B(n_2192),
.Y(n_2434)
);

INVx1_ASAP7_75t_L g2435 ( 
.A(n_2281),
.Y(n_2435)
);

AND2x2_ASAP7_75t_L g2436 ( 
.A(n_2246),
.B(n_2094),
.Y(n_2436)
);

INVx1_ASAP7_75t_SL g2437 ( 
.A(n_2329),
.Y(n_2437)
);

AND2x4_ASAP7_75t_L g2438 ( 
.A(n_2254),
.B(n_2185),
.Y(n_2438)
);

INVx2_ASAP7_75t_L g2439 ( 
.A(n_2381),
.Y(n_2439)
);

AND2x2_ASAP7_75t_L g2440 ( 
.A(n_2250),
.B(n_2134),
.Y(n_2440)
);

AOI221xp5_ASAP7_75t_L g2441 ( 
.A1(n_2252),
.A2(n_2263),
.B1(n_2288),
.B2(n_2279),
.C(n_2295),
.Y(n_2441)
);

AND2x2_ASAP7_75t_L g2442 ( 
.A(n_2250),
.B(n_2110),
.Y(n_2442)
);

NAND2xp5_ASAP7_75t_L g2443 ( 
.A(n_2268),
.B(n_2193),
.Y(n_2443)
);

NAND2xp5_ASAP7_75t_L g2444 ( 
.A(n_2268),
.B(n_2194),
.Y(n_2444)
);

OR2x2_ASAP7_75t_L g2445 ( 
.A(n_2290),
.B(n_2196),
.Y(n_2445)
);

INVx2_ASAP7_75t_L g2446 ( 
.A(n_2381),
.Y(n_2446)
);

INVx2_ASAP7_75t_L g2447 ( 
.A(n_2381),
.Y(n_2447)
);

NAND2xp5_ASAP7_75t_L g2448 ( 
.A(n_2270),
.B(n_2197),
.Y(n_2448)
);

INVx1_ASAP7_75t_L g2449 ( 
.A(n_2283),
.Y(n_2449)
);

AND2x2_ASAP7_75t_L g2450 ( 
.A(n_2297),
.B(n_2302),
.Y(n_2450)
);

INVxp67_ASAP7_75t_L g2451 ( 
.A(n_2391),
.Y(n_2451)
);

AND2x4_ASAP7_75t_L g2452 ( 
.A(n_2254),
.B(n_2287),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_2283),
.Y(n_2453)
);

NAND2xp5_ASAP7_75t_L g2454 ( 
.A(n_2270),
.B(n_2198),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2278),
.B(n_2201),
.Y(n_2455)
);

INVx2_ASAP7_75t_L g2456 ( 
.A(n_2381),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_L g2457 ( 
.A(n_2248),
.B(n_2205),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2292),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_2286),
.B(n_2210),
.Y(n_2459)
);

AOI22xp5_ASAP7_75t_L g2460 ( 
.A1(n_2280),
.A2(n_2185),
.B1(n_2164),
.B2(n_2096),
.Y(n_2460)
);

AND2x2_ASAP7_75t_L g2461 ( 
.A(n_2297),
.B(n_1993),
.Y(n_2461)
);

INVx1_ASAP7_75t_L g2462 ( 
.A(n_2292),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2306),
.Y(n_2463)
);

AND2x2_ASAP7_75t_L g2464 ( 
.A(n_2302),
.B(n_1993),
.Y(n_2464)
);

AOI22xp33_ASAP7_75t_L g2465 ( 
.A1(n_2285),
.A2(n_2187),
.B1(n_2118),
.B2(n_2044),
.Y(n_2465)
);

AND2x2_ASAP7_75t_L g2466 ( 
.A(n_2303),
.B(n_1996),
.Y(n_2466)
);

INVx1_ASAP7_75t_L g2467 ( 
.A(n_2301),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2378),
.B(n_2221),
.Y(n_2468)
);

INVxp67_ASAP7_75t_SL g2469 ( 
.A(n_2311),
.Y(n_2469)
);

OR2x2_ASAP7_75t_L g2470 ( 
.A(n_2278),
.B(n_2235),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2378),
.Y(n_2471)
);

AND2x2_ASAP7_75t_L g2472 ( 
.A(n_2303),
.B(n_2282),
.Y(n_2472)
);

INVx2_ASAP7_75t_L g2473 ( 
.A(n_2306),
.Y(n_2473)
);

OR2x2_ASAP7_75t_L g2474 ( 
.A(n_2309),
.B(n_2237),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_2301),
.Y(n_2475)
);

CKINVDCx20_ASAP7_75t_R g2476 ( 
.A(n_2366),
.Y(n_2476)
);

AND2x2_ASAP7_75t_L g2477 ( 
.A(n_2282),
.B(n_1996),
.Y(n_2477)
);

OR2x2_ASAP7_75t_L g2478 ( 
.A(n_2309),
.B(n_2241),
.Y(n_2478)
);

NAND2xp5_ASAP7_75t_L g2479 ( 
.A(n_2333),
.B(n_2242),
.Y(n_2479)
);

AND2x2_ASAP7_75t_L g2480 ( 
.A(n_2291),
.B(n_1849),
.Y(n_2480)
);

AND2x2_ASAP7_75t_L g2481 ( 
.A(n_2291),
.B(n_1849),
.Y(n_2481)
);

AND2x2_ASAP7_75t_L g2482 ( 
.A(n_2384),
.B(n_1865),
.Y(n_2482)
);

OAI21xp5_ASAP7_75t_L g2483 ( 
.A1(n_2322),
.A2(n_2217),
.B(n_2187),
.Y(n_2483)
);

NAND2xp5_ASAP7_75t_L g2484 ( 
.A(n_2333),
.B(n_2227),
.Y(n_2484)
);

OR2x2_ASAP7_75t_L g2485 ( 
.A(n_2305),
.B(n_2098),
.Y(n_2485)
);

OR2x2_ASAP7_75t_L g2486 ( 
.A(n_2305),
.B(n_2184),
.Y(n_2486)
);

NAND2xp5_ASAP7_75t_L g2487 ( 
.A(n_2344),
.B(n_2061),
.Y(n_2487)
);

BUFx2_ASAP7_75t_L g2488 ( 
.A(n_2287),
.Y(n_2488)
);

AND2x2_ASAP7_75t_L g2489 ( 
.A(n_2384),
.B(n_1865),
.Y(n_2489)
);

AND2x2_ASAP7_75t_L g2490 ( 
.A(n_2382),
.B(n_1975),
.Y(n_2490)
);

NAND3xp33_ASAP7_75t_L g2491 ( 
.A(n_2264),
.B(n_2215),
.C(n_2228),
.Y(n_2491)
);

OR2x2_ASAP7_75t_L g2492 ( 
.A(n_2320),
.B(n_2153),
.Y(n_2492)
);

NOR2x1p5_ASAP7_75t_L g2493 ( 
.A(n_2247),
.B(n_2180),
.Y(n_2493)
);

AND2x2_ASAP7_75t_L g2494 ( 
.A(n_2382),
.B(n_1975),
.Y(n_2494)
);

NAND2xp5_ASAP7_75t_L g2495 ( 
.A(n_2344),
.B(n_2216),
.Y(n_2495)
);

INVxp67_ASAP7_75t_SL g2496 ( 
.A(n_2311),
.Y(n_2496)
);

OR2x2_ASAP7_75t_L g2497 ( 
.A(n_2320),
.B(n_2207),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2314),
.Y(n_2498)
);

OR2x4_ASAP7_75t_L g2499 ( 
.A(n_2310),
.B(n_2099),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2325),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_2325),
.Y(n_2501)
);

AND2x2_ASAP7_75t_L g2502 ( 
.A(n_2382),
.B(n_2116),
.Y(n_2502)
);

INVx1_ASAP7_75t_L g2503 ( 
.A(n_2335),
.Y(n_2503)
);

AND2x2_ASAP7_75t_L g2504 ( 
.A(n_2400),
.B(n_2116),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2335),
.Y(n_2505)
);

AND2x2_ASAP7_75t_L g2506 ( 
.A(n_2400),
.B(n_2324),
.Y(n_2506)
);

INVx1_ASAP7_75t_L g2507 ( 
.A(n_2336),
.Y(n_2507)
);

AND2x2_ASAP7_75t_L g2508 ( 
.A(n_2400),
.B(n_2116),
.Y(n_2508)
);

AND2x4_ASAP7_75t_L g2509 ( 
.A(n_2262),
.B(n_2258),
.Y(n_2509)
);

AND2x2_ASAP7_75t_L g2510 ( 
.A(n_2324),
.B(n_2116),
.Y(n_2510)
);

NAND2xp5_ASAP7_75t_SL g2511 ( 
.A(n_2259),
.B(n_2209),
.Y(n_2511)
);

NAND2xp5_ASAP7_75t_L g2512 ( 
.A(n_2360),
.B(n_2233),
.Y(n_2512)
);

INVxp67_ASAP7_75t_L g2513 ( 
.A(n_2310),
.Y(n_2513)
);

INVx2_ASAP7_75t_L g2514 ( 
.A(n_2314),
.Y(n_2514)
);

INVx1_ASAP7_75t_L g2515 ( 
.A(n_2336),
.Y(n_2515)
);

OR2x2_ASAP7_75t_L g2516 ( 
.A(n_2350),
.B(n_2223),
.Y(n_2516)
);

NAND2xp5_ASAP7_75t_L g2517 ( 
.A(n_2360),
.B(n_2300),
.Y(n_2517)
);

INVx3_ASAP7_75t_L g2518 ( 
.A(n_2262),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2328),
.B(n_2130),
.Y(n_2519)
);

INVx1_ASAP7_75t_L g2520 ( 
.A(n_2346),
.Y(n_2520)
);

INVx1_ASAP7_75t_SL g2521 ( 
.A(n_2259),
.Y(n_2521)
);

INVx3_ASAP7_75t_L g2522 ( 
.A(n_2262),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2346),
.Y(n_2523)
);

INVx2_ASAP7_75t_L g2524 ( 
.A(n_2321),
.Y(n_2524)
);

AND2x2_ASAP7_75t_L g2525 ( 
.A(n_2328),
.B(n_2130),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2255),
.B(n_2130),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2255),
.B(n_2130),
.Y(n_2527)
);

BUFx2_ASAP7_75t_L g2528 ( 
.A(n_2321),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_L g2529 ( 
.A(n_2366),
.B(n_1922),
.Y(n_2529)
);

AND2x4_ASAP7_75t_L g2530 ( 
.A(n_2258),
.B(n_2168),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_L g2531 ( 
.A(n_2373),
.B(n_2000),
.Y(n_2531)
);

INVx1_ASAP7_75t_L g2532 ( 
.A(n_2347),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2528),
.Y(n_2533)
);

INVx2_ASAP7_75t_L g2534 ( 
.A(n_2488),
.Y(n_2534)
);

INVxp67_ASAP7_75t_SL g2535 ( 
.A(n_2422),
.Y(n_2535)
);

INVx3_ASAP7_75t_L g2536 ( 
.A(n_2452),
.Y(n_2536)
);

INVx1_ASAP7_75t_L g2537 ( 
.A(n_2528),
.Y(n_2537)
);

OAI21xp33_ASAP7_75t_L g2538 ( 
.A1(n_2441),
.A2(n_2256),
.B(n_2330),
.Y(n_2538)
);

NAND2xp5_ASAP7_75t_L g2539 ( 
.A(n_2521),
.B(n_2373),
.Y(n_2539)
);

AND2x2_ASAP7_75t_L g2540 ( 
.A(n_2450),
.B(n_2293),
.Y(n_2540)
);

OR2x2_ASAP7_75t_L g2541 ( 
.A(n_2434),
.B(n_2350),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_2488),
.Y(n_2542)
);

OAI32xp33_ASAP7_75t_L g2543 ( 
.A1(n_2432),
.A2(n_2317),
.A3(n_2245),
.B1(n_2331),
.B2(n_2313),
.Y(n_2543)
);

OAI21xp33_ASAP7_75t_L g2544 ( 
.A1(n_2483),
.A2(n_2388),
.B(n_2294),
.Y(n_2544)
);

INVx2_ASAP7_75t_L g2545 ( 
.A(n_2452),
.Y(n_2545)
);

AND2x2_ASAP7_75t_L g2546 ( 
.A(n_2450),
.B(n_2472),
.Y(n_2546)
);

NAND2x1_ASAP7_75t_L g2547 ( 
.A(n_2438),
.B(n_2326),
.Y(n_2547)
);

NOR2xp33_ASAP7_75t_L g2548 ( 
.A(n_2421),
.B(n_2385),
.Y(n_2548)
);

NAND2xp5_ASAP7_75t_L g2549 ( 
.A(n_2414),
.B(n_2310),
.Y(n_2549)
);

NAND2xp5_ASAP7_75t_L g2550 ( 
.A(n_2423),
.B(n_2310),
.Y(n_2550)
);

INVx1_ASAP7_75t_L g2551 ( 
.A(n_2419),
.Y(n_2551)
);

INVx2_ASAP7_75t_L g2552 ( 
.A(n_2452),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2419),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2431),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2472),
.B(n_2389),
.Y(n_2555)
);

HB1xp67_ASAP7_75t_L g2556 ( 
.A(n_2471),
.Y(n_2556)
);

AND2x2_ASAP7_75t_L g2557 ( 
.A(n_2402),
.B(n_2389),
.Y(n_2557)
);

OAI22xp33_ASAP7_75t_L g2558 ( 
.A1(n_2460),
.A2(n_2318),
.B1(n_2308),
.B2(n_2319),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2431),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_2516),
.B(n_2463),
.Y(n_2560)
);

OR2x2_ASAP7_75t_L g2561 ( 
.A(n_2516),
.B(n_2347),
.Y(n_2561)
);

INVx2_ASAP7_75t_L g2562 ( 
.A(n_2471),
.Y(n_2562)
);

BUFx2_ASAP7_75t_L g2563 ( 
.A(n_2499),
.Y(n_2563)
);

INVx2_ASAP7_75t_L g2564 ( 
.A(n_2476),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2435),
.Y(n_2565)
);

NOR3xp33_ASAP7_75t_L g2566 ( 
.A(n_2511),
.B(n_2397),
.C(n_2272),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2435),
.Y(n_2567)
);

HB1xp67_ASAP7_75t_L g2568 ( 
.A(n_2463),
.Y(n_2568)
);

HB1xp67_ASAP7_75t_L g2569 ( 
.A(n_2473),
.Y(n_2569)
);

NAND2xp5_ASAP7_75t_L g2570 ( 
.A(n_2437),
.B(n_2310),
.Y(n_2570)
);

INVx2_ASAP7_75t_SL g2571 ( 
.A(n_2499),
.Y(n_2571)
);

INVx1_ASAP7_75t_L g2572 ( 
.A(n_2449),
.Y(n_2572)
);

OAI21xp33_ASAP7_75t_L g2573 ( 
.A1(n_2420),
.A2(n_2392),
.B(n_2393),
.Y(n_2573)
);

OR2x2_ASAP7_75t_L g2574 ( 
.A(n_2473),
.B(n_2351),
.Y(n_2574)
);

INVx1_ASAP7_75t_L g2575 ( 
.A(n_2449),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2453),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2453),
.Y(n_2577)
);

NAND2xp5_ASAP7_75t_L g2578 ( 
.A(n_2451),
.B(n_2397),
.Y(n_2578)
);

NOR2x1_ASAP7_75t_L g2579 ( 
.A(n_2476),
.B(n_2326),
.Y(n_2579)
);

INVx1_ASAP7_75t_L g2580 ( 
.A(n_2458),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2458),
.Y(n_2581)
);

INVx2_ASAP7_75t_L g2582 ( 
.A(n_2518),
.Y(n_2582)
);

HB1xp67_ASAP7_75t_L g2583 ( 
.A(n_2498),
.Y(n_2583)
);

INVx1_ASAP7_75t_L g2584 ( 
.A(n_2462),
.Y(n_2584)
);

AND2x2_ASAP7_75t_L g2585 ( 
.A(n_2402),
.B(n_2257),
.Y(n_2585)
);

NAND2xp5_ASAP7_75t_L g2586 ( 
.A(n_2401),
.B(n_2257),
.Y(n_2586)
);

INVx1_ASAP7_75t_L g2587 ( 
.A(n_2462),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2401),
.B(n_2517),
.Y(n_2588)
);

AND2x2_ASAP7_75t_L g2589 ( 
.A(n_2506),
.B(n_2361),
.Y(n_2589)
);

INVx1_ASAP7_75t_L g2590 ( 
.A(n_2467),
.Y(n_2590)
);

INVx2_ASAP7_75t_L g2591 ( 
.A(n_2518),
.Y(n_2591)
);

INVx1_ASAP7_75t_L g2592 ( 
.A(n_2467),
.Y(n_2592)
);

INVx1_ASAP7_75t_L g2593 ( 
.A(n_2500),
.Y(n_2593)
);

INVxp67_ASAP7_75t_SL g2594 ( 
.A(n_2422),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2500),
.Y(n_2595)
);

AOI32xp33_ASAP7_75t_L g2596 ( 
.A1(n_2428),
.A2(n_2374),
.A3(n_2343),
.B1(n_2361),
.B2(n_2387),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2491),
.A2(n_2277),
.B1(n_2379),
.B2(n_2361),
.Y(n_2597)
);

NAND2xp5_ASAP7_75t_L g2598 ( 
.A(n_2498),
.B(n_2253),
.Y(n_2598)
);

AND2x2_ASAP7_75t_L g2599 ( 
.A(n_2506),
.B(n_2277),
.Y(n_2599)
);

NAND2xp5_ASAP7_75t_SL g2600 ( 
.A(n_2428),
.B(n_2277),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2404),
.B(n_2277),
.Y(n_2601)
);

AND2x2_ASAP7_75t_L g2602 ( 
.A(n_2404),
.B(n_2370),
.Y(n_2602)
);

AND2x2_ASAP7_75t_L g2603 ( 
.A(n_2407),
.B(n_2370),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2514),
.B(n_2390),
.Y(n_2604)
);

NAND2xp5_ASAP7_75t_L g2605 ( 
.A(n_2514),
.B(n_2340),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2407),
.B(n_2370),
.Y(n_2606)
);

INVxp67_ASAP7_75t_L g2607 ( 
.A(n_2438),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2501),
.Y(n_2608)
);

AND2x2_ASAP7_75t_L g2609 ( 
.A(n_2408),
.B(n_2343),
.Y(n_2609)
);

HB1xp67_ASAP7_75t_L g2610 ( 
.A(n_2524),
.Y(n_2610)
);

INVx2_ASAP7_75t_L g2611 ( 
.A(n_2518),
.Y(n_2611)
);

NAND2xp5_ASAP7_75t_L g2612 ( 
.A(n_2524),
.B(n_2340),
.Y(n_2612)
);

AND2x4_ASAP7_75t_L g2613 ( 
.A(n_2509),
.B(n_2258),
.Y(n_2613)
);

NAND3xp33_ASAP7_75t_L g2614 ( 
.A(n_2465),
.B(n_2425),
.C(n_2495),
.Y(n_2614)
);

AND2x2_ASAP7_75t_L g2615 ( 
.A(n_2408),
.B(n_2345),
.Y(n_2615)
);

AND2x2_ASAP7_75t_L g2616 ( 
.A(n_2427),
.B(n_2345),
.Y(n_2616)
);

INVx2_ASAP7_75t_L g2617 ( 
.A(n_2522),
.Y(n_2617)
);

INVx1_ASAP7_75t_L g2618 ( 
.A(n_2501),
.Y(n_2618)
);

INVx1_ASAP7_75t_L g2619 ( 
.A(n_2503),
.Y(n_2619)
);

INVx1_ASAP7_75t_L g2620 ( 
.A(n_2503),
.Y(n_2620)
);

OR2x2_ASAP7_75t_L g2621 ( 
.A(n_2455),
.B(n_2351),
.Y(n_2621)
);

INVx2_ASAP7_75t_L g2622 ( 
.A(n_2522),
.Y(n_2622)
);

INVx1_ASAP7_75t_L g2623 ( 
.A(n_2505),
.Y(n_2623)
);

NAND2xp5_ASAP7_75t_L g2624 ( 
.A(n_2438),
.B(n_2352),
.Y(n_2624)
);

BUFx2_ASAP7_75t_L g2625 ( 
.A(n_2499),
.Y(n_2625)
);

AND2x2_ASAP7_75t_L g2626 ( 
.A(n_2427),
.B(n_2332),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2505),
.Y(n_2627)
);

NAND2xp5_ASAP7_75t_L g2628 ( 
.A(n_2513),
.B(n_2353),
.Y(n_2628)
);

OR2x2_ASAP7_75t_L g2629 ( 
.A(n_2455),
.B(n_2359),
.Y(n_2629)
);

HB1xp67_ASAP7_75t_L g2630 ( 
.A(n_2522),
.Y(n_2630)
);

OR2x2_ASAP7_75t_L g2631 ( 
.A(n_2470),
.B(n_2359),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2507),
.Y(n_2632)
);

INVx1_ASAP7_75t_L g2633 ( 
.A(n_2507),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2515),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2416),
.B(n_2332),
.Y(n_2635)
);

INVx1_ASAP7_75t_L g2636 ( 
.A(n_2515),
.Y(n_2636)
);

OR2x2_ASAP7_75t_L g2637 ( 
.A(n_2470),
.B(n_2362),
.Y(n_2637)
);

AND2x2_ASAP7_75t_L g2638 ( 
.A(n_2416),
.B(n_2415),
.Y(n_2638)
);

INVx1_ASAP7_75t_L g2639 ( 
.A(n_2520),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2520),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2430),
.Y(n_2641)
);

AND2x2_ASAP7_75t_L g2642 ( 
.A(n_2415),
.B(n_2493),
.Y(n_2642)
);

AOI222xp33_ASAP7_75t_L g2643 ( 
.A1(n_2457),
.A2(n_2307),
.B1(n_2296),
.B2(n_2299),
.C1(n_2269),
.C2(n_2273),
.Y(n_2643)
);

BUFx3_ASAP7_75t_L g2644 ( 
.A(n_2509),
.Y(n_2644)
);

AND2x4_ASAP7_75t_L g2645 ( 
.A(n_2509),
.B(n_2258),
.Y(n_2645)
);

NAND2xp5_ASAP7_75t_L g2646 ( 
.A(n_2468),
.B(n_2398),
.Y(n_2646)
);

NOR2x1_ASAP7_75t_L g2647 ( 
.A(n_2430),
.B(n_2386),
.Y(n_2647)
);

INVx2_ASAP7_75t_L g2648 ( 
.A(n_2530),
.Y(n_2648)
);

INVx2_ASAP7_75t_L g2649 ( 
.A(n_2530),
.Y(n_2649)
);

INVx1_ASAP7_75t_L g2650 ( 
.A(n_2523),
.Y(n_2650)
);

OR2x2_ASAP7_75t_L g2651 ( 
.A(n_2445),
.B(n_2362),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2523),
.Y(n_2652)
);

INVx1_ASAP7_75t_L g2653 ( 
.A(n_2532),
.Y(n_2653)
);

AND2x2_ASAP7_75t_L g2654 ( 
.A(n_2482),
.B(n_2338),
.Y(n_2654)
);

AND2x2_ASAP7_75t_L g2655 ( 
.A(n_2482),
.B(n_2338),
.Y(n_2655)
);

INVx2_ASAP7_75t_L g2656 ( 
.A(n_2530),
.Y(n_2656)
);

AND2x2_ASAP7_75t_L g2657 ( 
.A(n_2489),
.B(n_2348),
.Y(n_2657)
);

AND2x4_ASAP7_75t_L g2658 ( 
.A(n_2439),
.B(n_2446),
.Y(n_2658)
);

NAND2xp5_ASAP7_75t_SL g2659 ( 
.A(n_2538),
.B(n_2469),
.Y(n_2659)
);

AND2x2_ASAP7_75t_L g2660 ( 
.A(n_2564),
.B(n_2489),
.Y(n_2660)
);

INVx2_ASAP7_75t_L g2661 ( 
.A(n_2536),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2564),
.B(n_2403),
.Y(n_2662)
);

INVx2_ASAP7_75t_L g2663 ( 
.A(n_2536),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2638),
.B(n_2409),
.Y(n_2664)
);

AND2x2_ASAP7_75t_L g2665 ( 
.A(n_2638),
.B(n_2409),
.Y(n_2665)
);

INVx2_ASAP7_75t_SL g2666 ( 
.A(n_2536),
.Y(n_2666)
);

INVx1_ASAP7_75t_L g2667 ( 
.A(n_2534),
.Y(n_2667)
);

NOR2x1p5_ASAP7_75t_L g2668 ( 
.A(n_2539),
.B(n_2487),
.Y(n_2668)
);

NOR2xp33_ASAP7_75t_L g2669 ( 
.A(n_2556),
.B(n_2459),
.Y(n_2669)
);

INVx2_ASAP7_75t_L g2670 ( 
.A(n_2547),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2534),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2542),
.Y(n_2672)
);

INVxp67_ASAP7_75t_SL g2673 ( 
.A(n_2579),
.Y(n_2673)
);

OR2x2_ASAP7_75t_L g2674 ( 
.A(n_2541),
.B(n_2411),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2542),
.Y(n_2675)
);

NAND2xp5_ASAP7_75t_L g2676 ( 
.A(n_2607),
.B(n_2479),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2568),
.Y(n_2677)
);

INVx1_ASAP7_75t_L g2678 ( 
.A(n_2569),
.Y(n_2678)
);

INVx1_ASAP7_75t_L g2679 ( 
.A(n_2583),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2546),
.B(n_2410),
.Y(n_2680)
);

AND2x2_ASAP7_75t_L g2681 ( 
.A(n_2546),
.B(n_2410),
.Y(n_2681)
);

OR2x2_ASAP7_75t_L g2682 ( 
.A(n_2541),
.B(n_2411),
.Y(n_2682)
);

INVxp67_ASAP7_75t_L g2683 ( 
.A(n_2563),
.Y(n_2683)
);

BUFx2_ASAP7_75t_L g2684 ( 
.A(n_2644),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2585),
.B(n_2442),
.Y(n_2685)
);

NOR2x1p5_ASAP7_75t_L g2686 ( 
.A(n_2570),
.B(n_2433),
.Y(n_2686)
);

AOI22xp5_ASAP7_75t_L g2687 ( 
.A1(n_2544),
.A2(n_2484),
.B1(n_2442),
.B2(n_2496),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2610),
.Y(n_2688)
);

NAND2xp5_ASAP7_75t_SL g2689 ( 
.A(n_2558),
.B(n_2258),
.Y(n_2689)
);

AND2x2_ASAP7_75t_L g2690 ( 
.A(n_2585),
.B(n_2413),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2547),
.Y(n_2691)
);

INVx3_ASAP7_75t_L g2692 ( 
.A(n_2644),
.Y(n_2692)
);

NAND2xp5_ASAP7_75t_L g2693 ( 
.A(n_2562),
.B(n_2439),
.Y(n_2693)
);

INVx2_ASAP7_75t_L g2694 ( 
.A(n_2545),
.Y(n_2694)
);

INVx2_ASAP7_75t_L g2695 ( 
.A(n_2545),
.Y(n_2695)
);

INVx1_ASAP7_75t_L g2696 ( 
.A(n_2560),
.Y(n_2696)
);

INVx1_ASAP7_75t_L g2697 ( 
.A(n_2560),
.Y(n_2697)
);

INVx1_ASAP7_75t_L g2698 ( 
.A(n_2537),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2557),
.B(n_2413),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2537),
.Y(n_2700)
);

NAND2xp5_ASAP7_75t_L g2701 ( 
.A(n_2562),
.B(n_2446),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2574),
.Y(n_2702)
);

NAND2xp5_ASAP7_75t_SL g2703 ( 
.A(n_2596),
.B(n_2447),
.Y(n_2703)
);

AOI221xp5_ASAP7_75t_L g2704 ( 
.A1(n_2543),
.A2(n_2614),
.B1(n_2573),
.B2(n_2566),
.C(n_2594),
.Y(n_2704)
);

NAND2xp5_ASAP7_75t_L g2705 ( 
.A(n_2552),
.B(n_2447),
.Y(n_2705)
);

INVx1_ASAP7_75t_L g2706 ( 
.A(n_2574),
.Y(n_2706)
);

NAND2xp5_ASAP7_75t_L g2707 ( 
.A(n_2552),
.B(n_2456),
.Y(n_2707)
);

INVx1_ASAP7_75t_L g2708 ( 
.A(n_2641),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2533),
.B(n_2474),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2587),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2557),
.B(n_2490),
.Y(n_2711)
);

OAI33xp33_ASAP7_75t_L g2712 ( 
.A1(n_2578),
.A2(n_2550),
.A3(n_2598),
.B1(n_2549),
.B2(n_2588),
.B3(n_2604),
.Y(n_2712)
);

NOR2xp33_ASAP7_75t_L g2713 ( 
.A(n_2548),
.B(n_2512),
.Y(n_2713)
);

AND2x2_ASAP7_75t_L g2714 ( 
.A(n_2635),
.B(n_2490),
.Y(n_2714)
);

INVx1_ASAP7_75t_SL g2715 ( 
.A(n_2555),
.Y(n_2715)
);

CKINVDCx16_ASAP7_75t_R g2716 ( 
.A(n_2599),
.Y(n_2716)
);

AND2x2_ASAP7_75t_L g2717 ( 
.A(n_2635),
.B(n_2494),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2587),
.Y(n_2718)
);

NAND2xp5_ASAP7_75t_L g2719 ( 
.A(n_2571),
.B(n_2456),
.Y(n_2719)
);

NAND2xp5_ASAP7_75t_L g2720 ( 
.A(n_2571),
.B(n_2555),
.Y(n_2720)
);

HB1xp67_ASAP7_75t_L g2721 ( 
.A(n_2630),
.Y(n_2721)
);

INVx2_ASAP7_75t_L g2722 ( 
.A(n_2589),
.Y(n_2722)
);

INVx3_ASAP7_75t_SL g2723 ( 
.A(n_2613),
.Y(n_2723)
);

OAI33xp33_ASAP7_75t_L g2724 ( 
.A1(n_2624),
.A2(n_2405),
.A3(n_2406),
.B1(n_2412),
.B2(n_2475),
.B3(n_2532),
.Y(n_2724)
);

INVx2_ASAP7_75t_L g2725 ( 
.A(n_2589),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2623),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2623),
.Y(n_2727)
);

NAND2xp5_ASAP7_75t_L g2728 ( 
.A(n_2563),
.B(n_2443),
.Y(n_2728)
);

NAND2xp5_ASAP7_75t_L g2729 ( 
.A(n_2625),
.B(n_2609),
.Y(n_2729)
);

INVx2_ASAP7_75t_L g2730 ( 
.A(n_2609),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2621),
.Y(n_2731)
);

OR2x2_ASAP7_75t_L g2732 ( 
.A(n_2605),
.B(n_2426),
.Y(n_2732)
);

OR2x2_ASAP7_75t_L g2733 ( 
.A(n_2612),
.B(n_2646),
.Y(n_2733)
);

INVx2_ASAP7_75t_L g2734 ( 
.A(n_2615),
.Y(n_2734)
);

INVx1_ASAP7_75t_L g2735 ( 
.A(n_2621),
.Y(n_2735)
);

AND2x4_ASAP7_75t_L g2736 ( 
.A(n_2613),
.B(n_2645),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2629),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2629),
.Y(n_2738)
);

OR2x2_ASAP7_75t_L g2739 ( 
.A(n_2561),
.B(n_2474),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2599),
.B(n_2494),
.Y(n_2740)
);

INVx1_ASAP7_75t_L g2741 ( 
.A(n_2631),
.Y(n_2741)
);

NAND2xp5_ASAP7_75t_L g2742 ( 
.A(n_2625),
.B(n_2444),
.Y(n_2742)
);

INVx2_ASAP7_75t_L g2743 ( 
.A(n_2615),
.Y(n_2743)
);

OA21x2_ASAP7_75t_L g2744 ( 
.A1(n_2535),
.A2(n_2418),
.B(n_2417),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2631),
.Y(n_2745)
);

AOI22xp33_ASAP7_75t_L g2746 ( 
.A1(n_2643),
.A2(n_2440),
.B1(n_2504),
.B2(n_2502),
.Y(n_2746)
);

NAND2xp5_ASAP7_75t_L g2747 ( 
.A(n_2586),
.B(n_2448),
.Y(n_2747)
);

NAND2xp5_ASAP7_75t_L g2748 ( 
.A(n_2540),
.B(n_2454),
.Y(n_2748)
);

CKINVDCx16_ASAP7_75t_R g2749 ( 
.A(n_2601),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2637),
.Y(n_2750)
);

INVx2_ASAP7_75t_L g2751 ( 
.A(n_2657),
.Y(n_2751)
);

AND2x2_ASAP7_75t_L g2752 ( 
.A(n_2601),
.B(n_2440),
.Y(n_2752)
);

AND2x2_ASAP7_75t_L g2753 ( 
.A(n_2642),
.B(n_2480),
.Y(n_2753)
);

NOR2xp33_ASAP7_75t_L g2754 ( 
.A(n_2543),
.B(n_2531),
.Y(n_2754)
);

OAI21x1_ASAP7_75t_L g2755 ( 
.A1(n_2647),
.A2(n_2363),
.B(n_2485),
.Y(n_2755)
);

HB1xp67_ASAP7_75t_L g2756 ( 
.A(n_2582),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2637),
.Y(n_2757)
);

AND2x2_ASAP7_75t_L g2758 ( 
.A(n_2642),
.B(n_2480),
.Y(n_2758)
);

INVx1_ASAP7_75t_SL g2759 ( 
.A(n_2540),
.Y(n_2759)
);

AOI221xp5_ASAP7_75t_L g2760 ( 
.A1(n_2600),
.A2(n_2597),
.B1(n_2628),
.B2(n_2554),
.C(n_2559),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2651),
.Y(n_2761)
);

INVx2_ASAP7_75t_L g2762 ( 
.A(n_2657),
.Y(n_2762)
);

AND2x4_ASAP7_75t_L g2763 ( 
.A(n_2613),
.B(n_2645),
.Y(n_2763)
);

INVx1_ASAP7_75t_L g2764 ( 
.A(n_2651),
.Y(n_2764)
);

INVx1_ASAP7_75t_L g2765 ( 
.A(n_2551),
.Y(n_2765)
);

NAND3xp33_ASAP7_75t_L g2766 ( 
.A(n_2600),
.B(n_2485),
.C(n_2478),
.Y(n_2766)
);

NAND4xp25_ASAP7_75t_SL g2767 ( 
.A(n_2616),
.B(n_2504),
.C(n_2508),
.D(n_2502),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2553),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2565),
.Y(n_2769)
);

INVx2_ASAP7_75t_L g2770 ( 
.A(n_2654),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2602),
.B(n_2481),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2561),
.B(n_2478),
.Y(n_2772)
);

NAND2xp5_ASAP7_75t_L g2773 ( 
.A(n_2715),
.B(n_2582),
.Y(n_2773)
);

NAND2xp5_ASAP7_75t_L g2774 ( 
.A(n_2660),
.B(n_2591),
.Y(n_2774)
);

NAND2xp5_ASAP7_75t_SL g2775 ( 
.A(n_2704),
.B(n_2645),
.Y(n_2775)
);

INVx3_ASAP7_75t_L g2776 ( 
.A(n_2692),
.Y(n_2776)
);

CKINVDCx16_ASAP7_75t_R g2777 ( 
.A(n_2716),
.Y(n_2777)
);

INVxp67_ASAP7_75t_L g2778 ( 
.A(n_2673),
.Y(n_2778)
);

OR2x2_ASAP7_75t_L g2779 ( 
.A(n_2759),
.B(n_2751),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2660),
.B(n_2591),
.Y(n_2780)
);

INVx1_ASAP7_75t_SL g2781 ( 
.A(n_2723),
.Y(n_2781)
);

INVx1_ASAP7_75t_SL g2782 ( 
.A(n_2723),
.Y(n_2782)
);

OR2x2_ASAP7_75t_L g2783 ( 
.A(n_2751),
.B(n_2426),
.Y(n_2783)
);

INVx2_ASAP7_75t_L g2784 ( 
.A(n_2692),
.Y(n_2784)
);

AOI33xp33_ASAP7_75t_L g2785 ( 
.A1(n_2746),
.A2(n_2575),
.A3(n_2590),
.B1(n_2567),
.B2(n_2572),
.B3(n_2653),
.Y(n_2785)
);

INVx1_ASAP7_75t_SL g2786 ( 
.A(n_2684),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2721),
.Y(n_2787)
);

NAND3xp33_ASAP7_75t_L g2788 ( 
.A(n_2754),
.B(n_2617),
.C(n_2611),
.Y(n_2788)
);

INVx2_ASAP7_75t_L g2789 ( 
.A(n_2692),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2739),
.Y(n_2790)
);

INVx2_ASAP7_75t_L g2791 ( 
.A(n_2666),
.Y(n_2791)
);

NAND2xp5_ASAP7_75t_L g2792 ( 
.A(n_2699),
.B(n_2611),
.Y(n_2792)
);

AND2x2_ASAP7_75t_L g2793 ( 
.A(n_2699),
.B(n_2602),
.Y(n_2793)
);

NAND2xp5_ASAP7_75t_L g2794 ( 
.A(n_2730),
.B(n_2617),
.Y(n_2794)
);

AND2x4_ASAP7_75t_L g2795 ( 
.A(n_2666),
.B(n_2622),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2670),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2690),
.B(n_2603),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2690),
.B(n_2603),
.Y(n_2798)
);

INVx1_ASAP7_75t_L g2799 ( 
.A(n_2739),
.Y(n_2799)
);

INVx2_ASAP7_75t_L g2800 ( 
.A(n_2670),
.Y(n_2800)
);

NAND2xp5_ASAP7_75t_L g2801 ( 
.A(n_2730),
.B(n_2622),
.Y(n_2801)
);

INVx2_ASAP7_75t_SL g2802 ( 
.A(n_2736),
.Y(n_2802)
);

INVx2_ASAP7_75t_L g2803 ( 
.A(n_2691),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2711),
.B(n_2606),
.Y(n_2804)
);

NOR2xp33_ASAP7_75t_L g2805 ( 
.A(n_2749),
.B(n_2658),
.Y(n_2805)
);

NOR2xp33_ASAP7_75t_L g2806 ( 
.A(n_2683),
.B(n_2658),
.Y(n_2806)
);

OR2x2_ASAP7_75t_L g2807 ( 
.A(n_2762),
.B(n_2616),
.Y(n_2807)
);

INVx2_ASAP7_75t_L g2808 ( 
.A(n_2691),
.Y(n_2808)
);

NOR2xp33_ASAP7_75t_L g2809 ( 
.A(n_2712),
.B(n_2658),
.Y(n_2809)
);

INVxp67_ASAP7_75t_L g2810 ( 
.A(n_2752),
.Y(n_2810)
);

NAND2xp5_ASAP7_75t_L g2811 ( 
.A(n_2711),
.B(n_2654),
.Y(n_2811)
);

INVx1_ASAP7_75t_L g2812 ( 
.A(n_2772),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2722),
.B(n_2655),
.Y(n_2813)
);

HB1xp67_ASAP7_75t_L g2814 ( 
.A(n_2661),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2772),
.Y(n_2815)
);

INVx1_ASAP7_75t_L g2816 ( 
.A(n_2694),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2694),
.Y(n_2817)
);

INVx2_ASAP7_75t_SL g2818 ( 
.A(n_2736),
.Y(n_2818)
);

OR2x2_ASAP7_75t_L g2819 ( 
.A(n_2762),
.B(n_2486),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2752),
.B(n_2685),
.Y(n_2820)
);

NAND2xp5_ASAP7_75t_L g2821 ( 
.A(n_2722),
.B(n_2655),
.Y(n_2821)
);

AND2x4_ASAP7_75t_L g2822 ( 
.A(n_2661),
.B(n_2648),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2664),
.B(n_2606),
.Y(n_2823)
);

OR2x2_ASAP7_75t_L g2824 ( 
.A(n_2770),
.B(n_2486),
.Y(n_2824)
);

NOR2x1_ASAP7_75t_L g2825 ( 
.A(n_2663),
.B(n_2648),
.Y(n_2825)
);

NAND2xp5_ASAP7_75t_L g2826 ( 
.A(n_2725),
.B(n_2626),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2695),
.Y(n_2827)
);

CKINVDCx20_ASAP7_75t_R g2828 ( 
.A(n_2662),
.Y(n_2828)
);

INVxp67_ASAP7_75t_L g2829 ( 
.A(n_2669),
.Y(n_2829)
);

AND2x2_ASAP7_75t_L g2830 ( 
.A(n_2664),
.B(n_2626),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2725),
.B(n_2649),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2695),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2756),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2665),
.B(n_2649),
.Y(n_2834)
);

NAND2xp5_ASAP7_75t_L g2835 ( 
.A(n_2685),
.B(n_2656),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2770),
.Y(n_2836)
);

AND2x2_ASAP7_75t_L g2837 ( 
.A(n_2665),
.B(n_2656),
.Y(n_2837)
);

AND2x2_ASAP7_75t_L g2838 ( 
.A(n_2753),
.B(n_2758),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2680),
.B(n_2461),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2663),
.Y(n_2840)
);

INVx1_ASAP7_75t_L g2841 ( 
.A(n_2667),
.Y(n_2841)
);

NAND2xp5_ASAP7_75t_L g2842 ( 
.A(n_2669),
.B(n_2576),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2754),
.B(n_2577),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2680),
.B(n_2461),
.Y(n_2844)
);

NAND2x1_ASAP7_75t_SL g2845 ( 
.A(n_2736),
.B(n_2508),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2671),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2672),
.Y(n_2847)
);

OR2x2_ASAP7_75t_L g2848 ( 
.A(n_2734),
.B(n_2445),
.Y(n_2848)
);

AND2x2_ASAP7_75t_L g2849 ( 
.A(n_2681),
.B(n_2464),
.Y(n_2849)
);

INVx2_ASAP7_75t_L g2850 ( 
.A(n_2763),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2675),
.Y(n_2851)
);

NAND2xp5_ASAP7_75t_L g2852 ( 
.A(n_2714),
.B(n_2580),
.Y(n_2852)
);

NAND2xp5_ASAP7_75t_L g2853 ( 
.A(n_2714),
.B(n_2581),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2734),
.Y(n_2854)
);

INVx2_ASAP7_75t_L g2855 ( 
.A(n_2763),
.Y(n_2855)
);

NAND2xp5_ASAP7_75t_L g2856 ( 
.A(n_2717),
.B(n_2584),
.Y(n_2856)
);

NAND2xp5_ASAP7_75t_L g2857 ( 
.A(n_2717),
.B(n_2592),
.Y(n_2857)
);

INVx1_ASAP7_75t_L g2858 ( 
.A(n_2743),
.Y(n_2858)
);

INVx1_ASAP7_75t_L g2859 ( 
.A(n_2743),
.Y(n_2859)
);

NAND2xp5_ASAP7_75t_L g2860 ( 
.A(n_2753),
.B(n_2593),
.Y(n_2860)
);

INVx1_ASAP7_75t_L g2861 ( 
.A(n_2709),
.Y(n_2861)
);

INVx1_ASAP7_75t_SL g2862 ( 
.A(n_2740),
.Y(n_2862)
);

NAND2xp5_ASAP7_75t_L g2863 ( 
.A(n_2758),
.B(n_2595),
.Y(n_2863)
);

OR2x2_ASAP7_75t_L g2864 ( 
.A(n_2729),
.B(n_2492),
.Y(n_2864)
);

NAND2xp5_ASAP7_75t_L g2865 ( 
.A(n_2809),
.B(n_2696),
.Y(n_2865)
);

OAI21xp33_ASAP7_75t_SL g2866 ( 
.A1(n_2845),
.A2(n_2746),
.B(n_2689),
.Y(n_2866)
);

INVx1_ASAP7_75t_L g2867 ( 
.A(n_2814),
.Y(n_2867)
);

OAI32xp33_ASAP7_75t_L g2868 ( 
.A1(n_2777),
.A2(n_2689),
.A3(n_2659),
.B1(n_2703),
.B2(n_2766),
.Y(n_2868)
);

OAI31xp33_ASAP7_75t_L g2869 ( 
.A1(n_2809),
.A2(n_2659),
.A3(n_2703),
.B(n_2678),
.Y(n_2869)
);

AOI21xp33_ASAP7_75t_L g2870 ( 
.A1(n_2829),
.A2(n_2760),
.B(n_2713),
.Y(n_2870)
);

OAI22xp33_ASAP7_75t_L g2871 ( 
.A1(n_2843),
.A2(n_2687),
.B1(n_2720),
.B2(n_2674),
.Y(n_2871)
);

INVxp67_ASAP7_75t_L g2872 ( 
.A(n_2805),
.Y(n_2872)
);

NOR2x1_ASAP7_75t_L g2873 ( 
.A(n_2776),
.B(n_2763),
.Y(n_2873)
);

OA21x2_ASAP7_75t_SL g2874 ( 
.A1(n_2775),
.A2(n_2719),
.B(n_2728),
.Y(n_2874)
);

OAI22xp33_ASAP7_75t_L g2875 ( 
.A1(n_2778),
.A2(n_2674),
.B1(n_2682),
.B2(n_2748),
.Y(n_2875)
);

NAND2xp5_ASAP7_75t_L g2876 ( 
.A(n_2862),
.B(n_2697),
.Y(n_2876)
);

AND2x2_ASAP7_75t_L g2877 ( 
.A(n_2793),
.B(n_2740),
.Y(n_2877)
);

INVx1_ASAP7_75t_L g2878 ( 
.A(n_2814),
.Y(n_2878)
);

AND2x2_ASAP7_75t_L g2879 ( 
.A(n_2793),
.B(n_2804),
.Y(n_2879)
);

NAND2xp5_ASAP7_75t_L g2880 ( 
.A(n_2786),
.B(n_2677),
.Y(n_2880)
);

AOI21xp5_ASAP7_75t_L g2881 ( 
.A1(n_2775),
.A2(n_2805),
.B(n_2842),
.Y(n_2881)
);

OAI21xp33_ASAP7_75t_L g2882 ( 
.A1(n_2838),
.A2(n_2713),
.B(n_2681),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2830),
.Y(n_2883)
);

AOI22xp33_ASAP7_75t_SL g2884 ( 
.A1(n_2828),
.A2(n_2771),
.B1(n_2679),
.B2(n_2688),
.Y(n_2884)
);

INVx1_ASAP7_75t_L g2885 ( 
.A(n_2830),
.Y(n_2885)
);

INVx1_ASAP7_75t_L g2886 ( 
.A(n_2776),
.Y(n_2886)
);

OAI222xp33_ASAP7_75t_L g2887 ( 
.A1(n_2781),
.A2(n_2682),
.B1(n_2742),
.B2(n_2709),
.C1(n_2708),
.C2(n_2676),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2802),
.B(n_2668),
.Y(n_2888)
);

OAI21xp33_ASAP7_75t_L g2889 ( 
.A1(n_2811),
.A2(n_2771),
.B(n_2747),
.Y(n_2889)
);

OAI21xp33_ASAP7_75t_L g2890 ( 
.A1(n_2820),
.A2(n_2733),
.B(n_2767),
.Y(n_2890)
);

AND2x2_ASAP7_75t_L g2891 ( 
.A(n_2804),
.B(n_2686),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2776),
.Y(n_2892)
);

INVx1_ASAP7_75t_L g2893 ( 
.A(n_2807),
.Y(n_2893)
);

OR2x2_ASAP7_75t_L g2894 ( 
.A(n_2792),
.B(n_2732),
.Y(n_2894)
);

INVx2_ASAP7_75t_L g2895 ( 
.A(n_2802),
.Y(n_2895)
);

OAI322xp33_ASAP7_75t_L g2896 ( 
.A1(n_2806),
.A2(n_2700),
.A3(n_2698),
.B1(n_2707),
.B2(n_2705),
.C1(n_2701),
.C2(n_2693),
.Y(n_2896)
);

AOI22xp5_ASAP7_75t_L g2897 ( 
.A1(n_2828),
.A2(n_2731),
.B1(n_2737),
.B2(n_2735),
.Y(n_2897)
);

INVx2_ASAP7_75t_L g2898 ( 
.A(n_2818),
.Y(n_2898)
);

NAND2xp5_ASAP7_75t_L g2899 ( 
.A(n_2810),
.B(n_2738),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2834),
.Y(n_2900)
);

INVx2_ASAP7_75t_L g2901 ( 
.A(n_2818),
.Y(n_2901)
);

OR2x2_ASAP7_75t_L g2902 ( 
.A(n_2774),
.B(n_2741),
.Y(n_2902)
);

NOR3xp33_ASAP7_75t_SL g2903 ( 
.A(n_2788),
.B(n_2773),
.C(n_2806),
.Y(n_2903)
);

INVx3_ASAP7_75t_L g2904 ( 
.A(n_2795),
.Y(n_2904)
);

AOI222xp33_ASAP7_75t_L g2905 ( 
.A1(n_2861),
.A2(n_2724),
.B1(n_2750),
.B2(n_2764),
.C1(n_2761),
.C2(n_2757),
.Y(n_2905)
);

OR2x2_ASAP7_75t_L g2906 ( 
.A(n_2780),
.B(n_2745),
.Y(n_2906)
);

AND2x2_ASAP7_75t_L g2907 ( 
.A(n_2797),
.B(n_2702),
.Y(n_2907)
);

AND2x2_ASAP7_75t_L g2908 ( 
.A(n_2797),
.B(n_2706),
.Y(n_2908)
);

AND2x2_ASAP7_75t_L g2909 ( 
.A(n_2798),
.B(n_2464),
.Y(n_2909)
);

OAI211xp5_ASAP7_75t_SL g2910 ( 
.A1(n_2782),
.A2(n_2768),
.B(n_2769),
.C(n_2765),
.Y(n_2910)
);

INVx1_ASAP7_75t_L g2911 ( 
.A(n_2834),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2798),
.B(n_2710),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2837),
.Y(n_2913)
);

INVx1_ASAP7_75t_L g2914 ( 
.A(n_2837),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2823),
.B(n_2850),
.Y(n_2915)
);

INVx1_ASAP7_75t_L g2916 ( 
.A(n_2822),
.Y(n_2916)
);

AOI21xp33_ASAP7_75t_L g2917 ( 
.A1(n_2779),
.A2(n_2787),
.B(n_2833),
.Y(n_2917)
);

INVx2_ASAP7_75t_L g2918 ( 
.A(n_2795),
.Y(n_2918)
);

OR2x2_ASAP7_75t_L g2919 ( 
.A(n_2813),
.B(n_2492),
.Y(n_2919)
);

OAI21xp33_ASAP7_75t_L g2920 ( 
.A1(n_2823),
.A2(n_2618),
.B(n_2608),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2850),
.B(n_2718),
.Y(n_2921)
);

OAI211xp5_ASAP7_75t_L g2922 ( 
.A1(n_2835),
.A2(n_2727),
.B(n_2726),
.C(n_2755),
.Y(n_2922)
);

AOI21xp5_ASAP7_75t_L g2923 ( 
.A1(n_2821),
.A2(n_2755),
.B(n_2744),
.Y(n_2923)
);

AOI222xp33_ASAP7_75t_L g2924 ( 
.A1(n_2790),
.A2(n_2812),
.B1(n_2815),
.B2(n_2799),
.C1(n_2841),
.C2(n_2846),
.Y(n_2924)
);

INVx1_ASAP7_75t_L g2925 ( 
.A(n_2822),
.Y(n_2925)
);

OR2x2_ASAP7_75t_L g2926 ( 
.A(n_2826),
.B(n_2497),
.Y(n_2926)
);

AND2x2_ASAP7_75t_L g2927 ( 
.A(n_2839),
.B(n_2466),
.Y(n_2927)
);

INVx1_ASAP7_75t_L g2928 ( 
.A(n_2822),
.Y(n_2928)
);

INVx1_ASAP7_75t_L g2929 ( 
.A(n_2825),
.Y(n_2929)
);

OR2x2_ASAP7_75t_L g2930 ( 
.A(n_2864),
.B(n_2497),
.Y(n_2930)
);

NOR4xp25_ASAP7_75t_L g2931 ( 
.A(n_2784),
.B(n_2620),
.C(n_2627),
.D(n_2619),
.Y(n_2931)
);

AOI22xp5_ASAP7_75t_L g2932 ( 
.A1(n_2839),
.A2(n_2529),
.B1(n_2633),
.B2(n_2632),
.Y(n_2932)
);

INVx2_ASAP7_75t_L g2933 ( 
.A(n_2795),
.Y(n_2933)
);

INVx1_ASAP7_75t_L g2934 ( 
.A(n_2784),
.Y(n_2934)
);

OR2x2_ASAP7_75t_L g2935 ( 
.A(n_2819),
.B(n_2634),
.Y(n_2935)
);

A2O1A1Ixp33_ASAP7_75t_L g2936 ( 
.A1(n_2785),
.A2(n_2636),
.B(n_2640),
.C(n_2639),
.Y(n_2936)
);

INVx1_ASAP7_75t_L g2937 ( 
.A(n_2789),
.Y(n_2937)
);

INVxp67_ASAP7_75t_L g2938 ( 
.A(n_2789),
.Y(n_2938)
);

AOI21xp5_ASAP7_75t_L g2939 ( 
.A1(n_2855),
.A2(n_2744),
.B(n_2652),
.Y(n_2939)
);

OR2x2_ASAP7_75t_L g2940 ( 
.A(n_2824),
.B(n_2650),
.Y(n_2940)
);

AND2x2_ASAP7_75t_L g2941 ( 
.A(n_2877),
.B(n_2855),
.Y(n_2941)
);

AOI22xp33_ASAP7_75t_L g2942 ( 
.A1(n_2869),
.A2(n_2844),
.B1(n_2849),
.B2(n_2836),
.Y(n_2942)
);

INVx1_ASAP7_75t_SL g2943 ( 
.A(n_2879),
.Y(n_2943)
);

INVx2_ASAP7_75t_L g2944 ( 
.A(n_2904),
.Y(n_2944)
);

NOR2xp33_ASAP7_75t_SL g2945 ( 
.A(n_2887),
.B(n_2791),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2904),
.Y(n_2946)
);

AND2x2_ASAP7_75t_L g2947 ( 
.A(n_2891),
.B(n_2844),
.Y(n_2947)
);

NAND2xp5_ASAP7_75t_L g2948 ( 
.A(n_2884),
.B(n_2791),
.Y(n_2948)
);

HB1xp67_ASAP7_75t_L g2949 ( 
.A(n_2873),
.Y(n_2949)
);

NOR2xp33_ASAP7_75t_L g2950 ( 
.A(n_2882),
.B(n_2863),
.Y(n_2950)
);

INVx1_ASAP7_75t_L g2951 ( 
.A(n_2916),
.Y(n_2951)
);

INVx1_ASAP7_75t_L g2952 ( 
.A(n_2925),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2928),
.Y(n_2953)
);

AND2x2_ASAP7_75t_L g2954 ( 
.A(n_2909),
.B(n_2849),
.Y(n_2954)
);

CKINVDCx14_ASAP7_75t_R g2955 ( 
.A(n_2895),
.Y(n_2955)
);

NOR2xp33_ASAP7_75t_L g2956 ( 
.A(n_2872),
.B(n_2860),
.Y(n_2956)
);

OAI21xp5_ASAP7_75t_SL g2957 ( 
.A1(n_2869),
.A2(n_2853),
.B(n_2852),
.Y(n_2957)
);

OAI22xp5_ASAP7_75t_L g2958 ( 
.A1(n_2865),
.A2(n_2881),
.B1(n_2897),
.B2(n_2903),
.Y(n_2958)
);

INVx2_ASAP7_75t_L g2959 ( 
.A(n_2918),
.Y(n_2959)
);

AND2x2_ASAP7_75t_SL g2960 ( 
.A(n_2865),
.B(n_2847),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2907),
.B(n_2854),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2933),
.Y(n_2962)
);

INVx1_ASAP7_75t_L g2963 ( 
.A(n_2867),
.Y(n_2963)
);

INVx2_ASAP7_75t_L g2964 ( 
.A(n_2929),
.Y(n_2964)
);

NAND2xp5_ASAP7_75t_L g2965 ( 
.A(n_2908),
.B(n_2858),
.Y(n_2965)
);

NAND2xp5_ASAP7_75t_L g2966 ( 
.A(n_2898),
.B(n_2859),
.Y(n_2966)
);

NAND2xp5_ASAP7_75t_L g2967 ( 
.A(n_2901),
.B(n_2840),
.Y(n_2967)
);

AND2x4_ASAP7_75t_L g2968 ( 
.A(n_2878),
.B(n_2796),
.Y(n_2968)
);

INVx1_ASAP7_75t_L g2969 ( 
.A(n_2886),
.Y(n_2969)
);

NAND2xp5_ASAP7_75t_L g2970 ( 
.A(n_2883),
.B(n_2796),
.Y(n_2970)
);

INVxp67_ASAP7_75t_L g2971 ( 
.A(n_2915),
.Y(n_2971)
);

INVx2_ASAP7_75t_L g2972 ( 
.A(n_2892),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2885),
.B(n_2800),
.Y(n_2973)
);

AND2x2_ASAP7_75t_L g2974 ( 
.A(n_2927),
.B(n_2900),
.Y(n_2974)
);

AND2x2_ASAP7_75t_L g2975 ( 
.A(n_2911),
.B(n_2800),
.Y(n_2975)
);

INVx2_ASAP7_75t_SL g2976 ( 
.A(n_2913),
.Y(n_2976)
);

INVx1_ASAP7_75t_L g2977 ( 
.A(n_2914),
.Y(n_2977)
);

NAND2xp33_ASAP7_75t_SL g2978 ( 
.A(n_2888),
.B(n_2785),
.Y(n_2978)
);

NAND2xp5_ASAP7_75t_L g2979 ( 
.A(n_2905),
.B(n_2803),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2880),
.Y(n_2980)
);

NAND2xp33_ASAP7_75t_L g2981 ( 
.A(n_2876),
.B(n_2794),
.Y(n_2981)
);

INVxp67_ASAP7_75t_L g2982 ( 
.A(n_2876),
.Y(n_2982)
);

INVx2_ASAP7_75t_L g2983 ( 
.A(n_2930),
.Y(n_2983)
);

AND2x2_ASAP7_75t_L g2984 ( 
.A(n_2893),
.B(n_2803),
.Y(n_2984)
);

AND2x2_ASAP7_75t_L g2985 ( 
.A(n_2938),
.B(n_2808),
.Y(n_2985)
);

NAND2x1p5_ASAP7_75t_L g2986 ( 
.A(n_2934),
.B(n_2808),
.Y(n_2986)
);

INVx1_ASAP7_75t_L g2987 ( 
.A(n_2880),
.Y(n_2987)
);

OR2x2_ASAP7_75t_L g2988 ( 
.A(n_2937),
.B(n_2848),
.Y(n_2988)
);

INVx2_ASAP7_75t_L g2989 ( 
.A(n_2935),
.Y(n_2989)
);

INVx2_ASAP7_75t_L g2990 ( 
.A(n_2940),
.Y(n_2990)
);

NAND2xp5_ASAP7_75t_SL g2991 ( 
.A(n_2870),
.B(n_2866),
.Y(n_2991)
);

NOR2xp33_ASAP7_75t_L g2992 ( 
.A(n_2868),
.B(n_2856),
.Y(n_2992)
);

INVx2_ASAP7_75t_L g2993 ( 
.A(n_2919),
.Y(n_2993)
);

OR2x2_ASAP7_75t_L g2994 ( 
.A(n_2912),
.B(n_2783),
.Y(n_2994)
);

NOR2xp67_ASAP7_75t_L g2995 ( 
.A(n_2939),
.B(n_2816),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2899),
.Y(n_2996)
);

INVx1_ASAP7_75t_SL g2997 ( 
.A(n_2894),
.Y(n_2997)
);

NAND2x1_ASAP7_75t_SL g2998 ( 
.A(n_2932),
.B(n_2817),
.Y(n_2998)
);

INVx1_ASAP7_75t_L g2999 ( 
.A(n_2899),
.Y(n_2999)
);

NAND2xp5_ASAP7_75t_SL g3000 ( 
.A(n_2870),
.B(n_2827),
.Y(n_3000)
);

INVxp67_ASAP7_75t_L g3001 ( 
.A(n_2924),
.Y(n_3001)
);

NAND2xp5_ASAP7_75t_L g3002 ( 
.A(n_2905),
.B(n_2801),
.Y(n_3002)
);

HB1xp67_ASAP7_75t_L g3003 ( 
.A(n_2926),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2871),
.B(n_2831),
.Y(n_3004)
);

NAND2xp5_ASAP7_75t_SL g3005 ( 
.A(n_2924),
.B(n_2832),
.Y(n_3005)
);

NOR4xp75_ASAP7_75t_L g3006 ( 
.A(n_2890),
.B(n_2857),
.C(n_2429),
.D(n_2436),
.Y(n_3006)
);

NAND2xp5_ASAP7_75t_L g3007 ( 
.A(n_2875),
.B(n_2851),
.Y(n_3007)
);

NOR2xp33_ASAP7_75t_L g3008 ( 
.A(n_2889),
.B(n_2316),
.Y(n_3008)
);

NAND2xp5_ASAP7_75t_L g3009 ( 
.A(n_2917),
.B(n_2481),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_SL g3010 ( 
.A(n_2923),
.B(n_2922),
.Y(n_3010)
);

OR2x2_ASAP7_75t_L g3011 ( 
.A(n_2943),
.B(n_2902),
.Y(n_3011)
);

OR4x1_ASAP7_75t_L g3012 ( 
.A(n_2976),
.B(n_2874),
.C(n_2917),
.D(n_2896),
.Y(n_3012)
);

OAI21xp5_ASAP7_75t_SL g3013 ( 
.A1(n_3001),
.A2(n_2910),
.B(n_2906),
.Y(n_3013)
);

AND2x2_ASAP7_75t_L g3014 ( 
.A(n_2947),
.B(n_2921),
.Y(n_3014)
);

NAND2xp5_ASAP7_75t_L g3015 ( 
.A(n_2947),
.B(n_2920),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2986),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2986),
.Y(n_3017)
);

NAND2xp5_ASAP7_75t_L g3018 ( 
.A(n_2941),
.B(n_2936),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2941),
.B(n_2954),
.Y(n_3019)
);

AND2x2_ASAP7_75t_L g3020 ( 
.A(n_2954),
.B(n_2931),
.Y(n_3020)
);

AOI22x1_ASAP7_75t_SL g3021 ( 
.A1(n_2997),
.A2(n_2931),
.B1(n_2424),
.B2(n_2418),
.Y(n_3021)
);

NAND2xp5_ASAP7_75t_L g3022 ( 
.A(n_2955),
.B(n_2466),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2961),
.B(n_2510),
.Y(n_3023)
);

HB1xp67_ASAP7_75t_L g3024 ( 
.A(n_2949),
.Y(n_3024)
);

INVx2_ASAP7_75t_L g3025 ( 
.A(n_2998),
.Y(n_3025)
);

INVxp67_ASAP7_75t_L g3026 ( 
.A(n_2945),
.Y(n_3026)
);

INVx2_ASAP7_75t_L g3027 ( 
.A(n_2968),
.Y(n_3027)
);

NAND2xp5_ASAP7_75t_L g3028 ( 
.A(n_2955),
.B(n_2477),
.Y(n_3028)
);

NOR3xp33_ASAP7_75t_L g3029 ( 
.A(n_2958),
.B(n_2424),
.C(n_2417),
.Y(n_3029)
);

INVx1_ASAP7_75t_L g3030 ( 
.A(n_2944),
.Y(n_3030)
);

NAND2xp5_ASAP7_75t_L g3031 ( 
.A(n_2960),
.B(n_2477),
.Y(n_3031)
);

NAND2xp5_ASAP7_75t_L g3032 ( 
.A(n_2960),
.B(n_2348),
.Y(n_3032)
);

A2O1A1Ixp33_ASAP7_75t_L g3033 ( 
.A1(n_2979),
.A2(n_2363),
.B(n_2251),
.C(n_2526),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2944),
.Y(n_3034)
);

OR2x2_ASAP7_75t_L g3035 ( 
.A(n_2983),
.B(n_3009),
.Y(n_3035)
);

NAND2xp5_ASAP7_75t_L g3036 ( 
.A(n_2961),
.B(n_2356),
.Y(n_3036)
);

NAND2xp5_ASAP7_75t_L g3037 ( 
.A(n_2942),
.B(n_2356),
.Y(n_3037)
);

OR2x2_ASAP7_75t_L g3038 ( 
.A(n_2983),
.B(n_2744),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2968),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2946),
.B(n_2365),
.Y(n_3040)
);

INVx1_ASAP7_75t_L g3041 ( 
.A(n_2968),
.Y(n_3041)
);

NAND2xp5_ASAP7_75t_L g3042 ( 
.A(n_2974),
.B(n_2369),
.Y(n_3042)
);

NAND2xp5_ASAP7_75t_SL g3043 ( 
.A(n_3002),
.B(n_2261),
.Y(n_3043)
);

AND2x2_ASAP7_75t_L g3044 ( 
.A(n_2974),
.B(n_3003),
.Y(n_3044)
);

INVx3_ASAP7_75t_L g3045 ( 
.A(n_2959),
.Y(n_3045)
);

AND2x2_ASAP7_75t_L g3046 ( 
.A(n_2984),
.B(n_2510),
.Y(n_3046)
);

INVxp33_ASAP7_75t_L g3047 ( 
.A(n_3005),
.Y(n_3047)
);

AND2x2_ASAP7_75t_L g3048 ( 
.A(n_2984),
.B(n_2519),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2959),
.B(n_2985),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2975),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2975),
.Y(n_3051)
);

NOR2xp33_ASAP7_75t_L g3052 ( 
.A(n_3005),
.B(n_2375),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2985),
.Y(n_3053)
);

NAND2xp5_ASAP7_75t_L g3054 ( 
.A(n_2976),
.B(n_2376),
.Y(n_3054)
);

NAND2xp5_ASAP7_75t_L g3055 ( 
.A(n_2962),
.B(n_2519),
.Y(n_3055)
);

NOR2xp33_ASAP7_75t_R g3056 ( 
.A(n_2981),
.B(n_2251),
.Y(n_3056)
);

NAND2xp5_ASAP7_75t_L g3057 ( 
.A(n_2992),
.B(n_2951),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2988),
.Y(n_3058)
);

NAND2xp5_ASAP7_75t_L g3059 ( 
.A(n_2952),
.B(n_2525),
.Y(n_3059)
);

NAND2xp5_ASAP7_75t_L g3060 ( 
.A(n_2953),
.B(n_2525),
.Y(n_3060)
);

NOR2xp33_ASAP7_75t_L g3061 ( 
.A(n_3010),
.B(n_2251),
.Y(n_3061)
);

NOR2x1_ASAP7_75t_R g3062 ( 
.A(n_2991),
.B(n_1936),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2988),
.Y(n_3063)
);

NAND2xp5_ASAP7_75t_L g3064 ( 
.A(n_2989),
.B(n_2526),
.Y(n_3064)
);

INVx1_ASAP7_75t_L g3065 ( 
.A(n_2965),
.Y(n_3065)
);

INVx1_ASAP7_75t_L g3066 ( 
.A(n_2970),
.Y(n_3066)
);

NAND2xp5_ASAP7_75t_L g3067 ( 
.A(n_2989),
.B(n_2527),
.Y(n_3067)
);

AOI21xp33_ASAP7_75t_SL g3068 ( 
.A1(n_3010),
.A2(n_2436),
.B(n_2429),
.Y(n_3068)
);

AND2x2_ASAP7_75t_L g3069 ( 
.A(n_2990),
.B(n_2527),
.Y(n_3069)
);

AOI32xp33_ASAP7_75t_L g3070 ( 
.A1(n_2978),
.A2(n_2261),
.A3(n_2265),
.B1(n_2387),
.B2(n_2358),
.Y(n_3070)
);

NOR2xp33_ASAP7_75t_L g3071 ( 
.A(n_3026),
.B(n_2982),
.Y(n_3071)
);

AND2x2_ASAP7_75t_L g3072 ( 
.A(n_3044),
.B(n_2993),
.Y(n_3072)
);

NOR2x1_ASAP7_75t_L g3073 ( 
.A(n_3045),
.B(n_3000),
.Y(n_3073)
);

NAND2x1_ASAP7_75t_L g3074 ( 
.A(n_3045),
.B(n_3027),
.Y(n_3074)
);

NAND4xp25_ASAP7_75t_SL g3075 ( 
.A(n_3037),
.B(n_2948),
.C(n_3004),
.D(n_3007),
.Y(n_3075)
);

NAND2xp5_ASAP7_75t_L g3076 ( 
.A(n_3049),
.B(n_2990),
.Y(n_3076)
);

NAND4xp25_ASAP7_75t_L g3077 ( 
.A(n_3022),
.B(n_2950),
.C(n_2956),
.D(n_2991),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_3049),
.B(n_2957),
.Y(n_3078)
);

NOR2xp33_ASAP7_75t_L g3079 ( 
.A(n_3028),
.B(n_2971),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_SL g3080 ( 
.A(n_3025),
.B(n_2993),
.Y(n_3080)
);

INVx2_ASAP7_75t_L g3081 ( 
.A(n_3027),
.Y(n_3081)
);

AND4x1_ASAP7_75t_L g3082 ( 
.A(n_3019),
.B(n_2980),
.C(n_2987),
.D(n_2967),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_3039),
.Y(n_3083)
);

INVx1_ASAP7_75t_L g3084 ( 
.A(n_3041),
.Y(n_3084)
);

HB1xp67_ASAP7_75t_L g3085 ( 
.A(n_3025),
.Y(n_3085)
);

NOR2xp33_ASAP7_75t_SL g3086 ( 
.A(n_3014),
.B(n_2994),
.Y(n_3086)
);

NOR2xp33_ASAP7_75t_L g3087 ( 
.A(n_3032),
.B(n_3000),
.Y(n_3087)
);

AND3x1_ASAP7_75t_L g3088 ( 
.A(n_3013),
.B(n_2966),
.C(n_2973),
.Y(n_3088)
);

NAND3xp33_ASAP7_75t_SL g3089 ( 
.A(n_3047),
.B(n_3006),
.C(n_2978),
.Y(n_3089)
);

NOR3xp33_ASAP7_75t_SL g3090 ( 
.A(n_3057),
.B(n_2999),
.C(n_2996),
.Y(n_3090)
);

AND2x2_ASAP7_75t_L g3091 ( 
.A(n_3053),
.B(n_2977),
.Y(n_3091)
);

NOR3xp33_ASAP7_75t_L g3092 ( 
.A(n_3058),
.B(n_2981),
.C(n_2995),
.Y(n_3092)
);

NOR3xp33_ASAP7_75t_L g3093 ( 
.A(n_3058),
.B(n_2963),
.C(n_2964),
.Y(n_3093)
);

NOR2xp67_ASAP7_75t_SL g3094 ( 
.A(n_3024),
.B(n_2964),
.Y(n_3094)
);

NOR3xp33_ASAP7_75t_L g3095 ( 
.A(n_3063),
.B(n_2972),
.C(n_2969),
.Y(n_3095)
);

AND2x2_ASAP7_75t_L g3096 ( 
.A(n_3069),
.B(n_2972),
.Y(n_3096)
);

NOR2xp33_ASAP7_75t_L g3097 ( 
.A(n_3031),
.B(n_3008),
.Y(n_3097)
);

AOI22xp33_ASAP7_75t_L g3098 ( 
.A1(n_3047),
.A2(n_2265),
.B1(n_2367),
.B2(n_2364),
.Y(n_3098)
);

INVx1_ASAP7_75t_L g3099 ( 
.A(n_3038),
.Y(n_3099)
);

NOR3xp33_ASAP7_75t_L g3100 ( 
.A(n_3020),
.B(n_3045),
.C(n_3017),
.Y(n_3100)
);

OR2x2_ASAP7_75t_L g3101 ( 
.A(n_3036),
.B(n_2372),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_3050),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_3051),
.Y(n_3103)
);

NAND4xp25_ASAP7_75t_L g3104 ( 
.A(n_3015),
.B(n_2209),
.C(n_2358),
.D(n_2372),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_3069),
.B(n_3011),
.Y(n_3105)
);

OAI211xp5_ASAP7_75t_L g3106 ( 
.A1(n_3070),
.A2(n_2371),
.B(n_2284),
.C(n_2337),
.Y(n_3106)
);

NOR3x1_ASAP7_75t_L g3107 ( 
.A(n_3018),
.B(n_2063),
.C(n_2371),
.Y(n_3107)
);

NOR2xp33_ASAP7_75t_L g3108 ( 
.A(n_3035),
.B(n_2399),
.Y(n_3108)
);

NAND2xp33_ASAP7_75t_SL g3109 ( 
.A(n_3020),
.B(n_2394),
.Y(n_3109)
);

NAND2xp5_ASAP7_75t_L g3110 ( 
.A(n_3030),
.B(n_2394),
.Y(n_3110)
);

NOR2xp33_ASAP7_75t_L g3111 ( 
.A(n_3062),
.B(n_2399),
.Y(n_3111)
);

AOI21xp5_ASAP7_75t_L g3112 ( 
.A1(n_3043),
.A2(n_3052),
.B(n_3061),
.Y(n_3112)
);

NAND2xp5_ASAP7_75t_L g3113 ( 
.A(n_3034),
.B(n_2395),
.Y(n_3113)
);

NOR3x1_ASAP7_75t_L g3114 ( 
.A(n_3055),
.B(n_2063),
.C(n_1845),
.Y(n_3114)
);

NAND2xp5_ASAP7_75t_L g3115 ( 
.A(n_3046),
.B(n_2395),
.Y(n_3115)
);

NAND4xp25_ASAP7_75t_L g3116 ( 
.A(n_3029),
.B(n_2398),
.C(n_2323),
.D(n_2349),
.Y(n_3116)
);

OAI21xp33_ASAP7_75t_SL g3117 ( 
.A1(n_3052),
.A2(n_2377),
.B(n_2284),
.Y(n_3117)
);

INVx1_ASAP7_75t_L g3118 ( 
.A(n_3016),
.Y(n_3118)
);

NAND2xp5_ASAP7_75t_SL g3119 ( 
.A(n_3068),
.B(n_2274),
.Y(n_3119)
);

OAI21xp5_ASAP7_75t_L g3120 ( 
.A1(n_3043),
.A2(n_2334),
.B(n_2274),
.Y(n_3120)
);

AOI21xp5_ASAP7_75t_L g3121 ( 
.A1(n_3073),
.A2(n_3061),
.B(n_3054),
.Y(n_3121)
);

OAI221xp5_ASAP7_75t_L g3122 ( 
.A1(n_3086),
.A2(n_3067),
.B1(n_3064),
.B2(n_3042),
.C(n_3066),
.Y(n_3122)
);

INVxp67_ASAP7_75t_L g3123 ( 
.A(n_3094),
.Y(n_3123)
);

AOI221xp5_ASAP7_75t_L g3124 ( 
.A1(n_3089),
.A2(n_3012),
.B1(n_3060),
.B2(n_3059),
.C(n_3065),
.Y(n_3124)
);

OAI22xp5_ASAP7_75t_L g3125 ( 
.A1(n_3078),
.A2(n_3033),
.B1(n_3023),
.B2(n_3040),
.Y(n_3125)
);

O2A1O1Ixp33_ASAP7_75t_L g3126 ( 
.A1(n_3092),
.A2(n_3012),
.B(n_3033),
.C(n_3021),
.Y(n_3126)
);

AOI221xp5_ASAP7_75t_L g3127 ( 
.A1(n_3100),
.A2(n_3048),
.B1(n_3046),
.B2(n_3023),
.C(n_3056),
.Y(n_3127)
);

AOI21xp5_ASAP7_75t_L g3128 ( 
.A1(n_3074),
.A2(n_3112),
.B(n_3080),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_3072),
.B(n_3048),
.Y(n_3129)
);

AOI32xp33_ASAP7_75t_L g3130 ( 
.A1(n_3088),
.A2(n_3056),
.A3(n_2377),
.B1(n_2368),
.B2(n_2367),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_3085),
.Y(n_3131)
);

AOI21xp5_ASAP7_75t_L g3132 ( 
.A1(n_3092),
.A2(n_2337),
.B(n_2334),
.Y(n_3132)
);

AOI322xp5_ASAP7_75t_L g3133 ( 
.A1(n_3100),
.A2(n_2368),
.A3(n_2364),
.B1(n_2355),
.B2(n_2354),
.C1(n_2342),
.C2(n_2341),
.Y(n_3133)
);

OAI21xp5_ASAP7_75t_SL g3134 ( 
.A1(n_3071),
.A2(n_1985),
.B(n_2339),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_3085),
.Y(n_3135)
);

AOI222xp33_ASAP7_75t_L g3136 ( 
.A1(n_3087),
.A2(n_2355),
.B1(n_2354),
.B2(n_2342),
.C1(n_2341),
.C2(n_2339),
.Y(n_3136)
);

AOI22xp5_ASAP7_75t_L g3137 ( 
.A1(n_3075),
.A2(n_2168),
.B1(n_1973),
.B2(n_1979),
.Y(n_3137)
);

BUFx8_ASAP7_75t_SL g3138 ( 
.A(n_3076),
.Y(n_3138)
);

NAND2xp5_ASAP7_75t_SL g3139 ( 
.A(n_3109),
.B(n_2100),
.Y(n_3139)
);

NAND5xp2_ASAP7_75t_L g3140 ( 
.A(n_3108),
.B(n_2215),
.C(n_2228),
.D(n_2222),
.E(n_2026),
.Y(n_3140)
);

AOI221x1_ASAP7_75t_L g3141 ( 
.A1(n_3093),
.A2(n_2112),
.B1(n_2113),
.B2(n_2218),
.C(n_2212),
.Y(n_3141)
);

AOI22xp5_ASAP7_75t_L g3142 ( 
.A1(n_3111),
.A2(n_1979),
.B1(n_2112),
.B2(n_2113),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_3081),
.B(n_2224),
.Y(n_3143)
);

AOI211xp5_ASAP7_75t_SL g3144 ( 
.A1(n_3079),
.A2(n_2044),
.B(n_2039),
.C(n_2236),
.Y(n_3144)
);

O2A1O1Ixp33_ASAP7_75t_L g3145 ( 
.A1(n_3093),
.A2(n_2232),
.B(n_2236),
.C(n_2224),
.Y(n_3145)
);

AOI222xp33_ASAP7_75t_L g3146 ( 
.A1(n_3083),
.A2(n_2140),
.B1(n_2131),
.B2(n_2208),
.C1(n_2144),
.C2(n_2159),
.Y(n_3146)
);

NOR3x1_ASAP7_75t_L g3147 ( 
.A(n_3077),
.B(n_2169),
.C(n_2179),
.Y(n_3147)
);

XOR2x2_ASAP7_75t_L g3148 ( 
.A(n_3082),
.B(n_2232),
.Y(n_3148)
);

NOR2xp33_ASAP7_75t_R g3149 ( 
.A(n_3105),
.B(n_1116),
.Y(n_3149)
);

AOI211x1_ASAP7_75t_SL g3150 ( 
.A1(n_3110),
.A2(n_2161),
.B(n_2159),
.C(n_2144),
.Y(n_3150)
);

AOI322xp5_ASAP7_75t_L g3151 ( 
.A1(n_3090),
.A2(n_3097),
.A3(n_3095),
.B1(n_3118),
.B2(n_3113),
.C1(n_3084),
.C2(n_3102),
.Y(n_3151)
);

OAI211xp5_ASAP7_75t_SL g3152 ( 
.A1(n_3090),
.A2(n_2222),
.B(n_2208),
.C(n_2161),
.Y(n_3152)
);

AOI211xp5_ASAP7_75t_SL g3153 ( 
.A1(n_3095),
.A2(n_2039),
.B(n_2140),
.C(n_2131),
.Y(n_3153)
);

AOI222xp33_ASAP7_75t_L g3154 ( 
.A1(n_3099),
.A2(n_1854),
.B1(n_2045),
.B2(n_2050),
.C1(n_2031),
.C2(n_2026),
.Y(n_3154)
);

OAI22xp5_ASAP7_75t_L g3155 ( 
.A1(n_3115),
.A2(n_2039),
.B1(n_2045),
.B2(n_2050),
.Y(n_3155)
);

OAI221xp5_ASAP7_75t_SL g3156 ( 
.A1(n_3117),
.A2(n_2031),
.B1(n_1868),
.B2(n_2045),
.C(n_2000),
.Y(n_3156)
);

NOR2x1_ASAP7_75t_L g3157 ( 
.A(n_3096),
.B(n_3103),
.Y(n_3157)
);

AOI21xp33_ASAP7_75t_L g3158 ( 
.A1(n_3091),
.A2(n_2220),
.B(n_2169),
.Y(n_3158)
);

AOI211xp5_ASAP7_75t_L g3159 ( 
.A1(n_3119),
.A2(n_2039),
.B(n_2179),
.C(n_2202),
.Y(n_3159)
);

OAI221xp5_ASAP7_75t_L g3160 ( 
.A1(n_3104),
.A2(n_2032),
.B1(n_2029),
.B2(n_2010),
.C(n_1997),
.Y(n_3160)
);

O2A1O1Ixp33_ASAP7_75t_L g3161 ( 
.A1(n_3126),
.A2(n_3123),
.B(n_3128),
.C(n_3121),
.Y(n_3161)
);

NOR3xp33_ASAP7_75t_L g3162 ( 
.A(n_3122),
.B(n_3116),
.C(n_3106),
.Y(n_3162)
);

NAND2xp5_ASAP7_75t_L g3163 ( 
.A(n_3131),
.B(n_3114),
.Y(n_3163)
);

OAI22xp5_ASAP7_75t_L g3164 ( 
.A1(n_3137),
.A2(n_3098),
.B1(n_3101),
.B2(n_3120),
.Y(n_3164)
);

OAI21xp33_ASAP7_75t_L g3165 ( 
.A1(n_3140),
.A2(n_3107),
.B(n_1868),
.Y(n_3165)
);

O2A1O1Ixp33_ASAP7_75t_L g3166 ( 
.A1(n_3135),
.A2(n_2220),
.B(n_1994),
.C(n_2024),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_3129),
.Y(n_3167)
);

BUFx2_ASAP7_75t_L g3168 ( 
.A(n_3157),
.Y(n_3168)
);

AOI222xp33_ASAP7_75t_L g3169 ( 
.A1(n_3124),
.A2(n_2029),
.B1(n_2032),
.B2(n_1997),
.C1(n_1994),
.C2(n_2001),
.Y(n_3169)
);

AOI221xp5_ASAP7_75t_L g3170 ( 
.A1(n_3125),
.A2(n_1857),
.B1(n_1864),
.B2(n_1869),
.C(n_1876),
.Y(n_3170)
);

NOR2x1_ASAP7_75t_L g3171 ( 
.A(n_3139),
.B(n_1173),
.Y(n_3171)
);

AOI221xp5_ASAP7_75t_L g3172 ( 
.A1(n_3127),
.A2(n_1857),
.B1(n_1864),
.B2(n_1869),
.C(n_1876),
.Y(n_3172)
);

AOI211xp5_ASAP7_75t_L g3173 ( 
.A1(n_3134),
.A2(n_2202),
.B(n_2125),
.C(n_2058),
.Y(n_3173)
);

INVx1_ASAP7_75t_L g3174 ( 
.A(n_3138),
.Y(n_3174)
);

OAI221xp5_ASAP7_75t_L g3175 ( 
.A1(n_3142),
.A2(n_2010),
.B1(n_2018),
.B2(n_2024),
.C(n_1994),
.Y(n_3175)
);

OAI221xp5_ASAP7_75t_SL g3176 ( 
.A1(n_3151),
.A2(n_2035),
.B1(n_2018),
.B2(n_2024),
.C(n_2001),
.Y(n_3176)
);

AOI21xp5_ASAP7_75t_L g3177 ( 
.A1(n_3148),
.A2(n_1932),
.B(n_2125),
.Y(n_3177)
);

AOI211xp5_ASAP7_75t_L g3178 ( 
.A1(n_3132),
.A2(n_2058),
.B(n_2055),
.C(n_2051),
.Y(n_3178)
);

AOI221xp5_ASAP7_75t_L g3179 ( 
.A1(n_3152),
.A2(n_2010),
.B1(n_2035),
.B2(n_1997),
.C(n_2001),
.Y(n_3179)
);

INVxp33_ASAP7_75t_SL g3180 ( 
.A(n_3149),
.Y(n_3180)
);

NOR2x1_ASAP7_75t_L g3181 ( 
.A(n_3143),
.B(n_1173),
.Y(n_3181)
);

AOI211xp5_ASAP7_75t_L g3182 ( 
.A1(n_3156),
.A2(n_3145),
.B(n_3158),
.C(n_3155),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3150),
.Y(n_3183)
);

OAI21xp5_ASAP7_75t_L g3184 ( 
.A1(n_3153),
.A2(n_3144),
.B(n_3133),
.Y(n_3184)
);

OAI221xp5_ASAP7_75t_SL g3185 ( 
.A1(n_3130),
.A2(n_2003),
.B1(n_2041),
.B2(n_2035),
.C(n_2018),
.Y(n_3185)
);

AOI22xp33_ASAP7_75t_L g3186 ( 
.A1(n_3154),
.A2(n_1932),
.B1(n_2191),
.B2(n_1165),
.Y(n_3186)
);

AOI221xp5_ASAP7_75t_L g3187 ( 
.A1(n_3159),
.A2(n_3160),
.B1(n_3147),
.B2(n_3153),
.C(n_3136),
.Y(n_3187)
);

NOR4xp25_ASAP7_75t_L g3188 ( 
.A(n_3141),
.B(n_3146),
.C(n_2041),
.D(n_2003),
.Y(n_3188)
);

BUFx8_ASAP7_75t_SL g3189 ( 
.A(n_3138),
.Y(n_3189)
);

AOI21xp5_ASAP7_75t_L g3190 ( 
.A1(n_3126),
.A2(n_2191),
.B(n_1932),
.Y(n_3190)
);

OAI211xp5_ASAP7_75t_SL g3191 ( 
.A1(n_3123),
.A2(n_1978),
.B(n_1984),
.C(n_2003),
.Y(n_3191)
);

INVx1_ASAP7_75t_L g3192 ( 
.A(n_3129),
.Y(n_3192)
);

NAND4xp25_ASAP7_75t_L g3193 ( 
.A(n_3124),
.B(n_1165),
.C(n_1151),
.D(n_1145),
.Y(n_3193)
);

AOI322xp5_ASAP7_75t_L g3194 ( 
.A1(n_3124),
.A2(n_2055),
.A3(n_2051),
.B1(n_2034),
.B2(n_2014),
.C1(n_2041),
.C2(n_1978),
.Y(n_3194)
);

A2O1A1Ixp33_ASAP7_75t_L g3195 ( 
.A1(n_3126),
.A2(n_2014),
.B(n_2034),
.C(n_1881),
.Y(n_3195)
);

NOR2xp67_ASAP7_75t_L g3196 ( 
.A(n_3174),
.B(n_2014),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3168),
.Y(n_3197)
);

OAI322xp33_ASAP7_75t_L g3198 ( 
.A1(n_3163),
.A2(n_2014),
.A3(n_2034),
.B1(n_1984),
.B2(n_1874),
.C1(n_1967),
.C2(n_1881),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_3161),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_SL g3200 ( 
.A(n_3187),
.B(n_2034),
.Y(n_3200)
);

NAND2xp5_ASAP7_75t_L g3201 ( 
.A(n_3165),
.B(n_1850),
.Y(n_3201)
);

AOI21xp5_ASAP7_75t_L g3202 ( 
.A1(n_3164),
.A2(n_2191),
.B(n_1932),
.Y(n_3202)
);

NAND2x1p5_ASAP7_75t_L g3203 ( 
.A(n_3167),
.B(n_1151),
.Y(n_3203)
);

A2O1A1Ixp33_ASAP7_75t_L g3204 ( 
.A1(n_3184),
.A2(n_1896),
.B(n_1892),
.C(n_1891),
.Y(n_3204)
);

NAND2xp5_ASAP7_75t_L g3205 ( 
.A(n_3162),
.B(n_1850),
.Y(n_3205)
);

AOI221xp5_ASAP7_75t_L g3206 ( 
.A1(n_3193),
.A2(n_1934),
.B1(n_1881),
.B2(n_1882),
.C(n_1883),
.Y(n_3206)
);

NOR2xp33_ASAP7_75t_L g3207 ( 
.A(n_3189),
.B(n_1159),
.Y(n_3207)
);

NOR2x1_ASAP7_75t_L g3208 ( 
.A(n_3192),
.B(n_1159),
.Y(n_3208)
);

INVx1_ASAP7_75t_L g3209 ( 
.A(n_3171),
.Y(n_3209)
);

OAI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_3183),
.A2(n_1968),
.B1(n_1882),
.B2(n_1883),
.Y(n_3210)
);

AOI22xp5_ASAP7_75t_L g3211 ( 
.A1(n_3180),
.A2(n_1931),
.B1(n_1980),
.B2(n_1976),
.Y(n_3211)
);

NAND3xp33_ASAP7_75t_SL g3212 ( 
.A(n_3182),
.B(n_1882),
.C(n_1980),
.Y(n_3212)
);

AOI321xp33_ASAP7_75t_L g3213 ( 
.A1(n_3195),
.A2(n_1165),
.A3(n_1980),
.B1(n_1976),
.B2(n_1972),
.C(n_1968),
.Y(n_3213)
);

OAI221xp5_ASAP7_75t_L g3214 ( 
.A1(n_3176),
.A2(n_1928),
.B1(n_1976),
.B2(n_1972),
.C(n_1968),
.Y(n_3214)
);

AOI221xp5_ASAP7_75t_L g3215 ( 
.A1(n_3188),
.A2(n_1928),
.B1(n_1874),
.B2(n_1883),
.C(n_1891),
.Y(n_3215)
);

AOI21xp5_ASAP7_75t_L g3216 ( 
.A1(n_3181),
.A2(n_1927),
.B(n_1972),
.Y(n_3216)
);

BUFx2_ASAP7_75t_L g3217 ( 
.A(n_3170),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3185),
.B(n_3186),
.Y(n_3218)
);

NOR2x1p5_ASAP7_75t_L g3219 ( 
.A(n_3194),
.B(n_1045),
.Y(n_3219)
);

AOI21xp5_ASAP7_75t_L g3220 ( 
.A1(n_3190),
.A2(n_1874),
.B(n_1967),
.Y(n_3220)
);

AOI221xp5_ASAP7_75t_L g3221 ( 
.A1(n_3191),
.A2(n_1931),
.B1(n_1891),
.B2(n_1892),
.C(n_1896),
.Y(n_3221)
);

NOR3xp33_ASAP7_75t_SL g3222 ( 
.A(n_3212),
.B(n_3172),
.C(n_3177),
.Y(n_3222)
);

NAND5xp2_ASAP7_75t_L g3223 ( 
.A(n_3197),
.B(n_3169),
.C(n_3173),
.D(n_3166),
.E(n_3177),
.Y(n_3223)
);

OR2x2_ASAP7_75t_L g3224 ( 
.A(n_3199),
.B(n_3209),
.Y(n_3224)
);

NAND2x1p5_ASAP7_75t_SL g3225 ( 
.A(n_3200),
.B(n_3178),
.Y(n_3225)
);

NOR3x2_ASAP7_75t_L g3226 ( 
.A(n_3218),
.B(n_3175),
.C(n_3179),
.Y(n_3226)
);

NOR3xp33_ASAP7_75t_L g3227 ( 
.A(n_3207),
.B(n_3217),
.C(n_3205),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_3219),
.A2(n_2036),
.B1(n_1059),
.B2(n_1073),
.Y(n_3228)
);

NAND4xp25_ASAP7_75t_L g3229 ( 
.A(n_3208),
.B(n_3201),
.C(n_3196),
.D(n_3204),
.Y(n_3229)
);

INVx2_ASAP7_75t_SL g3230 ( 
.A(n_3203),
.Y(n_3230)
);

NAND3xp33_ASAP7_75t_SL g3231 ( 
.A(n_3213),
.B(n_1896),
.C(n_1967),
.Y(n_3231)
);

INVx2_ASAP7_75t_L g3232 ( 
.A(n_3211),
.Y(n_3232)
);

INVx1_ASAP7_75t_L g3233 ( 
.A(n_3210),
.Y(n_3233)
);

AOI221xp5_ASAP7_75t_SL g3234 ( 
.A1(n_3198),
.A2(n_1966),
.B1(n_1892),
.B2(n_1903),
.C(n_1908),
.Y(n_3234)
);

NAND2xp5_ASAP7_75t_L g3235 ( 
.A(n_3216),
.B(n_1850),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3202),
.Y(n_3236)
);

OAI211xp5_ASAP7_75t_SL g3237 ( 
.A1(n_3220),
.A2(n_3215),
.B(n_3206),
.C(n_3214),
.Y(n_3237)
);

OAI221xp5_ASAP7_75t_L g3238 ( 
.A1(n_3221),
.A2(n_1931),
.B1(n_1966),
.B2(n_1949),
.C(n_1938),
.Y(n_3238)
);

NOR2x1_ASAP7_75t_L g3239 ( 
.A(n_3197),
.B(n_1903),
.Y(n_3239)
);

INVx1_ASAP7_75t_L g3240 ( 
.A(n_3197),
.Y(n_3240)
);

NAND5xp2_ASAP7_75t_L g3241 ( 
.A(n_3197),
.B(n_1431),
.C(n_1596),
.D(n_1589),
.E(n_1588),
.Y(n_3241)
);

CKINVDCx5p33_ASAP7_75t_R g3242 ( 
.A(n_3240),
.Y(n_3242)
);

AND2x2_ASAP7_75t_L g3243 ( 
.A(n_3227),
.B(n_1928),
.Y(n_3243)
);

NAND2xp33_ASAP7_75t_SL g3244 ( 
.A(n_3222),
.B(n_1045),
.Y(n_3244)
);

INVx1_ASAP7_75t_L g3245 ( 
.A(n_3224),
.Y(n_3245)
);

NOR3xp33_ASAP7_75t_L g3246 ( 
.A(n_3230),
.B(n_1511),
.C(n_1966),
.Y(n_3246)
);

CKINVDCx5p33_ASAP7_75t_R g3247 ( 
.A(n_3233),
.Y(n_3247)
);

BUFx6f_ASAP7_75t_L g3248 ( 
.A(n_3232),
.Y(n_3248)
);

CKINVDCx14_ASAP7_75t_R g3249 ( 
.A(n_3236),
.Y(n_3249)
);

HB1xp67_ASAP7_75t_L g3250 ( 
.A(n_3239),
.Y(n_3250)
);

OAI21xp33_ASAP7_75t_SL g3251 ( 
.A1(n_3229),
.A2(n_1908),
.B(n_1949),
.Y(n_3251)
);

INVx1_ASAP7_75t_SL g3252 ( 
.A(n_3226),
.Y(n_3252)
);

NOR2xp67_ASAP7_75t_L g3253 ( 
.A(n_3223),
.B(n_1903),
.Y(n_3253)
);

INVx1_ASAP7_75t_SL g3254 ( 
.A(n_3235),
.Y(n_3254)
);

NAND2xp33_ASAP7_75t_R g3255 ( 
.A(n_3225),
.B(n_2036),
.Y(n_3255)
);

INVx1_ASAP7_75t_L g3256 ( 
.A(n_3229),
.Y(n_3256)
);

INVx2_ASAP7_75t_L g3257 ( 
.A(n_3238),
.Y(n_3257)
);

OAI211xp5_ASAP7_75t_L g3258 ( 
.A1(n_3237),
.A2(n_1908),
.B(n_1916),
.C(n_1927),
.Y(n_3258)
);

INVx2_ASAP7_75t_L g3259 ( 
.A(n_3234),
.Y(n_3259)
);

CKINVDCx5p33_ASAP7_75t_R g3260 ( 
.A(n_3228),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_3250),
.Y(n_3261)
);

XOR2xp5_ASAP7_75t_L g3262 ( 
.A(n_3247),
.B(n_3231),
.Y(n_3262)
);

INVx4_ASAP7_75t_L g3263 ( 
.A(n_3248),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3245),
.Y(n_3264)
);

AOI221xp5_ASAP7_75t_L g3265 ( 
.A1(n_3244),
.A2(n_3241),
.B1(n_1949),
.B2(n_1938),
.C(n_1934),
.Y(n_3265)
);

AO21x2_ASAP7_75t_L g3266 ( 
.A1(n_3256),
.A2(n_1938),
.B(n_1934),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3248),
.Y(n_3267)
);

XOR2xp5_ASAP7_75t_L g3268 ( 
.A(n_3242),
.B(n_1045),
.Y(n_3268)
);

INVx1_ASAP7_75t_L g3269 ( 
.A(n_3248),
.Y(n_3269)
);

BUFx2_ASAP7_75t_L g3270 ( 
.A(n_3249),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3253),
.Y(n_3271)
);

INVx1_ASAP7_75t_L g3272 ( 
.A(n_3243),
.Y(n_3272)
);

AOI22x1_ASAP7_75t_L g3273 ( 
.A1(n_3252),
.A2(n_1045),
.B1(n_1059),
.B2(n_1073),
.Y(n_3273)
);

INVx1_ASAP7_75t_L g3274 ( 
.A(n_3259),
.Y(n_3274)
);

OAI22xp5_ASAP7_75t_L g3275 ( 
.A1(n_3260),
.A2(n_1927),
.B1(n_1916),
.B2(n_2036),
.Y(n_3275)
);

OAI22xp5_ASAP7_75t_SL g3276 ( 
.A1(n_3257),
.A2(n_1059),
.B1(n_1073),
.B2(n_1075),
.Y(n_3276)
);

AO21x2_ASAP7_75t_L g3277 ( 
.A1(n_3246),
.A2(n_1916),
.B(n_1595),
.Y(n_3277)
);

AND2x4_ASAP7_75t_L g3278 ( 
.A(n_3263),
.B(n_3254),
.Y(n_3278)
);

OAI22xp5_ASAP7_75t_SL g3279 ( 
.A1(n_3270),
.A2(n_3254),
.B1(n_3255),
.B2(n_3251),
.Y(n_3279)
);

BUFx2_ASAP7_75t_SL g3280 ( 
.A(n_3270),
.Y(n_3280)
);

AOI22xp5_ASAP7_75t_L g3281 ( 
.A1(n_3264),
.A2(n_3258),
.B1(n_2036),
.B2(n_1084),
.Y(n_3281)
);

OAI21xp5_ASAP7_75t_L g3282 ( 
.A1(n_3267),
.A2(n_1416),
.B(n_1414),
.Y(n_3282)
);

BUFx2_ASAP7_75t_L g3283 ( 
.A(n_3269),
.Y(n_3283)
);

OAI22xp5_ASAP7_75t_L g3284 ( 
.A1(n_3261),
.A2(n_1073),
.B1(n_1075),
.B2(n_1084),
.Y(n_3284)
);

OAI21xp5_ASAP7_75t_L g3285 ( 
.A1(n_3262),
.A2(n_1416),
.B(n_1414),
.Y(n_3285)
);

HB1xp67_ASAP7_75t_L g3286 ( 
.A(n_3271),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_3268),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_3266),
.Y(n_3288)
);

INVx2_ASAP7_75t_L g3289 ( 
.A(n_3273),
.Y(n_3289)
);

NAND2xp5_ASAP7_75t_L g3290 ( 
.A(n_3274),
.B(n_1850),
.Y(n_3290)
);

OAI22xp5_ASAP7_75t_L g3291 ( 
.A1(n_3272),
.A2(n_1073),
.B1(n_1075),
.B2(n_1084),
.Y(n_3291)
);

OAI22xp5_ASAP7_75t_L g3292 ( 
.A1(n_3276),
.A2(n_1075),
.B1(n_1084),
.B2(n_1095),
.Y(n_3292)
);

OR3x1_ASAP7_75t_L g3293 ( 
.A(n_3277),
.B(n_1431),
.C(n_1583),
.Y(n_3293)
);

INVx1_ASAP7_75t_L g3294 ( 
.A(n_3280),
.Y(n_3294)
);

HB1xp67_ASAP7_75t_L g3295 ( 
.A(n_3283),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_3279),
.Y(n_3296)
);

INVxp67_ASAP7_75t_SL g3297 ( 
.A(n_3286),
.Y(n_3297)
);

INVx1_ASAP7_75t_L g3298 ( 
.A(n_3278),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_3278),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3288),
.Y(n_3300)
);

INVx1_ASAP7_75t_L g3301 ( 
.A(n_3289),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3287),
.Y(n_3302)
);

INVx1_ASAP7_75t_L g3303 ( 
.A(n_3290),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3293),
.Y(n_3304)
);

OAI22xp5_ASAP7_75t_L g3305 ( 
.A1(n_3294),
.A2(n_3281),
.B1(n_3284),
.B2(n_3291),
.Y(n_3305)
);

NOR2x1p5_ASAP7_75t_L g3306 ( 
.A(n_3297),
.B(n_3292),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3295),
.Y(n_3307)
);

HB1xp67_ASAP7_75t_L g3308 ( 
.A(n_3297),
.Y(n_3308)
);

OAI22xp5_ASAP7_75t_L g3309 ( 
.A1(n_3298),
.A2(n_3265),
.B1(n_3285),
.B2(n_3282),
.Y(n_3309)
);

AOI22xp5_ASAP7_75t_L g3310 ( 
.A1(n_3299),
.A2(n_3275),
.B1(n_1084),
.B2(n_1095),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3296),
.Y(n_3311)
);

INVxp67_ASAP7_75t_SL g3312 ( 
.A(n_3308),
.Y(n_3312)
);

INVxp67_ASAP7_75t_L g3313 ( 
.A(n_3307),
.Y(n_3313)
);

OAI21x1_ASAP7_75t_SL g3314 ( 
.A1(n_3311),
.A2(n_3304),
.B(n_3301),
.Y(n_3314)
);

OAI221xp5_ASAP7_75t_L g3315 ( 
.A1(n_3312),
.A2(n_3300),
.B1(n_3302),
.B2(n_3309),
.C(n_3310),
.Y(n_3315)
);

O2A1O1Ixp33_ASAP7_75t_L g3316 ( 
.A1(n_3313),
.A2(n_3303),
.B(n_3305),
.C(n_3306),
.Y(n_3316)
);

AOI22xp33_ASAP7_75t_L g3317 ( 
.A1(n_3315),
.A2(n_3314),
.B1(n_1095),
.B2(n_1104),
.Y(n_3317)
);

AOI322xp5_ASAP7_75t_R g3318 ( 
.A1(n_3316),
.A2(n_1431),
.A3(n_1595),
.B1(n_1410),
.B2(n_1413),
.C1(n_1154),
.C2(n_1156),
.Y(n_3318)
);

AOI22xp5_ASAP7_75t_L g3319 ( 
.A1(n_3317),
.A2(n_1075),
.B1(n_1095),
.B2(n_1104),
.Y(n_3319)
);

AOI21xp5_ASAP7_75t_SL g3320 ( 
.A1(n_3319),
.A2(n_3318),
.B(n_1104),
.Y(n_3320)
);

AOI21xp5_ASAP7_75t_L g3321 ( 
.A1(n_3320),
.A2(n_1095),
.B(n_1104),
.Y(n_3321)
);

AOI211xp5_ASAP7_75t_L g3322 ( 
.A1(n_3321),
.A2(n_1104),
.B(n_1132),
.C(n_1154),
.Y(n_3322)
);


endmodule