module fake_netlist_5_2220_n_511 (n_137, n_91, n_82, n_122, n_142, n_10, n_140, n_24, n_124, n_86, n_136, n_146, n_143, n_83, n_132, n_61, n_90, n_127, n_75, n_101, n_65, n_78, n_74, n_144, n_114, n_57, n_96, n_37, n_111, n_108, n_129, n_31, n_13, n_66, n_98, n_60, n_155, n_152, n_16, n_43, n_107, n_0, n_58, n_9, n_69, n_18, n_116, n_42, n_22, n_1, n_45, n_117, n_46, n_21, n_94, n_113, n_38, n_123, n_139, n_105, n_80, n_4, n_125, n_35, n_128, n_73, n_17, n_92, n_19, n_149, n_120, n_135, n_30, n_156, n_5, n_33, n_126, n_14, n_84, n_23, n_130, n_157, n_29, n_79, n_131, n_151, n_47, n_25, n_53, n_8, n_158, n_44, n_40, n_34, n_100, n_62, n_138, n_148, n_71, n_154, n_109, n_112, n_85, n_95, n_119, n_59, n_26, n_133, n_55, n_99, n_2, n_3, n_49, n_20, n_6, n_39, n_54, n_147, n_12, n_67, n_121, n_36, n_76, n_87, n_150, n_27, n_64, n_77, n_102, n_106, n_81, n_118, n_28, n_89, n_70, n_115, n_68, n_93, n_72, n_134, n_32, n_41, n_104, n_103, n_56, n_51, n_63, n_97, n_141, n_11, n_153, n_7, n_15, n_145, n_48, n_50, n_52, n_88, n_110, n_511);

input n_137;
input n_91;
input n_82;
input n_122;
input n_142;
input n_10;
input n_140;
input n_24;
input n_124;
input n_86;
input n_136;
input n_146;
input n_143;
input n_83;
input n_132;
input n_61;
input n_90;
input n_127;
input n_75;
input n_101;
input n_65;
input n_78;
input n_74;
input n_144;
input n_114;
input n_57;
input n_96;
input n_37;
input n_111;
input n_108;
input n_129;
input n_31;
input n_13;
input n_66;
input n_98;
input n_60;
input n_155;
input n_152;
input n_16;
input n_43;
input n_107;
input n_0;
input n_58;
input n_9;
input n_69;
input n_18;
input n_116;
input n_42;
input n_22;
input n_1;
input n_45;
input n_117;
input n_46;
input n_21;
input n_94;
input n_113;
input n_38;
input n_123;
input n_139;
input n_105;
input n_80;
input n_4;
input n_125;
input n_35;
input n_128;
input n_73;
input n_17;
input n_92;
input n_19;
input n_149;
input n_120;
input n_135;
input n_30;
input n_156;
input n_5;
input n_33;
input n_126;
input n_14;
input n_84;
input n_23;
input n_130;
input n_157;
input n_29;
input n_79;
input n_131;
input n_151;
input n_47;
input n_25;
input n_53;
input n_8;
input n_158;
input n_44;
input n_40;
input n_34;
input n_100;
input n_62;
input n_138;
input n_148;
input n_71;
input n_154;
input n_109;
input n_112;
input n_85;
input n_95;
input n_119;
input n_59;
input n_26;
input n_133;
input n_55;
input n_99;
input n_2;
input n_3;
input n_49;
input n_20;
input n_6;
input n_39;
input n_54;
input n_147;
input n_12;
input n_67;
input n_121;
input n_36;
input n_76;
input n_87;
input n_150;
input n_27;
input n_64;
input n_77;
input n_102;
input n_106;
input n_81;
input n_118;
input n_28;
input n_89;
input n_70;
input n_115;
input n_68;
input n_93;
input n_72;
input n_134;
input n_32;
input n_41;
input n_104;
input n_103;
input n_56;
input n_51;
input n_63;
input n_97;
input n_141;
input n_11;
input n_153;
input n_7;
input n_15;
input n_145;
input n_48;
input n_50;
input n_52;
input n_88;
input n_110;

output n_511;

wire n_294;
wire n_431;
wire n_318;
wire n_380;
wire n_419;
wire n_444;
wire n_469;
wire n_194;
wire n_316;
wire n_389;
wire n_418;
wire n_248;
wire n_315;
wire n_268;
wire n_451;
wire n_408;
wire n_376;
wire n_503;
wire n_235;
wire n_226;
wire n_353;
wire n_351;
wire n_367;
wire n_452;
wire n_397;
wire n_493;
wire n_483;
wire n_467;
wire n_423;
wire n_284;
wire n_245;
wire n_501;
wire n_280;
wire n_378;
wire n_382;
wire n_254;
wire n_302;
wire n_265;
wire n_293;
wire n_372;
wire n_443;
wire n_244;
wire n_173;
wire n_198;
wire n_447;
wire n_247;
wire n_314;
wire n_368;
wire n_433;
wire n_321;
wire n_292;
wire n_455;
wire n_417;
wire n_212;
wire n_385;
wire n_498;
wire n_507;
wire n_497;
wire n_275;
wire n_252;
wire n_295;
wire n_330;
wire n_508;
wire n_506;
wire n_509;
wire n_373;
wire n_307;
wire n_439;
wire n_209;
wire n_259;
wire n_448;
wire n_375;
wire n_301;
wire n_186;
wire n_191;
wire n_492;
wire n_171;
wire n_399;
wire n_341;
wire n_204;
wire n_394;
wire n_250;
wire n_260;
wire n_298;
wire n_320;
wire n_505;
wire n_286;
wire n_282;
wire n_331;
wire n_406;
wire n_470;
wire n_325;
wire n_449;
wire n_281;
wire n_240;
wire n_381;
wire n_189;
wire n_220;
wire n_291;
wire n_231;
wire n_257;
wire n_390;
wire n_456;
wire n_371;
wire n_481;
wire n_317;
wire n_323;
wire n_195;
wire n_356;
wire n_227;
wire n_271;
wire n_335;
wire n_370;
wire n_167;
wire n_234;
wire n_343;
wire n_379;
wire n_308;
wire n_428;
wire n_267;
wire n_457;
wire n_297;
wire n_225;
wire n_377;
wire n_484;
wire n_219;
wire n_442;
wire n_192;
wire n_223;
wire n_392;
wire n_264;
wire n_472;
wire n_454;
wire n_387;
wire n_374;
wire n_163;
wire n_276;
wire n_339;
wire n_185;
wire n_183;
wire n_243;
wire n_398;
wire n_396;
wire n_347;
wire n_169;
wire n_255;
wire n_215;
wire n_350;
wire n_196;
wire n_459;
wire n_211;
wire n_218;
wire n_400;
wire n_181;
wire n_436;
wire n_290;
wire n_221;
wire n_178;
wire n_386;
wire n_287;
wire n_344;
wire n_473;
wire n_422;
wire n_475;
wire n_415;
wire n_485;
wire n_496;
wire n_355;
wire n_486;
wire n_336;
wire n_337;
wire n_430;
wire n_313;
wire n_479;
wire n_510;
wire n_216;
wire n_168;
wire n_395;
wire n_164;
wire n_432;
wire n_311;
wire n_208;
wire n_328;
wire n_214;
wire n_299;
wire n_303;
wire n_369;
wire n_296;
wire n_241;
wire n_357;
wire n_184;
wire n_446;
wire n_445;
wire n_165;
wire n_468;
wire n_499;
wire n_213;
wire n_342;
wire n_482;
wire n_361;
wire n_464;
wire n_363;
wire n_402;
wire n_413;
wire n_197;
wire n_236;
wire n_388;
wire n_249;
wire n_304;
wire n_329;
wire n_203;
wire n_274;
wire n_384;
wire n_460;
wire n_277;
wire n_338;
wire n_477;
wire n_461;
wire n_333;
wire n_309;
wire n_462;
wire n_322;
wire n_258;
wire n_306;
wire n_458;
wire n_288;
wire n_188;
wire n_190;
wire n_201;
wire n_263;
wire n_471;
wire n_224;
wire n_228;
wire n_283;
wire n_383;
wire n_474;
wire n_463;
wire n_488;
wire n_502;
wire n_239;
wire n_466;
wire n_420;
wire n_489;
wire n_310;
wire n_504;
wire n_465;
wire n_358;
wire n_362;
wire n_170;
wire n_332;
wire n_161;
wire n_273;
wire n_349;
wire n_270;
wire n_230;
wire n_279;
wire n_253;
wire n_261;
wire n_174;
wire n_289;
wire n_206;
wire n_172;
wire n_217;
wire n_440;
wire n_478;
wire n_441;
wire n_450;
wire n_312;
wire n_476;
wire n_429;
wire n_345;
wire n_210;
wire n_494;
wire n_365;
wire n_176;
wire n_182;
wire n_354;
wire n_480;
wire n_237;
wire n_425;
wire n_407;
wire n_180;
wire n_340;
wire n_207;
wire n_346;
wire n_393;
wire n_229;
wire n_487;
wire n_495;
wire n_437;
wire n_177;
wire n_403;
wire n_453;
wire n_421;
wire n_405;
wire n_359;
wire n_490;
wire n_326;
wire n_233;
wire n_404;
wire n_205;
wire n_366;
wire n_246;
wire n_179;
wire n_410;
wire n_269;
wire n_285;
wire n_412;
wire n_232;
wire n_327;
wire n_202;
wire n_266;
wire n_272;
wire n_491;
wire n_427;
wire n_193;
wire n_251;
wire n_352;
wire n_160;
wire n_426;
wire n_409;
wire n_500;
wire n_300;
wire n_435;
wire n_159;
wire n_334;
wire n_391;
wire n_434;
wire n_175;
wire n_262;
wire n_238;
wire n_411;
wire n_414;
wire n_319;
wire n_364;
wire n_242;
wire n_360;
wire n_200;
wire n_162;
wire n_222;
wire n_438;
wire n_324;
wire n_416;
wire n_199;
wire n_187;
wire n_401;
wire n_348;
wire n_166;
wire n_424;
wire n_256;
wire n_305;
wire n_278;

INVx2_ASAP7_75t_L g159 ( 
.A(n_146),
.Y(n_159)
);

INVx1_ASAP7_75t_SL g160 ( 
.A(n_77),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g161 ( 
.A(n_86),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_101),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_79),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_53),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g166 ( 
.A(n_60),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_23),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_115),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_125),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_102),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_17),
.Y(n_171)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_112),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_43),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_26),
.Y(n_174)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_74),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_58),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g177 ( 
.A(n_98),
.Y(n_177)
);

BUFx10_ASAP7_75t_L g178 ( 
.A(n_18),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g179 ( 
.A(n_88),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_49),
.Y(n_180)
);

BUFx5_ASAP7_75t_L g181 ( 
.A(n_113),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_122),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_118),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_34),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_54),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_148),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_132),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_92),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_127),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_130),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_129),
.Y(n_191)
);

BUFx6f_ASAP7_75t_L g192 ( 
.A(n_80),
.Y(n_192)
);

CKINVDCx5p33_ASAP7_75t_R g193 ( 
.A(n_105),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_48),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g195 ( 
.A(n_52),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_4),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g197 ( 
.A(n_69),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_27),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g199 ( 
.A(n_76),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_135),
.Y(n_200)
);

INVx1_ASAP7_75t_SL g201 ( 
.A(n_56),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_110),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_39),
.Y(n_203)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_111),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_95),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_158),
.Y(n_206)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_19),
.Y(n_207)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_89),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_96),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_82),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_5),
.Y(n_211)
);

INVx2_ASAP7_75t_SL g212 ( 
.A(n_156),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_119),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_104),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_9),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_30),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_25),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_6),
.Y(n_218)
);

INVx2_ASAP7_75t_L g219 ( 
.A(n_153),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_70),
.Y(n_220)
);

INVx2_ASAP7_75t_SL g221 ( 
.A(n_67),
.Y(n_221)
);

CKINVDCx5p33_ASAP7_75t_R g222 ( 
.A(n_90),
.Y(n_222)
);

BUFx10_ASAP7_75t_L g223 ( 
.A(n_123),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_84),
.Y(n_224)
);

INVxp67_ASAP7_75t_SL g225 ( 
.A(n_61),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_56),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_59),
.Y(n_227)
);

INVx2_ASAP7_75t_SL g228 ( 
.A(n_117),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_57),
.Y(n_229)
);

INVx1_ASAP7_75t_SL g230 ( 
.A(n_32),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_100),
.Y(n_231)
);

INVx2_ASAP7_75t_SL g232 ( 
.A(n_83),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_81),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_78),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_109),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_121),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_87),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_93),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_97),
.Y(n_239)
);

BUFx10_ASAP7_75t_L g240 ( 
.A(n_157),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_120),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_72),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_124),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_91),
.Y(n_244)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_75),
.Y(n_245)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_35),
.Y(n_246)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_85),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_11),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_107),
.Y(n_249)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

INVx2_ASAP7_75t_L g251 ( 
.A(n_64),
.Y(n_251)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_68),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_42),
.Y(n_253)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_128),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_31),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_106),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_103),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_150),
.Y(n_258)
);

INVx2_ASAP7_75t_L g259 ( 
.A(n_126),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_63),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_44),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_12),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_108),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_50),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_9),
.Y(n_265)
);

BUFx10_ASAP7_75t_L g266 ( 
.A(n_73),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_147),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_12),
.Y(n_268)
);

INVx2_ASAP7_75t_L g269 ( 
.A(n_52),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_141),
.Y(n_270)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_116),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_51),
.Y(n_272)
);

INVx1_ASAP7_75t_SL g273 ( 
.A(n_201),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_159),
.B(n_0),
.Y(n_274)
);

BUFx6f_ASAP7_75t_L g275 ( 
.A(n_161),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g276 ( 
.A(n_172),
.B(n_1),
.Y(n_276)
);

AND2x4_ASAP7_75t_L g277 ( 
.A(n_177),
.B(n_1),
.Y(n_277)
);

AND2x2_ASAP7_75t_L g278 ( 
.A(n_197),
.B(n_2),
.Y(n_278)
);

INVx2_ASAP7_75t_L g279 ( 
.A(n_181),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_159),
.B(n_3),
.Y(n_280)
);

INVx2_ASAP7_75t_SL g281 ( 
.A(n_178),
.Y(n_281)
);

BUFx6f_ASAP7_75t_L g282 ( 
.A(n_161),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_175),
.B(n_3),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_175),
.B(n_6),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_208),
.B(n_7),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_160),
.B(n_10),
.Y(n_286)
);

HB1xp67_ASAP7_75t_L g287 ( 
.A(n_207),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_208),
.B(n_10),
.Y(n_288)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_166),
.Y(n_289)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_219),
.B(n_62),
.Y(n_290)
);

AND2x2_ASAP7_75t_L g291 ( 
.A(n_179),
.B(n_271),
.Y(n_291)
);

BUFx6f_ASAP7_75t_L g292 ( 
.A(n_192),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g293 ( 
.A(n_247),
.B(n_13),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_185),
.Y(n_294)
);

AND2x4_ASAP7_75t_L g295 ( 
.A(n_251),
.B(n_14),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_223),
.B(n_14),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_SL g297 ( 
.A(n_223),
.B(n_15),
.Y(n_297)
);

AND2x4_ASAP7_75t_L g298 ( 
.A(n_252),
.B(n_16),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g299 ( 
.A(n_252),
.B(n_259),
.Y(n_299)
);

BUFx6f_ASAP7_75t_L g300 ( 
.A(n_259),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g301 ( 
.A(n_163),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_212),
.B(n_221),
.Y(n_302)
);

AND2x4_ASAP7_75t_L g303 ( 
.A(n_228),
.B(n_17),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_232),
.B(n_18),
.Y(n_304)
);

AND2x4_ASAP7_75t_L g305 ( 
.A(n_169),
.B(n_20),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_199),
.B(n_20),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_21),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g308 ( 
.A(n_269),
.B(n_22),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_225),
.B(n_22),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_226),
.B(n_24),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_170),
.B(n_24),
.Y(n_311)
);

BUFx2_ASAP7_75t_L g312 ( 
.A(n_165),
.Y(n_312)
);

BUFx12f_ASAP7_75t_L g313 ( 
.A(n_240),
.Y(n_313)
);

INVx4_ASAP7_75t_L g314 ( 
.A(n_266),
.Y(n_314)
);

BUFx12f_ASAP7_75t_L g315 ( 
.A(n_266),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_182),
.B(n_28),
.Y(n_316)
);

INVx5_ASAP7_75t_L g317 ( 
.A(n_167),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_183),
.B(n_29),
.Y(n_318)
);

AND2x4_ASAP7_75t_L g319 ( 
.A(n_188),
.B(n_31),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_202),
.B(n_205),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_210),
.Y(n_321)
);

AND2x2_ASAP7_75t_L g322 ( 
.A(n_230),
.B(n_32),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_213),
.B(n_33),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_224),
.B(n_237),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_239),
.B(n_34),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_243),
.B(n_36),
.Y(n_326)
);

INVx5_ASAP7_75t_L g327 ( 
.A(n_171),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_244),
.B(n_36),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_249),
.Y(n_329)
);

BUFx12f_ASAP7_75t_L g330 ( 
.A(n_173),
.Y(n_330)
);

BUFx12f_ASAP7_75t_L g331 ( 
.A(n_174),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_254),
.Y(n_332)
);

INVx5_ASAP7_75t_L g333 ( 
.A(n_176),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_180),
.B(n_37),
.Y(n_334)
);

INVx2_ASAP7_75t_SL g335 ( 
.A(n_194),
.Y(n_335)
);

INVx3_ASAP7_75t_L g336 ( 
.A(n_275),
.Y(n_336)
);

INVx2_ASAP7_75t_L g337 ( 
.A(n_275),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_275),
.Y(n_338)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_291),
.A2(n_204),
.B1(n_220),
.B2(n_162),
.Y(n_339)
);

INVx3_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g341 ( 
.A1(n_276),
.A2(n_198),
.B1(n_203),
.B2(n_196),
.Y(n_341)
);

AOI22xp5_ASAP7_75t_L g342 ( 
.A1(n_278),
.A2(n_234),
.B1(n_245),
.B2(n_164),
.Y(n_342)
);

OAI22xp33_ASAP7_75t_SL g343 ( 
.A1(n_276),
.A2(n_215),
.B1(n_216),
.B2(n_211),
.Y(n_343)
);

OAI22xp33_ASAP7_75t_L g344 ( 
.A1(n_273),
.A2(n_218),
.B1(n_227),
.B2(n_217),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_R g345 ( 
.A1(n_273),
.A2(n_246),
.B1(n_250),
.B2(n_229),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_314),
.B(n_234),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_306),
.A2(n_263),
.B1(n_248),
.B2(n_253),
.Y(n_347)
);

OAI22xp33_ASAP7_75t_SL g348 ( 
.A1(n_296),
.A2(n_261),
.B1(n_262),
.B2(n_255),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_286),
.A2(n_265),
.B1(n_268),
.B2(n_264),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_286),
.A2(n_272),
.B1(n_184),
.B2(n_195),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_312),
.B(n_168),
.Y(n_351)
);

OAI22xp33_ASAP7_75t_L g352 ( 
.A1(n_309),
.A2(n_187),
.B1(n_189),
.B2(n_186),
.Y(n_352)
);

OAI22xp33_ASAP7_75t_L g353 ( 
.A1(n_309),
.A2(n_191),
.B1(n_193),
.B2(n_190),
.Y(n_353)
);

OR2x6_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_37),
.Y(n_354)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_289),
.Y(n_355)
);

AND2x2_ASAP7_75t_L g356 ( 
.A(n_335),
.B(n_200),
.Y(n_356)
);

OAI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_297),
.A2(n_334),
.B1(n_304),
.B2(n_280),
.Y(n_357)
);

OAI22xp33_ASAP7_75t_L g358 ( 
.A1(n_304),
.A2(n_323),
.B1(n_328),
.B2(n_318),
.Y(n_358)
);

AO22x2_ASAP7_75t_L g359 ( 
.A1(n_277),
.A2(n_41),
.B1(n_38),
.B2(n_40),
.Y(n_359)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_331),
.A2(n_209),
.B1(n_214),
.B2(n_206),
.Y(n_360)
);

AOI22xp5_ASAP7_75t_L g361 ( 
.A1(n_322),
.A2(n_260),
.B1(n_270),
.B2(n_267),
.Y(n_361)
);

NOR2xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_222),
.Y(n_362)
);

OAI22xp33_ASAP7_75t_L g363 ( 
.A1(n_274),
.A2(n_283),
.B1(n_284),
.B2(n_280),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_281),
.A2(n_236),
.B1(n_257),
.B2(n_256),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_292),
.Y(n_365)
);

BUFx6f_ASAP7_75t_SL g366 ( 
.A(n_305),
.Y(n_366)
);

OAI22xp33_ASAP7_75t_L g367 ( 
.A1(n_284),
.A2(n_285),
.B1(n_293),
.B2(n_288),
.Y(n_367)
);

AO22x2_ASAP7_75t_L g368 ( 
.A1(n_303),
.A2(n_298),
.B1(n_295),
.B2(n_305),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_292),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_310),
.A2(n_258),
.B1(n_242),
.B2(n_241),
.Y(n_370)
);

AOI22xp5_ASAP7_75t_L g371 ( 
.A1(n_313),
.A2(n_235),
.B1(n_233),
.B2(n_231),
.Y(n_371)
);

OAI22xp33_ASAP7_75t_L g372 ( 
.A1(n_285),
.A2(n_238),
.B1(n_46),
.B2(n_47),
.Y(n_372)
);

INVx2_ASAP7_75t_SL g373 ( 
.A(n_317),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_315),
.A2(n_45),
.B1(n_46),
.B2(n_47),
.Y(n_374)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_317),
.B(n_65),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_368),
.A2(n_324),
.B(n_320),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_358),
.B(n_317),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_338),
.Y(n_378)
);

INVx2_ASAP7_75t_SL g379 ( 
.A(n_351),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_339),
.Y(n_380)
);

AOI21xp5_ASAP7_75t_L g381 ( 
.A1(n_368),
.A2(n_324),
.B(n_320),
.Y(n_381)
);

BUFx6f_ASAP7_75t_L g382 ( 
.A(n_337),
.Y(n_382)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_336),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_327),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_369),
.Y(n_385)
);

INVx2_ASAP7_75t_L g386 ( 
.A(n_340),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_340),
.Y(n_387)
);

INVxp33_ASAP7_75t_L g388 ( 
.A(n_350),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g389 ( 
.A(n_362),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_355),
.Y(n_390)
);

AND2x6_ASAP7_75t_L g391 ( 
.A(n_375),
.B(n_298),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_365),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_R g393 ( 
.A(n_354),
.B(n_319),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_L g394 ( 
.A(n_367),
.B(n_333),
.Y(n_394)
);

AND2x2_ASAP7_75t_SL g395 ( 
.A(n_342),
.B(n_319),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g396 ( 
.A(n_357),
.B(n_333),
.Y(n_396)
);

INVxp67_ASAP7_75t_SL g397 ( 
.A(n_372),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_366),
.Y(n_398)
);

NAND2xp33_ASAP7_75t_SL g399 ( 
.A(n_370),
.B(n_293),
.Y(n_399)
);

XOR2xp5_ASAP7_75t_L g400 ( 
.A(n_360),
.B(n_66),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_346),
.Y(n_401)
);

INVx2_ASAP7_75t_SL g402 ( 
.A(n_356),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_SL g403 ( 
.A(n_341),
.B(n_343),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g404 ( 
.A(n_347),
.Y(n_404)
);

INVxp33_ASAP7_75t_L g405 ( 
.A(n_349),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_359),
.Y(n_406)
);

INVx2_ASAP7_75t_L g407 ( 
.A(n_373),
.Y(n_407)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_361),
.Y(n_408)
);

AND2x2_ASAP7_75t_SL g409 ( 
.A(n_395),
.B(n_307),
.Y(n_409)
);

BUFx6f_ASAP7_75t_L g410 ( 
.A(n_382),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_378),
.Y(n_411)
);

AND2x2_ASAP7_75t_SL g412 ( 
.A(n_395),
.B(n_307),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_379),
.B(n_352),
.Y(n_413)
);

AND2x2_ASAP7_75t_L g414 ( 
.A(n_376),
.B(n_287),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_381),
.B(n_402),
.Y(n_415)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_399),
.A2(n_345),
.B1(n_316),
.B2(n_325),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_391),
.B(n_353),
.Y(n_417)
);

INVx2_ASAP7_75t_L g418 ( 
.A(n_385),
.Y(n_418)
);

BUFx6f_ASAP7_75t_L g419 ( 
.A(n_383),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g420 ( 
.A(n_377),
.B(n_348),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_396),
.B(n_299),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g422 ( 
.A(n_384),
.B(n_364),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_390),
.Y(n_423)
);

AND2x2_ASAP7_75t_L g424 ( 
.A(n_394),
.B(n_321),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g425 ( 
.A1(n_394),
.A2(n_325),
.B(n_311),
.Y(n_425)
);

AND2x2_ASAP7_75t_L g426 ( 
.A(n_397),
.B(n_329),
.Y(n_426)
);

AND2x4_ASAP7_75t_L g427 ( 
.A(n_392),
.B(n_290),
.Y(n_427)
);

INVx4_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

BUFx6f_ASAP7_75t_L g429 ( 
.A(n_387),
.Y(n_429)
);

NOR2xp33_ASAP7_75t_L g430 ( 
.A(n_405),
.B(n_371),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g431 ( 
.A(n_388),
.B(n_344),
.Y(n_431)
);

AND2x2_ASAP7_75t_SL g432 ( 
.A(n_403),
.B(n_308),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_406),
.B(n_332),
.Y(n_433)
);

HB1xp67_ASAP7_75t_L g434 ( 
.A(n_393),
.Y(n_434)
);

AND2x6_ASAP7_75t_L g435 ( 
.A(n_398),
.B(n_374),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_407),
.Y(n_436)
);

BUFx4f_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_415),
.B(n_401),
.Y(n_438)
);

INVx1_ASAP7_75t_L g439 ( 
.A(n_411),
.Y(n_439)
);

AND2x6_ASAP7_75t_L g440 ( 
.A(n_414),
.B(n_311),
.Y(n_440)
);

BUFx2_ASAP7_75t_L g441 ( 
.A(n_434),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g442 ( 
.A(n_414),
.B(n_300),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_L g443 ( 
.A(n_408),
.B(n_404),
.Y(n_443)
);

BUFx4f_ASAP7_75t_L g444 ( 
.A(n_435),
.Y(n_444)
);

NOR2xp33_ASAP7_75t_SL g445 ( 
.A(n_430),
.B(n_380),
.Y(n_445)
);

AND2x6_ASAP7_75t_L g446 ( 
.A(n_421),
.B(n_326),
.Y(n_446)
);

AND2x4_ASAP7_75t_L g447 ( 
.A(n_433),
.B(n_294),
.Y(n_447)
);

NOR2x1_ASAP7_75t_L g448 ( 
.A(n_417),
.B(n_400),
.Y(n_448)
);

NOR2xp33_ASAP7_75t_L g449 ( 
.A(n_422),
.B(n_301),
.Y(n_449)
);

BUFx6f_ASAP7_75t_L g450 ( 
.A(n_410),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_426),
.B(n_279),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_426),
.B(n_432),
.Y(n_452)
);

OAI22xp33_ASAP7_75t_SL g453 ( 
.A1(n_445),
.A2(n_420),
.B1(n_416),
.B2(n_431),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_439),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_438),
.B(n_409),
.Y(n_455)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_438),
.B(n_409),
.Y(n_456)
);

BUFx6f_ASAP7_75t_L g457 ( 
.A(n_450),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_441),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_452),
.B(n_424),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_451),
.B(n_424),
.Y(n_460)
);

AOI22xp33_ASAP7_75t_L g461 ( 
.A1(n_440),
.A2(n_425),
.B1(n_412),
.B2(n_416),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_L g462 ( 
.A(n_459),
.B(n_440),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_455),
.B(n_440),
.Y(n_463)
);

AOI22xp33_ASAP7_75t_SL g464 ( 
.A1(n_453),
.A2(n_445),
.B1(n_443),
.B2(n_444),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_454),
.Y(n_465)
);

INVx1_ASAP7_75t_SL g466 ( 
.A(n_458),
.Y(n_466)
);

AOI22xp33_ASAP7_75t_L g467 ( 
.A1(n_461),
.A2(n_448),
.B1(n_437),
.B2(n_446),
.Y(n_467)
);

AOI22xp33_ASAP7_75t_L g468 ( 
.A1(n_455),
.A2(n_446),
.B1(n_435),
.B2(n_413),
.Y(n_468)
);

AOI22xp33_ASAP7_75t_L g469 ( 
.A1(n_456),
.A2(n_446),
.B1(n_435),
.B2(n_447),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_L g470 ( 
.A(n_456),
.B(n_449),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_460),
.B(n_442),
.Y(n_471)
);

AOI22xp33_ASAP7_75t_L g472 ( 
.A1(n_464),
.A2(n_468),
.B1(n_463),
.B2(n_470),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_465),
.Y(n_473)
);

AOI22xp33_ASAP7_75t_L g474 ( 
.A1(n_471),
.A2(n_462),
.B1(n_467),
.B2(n_469),
.Y(n_474)
);

AND2x2_ASAP7_75t_L g475 ( 
.A(n_466),
.B(n_436),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_472),
.A2(n_418),
.B1(n_427),
.B2(n_423),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_474),
.A2(n_429),
.B1(n_419),
.B2(n_428),
.Y(n_477)
);

HB1xp67_ASAP7_75t_L g478 ( 
.A(n_475),
.Y(n_478)
);

NAND2xp5_ASAP7_75t_L g479 ( 
.A(n_473),
.B(n_457),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_478),
.B(n_55),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_479),
.B(n_71),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_L g482 ( 
.A(n_476),
.B(n_94),
.Y(n_482)
);

AND2x2_ASAP7_75t_L g483 ( 
.A(n_477),
.B(n_99),
.Y(n_483)
);

AND2x2_ASAP7_75t_L g484 ( 
.A(n_480),
.B(n_114),
.Y(n_484)
);

INVx1_ASAP7_75t_SL g485 ( 
.A(n_484),
.Y(n_485)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_485),
.Y(n_486)
);

BUFx2_ASAP7_75t_SL g487 ( 
.A(n_486),
.Y(n_487)
);

CKINVDCx16_ASAP7_75t_R g488 ( 
.A(n_487),
.Y(n_488)
);

INVx1_ASAP7_75t_SL g489 ( 
.A(n_488),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_489),
.Y(n_490)
);

INVx1_ASAP7_75t_L g491 ( 
.A(n_490),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_491),
.Y(n_492)
);

AO22x2_ASAP7_75t_L g493 ( 
.A1(n_492),
.A2(n_483),
.B1(n_481),
.B2(n_482),
.Y(n_493)
);

INVx2_ASAP7_75t_L g494 ( 
.A(n_493),
.Y(n_494)
);

BUFx2_ASAP7_75t_L g495 ( 
.A(n_493),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_495),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_494),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_495),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_496),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_498),
.Y(n_500)
);

INVx1_ASAP7_75t_L g501 ( 
.A(n_497),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g502 ( 
.A1(n_499),
.A2(n_131),
.B1(n_133),
.B2(n_134),
.Y(n_502)
);

OA22x2_ASAP7_75t_L g503 ( 
.A1(n_500),
.A2(n_137),
.B1(n_138),
.B2(n_139),
.Y(n_503)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_503),
.Y(n_504)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_502),
.Y(n_505)
);

OAI22xp33_ASAP7_75t_L g506 ( 
.A1(n_504),
.A2(n_501),
.B1(n_142),
.B2(n_143),
.Y(n_506)
);

OAI22xp33_ASAP7_75t_L g507 ( 
.A1(n_505),
.A2(n_140),
.B1(n_144),
.B2(n_145),
.Y(n_507)
);

INVx3_ASAP7_75t_L g508 ( 
.A(n_506),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_507),
.Y(n_509)
);

AOI221xp5_ASAP7_75t_L g510 ( 
.A1(n_509),
.A2(n_508),
.B1(n_149),
.B2(n_151),
.C(n_152),
.Y(n_510)
);

AOI211xp5_ASAP7_75t_L g511 ( 
.A1(n_510),
.A2(n_508),
.B(n_154),
.C(n_155),
.Y(n_511)
);


endmodule