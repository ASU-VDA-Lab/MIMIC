module fake_jpeg_6540_n_59 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_59);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_59;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_51;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx4f_ASAP7_75t_L g8 ( 
.A(n_1),
.Y(n_8)
);

BUFx12f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

OR2x2_ASAP7_75t_L g10 ( 
.A(n_1),
.B(n_3),
.Y(n_10)
);

BUFx3_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_3),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

INVx6_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

INVx8_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

INVx6_ASAP7_75t_SL g17 ( 
.A(n_9),
.Y(n_17)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_17),
.B(n_18),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

AND2x2_ASAP7_75t_L g21 ( 
.A(n_19),
.B(n_8),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_14),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g22 ( 
.A(n_20),
.B(n_10),
.Y(n_22)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_11),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_20),
.A2(n_15),
.B1(n_13),
.B2(n_12),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_23),
.A2(n_10),
.B1(n_16),
.B2(n_17),
.Y(n_29)
);

INVxp67_ASAP7_75t_L g27 ( 
.A(n_24),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g32 ( 
.A(n_27),
.B(n_29),
.Y(n_32)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_25),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_30),
.Y(n_33)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g37 ( 
.A1(n_31),
.A2(n_22),
.B(n_21),
.Y(n_37)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_31),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_34),
.B(n_35),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_29),
.B(n_23),
.Y(n_35)
);

OR2x2_ASAP7_75t_SL g36 ( 
.A(n_26),
.B(n_22),
.Y(n_36)
);

OAI21xp5_ASAP7_75t_SL g44 ( 
.A1(n_36),
.A2(n_38),
.B(n_18),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_28),
.B1(n_11),
.B2(n_18),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_L g38 ( 
.A1(n_26),
.A2(n_21),
.B(n_19),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_43),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_30),
.Y(n_40)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_40),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_44),
.C(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_45),
.B(n_40),
.C(n_2),
.Y(n_49)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_48),
.B(n_4),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_49),
.B(n_50),
.Y(n_52)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g53 ( 
.A(n_51),
.B(n_47),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_0),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_54),
.Y(n_56)
);

BUFx24_ASAP7_75t_SL g55 ( 
.A(n_52),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_56),
.B(n_55),
.C(n_2),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_57),
.B(n_0),
.Y(n_58)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_58),
.B(n_4),
.Y(n_59)
);


endmodule