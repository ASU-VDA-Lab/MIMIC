module fake_jpeg_26662_n_340 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g16 ( 
.A(n_5),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

INVx4_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_10),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_2),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_15),
.B(n_3),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_22),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_36),
.B(n_40),
.Y(n_50)
);

INVx6_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

INVx2_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_8),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_41),
.Y(n_66)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_30),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_42),
.Y(n_60)
);

INVx6_ASAP7_75t_L g43 ( 
.A(n_30),
.Y(n_43)
);

INVx3_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_32),
.Y(n_62)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_45),
.Y(n_56)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_46),
.Y(n_57)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_30),
.Y(n_47)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_40),
.B(n_34),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_51),
.B(n_59),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_24),
.B1(n_28),
.B2(n_18),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_52),
.A2(n_43),
.B1(n_18),
.B2(n_33),
.Y(n_87)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_64),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_63),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_38),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_39),
.B(n_32),
.Y(n_65)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

INVx11_ASAP7_75t_L g67 ( 
.A(n_42),
.Y(n_67)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_67),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_68),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_47),
.Y(n_69)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_69),
.Y(n_84)
);

CKINVDCx12_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_70),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_49),
.A2(n_37),
.B1(n_45),
.B2(n_39),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_71),
.A2(n_85),
.B1(n_87),
.B2(n_88),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_58),
.B(n_28),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_75),
.B(n_78),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_62),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_76),
.B(n_79),
.Y(n_101)
);

AND2x2_ASAP7_75t_SL g77 ( 
.A(n_64),
.B(n_38),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_77),
.B(n_83),
.C(n_66),
.Y(n_118)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_65),
.Y(n_79)
);

AND2x4_ASAP7_75t_L g81 ( 
.A(n_55),
.B(n_46),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g114 ( 
.A(n_81),
.B(n_57),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_50),
.B(n_28),
.Y(n_82)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_82),
.Y(n_116)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_55),
.B(n_46),
.C(n_38),
.Y(n_83)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_49),
.A2(n_37),
.B1(n_43),
.B2(n_45),
.Y(n_85)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_49),
.A2(n_43),
.B1(n_21),
.B2(n_20),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g89 ( 
.A(n_68),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_60),
.A2(n_19),
.B1(n_33),
.B2(n_29),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_92),
.A2(n_29),
.B1(n_33),
.B2(n_19),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_50),
.B(n_16),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_93),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_68),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_94),
.B(n_89),
.Y(n_121)
);

INVx2_ASAP7_75t_SL g95 ( 
.A(n_69),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_96),
.Y(n_113)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_79),
.A2(n_61),
.B1(n_48),
.B2(n_60),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_99),
.A2(n_103),
.B1(n_119),
.B2(n_85),
.Y(n_136)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_74),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_100),
.B(n_107),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_76),
.A2(n_61),
.B1(n_60),
.B2(n_63),
.Y(n_103)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_86),
.Y(n_105)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_77),
.A2(n_66),
.B(n_1),
.Y(n_106)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_106),
.A2(n_77),
.B(n_81),
.Y(n_129)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_74),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_108),
.Y(n_142)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx13_ASAP7_75t_L g130 ( 
.A(n_110),
.Y(n_130)
);

INVx3_ASAP7_75t_SL g111 ( 
.A(n_74),
.Y(n_111)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_111),
.A2(n_91),
.B1(n_95),
.B2(n_72),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_80),
.B(n_90),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_112),
.B(n_51),
.Y(n_154)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_114),
.B(n_118),
.Y(n_138)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_91),
.Y(n_117)
);

INVx13_ASAP7_75t_L g143 ( 
.A(n_117),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_121),
.Y(n_147)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_61),
.B1(n_53),
.B2(n_66),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_124),
.A2(n_125),
.B1(n_95),
.B2(n_91),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_81),
.A2(n_53),
.B1(n_67),
.B2(n_54),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_122),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_127),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_118),
.B(n_83),
.C(n_81),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_138),
.C(n_129),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g162 ( 
.A1(n_129),
.A2(n_131),
.B(n_139),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_114),
.A2(n_77),
.B(n_98),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_121),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g168 ( 
.A(n_132),
.B(n_134),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g188 ( 
.A(n_133),
.Y(n_188)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_101),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_112),
.B(n_97),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_135),
.B(n_146),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_136),
.A2(n_78),
.B1(n_72),
.B2(n_56),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_106),
.B(n_80),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_137),
.B(n_151),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g139 ( 
.A1(n_114),
.A2(n_96),
.B(n_94),
.Y(n_139)
);

INVx13_ASAP7_75t_L g141 ( 
.A(n_104),
.Y(n_141)
);

INVxp67_ASAP7_75t_SL g169 ( 
.A(n_141),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_115),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_144),
.Y(n_166)
);

AND2x2_ASAP7_75t_L g145 ( 
.A(n_109),
.B(n_71),
.Y(n_145)
);

OAI21xp33_ASAP7_75t_SL g186 ( 
.A1(n_145),
.A2(n_35),
.B(n_25),
.Y(n_186)
);

NAND3xp33_ASAP7_75t_L g146 ( 
.A(n_116),
.B(n_70),
.C(n_97),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_148),
.A2(n_19),
.B1(n_29),
.B2(n_27),
.Y(n_182)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_113),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g175 ( 
.A(n_149),
.B(n_153),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_113),
.A2(n_90),
.B1(n_73),
.B2(n_67),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_150),
.A2(n_117),
.B1(n_102),
.B2(n_104),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_56),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_56),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_155),
.Y(n_176)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_102),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g179 ( 
.A(n_154),
.B(n_17),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_123),
.B(n_105),
.Y(n_155)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_155),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_157),
.B(n_172),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_158),
.A2(n_161),
.B1(n_163),
.B2(n_167),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_136),
.A2(n_110),
.B1(n_108),
.B2(n_111),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_147),
.A2(n_111),
.B1(n_107),
.B2(n_100),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_164),
.B(n_165),
.C(n_173),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g165 ( 
.A(n_138),
.B(n_120),
.C(n_69),
.Y(n_165)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_132),
.A2(n_23),
.A3(n_17),
.B1(n_20),
.B2(n_21),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_SL g191 ( 
.A1(n_171),
.A2(n_186),
.B(n_148),
.Y(n_191)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_151),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g173 ( 
.A(n_138),
.B(n_21),
.C(n_31),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_152),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_174),
.B(n_180),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_128),
.B(n_21),
.C(n_31),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_177),
.B(n_179),
.C(n_185),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_137),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_178),
.B(n_139),
.Y(n_193)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_127),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_181),
.B(n_149),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_182),
.A2(n_184),
.B1(n_130),
.B2(n_142),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_154),
.B(n_17),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g198 ( 
.A1(n_183),
.A2(n_16),
.B(n_35),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_145),
.A2(n_27),
.B1(n_26),
.B2(n_25),
.Y(n_184)
);

XNOR2xp5_ASAP7_75t_L g185 ( 
.A(n_131),
.B(n_26),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_144),
.B(n_23),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_140),
.Y(n_189)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_189),
.Y(n_200)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_190),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_191),
.B(n_209),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_150),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g237 ( 
.A(n_192),
.B(n_130),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_193),
.B(n_196),
.Y(n_222)
);

OA22x2_ASAP7_75t_L g195 ( 
.A1(n_161),
.A2(n_145),
.B1(n_143),
.B2(n_153),
.Y(n_195)
);

INVx1_ASAP7_75t_SL g232 ( 
.A(n_195),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_176),
.B(n_140),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_198),
.B(n_8),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_176),
.B(n_159),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_201),
.B(n_202),
.Y(n_221)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_175),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_160),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_203),
.B(n_204),
.Y(n_235)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_205),
.B(n_208),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_166),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_206),
.A2(n_207),
.B(n_211),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g207 ( 
.A1(n_162),
.A2(n_143),
.B(n_1),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_159),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g209 ( 
.A(n_184),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g211 ( 
.A(n_189),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_178),
.B(n_141),
.Y(n_212)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_212),
.Y(n_231)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_213),
.B(n_214),
.Y(n_233)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_182),
.Y(n_214)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_162),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_217),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_188),
.A2(n_142),
.B(n_1),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g228 ( 
.A1(n_219),
.A2(n_0),
.B(n_2),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g220 ( 
.A(n_194),
.B(n_164),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_220),
.B(n_238),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g224 ( 
.A1(n_205),
.A2(n_188),
.B(n_185),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_224),
.B(n_240),
.Y(n_254)
);

OAI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_209),
.A2(n_183),
.B1(n_173),
.B2(n_177),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_225),
.A2(n_244),
.B1(n_217),
.B2(n_204),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_194),
.B(n_165),
.C(n_179),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_226),
.B(n_234),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_214),
.A2(n_170),
.B1(n_130),
.B2(n_141),
.Y(n_227)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_227),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_228),
.A2(n_192),
.B(n_191),
.Y(n_253)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_190),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_246),
.Y(n_258)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_210),
.B(n_23),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_203),
.Y(n_239)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_239),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_210),
.B(n_8),
.Y(n_241)
);

XOR2xp5_ASAP7_75t_L g259 ( 
.A(n_241),
.B(n_243),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_9),
.Y(n_243)
);

OAI22x1_ASAP7_75t_L g244 ( 
.A1(n_195),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_9),
.Y(n_245)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_241),
.Y(n_262)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_196),
.Y(n_246)
);

A2O1A1O1Ixp25_ASAP7_75t_L g247 ( 
.A1(n_224),
.A2(n_215),
.B(n_198),
.C(n_208),
.D(n_207),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_SL g276 ( 
.A(n_247),
.B(n_262),
.Y(n_276)
);

BUFx6f_ASAP7_75t_L g248 ( 
.A(n_244),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_248),
.B(n_266),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g249 ( 
.A(n_220),
.B(n_212),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_249),
.B(n_252),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_226),
.B(n_202),
.Y(n_252)
);

AO21x1_ASAP7_75t_L g269 ( 
.A1(n_253),
.A2(n_263),
.B(n_230),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g255 ( 
.A(n_239),
.B(n_206),
.Y(n_255)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_255),
.Y(n_272)
);

NAND3xp33_ASAP7_75t_L g260 ( 
.A(n_221),
.B(n_218),
.C(n_197),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g270 ( 
.A(n_260),
.B(n_261),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_235),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g263 ( 
.A(n_229),
.B(n_195),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_236),
.Y(n_264)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_264),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_265),
.A2(n_199),
.B1(n_231),
.B2(n_195),
.Y(n_280)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g267 ( 
.A(n_242),
.Y(n_267)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_267),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_245),
.B(n_213),
.Y(n_268)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_268),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_269),
.B(n_277),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_250),
.B(n_238),
.C(n_230),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_271),
.B(n_252),
.C(n_257),
.Y(n_286)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_250),
.B(n_222),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g278 ( 
.A1(n_251),
.A2(n_199),
.B1(n_233),
.B2(n_232),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g292 ( 
.A1(n_278),
.A2(n_282),
.B1(n_265),
.B2(n_248),
.Y(n_292)
);

FAx1_ASAP7_75t_L g279 ( 
.A(n_247),
.B(n_232),
.CI(n_219),
.CON(n_279),
.SN(n_279)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_279),
.A2(n_281),
.B(n_276),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_280),
.A2(n_281),
.B1(n_285),
.B2(n_254),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_263),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_267),
.A2(n_216),
.B1(n_228),
.B2(n_224),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g283 ( 
.A(n_258),
.Y(n_283)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_283),
.Y(n_291)
);

XOR2xp5_ASAP7_75t_L g308 ( 
.A(n_286),
.B(n_295),
.Y(n_308)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_272),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_293),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_288),
.A2(n_273),
.B1(n_11),
.B2(n_12),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_289),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_292),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_284),
.B(n_249),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_269),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_296),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_259),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_275),
.Y(n_296)
);

FAx1_ASAP7_75t_SL g297 ( 
.A(n_276),
.B(n_243),
.CI(n_240),
.CON(n_297),
.SN(n_297)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_298),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_279),
.A2(n_211),
.B(n_200),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_299),
.B(n_279),
.Y(n_301)
);

AOI221xp5_ASAP7_75t_L g300 ( 
.A1(n_274),
.A2(n_259),
.B1(n_262),
.B2(n_200),
.C(n_6),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_300),
.B(n_277),
.Y(n_304)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_301),
.Y(n_319)
);

INVx6_ASAP7_75t_L g302 ( 
.A(n_287),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_302),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_304),
.B(n_305),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g306 ( 
.A(n_290),
.B(n_273),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_306),
.B(n_312),
.Y(n_314)
);

OAI22xp5_ASAP7_75t_SL g320 ( 
.A1(n_307),
.A2(n_299),
.B1(n_291),
.B2(n_302),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_290),
.C(n_295),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_291),
.C(n_297),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_288),
.B(n_11),
.Y(n_312)
);

NOR2xp67_ASAP7_75t_SL g317 ( 
.A(n_310),
.B(n_294),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g329 ( 
.A(n_317),
.B(n_308),
.Y(n_329)
);

NAND3xp33_ASAP7_75t_L g318 ( 
.A(n_309),
.B(n_298),
.C(n_297),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g330 ( 
.A(n_318),
.B(n_320),
.Y(n_330)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_308),
.C(n_306),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_313),
.B(n_6),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_322),
.B(n_3),
.Y(n_327)
);

FAx1_ASAP7_75t_SL g323 ( 
.A(n_311),
.B(n_6),
.CI(n_9),
.CON(n_323),
.SN(n_323)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_323),
.B(n_15),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_L g333 ( 
.A1(n_324),
.A2(n_327),
.B1(n_319),
.B2(n_330),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_315),
.B(n_303),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g332 ( 
.A(n_325),
.B(n_323),
.Y(n_332)
);

INVxp33_ASAP7_75t_SL g326 ( 
.A(n_314),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_326),
.A2(n_328),
.B(n_329),
.Y(n_331)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_332),
.A2(n_333),
.B(n_316),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_334),
.B(n_331),
.Y(n_335)
);

OAI21xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_321),
.B(n_318),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g337 ( 
.A1(n_336),
.A2(n_12),
.B(n_13),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_13),
.Y(n_338)
);

OA21x2_ASAP7_75t_SL g339 ( 
.A1(n_338),
.A2(n_15),
.B(n_4),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_4),
.C(n_255),
.Y(n_340)
);


endmodule