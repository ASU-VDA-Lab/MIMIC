module fake_jpeg_12343_n_181 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_181);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_181;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_118;
wire n_100;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_3),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_8),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_2),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_5),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_11),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_5),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_5),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_16),
.B(n_24),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_33),
.B(n_39),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_25),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_34),
.Y(n_59)
);

INVx5_ASAP7_75t_L g35 ( 
.A(n_25),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_35),
.Y(n_65)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_37),
.Y(n_54)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_25),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_38),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g39 ( 
.A(n_16),
.B(n_13),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

CKINVDCx14_ASAP7_75t_R g67 ( 
.A(n_40),
.Y(n_67)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_28),
.Y(n_41)
);

INVx8_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_24),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_14),
.Y(n_43)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_43),
.Y(n_74)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_44),
.Y(n_76)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_24),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx6_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_47),
.B(n_31),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_20),
.B(n_0),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_52),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_19),
.B(n_0),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g71 ( 
.A(n_49),
.B(n_50),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_21),
.B(n_1),
.Y(n_50)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_22),
.Y(n_51)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_51),
.Y(n_78)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVxp67_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_55),
.B(n_57),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_26),
.B1(n_27),
.B2(n_30),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_56),
.A2(n_38),
.B1(n_36),
.B2(n_34),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_33),
.B(n_17),
.Y(n_57)
);

AO22x1_ASAP7_75t_SL g60 ( 
.A1(n_52),
.A2(n_26),
.B1(n_14),
.B2(n_30),
.Y(n_60)
);

AO22x1_ASAP7_75t_SL g80 ( 
.A1(n_60),
.A2(n_41),
.B1(n_40),
.B2(n_37),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_49),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_47),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_50),
.B(n_15),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_63),
.B(n_73),
.Y(n_100)
);

OAI22xp33_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_32),
.B1(n_29),
.B2(n_27),
.Y(n_72)
);

OAI22xp33_ASAP7_75t_L g98 ( 
.A1(n_72),
.A2(n_77),
.B1(n_38),
.B2(n_45),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_47),
.B(n_23),
.Y(n_73)
);

OAI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_46),
.A2(n_32),
.B1(n_29),
.B2(n_18),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_75),
.A2(n_47),
.B1(n_67),
.B2(n_54),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_48),
.A2(n_18),
.B1(n_21),
.B2(n_31),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_80),
.B(n_87),
.Y(n_111)
);

BUFx3_ASAP7_75t_L g81 ( 
.A(n_79),
.Y(n_81)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_81),
.Y(n_116)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_82),
.Y(n_106)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_84),
.Y(n_113)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_85),
.Y(n_105)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_86),
.Y(n_112)
);

NAND2xp33_ASAP7_75t_SL g87 ( 
.A(n_74),
.B(n_34),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_88),
.A2(n_91),
.B1(n_38),
.B2(n_65),
.Y(n_118)
);

OR2x2_ASAP7_75t_SL g89 ( 
.A(n_71),
.B(n_44),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_SL g121 ( 
.A(n_89),
.B(n_95),
.C(n_62),
.Y(n_121)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_64),
.Y(n_90)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_90),
.Y(n_114)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_64),
.Y(n_92)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_92),
.Y(n_115)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_72),
.Y(n_93)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_94),
.B(n_102),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g95 ( 
.A1(n_58),
.A2(n_35),
.B(n_42),
.Y(n_95)
);

A2O1A1Ixp33_ASAP7_75t_L g97 ( 
.A1(n_58),
.A2(n_23),
.B(n_15),
.C(n_43),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_97),
.B(n_62),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_74),
.B1(n_54),
.B2(n_60),
.Y(n_107)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_59),
.Y(n_99)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_99),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_59),
.Y(n_101)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_101),
.Y(n_122)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_66),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_77),
.B(n_13),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_70),
.Y(n_109)
);

INVxp33_ASAP7_75t_L g104 ( 
.A(n_88),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_104),
.B(n_80),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_107),
.A2(n_65),
.B1(n_83),
.B2(n_68),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g125 ( 
.A(n_109),
.B(n_110),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_96),
.B(n_60),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_117),
.B(n_69),
.Y(n_133)
);

AOI22x1_ASAP7_75t_L g127 ( 
.A1(n_118),
.A2(n_80),
.B1(n_87),
.B2(n_98),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_121),
.A2(n_83),
.B(n_65),
.Y(n_129)
);

XOR2x1_ASAP7_75t_L g123 ( 
.A(n_117),
.B(n_89),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g140 ( 
.A(n_123),
.B(n_126),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_108),
.B(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_124),
.B(n_128),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_95),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g146 ( 
.A1(n_127),
.A2(n_130),
.B1(n_137),
.B2(n_119),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_129),
.B(n_132),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_131),
.B(n_133),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_92),
.Y(n_132)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_105),
.Y(n_134)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_134),
.Y(n_139)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_112),
.Y(n_135)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g136 ( 
.A(n_106),
.B(n_12),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_136),
.B(n_12),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_111),
.A2(n_66),
.B1(n_101),
.B2(n_99),
.Y(n_137)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_118),
.B(n_69),
.Y(n_138)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_138),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_L g145 ( 
.A1(n_125),
.A2(n_119),
.B1(n_120),
.B2(n_122),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_145),
.A2(n_115),
.B1(n_114),
.B2(n_113),
.Y(n_158)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_146),
.B(n_138),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_137),
.Y(n_147)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_147),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_148),
.B(n_149),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_112),
.Y(n_149)
);

INVx2_ASAP7_75t_L g151 ( 
.A(n_139),
.Y(n_151)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_151),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g152 ( 
.A(n_142),
.B(n_129),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_152),
.B(n_157),
.Y(n_161)
);

NAND3xp33_ASAP7_75t_SL g153 ( 
.A(n_141),
.B(n_123),
.C(n_127),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_SL g164 ( 
.A(n_153),
.B(n_154),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_144),
.Y(n_154)
);

A2O1A1O1Ixp25_ASAP7_75t_L g156 ( 
.A1(n_140),
.A2(n_126),
.B(n_127),
.C(n_138),
.D(n_130),
.Y(n_156)
);

MAJx2_ASAP7_75t_L g166 ( 
.A(n_156),
.B(n_143),
.C(n_116),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g162 ( 
.A(n_158),
.B(n_150),
.C(n_115),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_165),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_154),
.B(n_140),
.C(n_141),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_163),
.B(n_159),
.C(n_158),
.Y(n_169)
);

AOI321xp33_ASAP7_75t_L g165 ( 
.A1(n_155),
.A2(n_149),
.A3(n_143),
.B1(n_147),
.B2(n_146),
.C(n_114),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_166),
.B(n_156),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_163),
.B(n_157),
.Y(n_168)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_168),
.B(n_169),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_170),
.B(n_79),
.C(n_68),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_164),
.A2(n_122),
.B1(n_120),
.B2(n_116),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_81),
.B1(n_2),
.B2(n_4),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_167),
.A2(n_161),
.B1(n_166),
.B2(n_160),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_172),
.B(n_174),
.C(n_175),
.Y(n_177)
);

AOI31xp67_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_169),
.A3(n_168),
.B(n_9),
.Y(n_176)
);

OAI21x1_ASAP7_75t_L g178 ( 
.A1(n_176),
.A2(n_9),
.B(n_177),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_178),
.A2(n_174),
.B(n_2),
.Y(n_179)
);

AOI321xp33_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_1),
.A3(n_4),
.B1(n_6),
.B2(n_7),
.C(n_173),
.Y(n_180)
);

XOR2xp5_ASAP7_75t_L g181 ( 
.A(n_180),
.B(n_7),
.Y(n_181)
);


endmodule