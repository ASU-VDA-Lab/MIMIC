module fake_jpeg_1836_n_578 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_578);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_578;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_14),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_5),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_2),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_18),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_7),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_3),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_17),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVxp33_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_4),
.Y(n_40)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_13),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_11),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_10),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_11),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_7),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_12),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_13),
.Y(n_51)
);

BUFx8_ASAP7_75t_L g52 ( 
.A(n_18),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_13),
.Y(n_53)
);

CKINVDCx16_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_5),
.Y(n_55)
);

BUFx12_ASAP7_75t_L g56 ( 
.A(n_52),
.Y(n_56)
);

INVx6_ASAP7_75t_SL g114 ( 
.A(n_56),
.Y(n_114)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_57),
.Y(n_135)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_59),
.Y(n_117)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_60),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_19),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_61),
.Y(n_137)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_52),
.Y(n_62)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_62),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_19),
.Y(n_63)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_63),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_27),
.B(n_18),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_64),
.B(n_85),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

INVx6_ASAP7_75t_L g169 ( 
.A(n_65),
.Y(n_169)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_66),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_30),
.Y(n_67)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_67),
.Y(n_116)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_34),
.Y(n_68)
);

INVx3_ASAP7_75t_L g139 ( 
.A(n_68),
.Y(n_139)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_26),
.Y(n_69)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_69),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_30),
.Y(n_70)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_70),
.Y(n_152)
);

HB1xp67_ASAP7_75t_L g71 ( 
.A(n_34),
.Y(n_71)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_71),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_72),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_SL g73 ( 
.A(n_20),
.B(n_8),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_73),
.B(n_78),
.Y(n_111)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_74),
.Y(n_132)
);

INVx11_ASAP7_75t_L g75 ( 
.A(n_52),
.Y(n_75)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_75),
.Y(n_121)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_27),
.Y(n_76)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_76),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g77 ( 
.A(n_52),
.Y(n_77)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_77),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g78 ( 
.A(n_27),
.B(n_8),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_30),
.Y(n_79)
);

INVx5_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

INVx11_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_33),
.Y(n_81)
);

INVx5_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx11_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

INVx4_ASAP7_75t_L g166 ( 
.A(n_82),
.Y(n_166)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_31),
.Y(n_83)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_83),
.Y(n_155)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_33),
.Y(n_84)
);

INVx5_ASAP7_75t_L g154 ( 
.A(n_84),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_20),
.B(n_7),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

BUFx3_ASAP7_75t_L g119 ( 
.A(n_86),
.Y(n_119)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_25),
.Y(n_87)
);

INVx3_ASAP7_75t_L g164 ( 
.A(n_87),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_88),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx4_ASAP7_75t_L g167 ( 
.A(n_89),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_90),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_21),
.B(n_9),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_97),
.Y(n_122)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_92),
.Y(n_158)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_35),
.Y(n_93)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_93),
.Y(n_162)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_25),
.Y(n_94)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_94),
.Y(n_165)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_31),
.Y(n_95)
);

AOI21xp33_ASAP7_75t_L g112 ( 
.A1(n_95),
.A2(n_105),
.B(n_35),
.Y(n_112)
);

BUFx4f_ASAP7_75t_SL g96 ( 
.A(n_43),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_108),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_31),
.B(n_50),
.Y(n_97)
);

INVx6_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_98),
.Y(n_172)
);

BUFx4f_ASAP7_75t_L g99 ( 
.A(n_50),
.Y(n_99)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_25),
.Y(n_100)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_50),
.Y(n_101)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_101),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_21),
.B(n_9),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_102),
.B(n_54),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_103),
.Y(n_148)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_44),
.Y(n_104)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_104),
.Y(n_160)
);

BUFx12_ASAP7_75t_L g105 ( 
.A(n_38),
.Y(n_105)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_23),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_106),
.B(n_107),
.Y(n_163)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_23),
.Y(n_107)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_23),
.Y(n_108)
);

AOI21xp33_ASAP7_75t_L g203 ( 
.A1(n_112),
.A2(n_146),
.B(n_45),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_78),
.B(n_39),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_123),
.B(n_127),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_81),
.A2(n_23),
.B1(n_46),
.B2(n_44),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_124),
.A2(n_151),
.B1(n_161),
.B2(n_171),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_68),
.A2(n_46),
.B1(n_54),
.B2(n_25),
.Y(n_126)
);

OA22x2_ASAP7_75t_L g193 ( 
.A1(n_126),
.A2(n_133),
.B1(n_147),
.B2(n_153),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_69),
.B(n_42),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_42),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_128),
.B(n_142),
.Y(n_195)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_62),
.A2(n_28),
.B1(n_36),
.B2(n_29),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_96),
.B(n_22),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_106),
.B(n_46),
.C(n_40),
.Y(n_144)
);

OAI32xp33_ASAP7_75t_L g191 ( 
.A1(n_144),
.A2(n_149),
.A3(n_56),
.B1(n_38),
.B2(n_45),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_100),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_145),
.B(n_156),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_75),
.A2(n_28),
.B1(n_36),
.B2(n_29),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_107),
.B(n_46),
.C(n_40),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g151 ( 
.A1(n_84),
.A2(n_22),
.B1(n_51),
.B2(n_48),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_74),
.A2(n_28),
.B1(n_29),
.B2(n_36),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_96),
.B(n_47),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_98),
.A2(n_32),
.B1(n_51),
.B2(n_47),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_24),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g210 ( 
.A(n_168),
.B(n_55),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_80),
.A2(n_55),
.B1(n_53),
.B2(n_49),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_SL g173 ( 
.A1(n_144),
.A2(n_53),
.B1(n_37),
.B2(n_49),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_173),
.Y(n_240)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_117),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g234 ( 
.A(n_174),
.Y(n_234)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_149),
.A2(n_37),
.B1(n_53),
.B2(n_49),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g266 ( 
.A(n_175),
.Y(n_266)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_114),
.Y(n_176)
);

BUFx3_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

INVx2_ASAP7_75t_L g177 ( 
.A(n_172),
.Y(n_177)
);

INVx2_ASAP7_75t_L g236 ( 
.A(n_177),
.Y(n_236)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_129),
.Y(n_179)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_179),
.Y(n_242)
);

INVx3_ASAP7_75t_L g180 ( 
.A(n_114),
.Y(n_180)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_180),
.Y(n_239)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

INVx2_ASAP7_75t_L g244 ( 
.A(n_181),
.Y(n_244)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_163),
.Y(n_182)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_182),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g183 ( 
.A(n_139),
.Y(n_183)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_183),
.Y(n_273)
);

INVx4_ASAP7_75t_L g184 ( 
.A(n_132),
.Y(n_184)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_184),
.Y(n_260)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_157),
.A2(n_45),
.B1(n_37),
.B2(n_82),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_185),
.A2(n_207),
.B1(n_216),
.B2(n_219),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g186 ( 
.A(n_132),
.Y(n_186)
);

INVx5_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_118),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_187),
.B(n_190),
.Y(n_267)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_117),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_188),
.Y(n_238)
);

INVx11_ASAP7_75t_L g189 ( 
.A(n_115),
.Y(n_189)
);

INVx8_ASAP7_75t_L g241 ( 
.A(n_189),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_113),
.Y(n_190)
);

AND2x2_ASAP7_75t_L g251 ( 
.A(n_191),
.B(n_198),
.Y(n_251)
);

INVx5_ASAP7_75t_L g192 ( 
.A(n_116),
.Y(n_192)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_192),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_122),
.A2(n_79),
.B1(n_61),
.B2(n_103),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g231 ( 
.A1(n_194),
.A2(n_206),
.B1(n_221),
.B2(n_147),
.Y(n_231)
);

CKINVDCx16_ASAP7_75t_R g196 ( 
.A(n_126),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_196),
.B(n_199),
.Y(n_246)
);

INVx4_ASAP7_75t_L g197 ( 
.A(n_115),
.Y(n_197)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_197),
.Y(n_278)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_116),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g199 ( 
.A(n_121),
.Y(n_199)
);

BUFx2_ASAP7_75t_L g200 ( 
.A(n_121),
.Y(n_200)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_200),
.Y(n_255)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_138),
.Y(n_201)
);

AND2x2_ASAP7_75t_L g253 ( 
.A(n_201),
.B(n_203),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_113),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_202),
.B(n_210),
.Y(n_262)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_131),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_204),
.B(n_209),
.Y(n_233)
);

INVx4_ASAP7_75t_L g205 ( 
.A(n_164),
.Y(n_205)
);

CKINVDCx14_ASAP7_75t_R g275 ( 
.A(n_205),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g206 ( 
.A1(n_109),
.A2(n_86),
.B1(n_59),
.B2(n_63),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_157),
.A2(n_48),
.B1(n_32),
.B2(n_24),
.Y(n_207)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_130),
.Y(n_209)
);

INVx6_ASAP7_75t_L g211 ( 
.A(n_137),
.Y(n_211)
);

INVx6_ASAP7_75t_L g257 ( 
.A(n_211),
.Y(n_257)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_148),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_212),
.B(n_222),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_140),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_213),
.B(n_214),
.Y(n_265)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_139),
.Y(n_214)
);

INVxp67_ASAP7_75t_L g215 ( 
.A(n_141),
.Y(n_215)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_215),
.Y(n_272)
);

INVx11_ASAP7_75t_L g216 ( 
.A(n_159),
.Y(n_216)
);

CKINVDCx20_ASAP7_75t_R g217 ( 
.A(n_134),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_218),
.Y(n_232)
);

INVx6_ASAP7_75t_L g218 ( 
.A(n_137),
.Y(n_218)
);

INVx3_ASAP7_75t_L g219 ( 
.A(n_164),
.Y(n_219)
);

INVx4_ASAP7_75t_SL g220 ( 
.A(n_141),
.Y(n_220)
);

NAND2x1_ASAP7_75t_SL g252 ( 
.A(n_220),
.B(n_176),
.Y(n_252)
);

AOI22xp33_ASAP7_75t_L g221 ( 
.A1(n_167),
.A2(n_55),
.B1(n_108),
.B2(n_88),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_111),
.B(n_104),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_135),
.A2(n_92),
.B1(n_94),
.B2(n_87),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_223),
.A2(n_225),
.B1(n_228),
.B2(n_229),
.Y(n_245)
);

INVx2_ASAP7_75t_L g225 ( 
.A(n_135),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_134),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_226),
.B(n_119),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_153),
.A2(n_67),
.B1(n_90),
.B2(n_89),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_227),
.A2(n_38),
.B1(n_35),
.B2(n_105),
.Y(n_276)
);

INVx5_ASAP7_75t_L g228 ( 
.A(n_152),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_158),
.A2(n_162),
.B1(n_165),
.B2(n_160),
.Y(n_229)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_110),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_SL g249 ( 
.A1(n_230),
.A2(n_166),
.B1(n_119),
.B2(n_167),
.Y(n_249)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_231),
.A2(n_256),
.B1(n_268),
.B2(n_269),
.Y(n_280)
);

AO22x2_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_133),
.B1(n_171),
.B2(n_159),
.Y(n_237)
);

AO22x1_ASAP7_75t_SL g315 ( 
.A1(n_237),
.A2(n_38),
.B1(n_1),
.B2(n_2),
.Y(n_315)
);

AND2x4_ASAP7_75t_SL g247 ( 
.A(n_182),
.B(n_136),
.Y(n_247)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_247),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g293 ( 
.A(n_249),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_195),
.B(n_155),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_250),
.B(n_254),
.Y(n_287)
);

INVx11_ASAP7_75t_L g319 ( 
.A(n_252),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_187),
.B(n_208),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_194),
.A2(n_150),
.B1(n_125),
.B2(n_65),
.Y(n_256)
);

AOI22xp33_ASAP7_75t_L g258 ( 
.A1(n_224),
.A2(n_170),
.B1(n_143),
.B2(n_154),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_SL g296 ( 
.A1(n_258),
.A2(n_261),
.B1(n_271),
.B2(n_220),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_170),
.B1(n_143),
.B2(n_154),
.Y(n_261)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_206),
.A2(n_191),
.B1(n_193),
.B2(n_178),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_193),
.A2(n_169),
.B1(n_120),
.B2(n_72),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g270 ( 
.A1(n_193),
.A2(n_120),
.B1(n_169),
.B2(n_70),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_270),
.A2(n_276),
.B1(n_277),
.B2(n_184),
.Y(n_294)
);

AOI22xp33_ASAP7_75t_L g271 ( 
.A1(n_204),
.A2(n_166),
.B1(n_56),
.B2(n_152),
.Y(n_271)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_193),
.A2(n_105),
.B1(n_38),
.B2(n_2),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_SL g279 ( 
.A1(n_240),
.A2(n_202),
.B1(n_190),
.B2(n_217),
.Y(n_279)
);

INVxp67_ASAP7_75t_L g332 ( 
.A(n_279),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_SL g281 ( 
.A(n_267),
.B(n_230),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g321 ( 
.A(n_281),
.B(n_284),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_248),
.Y(n_282)
);

BUFx3_ASAP7_75t_L g341 ( 
.A(n_282),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_267),
.B(n_179),
.Y(n_284)
);

INVx3_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g342 ( 
.A(n_285),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g286 ( 
.A(n_252),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_286),
.B(n_298),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_254),
.B(n_213),
.Y(n_288)
);

INVxp67_ASAP7_75t_L g356 ( 
.A(n_288),
.Y(n_356)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_242),
.Y(n_289)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_289),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g290 ( 
.A(n_253),
.B(n_209),
.C(n_180),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_290),
.B(n_313),
.C(n_320),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_SL g291 ( 
.A1(n_251),
.A2(n_229),
.B1(n_226),
.B2(n_219),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_291),
.A2(n_294),
.B1(n_304),
.B2(n_312),
.Y(n_337)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_242),
.Y(n_295)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_295),
.Y(n_325)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_296),
.A2(n_307),
.B1(n_317),
.B2(n_231),
.Y(n_331)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_232),
.Y(n_297)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_297),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_262),
.B(n_215),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_232),
.Y(n_299)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g300 ( 
.A1(n_240),
.A2(n_186),
.B1(n_198),
.B2(n_228),
.Y(n_300)
);

OAI21xp5_ASAP7_75t_L g330 ( 
.A1(n_300),
.A2(n_310),
.B(n_245),
.Y(n_330)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_233),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g334 ( 
.A(n_301),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_201),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_302),
.B(n_309),
.Y(n_326)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_233),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_303),
.B(n_311),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g304 ( 
.A1(n_251),
.A2(n_174),
.B1(n_218),
.B2(n_211),
.Y(n_304)
);

INVx6_ASAP7_75t_L g305 ( 
.A(n_234),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g340 ( 
.A(n_305),
.Y(n_340)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_278),
.Y(n_306)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_306),
.Y(n_344)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_238),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_268),
.A2(n_205),
.B1(n_181),
.B2(n_225),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_L g336 ( 
.A1(n_308),
.A2(n_275),
.B1(n_244),
.B2(n_255),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_252),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_266),
.A2(n_177),
.B(n_214),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_263),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g312 ( 
.A1(n_276),
.A2(n_188),
.B1(n_192),
.B2(n_220),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_253),
.B(n_197),
.C(n_200),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_236),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_314),
.B(n_316),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_315),
.B(n_318),
.Y(n_350)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_236),
.Y(n_316)
);

AOI22xp33_ASAP7_75t_SL g317 ( 
.A1(n_266),
.A2(n_246),
.B1(n_277),
.B2(n_269),
.Y(n_317)
);

INVx2_ASAP7_75t_SL g318 ( 
.A(n_257),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_259),
.B(n_216),
.Y(n_320)
);

XNOR2x1_ASAP7_75t_SL g324 ( 
.A(n_287),
.B(n_253),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_324),
.A2(n_346),
.B(n_357),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_280),
.A2(n_270),
.B1(n_259),
.B2(n_237),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g363 ( 
.A1(n_327),
.A2(n_336),
.B1(n_338),
.B2(n_353),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_SL g392 ( 
.A1(n_330),
.A2(n_331),
.B(n_339),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g338 ( 
.A1(n_280),
.A2(n_237),
.B1(n_250),
.B2(n_235),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_L g339 ( 
.A1(n_286),
.A2(n_243),
.B(n_237),
.Y(n_339)
);

AOI32xp33_ASAP7_75t_L g343 ( 
.A1(n_302),
.A2(n_247),
.A3(n_237),
.B1(n_243),
.B2(n_265),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g388 ( 
.A(n_343),
.B(n_264),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_287),
.B(n_247),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_345),
.B(n_347),
.C(n_348),
.Y(n_381)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_309),
.A2(n_292),
.B(n_297),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g347 ( 
.A(n_290),
.B(n_247),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g349 ( 
.A(n_301),
.B(n_239),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_SL g360 ( 
.A(n_349),
.B(n_355),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_L g351 ( 
.A1(n_294),
.A2(n_256),
.B1(n_257),
.B2(n_274),
.Y(n_351)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_351),
.A2(n_295),
.B1(n_289),
.B2(n_279),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_299),
.B(n_274),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_352),
.B(n_358),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_SL g353 ( 
.A1(n_308),
.A2(n_234),
.B1(n_238),
.B2(n_239),
.Y(n_353)
);

OAI21x1_ASAP7_75t_L g354 ( 
.A1(n_319),
.A2(n_273),
.B(n_278),
.Y(n_354)
);

OA21x2_ASAP7_75t_L g384 ( 
.A1(n_354),
.A2(n_315),
.B(n_260),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g355 ( 
.A(n_303),
.B(n_283),
.Y(n_355)
);

AOI22xp33_ASAP7_75t_SL g357 ( 
.A1(n_293),
.A2(n_264),
.B1(n_260),
.B2(n_273),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_283),
.B(n_244),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_SL g359 ( 
.A(n_284),
.B(n_313),
.Y(n_359)
);

MAJx2_ASAP7_75t_L g373 ( 
.A(n_359),
.B(n_320),
.C(n_281),
.Y(n_373)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_352),
.Y(n_361)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_361),
.Y(n_409)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_333),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_362),
.B(n_366),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_324),
.B(n_311),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_364),
.B(n_376),
.Y(n_412)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_365),
.A2(n_382),
.B1(n_383),
.B2(n_384),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_333),
.Y(n_366)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_322),
.Y(n_368)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_368),
.Y(n_411)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_322),
.Y(n_369)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_369),
.Y(n_414)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_325),
.Y(n_370)
);

INVx2_ASAP7_75t_L g422 ( 
.A(n_370),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_358),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_387),
.Y(n_425)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_325),
.Y(n_372)
);

INVxp67_ASAP7_75t_L g415 ( 
.A(n_372),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_SL g396 ( 
.A(n_373),
.B(n_345),
.Y(n_396)
);

INVx2_ASAP7_75t_L g374 ( 
.A(n_342),
.Y(n_374)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_374),
.Y(n_426)
);

OAI21xp5_ASAP7_75t_L g375 ( 
.A1(n_339),
.A2(n_323),
.B(n_326),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_375),
.A2(n_380),
.B(n_384),
.Y(n_398)
);

XOR2xp5_ASAP7_75t_L g376 ( 
.A(n_359),
.B(n_291),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g378 ( 
.A(n_323),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_378),
.B(n_386),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_348),
.B(n_304),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_379),
.B(n_381),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g380 ( 
.A1(n_326),
.A2(n_319),
.B(n_310),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_327),
.A2(n_312),
.B1(n_315),
.B2(n_293),
.Y(n_382)
);

AOI22xp5_ASAP7_75t_L g383 ( 
.A1(n_338),
.A2(n_315),
.B1(n_318),
.B2(n_285),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_347),
.B(n_316),
.C(n_314),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_385),
.B(n_391),
.Y(n_418)
);

CKINVDCx16_ASAP7_75t_R g386 ( 
.A(n_342),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g387 ( 
.A(n_329),
.B(n_318),
.Y(n_387)
);

AOI21xp5_ASAP7_75t_SL g402 ( 
.A1(n_388),
.A2(n_355),
.B(n_329),
.Y(n_402)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_328),
.Y(n_389)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_389),
.Y(n_427)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_328),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_390),
.B(n_393),
.Y(n_428)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_346),
.B(n_300),
.C(n_282),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_349),
.Y(n_393)
);

AOI21xp5_ASAP7_75t_L g394 ( 
.A1(n_354),
.A2(n_272),
.B(n_305),
.Y(n_394)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_394),
.A2(n_330),
.B(n_332),
.Y(n_399)
);

NAND3xp33_ASAP7_75t_L g395 ( 
.A(n_356),
.B(n_272),
.C(n_234),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_395),
.B(n_342),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g458 ( 
.A(n_396),
.B(n_421),
.Y(n_458)
);

OAI21xp5_ASAP7_75t_L g440 ( 
.A1(n_399),
.A2(n_402),
.B(n_367),
.Y(n_440)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_383),
.A2(n_350),
.B1(n_335),
.B2(n_337),
.Y(n_400)
);

OAI22xp5_ASAP7_75t_L g443 ( 
.A1(n_400),
.A2(n_413),
.B1(n_420),
.B2(n_365),
.Y(n_443)
);

AND2x2_ASAP7_75t_L g401 ( 
.A(n_394),
.B(n_350),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_401),
.Y(n_433)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_387),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_403),
.B(n_407),
.Y(n_438)
);

AOI22xp5_ASAP7_75t_L g446 ( 
.A1(n_405),
.A2(n_419),
.B1(n_430),
.B2(n_380),
.Y(n_446)
);

HB1xp67_ASAP7_75t_L g453 ( 
.A(n_406),
.Y(n_453)
);

CKINVDCx20_ASAP7_75t_R g407 ( 
.A(n_375),
.Y(n_407)
);

INVx3_ASAP7_75t_L g408 ( 
.A(n_374),
.Y(n_408)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_408),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_SL g410 ( 
.A(n_378),
.B(n_321),
.Y(n_410)
);

NOR2xp33_ASAP7_75t_SL g439 ( 
.A(n_410),
.B(n_393),
.Y(n_439)
);

AOI22xp5_ASAP7_75t_L g413 ( 
.A1(n_363),
.A2(n_335),
.B1(n_337),
.B2(n_351),
.Y(n_413)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_361),
.Y(n_416)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_416),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g419 ( 
.A1(n_363),
.A2(n_334),
.B1(n_343),
.B2(n_321),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_384),
.A2(n_334),
.B1(n_353),
.B2(n_336),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_381),
.B(n_334),
.Y(n_421)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_360),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_423),
.B(n_360),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g424 ( 
.A(n_376),
.B(n_344),
.Y(n_424)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_424),
.B(n_379),
.Y(n_434)
);

CKINVDCx14_ASAP7_75t_R g429 ( 
.A(n_377),
.Y(n_429)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_429),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_SL g430 ( 
.A1(n_382),
.A2(n_344),
.B1(n_340),
.B2(n_341),
.Y(n_430)
);

AOI22xp33_ASAP7_75t_L g466 ( 
.A1(n_432),
.A2(n_443),
.B1(n_445),
.B2(n_447),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_404),
.Y(n_464)
);

NAND2xp5_ASAP7_75t_L g435 ( 
.A(n_415),
.B(n_362),
.Y(n_435)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_435),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_415),
.B(n_366),
.Y(n_436)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_436),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g468 ( 
.A(n_439),
.B(n_442),
.Y(n_468)
);

AOI21xp5_ASAP7_75t_L g479 ( 
.A1(n_440),
.A2(n_408),
.B(n_241),
.Y(n_479)
);

CKINVDCx16_ASAP7_75t_R g442 ( 
.A(n_397),
.Y(n_442)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_417),
.Y(n_444)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_444),
.Y(n_482)
);

CKINVDCx20_ASAP7_75t_R g445 ( 
.A(n_417),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_446),
.A2(n_398),
.B1(n_414),
.B2(n_372),
.Y(n_470)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_425),
.Y(n_447)
);

AO21x2_ASAP7_75t_SL g448 ( 
.A1(n_401),
.A2(n_392),
.B(n_371),
.Y(n_448)
);

CKINVDCx20_ASAP7_75t_R g474 ( 
.A(n_448),
.Y(n_474)
);

OAI22xp5_ASAP7_75t_L g449 ( 
.A1(n_400),
.A2(n_367),
.B1(n_377),
.B2(n_391),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_449),
.A2(n_454),
.B1(n_459),
.B2(n_461),
.Y(n_471)
);

INVxp67_ASAP7_75t_SL g450 ( 
.A(n_428),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_450),
.B(n_452),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_L g451 ( 
.A(n_427),
.B(n_390),
.Y(n_451)
);

INVxp67_ASAP7_75t_L g476 ( 
.A(n_451),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_L g452 ( 
.A(n_421),
.B(n_341),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_L g454 ( 
.A1(n_413),
.A2(n_364),
.B1(n_389),
.B2(n_392),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_402),
.B(n_341),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g483 ( 
.A(n_455),
.B(n_457),
.Y(n_483)
);

BUFx12_ASAP7_75t_L g456 ( 
.A(n_426),
.Y(n_456)
);

CKINVDCx16_ASAP7_75t_R g477 ( 
.A(n_456),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_SL g457 ( 
.A(n_409),
.B(n_369),
.Y(n_457)
);

OAI22xp5_ASAP7_75t_L g459 ( 
.A1(n_420),
.A2(n_425),
.B1(n_428),
.B2(n_401),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_422),
.Y(n_460)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_460),
.A2(n_426),
.B1(n_427),
.B2(n_422),
.Y(n_463)
);

NOR2xp33_ASAP7_75t_SL g461 ( 
.A(n_411),
.B(n_368),
.Y(n_461)
);

FAx1_ASAP7_75t_SL g462 ( 
.A(n_448),
.B(n_419),
.CI(n_373),
.CON(n_462),
.SN(n_462)
);

FAx1_ASAP7_75t_SL g504 ( 
.A(n_462),
.B(n_457),
.CI(n_461),
.CON(n_504),
.SN(n_504)
);

INVx1_ASAP7_75t_L g490 ( 
.A(n_463),
.Y(n_490)
);

XNOR2xp5_ASAP7_75t_L g488 ( 
.A(n_464),
.B(n_458),
.Y(n_488)
);

AOI22xp5_ASAP7_75t_L g465 ( 
.A1(n_443),
.A2(n_430),
.B1(n_399),
.B2(n_418),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g505 ( 
.A1(n_465),
.A2(n_469),
.B1(n_431),
.B2(n_456),
.Y(n_505)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_459),
.A2(n_418),
.B1(n_424),
.B2(n_398),
.Y(n_469)
);

AOI22xp5_ASAP7_75t_L g487 ( 
.A1(n_470),
.A2(n_473),
.B1(n_485),
.B2(n_486),
.Y(n_487)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_446),
.A2(n_370),
.B1(n_412),
.B2(n_396),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_434),
.B(n_404),
.C(n_385),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g502 ( 
.A(n_475),
.B(n_478),
.C(n_437),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_458),
.B(n_412),
.C(n_340),
.Y(n_478)
);

OAI21xp33_ASAP7_75t_L g492 ( 
.A1(n_479),
.A2(n_481),
.B(n_448),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g481 ( 
.A1(n_448),
.A2(n_241),
.B(n_307),
.Y(n_481)
);

OAI22xp5_ASAP7_75t_L g484 ( 
.A1(n_445),
.A2(n_307),
.B1(n_238),
.B2(n_241),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_L g497 ( 
.A1(n_484),
.A2(n_437),
.B1(n_431),
.B2(n_460),
.Y(n_497)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_444),
.A2(n_38),
.B1(n_189),
.B2(n_10),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g486 ( 
.A1(n_447),
.A2(n_9),
.B1(n_15),
.B2(n_14),
.Y(n_486)
);

XNOR2xp5_ASAP7_75t_L g510 ( 
.A(n_488),
.B(n_491),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g489 ( 
.A1(n_471),
.A2(n_438),
.B1(n_449),
.B2(n_454),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_489),
.B(n_494),
.Y(n_522)
);

XNOR2xp5_ASAP7_75t_L g491 ( 
.A(n_464),
.B(n_440),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_SL g523 ( 
.A1(n_492),
.A2(n_504),
.B(n_462),
.Y(n_523)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_436),
.Y(n_493)
);

XNOR2xp5_ASAP7_75t_L g514 ( 
.A(n_493),
.B(n_495),
.Y(n_514)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_468),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_471),
.A2(n_441),
.B1(n_433),
.B2(n_435),
.Y(n_495)
);

XNOR2xp5_ASAP7_75t_SL g496 ( 
.A(n_473),
.B(n_453),
.Y(n_496)
);

XNOR2xp5_ASAP7_75t_L g519 ( 
.A(n_496),
.B(n_499),
.Y(n_519)
);

NOR2xp33_ASAP7_75t_L g509 ( 
.A(n_497),
.B(n_498),
.Y(n_509)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_472),
.Y(n_498)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_478),
.B(n_439),
.Y(n_499)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_466),
.A2(n_441),
.B1(n_467),
.B2(n_480),
.Y(n_500)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_500),
.B(n_501),
.Y(n_515)
);

INVx2_ASAP7_75t_SL g501 ( 
.A(n_482),
.Y(n_501)
);

OAI21xp5_ASAP7_75t_L g511 ( 
.A1(n_502),
.A2(n_465),
.B(n_477),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_475),
.B(n_433),
.C(n_451),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_503),
.B(n_476),
.C(n_477),
.Y(n_512)
);

NOR2xp33_ASAP7_75t_L g516 ( 
.A(n_505),
.B(n_506),
.Y(n_516)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_483),
.Y(n_506)
);

OAI321xp33_ASAP7_75t_L g507 ( 
.A1(n_490),
.A2(n_480),
.A3(n_467),
.B1(n_482),
.B2(n_481),
.C(n_479),
.Y(n_507)
);

AOI22xp5_ASAP7_75t_L g533 ( 
.A1(n_507),
.A2(n_486),
.B1(n_9),
.B2(n_10),
.Y(n_533)
);

CKINVDCx20_ASAP7_75t_R g508 ( 
.A(n_495),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_508),
.B(n_511),
.Y(n_528)
);

NOR2xp67_ASAP7_75t_SL g535 ( 
.A(n_512),
.B(n_518),
.Y(n_535)
);

BUFx24_ASAP7_75t_SL g513 ( 
.A(n_504),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g536 ( 
.A(n_513),
.B(n_517),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_503),
.B(n_470),
.Y(n_517)
);

MAJIxp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_474),
.C(n_463),
.Y(n_518)
);

FAx1_ASAP7_75t_SL g520 ( 
.A(n_504),
.B(n_462),
.CI(n_474),
.CON(n_520),
.SN(n_520)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_520),
.B(n_6),
.Y(n_534)
);

CKINVDCx16_ASAP7_75t_R g521 ( 
.A(n_487),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_SL g526 ( 
.A(n_521),
.B(n_524),
.Y(n_526)
);

OAI21xp5_ASAP7_75t_SL g530 ( 
.A1(n_523),
.A2(n_496),
.B(n_487),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_499),
.B(n_476),
.C(n_484),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g525 ( 
.A(n_493),
.B(n_456),
.C(n_485),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_525),
.B(n_6),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g527 ( 
.A(n_518),
.B(n_489),
.C(n_488),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_527),
.B(n_529),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g529 ( 
.A(n_512),
.B(n_524),
.C(n_510),
.Y(n_529)
);

AOI21xp5_ASAP7_75t_L g545 ( 
.A1(n_530),
.A2(n_523),
.B(n_516),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_510),
.B(n_491),
.C(n_501),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_531),
.B(n_532),
.Y(n_549)
);

MAJIxp5_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_492),
.C(n_456),
.Y(n_532)
);

OR2x2_ASAP7_75t_L g544 ( 
.A(n_533),
.B(n_534),
.Y(n_544)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_519),
.B(n_6),
.Y(n_537)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_537),
.Y(n_547)
);

CKINVDCx20_ASAP7_75t_R g538 ( 
.A(n_515),
.Y(n_538)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_538),
.B(n_540),
.Y(n_554)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_539),
.Y(n_548)
);

XOR2xp5_ASAP7_75t_L g540 ( 
.A(n_519),
.B(n_514),
.Y(n_540)
);

CKINVDCx20_ASAP7_75t_R g541 ( 
.A(n_509),
.Y(n_541)
);

CKINVDCx20_ASAP7_75t_R g551 ( 
.A(n_541),
.Y(n_551)
);

OAI22xp5_ASAP7_75t_SL g542 ( 
.A1(n_522),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_SL g550 ( 
.A1(n_542),
.A2(n_520),
.B1(n_525),
.B2(n_11),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_529),
.B(n_535),
.C(n_527),
.Y(n_543)
);

NOR2xp67_ASAP7_75t_SL g560 ( 
.A(n_543),
.B(n_542),
.Y(n_560)
);

AOI22xp5_ASAP7_75t_L g561 ( 
.A1(n_545),
.A2(n_552),
.B1(n_0),
.B2(n_1),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g559 ( 
.A(n_550),
.B(n_533),
.Y(n_559)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_526),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_552)
);

AOI22xp33_ASAP7_75t_SL g553 ( 
.A1(n_528),
.A2(n_16),
.B1(n_12),
.B2(n_2),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g557 ( 
.A1(n_553),
.A2(n_555),
.B(n_530),
.Y(n_557)
);

OR2x2_ASAP7_75t_L g555 ( 
.A(n_534),
.B(n_532),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g556 ( 
.A(n_543),
.B(n_531),
.C(n_540),
.Y(n_556)
);

NAND2xp5_ASAP7_75t_L g565 ( 
.A(n_556),
.B(n_557),
.Y(n_565)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_546),
.B(n_536),
.C(n_537),
.Y(n_558)
);

AND2x2_ASAP7_75t_L g568 ( 
.A(n_558),
.B(n_563),
.Y(n_568)
);

NOR2xp33_ASAP7_75t_L g566 ( 
.A(n_559),
.B(n_555),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_560),
.B(n_549),
.C(n_550),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_SL g564 ( 
.A(n_561),
.B(n_562),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_554),
.B(n_5),
.Y(n_562)
);

AOI21xp5_ASAP7_75t_L g563 ( 
.A1(n_551),
.A2(n_5),
.B(n_1),
.Y(n_563)
);

OAI211xp5_ASAP7_75t_L g570 ( 
.A1(n_566),
.A2(n_567),
.B(n_547),
.C(n_548),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g569 ( 
.A(n_568),
.B(n_556),
.Y(n_569)
);

OAI21xp5_ASAP7_75t_SL g572 ( 
.A1(n_569),
.A2(n_570),
.B(n_571),
.Y(n_572)
);

OAI21xp5_ASAP7_75t_SL g571 ( 
.A1(n_565),
.A2(n_544),
.B(n_553),
.Y(n_571)
);

OAI311xp33_ASAP7_75t_L g573 ( 
.A1(n_570),
.A2(n_544),
.A3(n_564),
.B1(n_3),
.C1(n_4),
.Y(n_573)
);

AOI21xp5_ASAP7_75t_L g574 ( 
.A1(n_573),
.A2(n_0),
.B(n_1),
.Y(n_574)
);

AOI211x1_ASAP7_75t_L g575 ( 
.A1(n_574),
.A2(n_572),
.B(n_3),
.C(n_4),
.Y(n_575)
);

AOI21xp5_ASAP7_75t_SL g576 ( 
.A1(n_575),
.A2(n_0),
.B(n_3),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_576),
.B(n_3),
.Y(n_577)
);

AOI21xp5_ASAP7_75t_L g578 ( 
.A1(n_577),
.A2(n_4),
.B(n_5),
.Y(n_578)
);


endmodule