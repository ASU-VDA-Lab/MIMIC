module fake_jpeg_6317_n_102 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_35, n_4, n_34, n_30, n_39, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_12, n_32, n_8, n_15, n_7, n_102);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_35;
input n_4;
input n_34;
input n_30;
input n_39;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_102;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_43;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_30),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_27),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_24),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_1),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_15),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_18),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_32),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_33),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_26),
.Y(n_57)
);

BUFx10_ASAP7_75t_L g58 ( 
.A(n_2),
.Y(n_58)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_16),
.Y(n_59)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_58),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_60),
.Y(n_67)
);

AND2x2_ASAP7_75t_SL g61 ( 
.A(n_41),
.B(n_0),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_65),
.B(n_44),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_1),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_48),
.Y(n_66)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_58),
.Y(n_63)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_47),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_64),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_5),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_66),
.B(n_45),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_65),
.A2(n_59),
.B1(n_42),
.B2(n_56),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g74 ( 
.A1(n_68),
.A2(n_72),
.B1(n_40),
.B2(n_46),
.Y(n_74)
);

OAI21xp33_ASAP7_75t_L g73 ( 
.A1(n_70),
.A2(n_57),
.B(n_50),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g72 ( 
.A1(n_61),
.A2(n_55),
.B1(n_43),
.B2(n_53),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g84 ( 
.A1(n_73),
.A2(n_67),
.B(n_9),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_74),
.B(n_75),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_71),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_76),
.B(n_77),
.Y(n_81)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_69),
.Y(n_77)
);

O2A1O1Ixp33_ASAP7_75t_L g78 ( 
.A1(n_73),
.A2(n_67),
.B(n_54),
.C(n_52),
.Y(n_78)
);

AO22x1_ASAP7_75t_SL g86 ( 
.A1(n_78),
.A2(n_80),
.B1(n_6),
.B2(n_11),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_73),
.A2(n_51),
.B1(n_7),
.B2(n_8),
.Y(n_80)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_82),
.B(n_83),
.Y(n_88)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_84),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g85 ( 
.A(n_74),
.Y(n_85)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_85),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_86),
.A2(n_79),
.B(n_85),
.Y(n_90)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_90),
.B(n_91),
.C(n_89),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g91 ( 
.A(n_88),
.B(n_81),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_87),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_93),
.Y(n_94)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_12),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_13),
.B1(n_14),
.B2(n_17),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_96),
.A2(n_39),
.B1(n_20),
.B2(n_21),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g98 ( 
.A(n_97),
.B(n_19),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g99 ( 
.A1(n_98),
.A2(n_37),
.B(n_25),
.Y(n_99)
);

FAx1_ASAP7_75t_SL g100 ( 
.A(n_99),
.B(n_23),
.CI(n_28),
.CON(n_100),
.SN(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_100),
.B(n_36),
.Y(n_101)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_101),
.B(n_31),
.Y(n_102)
);


endmodule