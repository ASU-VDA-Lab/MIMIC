module fake_jpeg_32118_n_350 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_350);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_350;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_7),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_9),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_11),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx24_ASAP7_75t_L g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_1),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx12_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_8),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx16f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_8),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_39),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_40),
.B(n_47),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_41),
.Y(n_85)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx11_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_43),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_14),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_44),
.Y(n_98)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_35),
.Y(n_45)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_45),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_14),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_46),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_15),
.B(n_13),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_48),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g49 ( 
.A(n_15),
.B(n_13),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_56),
.Y(n_105)
);

BUFx5_ASAP7_75t_L g50 ( 
.A(n_25),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_50),
.Y(n_104)
);

INVx6_ASAP7_75t_SL g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g80 ( 
.A(n_51),
.Y(n_80)
);

BUFx5_ASAP7_75t_L g52 ( 
.A(n_25),
.Y(n_52)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_52),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g53 ( 
.A(n_18),
.B(n_13),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_53),
.B(n_57),
.Y(n_117)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_25),
.Y(n_54)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_25),
.Y(n_55)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_55),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_39),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_30),
.B(n_0),
.Y(n_57)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_14),
.Y(n_58)
);

INVx4_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

NAND2x1_ASAP7_75t_L g59 ( 
.A(n_32),
.B(n_0),
.Y(n_59)
);

MAJIxp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_16),
.C(n_38),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_31),
.B(n_0),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_60),
.B(n_61),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_39),
.Y(n_61)
);

BUFx5_ASAP7_75t_L g62 ( 
.A(n_25),
.Y(n_62)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_32),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_63),
.B(n_68),
.Y(n_125)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_26),
.Y(n_64)
);

BUFx8_ASAP7_75t_L g91 ( 
.A(n_64),
.Y(n_91)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_35),
.Y(n_65)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_66),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g67 ( 
.A(n_21),
.Y(n_67)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_18),
.B(n_0),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_69),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_26),
.Y(n_70)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_22),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_71),
.B(n_29),
.Y(n_126)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_17),
.Y(n_72)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_72),
.Y(n_121)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_73),
.Y(n_124)
);

INVx11_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx6_ASAP7_75t_L g113 ( 
.A(n_74),
.Y(n_113)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_75),
.Y(n_100)
);

INVx1_ASAP7_75t_SL g76 ( 
.A(n_20),
.Y(n_76)
);

CKINVDCx14_ASAP7_75t_R g88 ( 
.A(n_76),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_77),
.B(n_93),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_73),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_82),
.A2(n_84),
.B1(n_101),
.B2(n_107),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_41),
.A2(n_21),
.B1(n_28),
.B2(n_23),
.Y(n_84)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_45),
.A2(n_28),
.B1(n_23),
.B2(n_19),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_57),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g145 ( 
.A(n_95),
.B(n_112),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_71),
.A2(n_22),
.B1(n_33),
.B2(n_19),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_106),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_64),
.A2(n_24),
.B1(n_19),
.B2(n_33),
.Y(n_101)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

HB1xp67_ASAP7_75t_L g141 ( 
.A(n_103),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_48),
.A2(n_33),
.B1(n_24),
.B2(n_38),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_64),
.A2(n_24),
.B1(n_37),
.B2(n_20),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_66),
.A2(n_37),
.B1(n_36),
.B2(n_34),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_108),
.A2(n_123),
.B1(n_75),
.B2(n_70),
.Y(n_156)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_109),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g110 ( 
.A1(n_72),
.A2(n_30),
.B1(n_34),
.B2(n_36),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_110),
.B(n_118),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_63),
.B(n_27),
.C(n_16),
.Y(n_112)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_61),
.Y(n_114)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_114),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_76),
.B(n_27),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_44),
.A2(n_29),
.B1(n_2),
.B2(n_3),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_120),
.B(n_1),
.Y(n_144)
);

INVx6_ASAP7_75t_L g122 ( 
.A(n_46),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_122),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_65),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_126),
.B(n_29),
.Y(n_149)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_128),
.Y(n_173)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_121),
.Y(n_129)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_129),
.Y(n_175)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_78),
.Y(n_130)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_130),
.Y(n_180)
);

INVx4_ASAP7_75t_SL g131 ( 
.A(n_80),
.Y(n_131)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_100),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_138),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_117),
.B(n_59),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_SL g183 ( 
.A(n_134),
.B(n_149),
.Y(n_183)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_59),
.C(n_69),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx5_ASAP7_75t_L g185 ( 
.A(n_139),
.Y(n_185)
);

INVx6_ASAP7_75t_L g140 ( 
.A(n_85),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g172 ( 
.A(n_140),
.Y(n_172)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_81),
.Y(n_143)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_143),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g196 ( 
.A(n_144),
.B(n_123),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_105),
.B(n_51),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_160),
.Y(n_204)
);

A2O1A1Ixp33_ASAP7_75t_L g147 ( 
.A1(n_116),
.A2(n_75),
.B(n_70),
.C(n_66),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_147),
.B(n_91),
.Y(n_199)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_115),
.Y(n_148)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_148),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_125),
.B(n_29),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_150),
.B(n_154),
.Y(n_188)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_85),
.Y(n_151)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_151),
.Y(n_179)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_113),
.Y(n_153)
);

INVx3_ASAP7_75t_L g176 ( 
.A(n_153),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_88),
.B(n_54),
.Y(n_154)
);

BUFx12f_ASAP7_75t_L g155 ( 
.A(n_80),
.Y(n_155)
);

BUFx4f_ASAP7_75t_SL g201 ( 
.A(n_155),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_156),
.A2(n_58),
.B1(n_87),
.B2(n_62),
.Y(n_198)
);

AND2x6_ASAP7_75t_L g157 ( 
.A(n_108),
.B(n_75),
.Y(n_157)
);

AND2x6_ASAP7_75t_L g192 ( 
.A(n_157),
.B(n_101),
.Y(n_192)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_158),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_119),
.B(n_93),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_159),
.B(n_161),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_122),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_102),
.B(n_29),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_124),
.B(n_42),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_162),
.B(n_169),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_98),
.Y(n_163)
);

INVx8_ASAP7_75t_L g178 ( 
.A(n_163),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_91),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_165),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_83),
.B(n_43),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_83),
.B(n_52),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_166),
.B(n_167),
.Y(n_205)
);

INVx5_ASAP7_75t_L g167 ( 
.A(n_79),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_89),
.B(n_50),
.Y(n_168)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_96),
.B(n_3),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_104),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g200 ( 
.A(n_170),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g171 ( 
.A(n_107),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_171),
.B(n_55),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_86),
.B1(n_94),
.B2(n_90),
.Y(n_177)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_177),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_145),
.B(n_133),
.C(n_147),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_181),
.B(n_196),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_L g182 ( 
.A1(n_135),
.A2(n_142),
.B1(n_137),
.B2(n_156),
.Y(n_182)
);

INVxp67_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_157),
.A2(n_74),
.B(n_91),
.Y(n_184)
);

OAI21xp5_ASAP7_75t_L g238 ( 
.A1(n_184),
.A2(n_207),
.B(n_196),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_L g189 ( 
.A1(n_142),
.A2(n_111),
.B1(n_98),
.B2(n_96),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_189),
.A2(n_131),
.B1(n_170),
.B2(n_139),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_141),
.A2(n_94),
.B(n_86),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_190),
.A2(n_192),
.B(n_207),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_143),
.A2(n_84),
.B1(n_82),
.B2(n_111),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_193),
.A2(n_197),
.B1(n_163),
.B2(n_158),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_127),
.A2(n_67),
.B1(n_136),
.B2(n_152),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_198),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_233)
);

OR2x2_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_4),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g208 ( 
.A(n_202),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_208),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_206),
.B(n_204),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_209),
.B(n_211),
.Y(n_265)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_187),
.Y(n_210)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_210),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_206),
.B(n_204),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_188),
.B(n_183),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_214),
.B(n_222),
.Y(n_255)
);

AO22x2_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_151),
.B1(n_140),
.B2(n_152),
.Y(n_215)
);

AO22x1_ASAP7_75t_SL g243 ( 
.A1(n_215),
.A2(n_172),
.B1(n_176),
.B2(n_185),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_181),
.B(n_199),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g252 ( 
.A(n_216),
.B(n_217),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_195),
.B(n_127),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_226),
.Y(n_251)
);

OAI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_220),
.A2(n_233),
.B1(n_200),
.B2(n_178),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_136),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g256 ( 
.A(n_221),
.B(n_231),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_173),
.B(n_155),
.Y(n_222)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_187),
.Y(n_224)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_224),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_SL g225 ( 
.A1(n_185),
.A2(n_155),
.B1(n_87),
.B2(n_153),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_225),
.A2(n_230),
.B(n_200),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_175),
.B(n_130),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_186),
.B(n_167),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_227),
.B(n_228),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_191),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_229),
.A2(n_193),
.B1(n_179),
.B2(n_178),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_174),
.B(n_132),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_190),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_232),
.B(n_236),
.Y(n_260)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_180),
.Y(n_234)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_234),
.Y(n_250)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_203),
.Y(n_235)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_235),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_197),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_196),
.B(n_4),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_SL g257 ( 
.A(n_237),
.B(n_6),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_238),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_176),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_L g258 ( 
.A1(n_239),
.A2(n_201),
.B(n_7),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g242 ( 
.A1(n_232),
.A2(n_184),
.B(n_198),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g270 ( 
.A(n_242),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_243),
.B(n_247),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g284 ( 
.A1(n_244),
.A2(n_245),
.B1(n_220),
.B2(n_227),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_219),
.A2(n_179),
.B1(n_172),
.B2(n_194),
.Y(n_247)
);

AO21x1_ASAP7_75t_L g276 ( 
.A1(n_249),
.A2(n_258),
.B(n_225),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_212),
.A2(n_201),
.B(n_194),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g282 ( 
.A(n_253),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g267 ( 
.A(n_257),
.B(n_237),
.Y(n_267)
);

AND2x2_ASAP7_75t_L g275 ( 
.A(n_258),
.B(n_222),
.Y(n_275)
);

AOI21xp5_ASAP7_75t_L g261 ( 
.A1(n_212),
.A2(n_238),
.B(n_213),
.Y(n_261)
);

NAND2x1_ASAP7_75t_L g281 ( 
.A(n_261),
.B(n_223),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g262 ( 
.A(n_216),
.B(n_201),
.C(n_7),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_262),
.B(n_230),
.C(n_209),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_229),
.A2(n_6),
.B1(n_8),
.B2(n_236),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_263),
.B(n_233),
.Y(n_269)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_210),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_264),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_267),
.B(n_277),
.Y(n_302)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_269),
.Y(n_293)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_259),
.Y(n_271)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_271),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_211),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_272),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_246),
.B(n_214),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g304 ( 
.A(n_273),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_255),
.B(n_254),
.Y(n_274)
);

HB1xp67_ASAP7_75t_L g303 ( 
.A(n_274),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_275),
.A2(n_279),
.B1(n_280),
.B2(n_283),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_276),
.A2(n_249),
.B(n_233),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_251),
.B(n_208),
.Y(n_277)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_252),
.B(n_223),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_278),
.B(n_285),
.C(n_252),
.Y(n_297)
);

INVx13_ASAP7_75t_L g279 ( 
.A(n_259),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_265),
.B(n_218),
.Y(n_280)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_281),
.A2(n_287),
.B(n_231),
.Y(n_300)
);

CKINVDCx20_ASAP7_75t_R g283 ( 
.A(n_260),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_284),
.A2(n_286),
.B1(n_240),
.B2(n_244),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_256),
.B(n_221),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_288),
.A2(n_292),
.B1(n_295),
.B2(n_299),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_282),
.A2(n_245),
.B1(n_253),
.B2(n_270),
.Y(n_289)
);

OAI22xp5_ASAP7_75t_SL g311 ( 
.A1(n_289),
.A2(n_291),
.B1(n_294),
.B2(n_293),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_282),
.A2(n_242),
.B1(n_261),
.B2(n_240),
.Y(n_291)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_284),
.A2(n_270),
.B1(n_268),
.B2(n_269),
.Y(n_292)
);

AOI21x1_ASAP7_75t_SL g294 ( 
.A1(n_276),
.A2(n_243),
.B(n_215),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_268),
.A2(n_263),
.B1(n_215),
.B2(n_243),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_297),
.B(n_298),
.C(n_267),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_256),
.C(n_262),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g308 ( 
.A(n_300),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_297),
.B(n_286),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_305),
.B(n_306),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_302),
.B(n_285),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_307),
.B(n_313),
.C(n_314),
.Y(n_324)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_303),
.Y(n_309)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_309),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_293),
.A2(n_275),
.B1(n_266),
.B2(n_287),
.Y(n_310)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_310),
.B(n_315),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_311),
.A2(n_292),
.B1(n_299),
.B2(n_294),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_302),
.B(n_272),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_298),
.B(n_215),
.C(n_281),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_288),
.A2(n_275),
.B1(n_215),
.B2(n_281),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_300),
.B(n_215),
.C(n_271),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_317),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_295),
.A2(n_266),
.B1(n_241),
.B2(n_264),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_318),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_304),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_321),
.B(n_326),
.Y(n_333)
);

OAI21xp5_ASAP7_75t_L g322 ( 
.A1(n_312),
.A2(n_291),
.B(n_289),
.Y(n_322)
);

OAI21xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_301),
.B(n_307),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_323),
.A2(n_315),
.B1(n_290),
.B2(n_247),
.Y(n_331)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_306),
.B(n_296),
.Y(n_326)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_314),
.B(n_296),
.Y(n_327)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_327),
.A2(n_313),
.B(n_305),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_320),
.A2(n_290),
.B1(n_312),
.B2(n_316),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_330),
.B(n_335),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_334),
.Y(n_340)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_332),
.A2(n_322),
.B(n_328),
.Y(n_338)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_325),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_319),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_336),
.A2(n_324),
.B(n_329),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_332),
.B(n_324),
.C(n_329),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_337),
.B(n_333),
.Y(n_344)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_338),
.B(n_339),
.Y(n_343)
);

OR2x2_ASAP7_75t_L g342 ( 
.A(n_340),
.B(n_304),
.Y(n_342)
);

AOI322xp5_ASAP7_75t_L g345 ( 
.A1(n_342),
.A2(n_344),
.A3(n_279),
.B1(n_248),
.B2(n_250),
.C1(n_341),
.C2(n_228),
.Y(n_345)
);

OAI22xp5_ASAP7_75t_L g347 ( 
.A1(n_345),
.A2(n_346),
.B1(n_217),
.B2(n_224),
.Y(n_347)
);

AOI322xp5_ASAP7_75t_L g346 ( 
.A1(n_343),
.A2(n_330),
.A3(n_327),
.B1(n_323),
.B2(n_326),
.C1(n_250),
.C2(n_239),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_347),
.B(n_226),
.C(n_234),
.Y(n_348)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_235),
.B1(n_230),
.B2(n_257),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_6),
.Y(n_350)
);


endmodule