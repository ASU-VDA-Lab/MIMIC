module fake_jpeg_5825_n_331 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_331);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_331;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_27;
wire n_179;
wire n_185;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_2),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_7),
.B(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_9),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_6),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx3_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_23),
.Y(n_36)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_39),
.Y(n_59)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_38),
.B(n_34),
.Y(n_72)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx11_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_23),
.Y(n_41)
);

OR2x2_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

BUFx2_ASAP7_75t_R g42 ( 
.A(n_23),
.Y(n_42)
);

INVx2_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_43),
.B(n_21),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_24),
.B(n_0),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_44),
.B(n_45),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_0),
.Y(n_45)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_48),
.Y(n_74)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_47),
.B(n_60),
.Y(n_77)
);

INVx2_ASAP7_75t_SL g48 ( 
.A(n_41),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

HB1xp67_ASAP7_75t_L g97 ( 
.A(n_49),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_42),
.A2(n_29),
.B1(n_32),
.B2(n_27),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_51),
.A2(n_52),
.B1(n_56),
.B2(n_64),
.Y(n_94)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_42),
.A2(n_27),
.B1(n_22),
.B2(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_53),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_42),
.A2(n_22),
.B1(n_19),
.B2(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_57),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_41),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g87 ( 
.A(n_58),
.Y(n_87)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_61),
.B(n_71),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_35),
.Y(n_63)
);

INVx5_ASAP7_75t_L g78 ( 
.A(n_63),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_42),
.A2(n_25),
.B1(n_17),
.B2(n_24),
.Y(n_64)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_66),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_39),
.A2(n_18),
.B1(n_25),
.B2(n_30),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

AO22x1_ASAP7_75t_SL g68 ( 
.A1(n_44),
.A2(n_34),
.B1(n_30),
.B2(n_26),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_68),
.A2(n_70),
.B1(n_18),
.B2(n_43),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx5_ASAP7_75t_L g83 ( 
.A(n_69),
.Y(n_83)
);

AOI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_39),
.A2(n_24),
.B1(n_30),
.B2(n_26),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_44),
.B(n_31),
.Y(n_71)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_65),
.B(n_45),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_73),
.B(n_75),
.Y(n_121)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_65),
.B(n_62),
.Y(n_75)
);

OAI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_68),
.A2(n_39),
.B1(n_40),
.B2(n_43),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_76),
.A2(n_54),
.B1(n_40),
.B2(n_61),
.Y(n_105)
);

INVx13_ASAP7_75t_L g79 ( 
.A(n_47),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_79),
.B(n_92),
.Y(n_107)
);

O2A1O1Ixp33_ASAP7_75t_L g80 ( 
.A1(n_68),
.A2(n_45),
.B(n_44),
.C(n_35),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g106 ( 
.A1(n_80),
.A2(n_93),
.B1(n_66),
.B2(n_48),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g82 ( 
.A(n_62),
.B(n_38),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_82),
.B(n_99),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_45),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_86),
.B(n_90),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_68),
.B(n_37),
.Y(n_90)
);

NAND3xp33_ASAP7_75t_L g91 ( 
.A(n_62),
.B(n_50),
.C(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_91),
.A2(n_55),
.B1(n_57),
.B2(n_49),
.Y(n_124)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_59),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_96),
.B(n_46),
.Y(n_113)
);

CKINVDCx6p67_ASAP7_75t_R g98 ( 
.A(n_50),
.Y(n_98)
);

INVx5_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_48),
.B(n_43),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_72),
.B(n_37),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g108 ( 
.A(n_100),
.B(n_73),
.Y(n_108)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_77),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_102),
.B(n_104),
.Y(n_136)
);

CKINVDCx5p33_ASAP7_75t_R g104 ( 
.A(n_98),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_105),
.A2(n_106),
.B1(n_110),
.B2(n_112),
.Y(n_130)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_108),
.B(n_129),
.Y(n_144)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_77),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_109),
.B(n_111),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g110 ( 
.A1(n_93),
.A2(n_54),
.B1(n_40),
.B2(n_38),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_100),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_90),
.A2(n_40),
.B1(n_54),
.B2(n_38),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_113),
.B(n_116),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_73),
.B(n_60),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_114),
.B(n_115),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_75),
.B(n_37),
.Y(n_115)
);

INVx2_ASAP7_75t_R g116 ( 
.A(n_98),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g117 ( 
.A1(n_95),
.A2(n_38),
.B1(n_61),
.B2(n_55),
.Y(n_117)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_117),
.Y(n_131)
);

INVx4_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_75),
.B(n_20),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_125),
.Y(n_143)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_74),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_120),
.B(n_123),
.Y(n_155)
);

AOI22x1_ASAP7_75t_SL g122 ( 
.A1(n_94),
.A2(n_53),
.B1(n_58),
.B2(n_46),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_122),
.A2(n_95),
.B1(n_88),
.B2(n_84),
.Y(n_132)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_78),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g135 ( 
.A1(n_124),
.A2(n_85),
.B(n_84),
.Y(n_135)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_74),
.Y(n_125)
);

INVx13_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

INVx3_ASAP7_75t_L g154 ( 
.A(n_127),
.Y(n_154)
);

HB1xp67_ASAP7_75t_L g128 ( 
.A(n_78),
.Y(n_128)
);

INVxp33_ASAP7_75t_SL g141 ( 
.A(n_128),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g129 ( 
.A(n_82),
.B(n_58),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_132),
.A2(n_124),
.B1(n_122),
.B2(n_106),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_107),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_134),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_135),
.A2(n_158),
.B(n_98),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_107),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_139),
.Y(n_184)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_113),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_140),
.B(n_142),
.Y(n_181)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_112),
.Y(n_142)
);

CKINVDCx14_ASAP7_75t_R g145 ( 
.A(n_126),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_145),
.B(n_149),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g146 ( 
.A(n_108),
.B(n_114),
.Y(n_146)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_146),
.B(n_153),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_88),
.B1(n_80),
.B2(n_82),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

OR2x2_ASAP7_75t_L g148 ( 
.A(n_101),
.B(n_99),
.Y(n_148)
);

AOI21xp5_ASAP7_75t_SL g192 ( 
.A1(n_148),
.A2(n_28),
.B(n_21),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_103),
.B(n_86),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_151),
.B(n_111),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_126),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_152),
.B(n_157),
.Y(n_167)
);

MAJx2_ASAP7_75t_L g153 ( 
.A(n_121),
.B(n_85),
.C(n_99),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g156 ( 
.A(n_103),
.B(n_96),
.Y(n_156)
);

XNOR2xp5_ASAP7_75t_L g172 ( 
.A(n_156),
.B(n_129),
.Y(n_172)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_115),
.Y(n_157)
);

OAI21xp5_ASAP7_75t_SL g158 ( 
.A1(n_101),
.A2(n_92),
.B(n_81),
.Y(n_158)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_121),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_159),
.B(n_160),
.Y(n_179)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_116),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_161),
.B(n_188),
.Y(n_194)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_141),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_162),
.B(n_163),
.Y(n_215)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_136),
.Y(n_163)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_164),
.A2(n_173),
.B1(n_183),
.B2(n_185),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g165 ( 
.A(n_146),
.B(n_119),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_165),
.B(n_175),
.C(n_178),
.Y(n_212)
);

NAND2xp33_ASAP7_75t_SL g166 ( 
.A(n_148),
.B(n_101),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g201 ( 
.A1(n_166),
.A2(n_192),
.B(n_143),
.Y(n_201)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_155),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g208 ( 
.A(n_168),
.B(n_174),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_137),
.A2(n_147),
.B(n_158),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_171),
.A2(n_186),
.B(n_143),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g218 ( 
.A(n_172),
.B(n_169),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_142),
.A2(n_129),
.B1(n_120),
.B2(n_125),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_133),
.Y(n_174)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_135),
.B(n_109),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_130),
.A2(n_102),
.B1(n_116),
.B2(n_83),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_176),
.A2(n_154),
.B1(n_69),
.B2(n_63),
.Y(n_214)
);

OAI21xp5_ASAP7_75t_SL g217 ( 
.A1(n_177),
.A2(n_87),
.B(n_1),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g178 ( 
.A(n_156),
.B(n_83),
.Y(n_178)
);

OAI22xp33_ASAP7_75t_SL g180 ( 
.A1(n_159),
.A2(n_97),
.B1(n_128),
.B2(n_104),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_180),
.A2(n_160),
.B1(n_140),
.B2(n_131),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_132),
.A2(n_55),
.B1(n_53),
.B2(n_118),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_130),
.A2(n_118),
.B1(n_89),
.B2(n_26),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_144),
.A2(n_127),
.B(n_79),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_151),
.B(n_127),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_134),
.B(n_139),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_189),
.B(n_191),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_138),
.Y(n_190)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_190),
.Y(n_193)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_138),
.Y(n_191)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_188),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_196),
.Y(n_225)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_187),
.Y(n_196)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_197),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_R g198 ( 
.A(n_166),
.B(n_153),
.Y(n_198)
);

AOI21xp5_ASAP7_75t_L g222 ( 
.A1(n_198),
.A2(n_199),
.B(n_201),
.Y(n_222)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_161),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_200),
.B(n_205),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_182),
.A2(n_157),
.B1(n_177),
.B2(n_131),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_202),
.A2(n_203),
.B1(n_209),
.B2(n_217),
.Y(n_240)
);

OAI22x1_ASAP7_75t_SL g203 ( 
.A1(n_182),
.A2(n_144),
.B1(n_137),
.B2(n_152),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_181),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_191),
.B(n_144),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_206),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_190),
.B(n_149),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_207),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_192),
.A2(n_154),
.B1(n_28),
.B2(n_63),
.Y(n_209)
);

BUFx12f_ASAP7_75t_SL g211 ( 
.A(n_163),
.Y(n_211)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_211),
.Y(n_226)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_167),
.Y(n_213)
);

BUFx24_ASAP7_75t_SL g235 ( 
.A(n_213),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_185),
.B1(n_162),
.B2(n_183),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_178),
.B(n_69),
.C(n_79),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_212),
.C(n_207),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_218),
.B(n_150),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_186),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_172),
.B(n_0),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g237 ( 
.A(n_220),
.Y(n_237)
);

NAND4xp25_ASAP7_75t_L g257 ( 
.A(n_223),
.B(n_246),
.C(n_217),
.D(n_209),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_203),
.A2(n_164),
.B1(n_171),
.B2(n_173),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g264 ( 
.A1(n_224),
.A2(n_228),
.B1(n_229),
.B2(n_230),
.Y(n_264)
);

AOI211xp5_ASAP7_75t_L g227 ( 
.A1(n_198),
.A2(n_175),
.B(n_170),
.C(n_184),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_227),
.A2(n_10),
.B(n_15),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_214),
.A2(n_184),
.B1(n_170),
.B2(n_176),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_206),
.A2(n_174),
.B1(n_179),
.B2(n_169),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_201),
.A2(n_165),
.B1(n_150),
.B2(n_89),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_231),
.B(n_212),
.C(n_220),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_200),
.A2(n_195),
.B1(n_193),
.B2(n_204),
.Y(n_233)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_204),
.A2(n_89),
.B1(n_150),
.B2(n_3),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g247 ( 
.A1(n_234),
.A2(n_205),
.B1(n_213),
.B2(n_196),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_238),
.B(n_245),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_193),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_241)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_241),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_202),
.A2(n_15),
.B1(n_14),
.B2(n_13),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_242),
.B(n_244),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_211),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_16),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_194),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_246)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_247),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_236),
.B(n_194),
.Y(n_249)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_249),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g250 ( 
.A1(n_221),
.A2(n_240),
.B1(n_234),
.B2(n_232),
.Y(n_250)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_250),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_239),
.B(n_210),
.Y(n_251)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_251),
.Y(n_281)
);

BUFx2_ASAP7_75t_L g252 ( 
.A(n_239),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_252),
.B(n_256),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g253 ( 
.A1(n_226),
.A2(n_199),
.B1(n_216),
.B2(n_219),
.Y(n_253)
);

OA22x2_ASAP7_75t_L g278 ( 
.A1(n_253),
.A2(n_257),
.B1(n_246),
.B2(n_241),
.Y(n_278)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_255),
.B(n_258),
.C(n_266),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_225),
.B(n_208),
.Y(n_256)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_231),
.B(n_215),
.C(n_3),
.Y(n_258)
);

CKINVDCx14_ASAP7_75t_R g279 ( 
.A(n_259),
.Y(n_279)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_226),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_260),
.A2(n_261),
.B(n_262),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_233),
.B(n_2),
.Y(n_261)
);

CKINVDCx20_ASAP7_75t_R g262 ( 
.A(n_243),
.Y(n_262)
);

BUFx12_ASAP7_75t_L g263 ( 
.A(n_238),
.Y(n_263)
);

INVxp67_ASAP7_75t_L g283 ( 
.A(n_263),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_230),
.B(n_5),
.C(n_6),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_254),
.B(n_222),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g291 ( 
.A(n_268),
.B(n_271),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_267),
.A2(n_227),
.B1(n_224),
.B2(n_228),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_269),
.A2(n_267),
.B1(n_250),
.B2(n_253),
.Y(n_287)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_245),
.Y(n_271)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_263),
.B(n_229),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_273),
.B(n_5),
.C(n_6),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_223),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_275),
.B(n_264),
.Y(n_289)
);

AO21x1_ASAP7_75t_L g284 ( 
.A1(n_278),
.A2(n_259),
.B(n_257),
.Y(n_284)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_260),
.A2(n_237),
.B(n_235),
.Y(n_282)
);

AOI21xp5_ASAP7_75t_L g286 ( 
.A1(n_282),
.A2(n_248),
.B(n_249),
.Y(n_286)
);

AO21x1_ASAP7_75t_L g302 ( 
.A1(n_284),
.A2(n_279),
.B(n_273),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g285 ( 
.A(n_280),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_L g301 ( 
.A1(n_285),
.A2(n_292),
.B(n_294),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_286),
.B(n_276),
.Y(n_306)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_278),
.B1(n_283),
.B2(n_269),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_258),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g300 ( 
.A(n_288),
.B(n_290),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_289),
.B(n_297),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_275),
.B(n_265),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_252),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_274),
.A2(n_247),
.B1(n_266),
.B2(n_261),
.Y(n_293)
);

INVxp67_ASAP7_75t_L g303 ( 
.A(n_293),
.Y(n_303)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_277),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_270),
.B(n_255),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g307 ( 
.A(n_295),
.B(n_271),
.Y(n_307)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_278),
.A2(n_263),
.B1(n_6),
.B2(n_7),
.Y(n_296)
);

CKINVDCx16_ASAP7_75t_R g309 ( 
.A(n_296),
.Y(n_309)
);

OR2x2_ASAP7_75t_L g298 ( 
.A(n_284),
.B(n_278),
.Y(n_298)
);

AND2x4_ASAP7_75t_L g317 ( 
.A(n_298),
.B(n_302),
.Y(n_317)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_299),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g304 ( 
.A1(n_287),
.A2(n_283),
.B(n_276),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g311 ( 
.A(n_304),
.B(n_307),
.C(n_308),
.Y(n_311)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_306),
.B(n_305),
.Y(n_310)
);

AOI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_289),
.A2(n_268),
.B1(n_12),
.B2(n_13),
.Y(n_308)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_310),
.Y(n_319)
);

AOI21xp5_ASAP7_75t_SL g312 ( 
.A1(n_303),
.A2(n_298),
.B(n_302),
.Y(n_312)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_312),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_303),
.B(n_293),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_314),
.B(n_315),
.C(n_316),
.Y(n_321)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_291),
.C(n_296),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_309),
.B(n_297),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_291),
.Y(n_318)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_318),
.B(n_10),
.Y(n_322)
);

AOI322xp5_ASAP7_75t_L g320 ( 
.A1(n_317),
.A2(n_285),
.A3(n_12),
.B1(n_14),
.B2(n_10),
.C1(n_11),
.C2(n_16),
.Y(n_320)
);

BUFx24_ASAP7_75t_SL g327 ( 
.A(n_320),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_SL g326 ( 
.A(n_322),
.B(n_323),
.Y(n_326)
);

HB1xp67_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

OAI321xp33_ASAP7_75t_L g328 ( 
.A1(n_324),
.A2(n_325),
.A3(n_7),
.B1(n_8),
.B2(n_9),
.C(n_321),
.Y(n_328)
);

AOI322xp5_ASAP7_75t_L g325 ( 
.A1(n_313),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_11),
.C1(n_15),
.C2(n_311),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g329 ( 
.A1(n_326),
.A2(n_328),
.B(n_324),
.Y(n_329)
);

MAJIxp5_ASAP7_75t_L g330 ( 
.A(n_329),
.B(n_319),
.C(n_327),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_330),
.B(n_8),
.Y(n_331)
);


endmodule