module fake_ariane_884_n_185 (n_8, n_24, n_7, n_22, n_1, n_6, n_13, n_20, n_27, n_29, n_17, n_4, n_2, n_18, n_28, n_9, n_11, n_26, n_3, n_14, n_0, n_19, n_30, n_31, n_16, n_5, n_12, n_15, n_21, n_23, n_10, n_25, n_185);

input n_8;
input n_24;
input n_7;
input n_22;
input n_1;
input n_6;
input n_13;
input n_20;
input n_27;
input n_29;
input n_17;
input n_4;
input n_2;
input n_18;
input n_28;
input n_9;
input n_11;
input n_26;
input n_3;
input n_14;
input n_0;
input n_19;
input n_30;
input n_31;
input n_16;
input n_5;
input n_12;
input n_15;
input n_21;
input n_23;
input n_10;
input n_25;

output n_185;

wire n_83;
wire n_56;
wire n_60;
wire n_170;
wire n_160;
wire n_64;
wire n_180;
wire n_179;
wire n_119;
wire n_124;
wire n_167;
wire n_90;
wire n_38;
wire n_47;
wire n_110;
wire n_153;
wire n_86;
wire n_75;
wire n_89;
wire n_67;
wire n_176;
wire n_149;
wire n_34;
wire n_158;
wire n_172;
wire n_69;
wire n_95;
wire n_175;
wire n_92;
wire n_143;
wire n_183;
wire n_150;
wire n_98;
wire n_74;
wire n_113;
wire n_114;
wire n_33;
wire n_40;
wire n_181;
wire n_152;
wire n_120;
wire n_169;
wire n_106;
wire n_53;
wire n_173;
wire n_111;
wire n_115;
wire n_133;
wire n_66;
wire n_71;
wire n_109;
wire n_96;
wire n_156;
wire n_49;
wire n_174;
wire n_100;
wire n_50;
wire n_132;
wire n_62;
wire n_147;
wire n_51;
wire n_166;
wire n_76;
wire n_103;
wire n_79;
wire n_46;
wire n_84;
wire n_36;
wire n_91;
wire n_159;
wire n_107;
wire n_72;
wire n_105;
wire n_128;
wire n_44;
wire n_82;
wire n_178;
wire n_42;
wire n_57;
wire n_131;
wire n_70;
wire n_117;
wire n_139;
wire n_165;
wire n_85;
wire n_130;
wire n_144;
wire n_48;
wire n_94;
wire n_101;
wire n_134;
wire n_32;
wire n_58;
wire n_37;
wire n_65;
wire n_123;
wire n_138;
wire n_112;
wire n_45;
wire n_162;
wire n_129;
wire n_126;
wire n_137;
wire n_122;
wire n_148;
wire n_164;
wire n_52;
wire n_157;
wire n_184;
wire n_177;
wire n_135;
wire n_73;
wire n_77;
wire n_171;
wire n_118;
wire n_93;
wire n_121;
wire n_61;
wire n_108;
wire n_102;
wire n_182;
wire n_125;
wire n_168;
wire n_43;
wire n_81;
wire n_87;
wire n_41;
wire n_140;
wire n_55;
wire n_151;
wire n_136;
wire n_80;
wire n_146;
wire n_97;
wire n_154;
wire n_142;
wire n_161;
wire n_163;
wire n_88;
wire n_141;
wire n_68;
wire n_116;
wire n_104;
wire n_145;
wire n_78;
wire n_39;
wire n_63;
wire n_59;
wire n_99;
wire n_155;
wire n_127;
wire n_35;
wire n_54;

INVx1_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g35 ( 
.A(n_23),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g37 ( 
.A(n_11),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_0),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_13),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

HB1xp67_ASAP7_75t_L g43 ( 
.A(n_1),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_9),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_1),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_17),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_6),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_18),
.Y(n_49)
);

INVxp33_ASAP7_75t_L g50 ( 
.A(n_8),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_21),
.Y(n_51)
);

CKINVDCx5p33_ASAP7_75t_R g52 ( 
.A(n_26),
.Y(n_52)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

BUFx6f_ASAP7_75t_SL g54 ( 
.A(n_40),
.Y(n_54)
);

AND2x6_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_15),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_34),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_34),
.Y(n_57)
);

INVx2_ASAP7_75t_SL g58 ( 
.A(n_43),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_45),
.B(n_2),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx10_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_41),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_39),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_50),
.B(n_2),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_32),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_67)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_32),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_49),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_51),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_51),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g73 ( 
.A(n_33),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_38),
.B(n_3),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_73),
.A2(n_53),
.B1(n_46),
.B2(n_48),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g76 ( 
.A(n_61),
.B(n_58),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_58),
.Y(n_77)
);

AOI221xp5_ASAP7_75t_L g78 ( 
.A1(n_67),
.A2(n_37),
.B1(n_48),
.B2(n_46),
.C(n_44),
.Y(n_78)
);

HB1xp67_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_61),
.B(n_47),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_52),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_57),
.B(n_64),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_62),
.B(n_35),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_56),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_61),
.B(n_62),
.Y(n_86)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_60),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_64),
.B(n_44),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_60),
.Y(n_89)
);

NAND3xp33_ASAP7_75t_SL g90 ( 
.A(n_66),
.B(n_42),
.C(n_5),
.Y(n_90)
);

AND2x2_ASAP7_75t_L g91 ( 
.A(n_68),
.B(n_4),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_86),
.B(n_83),
.Y(n_92)
);

OAI21x1_ASAP7_75t_L g93 ( 
.A1(n_82),
.A2(n_71),
.B(n_65),
.Y(n_93)
);

BUFx10_ASAP7_75t_L g94 ( 
.A(n_84),
.Y(n_94)
);

CKINVDCx5p33_ASAP7_75t_R g95 ( 
.A(n_79),
.Y(n_95)
);

NAND3xp33_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_71),
.C(n_74),
.Y(n_96)
);

INVxp67_ASAP7_75t_SL g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx4f_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_81),
.A2(n_70),
.B(n_69),
.Y(n_100)
);

A2O1A1Ixp33_ASAP7_75t_L g101 ( 
.A1(n_91),
.A2(n_74),
.B(n_65),
.C(n_70),
.Y(n_101)
);

AO21x1_ASAP7_75t_L g102 ( 
.A1(n_91),
.A2(n_59),
.B(n_69),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_81),
.A2(n_72),
.B(n_68),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_94),
.B(n_80),
.Y(n_105)
);

OA21x2_ASAP7_75t_L g106 ( 
.A1(n_93),
.A2(n_83),
.B(n_89),
.Y(n_106)
);

O2A1O1Ixp5_ASAP7_75t_L g107 ( 
.A1(n_102),
.A2(n_92),
.B(n_101),
.C(n_98),
.Y(n_107)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_97),
.B(n_77),
.Y(n_108)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_96),
.A2(n_90),
.B(n_76),
.C(n_87),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_103),
.A2(n_88),
.B(n_68),
.C(n_72),
.Y(n_110)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_95),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g112 ( 
.A(n_111),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_L g113 ( 
.A1(n_107),
.A2(n_96),
.B(n_100),
.C(n_98),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_108),
.B(n_102),
.Y(n_114)
);

AND2x2_ASAP7_75t_L g115 ( 
.A(n_111),
.B(n_95),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_108),
.B(n_75),
.Y(n_116)
);

HB1xp67_ASAP7_75t_L g117 ( 
.A(n_109),
.Y(n_117)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_104),
.Y(n_118)
);

INVx5_ASAP7_75t_L g119 ( 
.A(n_118),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_117),
.Y(n_120)
);

AND2x4_ASAP7_75t_L g121 ( 
.A(n_116),
.B(n_105),
.Y(n_121)
);

AOI21xp33_ASAP7_75t_L g122 ( 
.A1(n_114),
.A2(n_107),
.B(n_98),
.Y(n_122)
);

AO21x1_ASAP7_75t_L g123 ( 
.A1(n_114),
.A2(n_93),
.B(n_104),
.Y(n_123)
);

AND2x2_ASAP7_75t_L g124 ( 
.A(n_121),
.B(n_85),
.Y(n_124)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_85),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_120),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_115),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g128 ( 
.A(n_119),
.B(n_121),
.Y(n_128)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_119),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_119),
.B(n_87),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g131 ( 
.A(n_119),
.Y(n_131)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_119),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_123),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_122),
.B(n_112),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_133),
.A2(n_113),
.B(n_123),
.Y(n_135)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_126),
.Y(n_136)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_124),
.B(n_106),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_127),
.B(n_89),
.Y(n_138)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_124),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_134),
.A2(n_110),
.B(n_106),
.Y(n_140)
);

NAND2xp33_ASAP7_75t_SL g141 ( 
.A(n_129),
.B(n_94),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g142 ( 
.A(n_126),
.B(n_106),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_135),
.A2(n_133),
.B(n_130),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_125),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g145 ( 
.A(n_138),
.B(n_125),
.C(n_130),
.Y(n_145)
);

AOI211xp5_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_128),
.B(n_110),
.C(n_129),
.Y(n_146)
);

NAND2xp67_ASAP7_75t_SL g147 ( 
.A(n_137),
.B(n_106),
.Y(n_147)
);

O2A1O1Ixp33_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_129),
.B(n_132),
.C(n_131),
.Y(n_148)
);

NAND2x1_ASAP7_75t_L g149 ( 
.A(n_137),
.B(n_132),
.Y(n_149)
);

AOI21xp5_ASAP7_75t_L g150 ( 
.A1(n_141),
.A2(n_131),
.B(n_106),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_131),
.B1(n_55),
.B2(n_54),
.Y(n_151)
);

AND2x2_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_136),
.Y(n_152)
);

AOI32xp33_ASAP7_75t_L g153 ( 
.A1(n_144),
.A2(n_7),
.A3(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_153)
);

OAI21xp33_ASAP7_75t_L g154 ( 
.A1(n_143),
.A2(n_146),
.B(n_145),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_143),
.B(n_136),
.Y(n_155)
);

INVx1_ASAP7_75t_SL g156 ( 
.A(n_150),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_148),
.B(n_7),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g158 ( 
.A(n_147),
.B(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_SL g159 ( 
.A(n_151),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_144),
.Y(n_160)
);

AOI21xp33_ASAP7_75t_SL g161 ( 
.A1(n_154),
.A2(n_153),
.B(n_157),
.Y(n_161)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g163 ( 
.A1(n_156),
.A2(n_99),
.B(n_94),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_158),
.Y(n_164)
);

AND2x4_ASAP7_75t_L g165 ( 
.A(n_152),
.B(n_19),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g166 ( 
.A(n_155),
.B(n_54),
.C(n_25),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_160),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_158),
.B(n_22),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_167),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_167),
.Y(n_170)
);

AOI322xp5_ASAP7_75t_L g171 ( 
.A1(n_161),
.A2(n_159),
.A3(n_54),
.B1(n_55),
.B2(n_30),
.C1(n_27),
.C2(n_29),
.Y(n_171)
);

AOI22x1_ASAP7_75t_L g172 ( 
.A1(n_164),
.A2(n_28),
.B1(n_31),
.B2(n_55),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

INVx2_ASAP7_75t_SL g174 ( 
.A(n_164),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_171),
.A2(n_164),
.B(n_168),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_173),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_173),
.Y(n_177)
);

NAND3xp33_ASAP7_75t_L g178 ( 
.A(n_169),
.B(n_166),
.C(n_163),
.Y(n_178)
);

INVxp67_ASAP7_75t_L g179 ( 
.A(n_170),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_174),
.Y(n_180)
);

AND2x4_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_176),
.Y(n_181)
);

NAND4xp25_ASAP7_75t_L g182 ( 
.A(n_175),
.B(n_165),
.C(n_162),
.D(n_174),
.Y(n_182)
);

AOI22x1_ASAP7_75t_L g183 ( 
.A1(n_180),
.A2(n_172),
.B1(n_55),
.B2(n_94),
.Y(n_183)
);

AO22x1_ASAP7_75t_L g184 ( 
.A1(n_181),
.A2(n_179),
.B1(n_177),
.B2(n_172),
.Y(n_184)
);

AOI221xp5_ASAP7_75t_L g185 ( 
.A1(n_184),
.A2(n_55),
.B1(n_182),
.B2(n_183),
.C(n_161),
.Y(n_185)
);


endmodule