module fake_jpeg_31364_n_182 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_182);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_182;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_175;
wire n_57;
wire n_171;
wire n_119;
wire n_69;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_11),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_3),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_6),
.Y(n_56)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_13),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

HB1xp67_ASAP7_75t_L g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_3),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_29),
.B(n_0),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_6),
.Y(n_63)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_16),
.Y(n_64)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_5),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_50),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_1),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_8),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_24),
.Y(n_70)
);

BUFx4f_ASAP7_75t_L g71 ( 
.A(n_43),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_9),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_SL g75 ( 
.A(n_32),
.B(n_10),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_11),
.B(n_47),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_51),
.Y(n_78)
);

INVx6_ASAP7_75t_L g79 ( 
.A(n_33),
.Y(n_79)
);

INVx6_ASAP7_75t_L g80 ( 
.A(n_71),
.Y(n_80)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_80),
.Y(n_92)
);

BUFx12_ASAP7_75t_L g81 ( 
.A(n_71),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_81),
.B(n_82),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_73),
.B(n_0),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_75),
.B(n_1),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_88),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx4_ASAP7_75t_L g97 ( 
.A(n_84),
.Y(n_97)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

INVx4_ASAP7_75t_L g100 ( 
.A(n_85),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_86),
.B(n_87),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_27),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g88 ( 
.A(n_62),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g90 ( 
.A1(n_80),
.A2(n_53),
.B1(n_76),
.B2(n_68),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g119 ( 
.A1(n_90),
.A2(n_54),
.B1(n_70),
.B2(n_78),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_87),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_91),
.B(n_95),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_85),
.B(n_66),
.C(n_60),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_93),
.B(n_57),
.Y(n_113)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_81),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_86),
.B(n_75),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_98),
.B(n_99),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_53),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_81),
.B(n_61),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_102),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_88),
.B(n_55),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_88),
.B(n_69),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_74),
.Y(n_114)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_100),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_105),
.Y(n_124)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_100),
.Y(n_106)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_106),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g108 ( 
.A(n_92),
.Y(n_108)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_108),
.Y(n_133)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_92),
.Y(n_109)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_109),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_97),
.A2(n_76),
.B1(n_59),
.B2(n_56),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_110),
.A2(n_111),
.B1(n_121),
.B2(n_77),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_90),
.A2(n_63),
.B1(n_60),
.B2(n_64),
.Y(n_111)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_2),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_114),
.B(n_117),
.Y(n_136)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_99),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_115),
.B(n_116),
.Y(n_143)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g117 ( 
.A(n_89),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_96),
.B(n_62),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_118),
.B(n_120),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_119),
.A2(n_2),
.B1(n_4),
.B2(n_7),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_93),
.B(n_77),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g121 ( 
.A1(n_97),
.A2(n_58),
.B1(n_4),
.B2(n_5),
.Y(n_121)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_100),
.Y(n_122)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_101),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_123),
.B(n_7),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_108),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_125),
.B(n_128),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_SL g145 ( 
.A1(n_126),
.A2(n_19),
.B(n_20),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_127),
.A2(n_144),
.B1(n_22),
.B2(n_23),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_104),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_122),
.Y(n_129)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_129),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_110),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g134 ( 
.A(n_112),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_138),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g135 ( 
.A(n_121),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_135),
.B(n_140),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g152 ( 
.A(n_137),
.B(n_141),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_107),
.B(n_9),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_113),
.B(n_12),
.Y(n_141)
);

NOR2x1_ASAP7_75t_L g142 ( 
.A(n_111),
.B(n_14),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_142),
.B(n_34),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_117),
.A2(n_15),
.B1(n_17),
.B2(n_18),
.Y(n_144)
);

AOI21xp5_ASAP7_75t_L g166 ( 
.A1(n_145),
.A2(n_154),
.B(n_48),
.Y(n_166)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_139),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_146),
.B(n_149),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g149 ( 
.A(n_133),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_155),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g151 ( 
.A1(n_130),
.A2(n_25),
.B(n_30),
.C(n_31),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_SL g165 ( 
.A1(n_151),
.A2(n_154),
.B(n_159),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_SL g155 ( 
.A(n_143),
.B(n_52),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_136),
.B(n_35),
.Y(n_156)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_156),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g158 ( 
.A(n_137),
.B(n_36),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_158),
.B(n_160),
.C(n_132),
.Y(n_164)
);

AO22x1_ASAP7_75t_L g159 ( 
.A1(n_135),
.A2(n_37),
.B1(n_38),
.B2(n_39),
.Y(n_159)
);

OAI21xp33_ASAP7_75t_L g168 ( 
.A1(n_159),
.A2(n_157),
.B(n_142),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_124),
.B(n_42),
.C(n_44),
.Y(n_160)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_152),
.B(n_147),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_162),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_164),
.B(n_165),
.Y(n_170)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_166),
.Y(n_172)
);

INVx1_ASAP7_75t_SL g171 ( 
.A(n_168),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_170),
.B(n_162),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_SL g175 ( 
.A1(n_173),
.A2(n_174),
.B(n_169),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_171),
.A2(n_127),
.B1(n_168),
.B2(n_163),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_SL g176 ( 
.A(n_175),
.B(n_172),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_176),
.A2(n_167),
.B1(n_151),
.B2(n_153),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_177),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_178),
.B(n_149),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_179),
.A2(n_131),
.B(n_49),
.Y(n_180)
);

OAI21xp5_ASAP7_75t_L g181 ( 
.A1(n_180),
.A2(n_45),
.B(n_148),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_181),
.B(n_148),
.Y(n_182)
);


endmodule