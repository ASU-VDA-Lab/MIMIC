module fake_jpeg_8982_n_104 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_104);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_104;

wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_49;
wire n_76;
wire n_88;
wire n_74;
wire n_103;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_93;
wire n_91;
wire n_101;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_62;
wire n_100;
wire n_82;
wire n_96;

INVx8_ASAP7_75t_L g44 ( 
.A(n_32),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_37),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_27),
.Y(n_47)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_38),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_35),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_33),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_30),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_3),
.Y(n_54)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_22),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

INVx8_ASAP7_75t_SL g57 ( 
.A(n_1),
.Y(n_57)
);

BUFx4f_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx2_ASAP7_75t_L g59 ( 
.A(n_10),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_28),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_8),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_15),
.Y(n_63)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_57),
.Y(n_64)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_65),
.Y(n_85)
);

AOI21xp33_ASAP7_75t_L g66 ( 
.A1(n_55),
.A2(n_0),
.B(n_1),
.Y(n_66)
);

NAND3xp33_ASAP7_75t_L g78 ( 
.A(n_66),
.B(n_74),
.C(n_0),
.Y(n_78)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_48),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_67),
.Y(n_76)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_68),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_60),
.Y(n_69)
);

AND2x4_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_2),
.Y(n_82)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_54),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_70),
.Y(n_84)
);

INVx4_ASAP7_75t_SL g71 ( 
.A(n_61),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_71),
.A2(n_50),
.B1(n_52),
.B2(n_63),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI21xp33_ASAP7_75t_SL g79 ( 
.A1(n_72),
.A2(n_73),
.B(n_25),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_56),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_SL g75 ( 
.A1(n_71),
.A2(n_44),
.B1(n_56),
.B2(n_60),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_75),
.B(n_78),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g90 ( 
.A1(n_79),
.A2(n_80),
.B1(n_46),
.B2(n_45),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_69),
.A2(n_49),
.B1(n_62),
.B2(n_47),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_81),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g87 ( 
.A(n_82),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_88),
.Y(n_91)
);

BUFx12f_ASAP7_75t_L g88 ( 
.A(n_83),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_82),
.B1(n_85),
.B2(n_84),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_92),
.A2(n_86),
.B1(n_82),
.B2(n_89),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g94 ( 
.A(n_93),
.B(n_91),
.Y(n_94)
);

XOR2xp5_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_77),
.Y(n_95)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_95),
.A2(n_76),
.B(n_88),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_96),
.B(n_4),
.C(n_5),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_6),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_98),
.B(n_7),
.C(n_12),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_99),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_100)
);

AOI22x1_ASAP7_75t_L g101 ( 
.A1(n_100),
.A2(n_18),
.B1(n_19),
.B2(n_20),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g102 ( 
.A1(n_101),
.A2(n_21),
.A3(n_23),
.B1(n_24),
.B2(n_29),
.C1(n_31),
.C2(n_34),
.Y(n_102)
);

AOI21xp5_ASAP7_75t_SL g103 ( 
.A1(n_102),
.A2(n_43),
.B(n_39),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_41),
.Y(n_104)
);


endmodule