module fake_jpeg_26586_n_247 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_247);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_247;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_96;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_11),
.Y(n_17)
);

INVx6_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_15),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_16),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx5_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_0),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_19),
.Y(n_35)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_36),
.Y(n_60)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_17),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_38),
.B(n_39),
.Y(n_58)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_40),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_41),
.B(n_42),
.Y(n_62)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx3_ASAP7_75t_L g43 ( 
.A(n_19),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_43),
.Y(n_48)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_21),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_45),
.Y(n_63)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_19),
.Y(n_45)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_27),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_42),
.A2(n_18),
.B1(n_34),
.B2(n_22),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_49),
.A2(n_51),
.B1(n_26),
.B2(n_23),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_50),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_27),
.C(n_30),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_52),
.B(n_61),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_36),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_55),
.B(n_59),
.Y(n_74)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_45),
.A2(n_18),
.B1(n_43),
.B2(n_46),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_67),
.B1(n_22),
.B2(n_26),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_43),
.A2(n_18),
.B1(n_27),
.B2(n_29),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_57),
.A2(n_22),
.B1(n_26),
.B2(n_30),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_25),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_44),
.B(n_27),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_36),
.B(n_29),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_40),
.B(n_21),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_46),
.A2(n_18),
.B1(n_25),
.B2(n_24),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_37),
.A2(n_24),
.B1(n_25),
.B2(n_30),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_68),
.A2(n_33),
.B1(n_28),
.B2(n_31),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_23),
.Y(n_69)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_69),
.A2(n_33),
.B(n_28),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_70),
.B(n_75),
.Y(n_114)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_71),
.Y(n_95)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_47),
.Y(n_76)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_76),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_50),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_77),
.Y(n_104)
);

NAND2xp33_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_28),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_SL g99 ( 
.A(n_78),
.B(n_52),
.Y(n_99)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx3_ASAP7_75t_L g115 ( 
.A(n_79),
.Y(n_115)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_62),
.Y(n_80)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_80),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_81),
.A2(n_84),
.B1(n_51),
.B2(n_69),
.Y(n_100)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_47),
.Y(n_82)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_82),
.Y(n_105)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_47),
.Y(n_85)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_85),
.Y(n_108)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_86),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_87),
.B(n_91),
.Y(n_94)
);

AO22x2_ASAP7_75t_SL g88 ( 
.A1(n_57),
.A2(n_40),
.B1(n_41),
.B2(n_33),
.Y(n_88)
);

O2A1O1Ixp33_ASAP7_75t_SL g97 ( 
.A1(n_88),
.A2(n_63),
.B(n_49),
.C(n_54),
.Y(n_97)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_48),
.Y(n_89)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_89),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_58),
.B(n_32),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g102 ( 
.A(n_90),
.B(n_69),
.Y(n_102)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_63),
.Y(n_92)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_92),
.Y(n_118)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_55),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_97),
.A2(n_103),
.B1(n_88),
.B2(n_84),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_77),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_79),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_100),
.A2(n_106),
.B1(n_88),
.B2(n_80),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_102),
.B(n_74),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_93),
.A2(n_53),
.B1(n_64),
.B2(n_60),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g107 ( 
.A(n_73),
.B(n_54),
.C(n_48),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_107),
.B(n_116),
.C(n_72),
.Y(n_121)
);

OAI32xp33_ASAP7_75t_L g109 ( 
.A1(n_73),
.A2(n_58),
.A3(n_65),
.B1(n_66),
.B2(n_60),
.Y(n_109)
);

OAI32xp33_ASAP7_75t_L g140 ( 
.A1(n_109),
.A2(n_31),
.A3(n_20),
.B1(n_89),
.B2(n_86),
.Y(n_140)
);

BUFx24_ASAP7_75t_SL g111 ( 
.A(n_70),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_111),
.B(n_31),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_92),
.B(n_54),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_117),
.Y(n_127)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_75),
.B(n_64),
.C(n_32),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_83),
.B(n_32),
.Y(n_117)
);

MAJx2_ASAP7_75t_L g119 ( 
.A(n_107),
.B(n_78),
.C(n_87),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_119),
.B(n_135),
.C(n_101),
.Y(n_143)
);

BUFx5_ASAP7_75t_L g120 ( 
.A(n_115),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_130),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_121),
.B(n_136),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_122),
.A2(n_94),
.B1(n_97),
.B2(n_95),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g124 ( 
.A(n_98),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_113),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_125),
.B(n_129),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_126),
.B(n_139),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g149 ( 
.A1(n_128),
.A2(n_133),
.B1(n_130),
.B2(n_137),
.Y(n_149)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_100),
.Y(n_130)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_103),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_131),
.B(n_137),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_104),
.Y(n_132)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_132),
.Y(n_146)
);

NOR2x1_ASAP7_75t_L g133 ( 
.A(n_109),
.B(n_88),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_99),
.B(n_83),
.C(n_72),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_116),
.Y(n_137)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_117),
.Y(n_138)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_138),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_L g160 ( 
.A1(n_140),
.A2(n_105),
.B(n_110),
.Y(n_160)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_141),
.Y(n_145)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_143),
.B(n_148),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g178 ( 
.A1(n_147),
.A2(n_156),
.B1(n_76),
.B2(n_115),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g171 ( 
.A1(n_149),
.A2(n_160),
.B1(n_110),
.B2(n_82),
.Y(n_171)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_122),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_151),
.B(n_152),
.Y(n_166)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_127),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_123),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_153),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_136),
.B(n_101),
.C(n_118),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_154),
.B(n_157),
.C(n_20),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_129),
.A2(n_97),
.B1(n_95),
.B2(n_94),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_121),
.B(n_118),
.C(n_96),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_128),
.A2(n_96),
.B1(n_112),
.B2(n_105),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_159),
.A2(n_131),
.B1(n_138),
.B2(n_140),
.Y(n_169)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_127),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_161),
.B(n_163),
.Y(n_174)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_150),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_165),
.B(n_168),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_SL g167 ( 
.A(n_164),
.B(n_119),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_167),
.B(n_170),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_159),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_169),
.A2(n_171),
.B1(n_172),
.B2(n_156),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_148),
.B(n_135),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_149),
.A2(n_108),
.B1(n_76),
.B2(n_85),
.Y(n_172)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_145),
.Y(n_173)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_173),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_151),
.A2(n_108),
.B(n_120),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_175),
.A2(n_176),
.B(n_181),
.Y(n_193)
);

OAI21xp5_ASAP7_75t_L g176 ( 
.A1(n_160),
.A2(n_1),
.B(n_2),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_177),
.B(n_180),
.C(n_157),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_178),
.A2(n_179),
.B1(n_142),
.B2(n_144),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_147),
.A2(n_20),
.B1(n_15),
.B2(n_14),
.Y(n_179)
);

XOR2x2_ASAP7_75t_SL g181 ( 
.A(n_143),
.B(n_1),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g182 ( 
.A(n_155),
.Y(n_182)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_182),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g184 ( 
.A1(n_153),
.A2(n_1),
.B(n_2),
.Y(n_184)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_184),
.A2(n_176),
.B(n_4),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_185),
.B(n_186),
.Y(n_209)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_167),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_187),
.B(n_200),
.C(n_180),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_188),
.A2(n_191),
.B1(n_163),
.B2(n_145),
.Y(n_212)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_174),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_189),
.B(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_166),
.B(n_152),
.Y(n_190)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_190),
.Y(n_207)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_194),
.Y(n_211)
);

AOI21xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_162),
.B(n_146),
.Y(n_195)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_195),
.A2(n_142),
.B(n_173),
.C(n_184),
.Y(n_210)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_172),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_177),
.B(n_154),
.C(n_162),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_175),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_201),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_202),
.B(n_205),
.C(n_214),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_192),
.B(n_158),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_203),
.B(n_213),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g205 ( 
.A(n_187),
.B(n_170),
.C(n_161),
.Y(n_205)
);

OAI21x1_ASAP7_75t_L g206 ( 
.A1(n_197),
.A2(n_181),
.B(n_179),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_206),
.A2(n_193),
.B(n_190),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_200),
.B(n_169),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g223 ( 
.A(n_208),
.B(n_3),
.Y(n_223)
);

A2O1A1Ixp33_ASAP7_75t_SL g218 ( 
.A1(n_210),
.A2(n_195),
.B(n_191),
.C(n_193),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_212),
.A2(n_198),
.B1(n_201),
.B2(n_196),
.Y(n_217)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_199),
.B(n_13),
.C(n_5),
.Y(n_214)
);

BUFx24_ASAP7_75t_SL g215 ( 
.A(n_209),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_215),
.B(n_220),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_207),
.B(n_192),
.Y(n_216)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_216),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g225 ( 
.A1(n_217),
.A2(n_219),
.B1(n_210),
.B2(n_214),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_218),
.A2(n_210),
.B(n_6),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_211),
.A2(n_188),
.B1(n_186),
.B2(n_199),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_204),
.A2(n_186),
.B1(n_13),
.B2(n_6),
.Y(n_222)
);

AND2x2_ASAP7_75t_L g231 ( 
.A(n_222),
.B(n_5),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_223),
.B(n_205),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_225),
.B(n_226),
.Y(n_234)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_229),
.B(n_12),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g235 ( 
.A1(n_230),
.A2(n_12),
.B1(n_7),
.B2(n_8),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_231),
.A2(n_224),
.B(n_218),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_232),
.B(n_233),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_221),
.C(n_218),
.Y(n_233)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_235),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g239 ( 
.A(n_236),
.B(n_237),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_227),
.B(n_6),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_234),
.B(n_230),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_241),
.B(n_233),
.C(n_231),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_242),
.Y(n_245)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_238),
.Y(n_243)
);

OAI321xp33_ASAP7_75t_L g244 ( 
.A1(n_243),
.A2(n_240),
.A3(n_239),
.B1(n_11),
.B2(n_10),
.C(n_9),
.Y(n_244)
);

OAI21xp5_ASAP7_75t_SL g246 ( 
.A1(n_244),
.A2(n_9),
.B(n_10),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_246),
.B(n_245),
.Y(n_247)
);


endmodule