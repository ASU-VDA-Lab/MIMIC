module fake_jpeg_21410_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_121;
wire n_99;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_49),
.Y(n_50)
);

INVxp67_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_25),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_27),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_44),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

BUFx12_ASAP7_75t_L g58 ( 
.A(n_23),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_14),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_18),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_46),
.Y(n_61)
);

INVx1_ASAP7_75t_SL g62 ( 
.A(n_6),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_SL g64 ( 
.A(n_35),
.B(n_32),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_48),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_24),
.B(n_47),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_20),
.Y(n_69)
);

INVx4_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_9),
.Y(n_71)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_12),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_2),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_36),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_15),
.Y(n_75)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_16),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_11),
.Y(n_78)
);

BUFx24_ASAP7_75t_L g79 ( 
.A(n_10),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_55),
.Y(n_80)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_80),
.Y(n_95)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_76),
.Y(n_81)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_81),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_82),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_59),
.Y(n_83)
);

INVx1_ASAP7_75t_SL g92 ( 
.A(n_83),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_79),
.Y(n_84)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_84),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_65),
.B(n_0),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_85),
.B(n_1),
.Y(n_91)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_76),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_86),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_62),
.B(n_0),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_87),
.B(n_58),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_90),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_81),
.B(n_72),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_91),
.B(n_1),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_80),
.A2(n_66),
.B1(n_70),
.B2(n_79),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_93),
.A2(n_51),
.B1(n_66),
.B2(n_58),
.Y(n_103)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_82),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g112 ( 
.A(n_97),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g100 ( 
.A(n_89),
.B(n_50),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_100),
.B(n_105),
.Y(n_122)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_94),
.Y(n_101)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_101),
.Y(n_119)
);

AOI21xp5_ASAP7_75t_L g102 ( 
.A1(n_92),
.A2(n_51),
.B(n_76),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_102),
.A2(n_63),
.B(n_61),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_103),
.A2(n_56),
.B1(n_3),
.B2(n_4),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_95),
.B(n_83),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_104),
.B(n_75),
.Y(n_116)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_98),
.Y(n_105)
);

INVx11_ASAP7_75t_L g106 ( 
.A(n_96),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g129 ( 
.A(n_106),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_107),
.B(n_2),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_94),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_108),
.B(n_110),
.Y(n_128)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_95),
.A2(n_71),
.B1(n_73),
.B2(n_59),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_109),
.A2(n_111),
.B1(n_74),
.B2(n_67),
.Y(n_124)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_97),
.A2(n_71),
.B1(n_73),
.B2(n_78),
.Y(n_111)
);

CKINVDCx20_ASAP7_75t_R g113 ( 
.A(n_100),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_113),
.B(n_114),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_102),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_92),
.B1(n_93),
.B2(n_77),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_118),
.B1(n_120),
.B2(n_60),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_116),
.B(n_125),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_117),
.A2(n_121),
.B(n_64),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_L g118 ( 
.A1(n_99),
.A2(n_53),
.B1(n_69),
.B2(n_54),
.Y(n_118)
);

AND2x2_ASAP7_75t_L g121 ( 
.A(n_103),
.B(n_68),
.Y(n_121)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_123),
.B(n_124),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_112),
.B(n_68),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_126),
.B(n_127),
.Y(n_140)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_110),
.Y(n_127)
);

NAND3xp33_ASAP7_75t_L g148 ( 
.A(n_131),
.B(n_4),
.C(n_5),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_132),
.A2(n_136),
.B1(n_123),
.B2(n_5),
.Y(n_146)
);

BUFx24_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_133),
.Y(n_143)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_135),
.B(n_137),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_114),
.A2(n_57),
.B1(n_52),
.B2(n_106),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_119),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_139),
.B(n_141),
.Y(n_144)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_115),
.Y(n_141)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_3),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_6),
.C(n_7),
.Y(n_149)
);

MAJx2_ASAP7_75t_L g145 ( 
.A(n_134),
.B(n_142),
.C(n_117),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_148),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_146),
.A2(n_130),
.B1(n_138),
.B2(n_140),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_149),
.A2(n_140),
.B1(n_8),
.B2(n_9),
.Y(n_151)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_153),
.B(n_147),
.Y(n_154)
);

BUFx24_ASAP7_75t_SL g155 ( 
.A(n_154),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_143),
.C(n_147),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_144),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_157),
.B(n_144),
.Y(n_158)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_158),
.A2(n_150),
.B(n_130),
.Y(n_159)
);

AOI21xp5_ASAP7_75t_L g160 ( 
.A1(n_159),
.A2(n_150),
.B(n_33),
.Y(n_160)
);

OAI311xp33_ASAP7_75t_L g161 ( 
.A1(n_160),
.A2(n_133),
.A3(n_31),
.B1(n_34),
.C1(n_17),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_28),
.A3(n_43),
.B1(n_39),
.B2(n_19),
.C1(n_22),
.C2(n_26),
.Y(n_162)
);

OAI321xp33_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_37),
.A3(n_38),
.B1(n_45),
.B2(n_7),
.C(n_11),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_163),
.B(n_12),
.Y(n_164)
);


endmodule