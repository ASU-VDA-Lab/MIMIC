module fake_netlist_1_8606_n_728 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_80, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_728);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_80;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_728;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_724;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_141;
wire n_119;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g81 ( .A(n_41), .Y(n_81) );
BUFx3_ASAP7_75t_L g82 ( .A(n_42), .Y(n_82) );
BUFx6f_ASAP7_75t_L g83 ( .A(n_2), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_69), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_70), .Y(n_85) );
CKINVDCx16_ASAP7_75t_R g86 ( .A(n_64), .Y(n_86) );
BUFx3_ASAP7_75t_L g87 ( .A(n_9), .Y(n_87) );
INVx1_ASAP7_75t_L g88 ( .A(n_17), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_48), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_74), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_66), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_67), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_44), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_19), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_28), .Y(n_95) );
HB1xp67_ASAP7_75t_L g96 ( .A(n_63), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_0), .Y(n_97) );
INVx2_ASAP7_75t_L g98 ( .A(n_78), .Y(n_98) );
INVx1_ASAP7_75t_L g99 ( .A(n_40), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_0), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_11), .Y(n_101) );
INVx1_ASAP7_75t_L g102 ( .A(n_14), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_50), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_4), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_18), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_25), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_1), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_23), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_24), .Y(n_109) );
INVxp67_ASAP7_75t_SL g110 ( .A(n_16), .Y(n_110) );
INVxp33_ASAP7_75t_L g111 ( .A(n_57), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_11), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_8), .Y(n_113) );
BUFx3_ASAP7_75t_L g114 ( .A(n_54), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_29), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_35), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_61), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_73), .Y(n_118) );
INVxp67_ASAP7_75t_SL g119 ( .A(n_51), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_9), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_45), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_59), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_37), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_22), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_4), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_15), .Y(n_126) );
INVx2_ASAP7_75t_L g127 ( .A(n_68), .Y(n_127) );
INVx1_ASAP7_75t_SL g128 ( .A(n_49), .Y(n_128) );
INVxp67_ASAP7_75t_SL g129 ( .A(n_15), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_81), .Y(n_130) );
OR2x2_ASAP7_75t_L g131 ( .A(n_100), .B(n_1), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_81), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_96), .B(n_2), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx2_ASAP7_75t_L g135 ( .A(n_98), .Y(n_135) );
INVx2_ASAP7_75t_L g136 ( .A(n_98), .Y(n_136) );
CKINVDCx5p33_ASAP7_75t_R g137 ( .A(n_86), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_84), .Y(n_138) );
NAND2xp5_ASAP7_75t_L g139 ( .A(n_104), .B(n_3), .Y(n_139) );
BUFx8_ASAP7_75t_L g140 ( .A(n_127), .Y(n_140) );
INVx2_ASAP7_75t_L g141 ( .A(n_127), .Y(n_141) );
NOR2x1_ASAP7_75t_L g142 ( .A(n_87), .B(n_3), .Y(n_142) );
INVx5_ASAP7_75t_L g143 ( .A(n_82), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_85), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_85), .Y(n_145) );
HB1xp67_ASAP7_75t_L g146 ( .A(n_87), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_88), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_88), .Y(n_148) );
HB1xp67_ASAP7_75t_L g149 ( .A(n_100), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_89), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_89), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_91), .Y(n_152) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_107), .B(n_5), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_112), .B(n_5), .Y(n_154) );
NAND3xp33_ASAP7_75t_L g155 ( .A(n_101), .B(n_39), .C(n_79), .Y(n_155) );
INVx1_ASAP7_75t_L g156 ( .A(n_91), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_92), .Y(n_157) );
OAI22xp33_ASAP7_75t_L g158 ( .A1(n_101), .A2(n_6), .B1(n_7), .B2(n_8), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_92), .Y(n_159) );
AND2x2_ASAP7_75t_L g160 ( .A(n_111), .B(n_6), .Y(n_160) );
INVx2_ASAP7_75t_L g161 ( .A(n_93), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_93), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_113), .B(n_7), .Y(n_163) );
INVx3_ASAP7_75t_L g164 ( .A(n_83), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_94), .Y(n_165) );
AND2x4_ASAP7_75t_L g166 ( .A(n_102), .B(n_10), .Y(n_166) );
INVx3_ASAP7_75t_L g167 ( .A(n_83), .Y(n_167) );
OAI21x1_ASAP7_75t_L g168 ( .A1(n_94), .A2(n_43), .B(n_77), .Y(n_168) );
INVx2_ASAP7_75t_L g169 ( .A(n_99), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_99), .Y(n_170) );
NAND2xp33_ASAP7_75t_SL g171 ( .A(n_90), .B(n_10), .Y(n_171) );
AND2x2_ASAP7_75t_L g172 ( .A(n_102), .B(n_12), .Y(n_172) );
INVx2_ASAP7_75t_L g173 ( .A(n_103), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_120), .B(n_12), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_146), .B(n_106), .Y(n_175) );
NAND2x1p5_ASAP7_75t_L g176 ( .A(n_166), .B(n_122), .Y(n_176) );
INVx2_ASAP7_75t_L g177 ( .A(n_164), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_166), .Y(n_178) );
AOI22xp5_ASAP7_75t_L g179 ( .A1(n_160), .A2(n_126), .B1(n_125), .B2(n_129), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_149), .B(n_125), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_137), .B(n_105), .Y(n_182) );
BUFx6f_ASAP7_75t_L g183 ( .A(n_168), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_164), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_168), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_166), .Y(n_186) );
AND2x4_ASAP7_75t_L g187 ( .A(n_130), .B(n_126), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_164), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_130), .B(n_109), .Y(n_189) );
INVx2_ASAP7_75t_SL g190 ( .A(n_140), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_132), .B(n_90), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_164), .Y(n_192) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_167), .Y(n_193) );
CKINVDCx20_ASAP7_75t_R g194 ( .A(n_160), .Y(n_194) );
NAND2x1p5_ASAP7_75t_L g195 ( .A(n_172), .B(n_108), .Y(n_195) );
INVx2_ASAP7_75t_L g196 ( .A(n_167), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_132), .B(n_95), .Y(n_197) );
AND2x4_ASAP7_75t_L g198 ( .A(n_134), .B(n_124), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_134), .B(n_95), .Y(n_199) );
INVx4_ASAP7_75t_L g200 ( .A(n_143), .Y(n_200) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_138), .B(n_123), .Y(n_201) );
INVx1_ASAP7_75t_L g202 ( .A(n_172), .Y(n_202) );
AND2x2_ASAP7_75t_L g203 ( .A(n_138), .B(n_123), .Y(n_203) );
INVx1_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
NAND2x1p5_ASAP7_75t_L g205 ( .A(n_147), .B(n_103), .Y(n_205) );
INVx3_ASAP7_75t_L g206 ( .A(n_135), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_147), .B(n_106), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_167), .Y(n_208) );
INVx2_ASAP7_75t_L g209 ( .A(n_167), .Y(n_209) );
CKINVDCx20_ASAP7_75t_R g210 ( .A(n_171), .Y(n_210) );
BUFx6f_ASAP7_75t_L g211 ( .A(n_145), .Y(n_211) );
BUFx6f_ASAP7_75t_L g212 ( .A(n_145), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_148), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_148), .Y(n_214) );
INVx4_ASAP7_75t_L g215 ( .A(n_143), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_150), .B(n_116), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_148), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_152), .Y(n_218) );
AND2x2_ASAP7_75t_L g219 ( .A(n_150), .B(n_97), .Y(n_219) );
AND2x4_ASAP7_75t_L g220 ( .A(n_156), .B(n_124), .Y(n_220) );
AND2x4_ASAP7_75t_L g221 ( .A(n_156), .B(n_122), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_152), .Y(n_222) );
INVx1_ASAP7_75t_L g223 ( .A(n_152), .Y(n_223) );
INVx2_ASAP7_75t_SL g224 ( .A(n_140), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_173), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_140), .B(n_115), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_173), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_157), .B(n_118), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_173), .Y(n_229) );
INVx8_ASAP7_75t_L g230 ( .A(n_143), .Y(n_230) );
INVx4_ASAP7_75t_SL g231 ( .A(n_157), .Y(n_231) );
INVx2_ASAP7_75t_L g232 ( .A(n_135), .Y(n_232) );
NAND2xp5_ASAP7_75t_L g233 ( .A(n_159), .B(n_121), .Y(n_233) );
NAND2xp5_ASAP7_75t_SL g234 ( .A(n_140), .B(n_108), .Y(n_234) );
AND2x4_ASAP7_75t_L g235 ( .A(n_159), .B(n_110), .Y(n_235) );
INVx2_ASAP7_75t_L g236 ( .A(n_136), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_136), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_211), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
INVx1_ASAP7_75t_L g240 ( .A(n_205), .Y(n_240) );
AND2x4_ASAP7_75t_L g241 ( .A(n_203), .B(n_131), .Y(n_241) );
INVx1_ASAP7_75t_SL g242 ( .A(n_203), .Y(n_242) );
HB1xp67_ASAP7_75t_L g243 ( .A(n_207), .Y(n_243) );
NOR2xp33_ASAP7_75t_SL g244 ( .A(n_190), .B(n_158), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_175), .B(n_133), .Y(n_245) );
BUFx6f_ASAP7_75t_L g246 ( .A(n_190), .Y(n_246) );
AND2x4_ASAP7_75t_L g247 ( .A(n_207), .B(n_131), .Y(n_247) );
BUFx6f_ASAP7_75t_L g248 ( .A(n_224), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g249 ( .A(n_191), .B(n_165), .Y(n_249) );
INVx3_ASAP7_75t_L g250 ( .A(n_186), .Y(n_250) );
NOR2xp33_ASAP7_75t_L g251 ( .A(n_202), .B(n_170), .Y(n_251) );
INVx5_ASAP7_75t_L g252 ( .A(n_230), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g253 ( .A(n_197), .B(n_165), .Y(n_253) );
BUFx4f_ASAP7_75t_L g254 ( .A(n_176), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_204), .Y(n_255) );
BUFx4f_ASAP7_75t_L g256 ( .A(n_176), .Y(n_256) );
BUFx2_ASAP7_75t_L g257 ( .A(n_194), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_194), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_205), .Y(n_259) );
BUFx3_ASAP7_75t_L g260 ( .A(n_224), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_204), .Y(n_261) );
INVx1_ASAP7_75t_L g262 ( .A(n_213), .Y(n_262) );
NAND2xp5_ASAP7_75t_SL g263 ( .A(n_183), .B(n_170), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_213), .Y(n_264) );
AND2x2_ASAP7_75t_SL g265 ( .A(n_198), .B(n_174), .Y(n_265) );
INVx3_ASAP7_75t_L g266 ( .A(n_186), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g267 ( .A(n_199), .B(n_169), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_187), .Y(n_268) );
INVx2_ASAP7_75t_L g269 ( .A(n_211), .Y(n_269) );
HB1xp67_ASAP7_75t_L g270 ( .A(n_195), .Y(n_270) );
INVx2_ASAP7_75t_L g271 ( .A(n_211), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_187), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_201), .B(n_169), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_235), .B(n_142), .Y(n_274) );
CKINVDCx5p33_ASAP7_75t_R g275 ( .A(n_210), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_187), .Y(n_276) );
INVx2_ASAP7_75t_L g277 ( .A(n_211), .Y(n_277) );
BUFx3_ASAP7_75t_L g278 ( .A(n_230), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_195), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_195), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g281 ( .A1(n_235), .A2(n_142), .B1(n_163), .B2(n_139), .Y(n_281) );
BUFx3_ASAP7_75t_L g282 ( .A(n_230), .Y(n_282) );
INVx2_ASAP7_75t_L g283 ( .A(n_211), .Y(n_283) );
AND2x2_ASAP7_75t_L g284 ( .A(n_235), .B(n_162), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_198), .B(n_162), .Y(n_285) );
NAND2xp5_ASAP7_75t_SL g286 ( .A(n_183), .B(n_155), .Y(n_286) );
NAND2xp5_ASAP7_75t_L g287 ( .A(n_198), .B(n_161), .Y(n_287) );
AO21x2_ASAP7_75t_L g288 ( .A1(n_234), .A2(n_155), .B(n_153), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_220), .A2(n_154), .B1(n_161), .B2(n_151), .Y(n_289) );
AND2x2_ASAP7_75t_L g290 ( .A(n_219), .B(n_144), .Y(n_290) );
HB1xp67_ASAP7_75t_L g291 ( .A(n_180), .Y(n_291) );
INVx1_ASAP7_75t_L g292 ( .A(n_206), .Y(n_292) );
NAND2xp5_ASAP7_75t_L g293 ( .A(n_220), .B(n_221), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_183), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_206), .Y(n_295) );
O2A1O1Ixp33_ASAP7_75t_L g296 ( .A1(n_180), .A2(n_151), .B(n_144), .C(n_141), .Y(n_296) );
INVx2_ASAP7_75t_SL g297 ( .A(n_176), .Y(n_297) );
AOI22xp33_ASAP7_75t_SL g298 ( .A1(n_210), .A2(n_83), .B1(n_117), .B2(n_119), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_220), .B(n_221), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_221), .B(n_141), .Y(n_300) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_219), .B(n_143), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_206), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_186), .B(n_143), .Y(n_303) );
BUFx6f_ASAP7_75t_SL g304 ( .A(n_178), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_181), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_232), .Y(n_306) );
OAI22xp5_ASAP7_75t_L g307 ( .A1(n_254), .A2(n_216), .B1(n_233), .B2(n_228), .Y(n_307) );
AOI21xp5_ASAP7_75t_L g308 ( .A1(n_263), .A2(n_226), .B(n_185), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_268), .Y(n_309) );
O2A1O1Ixp33_ASAP7_75t_L g310 ( .A1(n_243), .A2(n_189), .B(n_223), .C(n_225), .Y(n_310) );
INVxp67_ASAP7_75t_SL g311 ( .A(n_297), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_263), .A2(n_185), .B(n_183), .Y(n_312) );
INVx2_ASAP7_75t_SL g313 ( .A(n_254), .Y(n_313) );
INVx4_ASAP7_75t_L g314 ( .A(n_252), .Y(n_314) );
AND2x4_ASAP7_75t_L g315 ( .A(n_279), .B(n_179), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_280), .B(n_182), .Y(n_316) );
INVx4_ASAP7_75t_SL g317 ( .A(n_304), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_272), .Y(n_318) );
AND2x4_ASAP7_75t_L g319 ( .A(n_270), .B(n_231), .Y(n_319) );
AOI22xp33_ASAP7_75t_L g320 ( .A1(n_274), .A2(n_227), .B1(n_218), .B2(n_229), .Y(n_320) );
AOI22xp5_ASAP7_75t_L g321 ( .A1(n_293), .A2(n_222), .B1(n_214), .B2(n_217), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_254), .Y(n_322) );
AND2x4_ASAP7_75t_L g323 ( .A(n_241), .B(n_231), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_241), .B(n_222), .Y(n_324) );
NOR2x1_ASAP7_75t_L g325 ( .A(n_274), .B(n_237), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_252), .Y(n_326) );
INVx1_ASAP7_75t_L g327 ( .A(n_276), .Y(n_327) );
INVx2_ASAP7_75t_L g328 ( .A(n_250), .Y(n_328) );
INVx4_ASAP7_75t_SL g329 ( .A(n_304), .Y(n_329) );
INVx2_ASAP7_75t_L g330 ( .A(n_250), .Y(n_330) );
AND2x2_ASAP7_75t_SL g331 ( .A(n_256), .B(n_183), .Y(n_331) );
BUFx6f_ASAP7_75t_L g332 ( .A(n_252), .Y(n_332) );
INVx5_ASAP7_75t_L g333 ( .A(n_252), .Y(n_333) );
OR2x6_ASAP7_75t_L g334 ( .A(n_297), .B(n_230), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_290), .Y(n_335) );
HB1xp67_ASAP7_75t_L g336 ( .A(n_242), .Y(n_336) );
INVx2_ASAP7_75t_L g337 ( .A(n_250), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_290), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_266), .Y(n_339) );
NAND2x1p5_ASAP7_75t_L g340 ( .A(n_256), .B(n_218), .Y(n_340) );
BUFx12f_ASAP7_75t_L g341 ( .A(n_275), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g342 ( .A1(n_299), .A2(n_217), .B1(n_214), .B2(n_229), .Y(n_342) );
INVx1_ASAP7_75t_L g343 ( .A(n_266), .Y(n_343) );
BUFx10_ASAP7_75t_L g344 ( .A(n_241), .Y(n_344) );
BUFx2_ASAP7_75t_R g345 ( .A(n_275), .Y(n_345) );
INVx3_ASAP7_75t_L g346 ( .A(n_252), .Y(n_346) );
OR2x6_ASAP7_75t_SL g347 ( .A(n_239), .B(n_240), .Y(n_347) );
NOR2xp33_ASAP7_75t_L g348 ( .A(n_291), .B(n_185), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_256), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_266), .Y(n_350) );
HB1xp67_ASAP7_75t_L g351 ( .A(n_257), .Y(n_351) );
INVx1_ASAP7_75t_L g352 ( .A(n_300), .Y(n_352) );
INVx1_ASAP7_75t_L g353 ( .A(n_284), .Y(n_353) );
AOI21xp33_ASAP7_75t_L g354 ( .A1(n_288), .A2(n_185), .B(n_236), .Y(n_354) );
HB1xp67_ASAP7_75t_L g355 ( .A(n_257), .Y(n_355) );
AND2x4_ASAP7_75t_L g356 ( .A(n_247), .B(n_231), .Y(n_356) );
AND2x4_ASAP7_75t_L g357 ( .A(n_247), .B(n_231), .Y(n_357) );
BUFx3_ASAP7_75t_L g358 ( .A(n_258), .Y(n_358) );
INVx2_ASAP7_75t_L g359 ( .A(n_255), .Y(n_359) );
OAI221xp5_ASAP7_75t_L g360 ( .A1(n_281), .A2(n_237), .B1(n_236), .B2(n_232), .C(n_128), .Y(n_360) );
INVx1_ASAP7_75t_SL g361 ( .A(n_259), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_359), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_333), .Y(n_363) );
INVx3_ASAP7_75t_SL g364 ( .A(n_333), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_361), .B(n_247), .Y(n_365) );
NAND2xp5_ASAP7_75t_SL g366 ( .A(n_333), .B(n_260), .Y(n_366) );
INVx1_ASAP7_75t_SL g367 ( .A(n_361), .Y(n_367) );
INVx2_ASAP7_75t_SL g368 ( .A(n_334), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_314), .Y(n_369) );
NAND2x1_ASAP7_75t_L g370 ( .A(n_314), .B(n_255), .Y(n_370) );
AOI222xp33_ASAP7_75t_L g371 ( .A1(n_335), .A2(n_258), .B1(n_274), .B2(n_244), .C1(n_251), .C2(n_284), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_322), .B(n_278), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_309), .Y(n_373) );
OAI222xp33_ASAP7_75t_L g374 ( .A1(n_307), .A2(n_298), .B1(n_289), .B2(n_253), .C1(n_249), .C2(n_287), .Y(n_374) );
CKINVDCx12_ASAP7_75t_R g375 ( .A(n_334), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_328), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_318), .Y(n_377) );
CKINVDCx5p33_ASAP7_75t_R g378 ( .A(n_341), .Y(n_378) );
CKINVDCx6p67_ASAP7_75t_R g379 ( .A(n_347), .Y(n_379) );
AND2x4_ASAP7_75t_L g380 ( .A(n_349), .B(n_278), .Y(n_380) );
O2A1O1Ixp33_ASAP7_75t_SL g381 ( .A1(n_354), .A2(n_286), .B(n_261), .C(n_262), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g382 ( .A(n_336), .B(n_265), .Y(n_382) );
AO21x2_ASAP7_75t_L g383 ( .A1(n_354), .A2(n_286), .B(n_288), .Y(n_383) );
AOI21xp5_ASAP7_75t_L g384 ( .A1(n_312), .A2(n_305), .B(n_260), .Y(n_384) );
INVx1_ASAP7_75t_L g385 ( .A(n_327), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_338), .B(n_265), .Y(n_386) );
INVx1_ASAP7_75t_L g387 ( .A(n_352), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_330), .Y(n_388) );
INVx4_ASAP7_75t_L g389 ( .A(n_326), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_324), .B(n_285), .Y(n_390) );
AND2x2_ASAP7_75t_L g391 ( .A(n_344), .B(n_264), .Y(n_391) );
AOI22xp33_ASAP7_75t_SL g392 ( .A1(n_358), .A2(n_304), .B1(n_245), .B2(n_246), .Y(n_392) );
INVx2_ASAP7_75t_L g393 ( .A(n_337), .Y(n_393) );
INVx3_ASAP7_75t_L g394 ( .A(n_326), .Y(n_394) );
NAND2xp5_ASAP7_75t_L g395 ( .A(n_315), .B(n_267), .Y(n_395) );
INVx1_ASAP7_75t_SL g396 ( .A(n_351), .Y(n_396) );
AOI22xp33_ASAP7_75t_L g397 ( .A1(n_371), .A2(n_307), .B1(n_360), .B2(n_355), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
OAI211xp5_ASAP7_75t_L g399 ( .A1(n_367), .A2(n_360), .B(n_310), .C(n_324), .Y(n_399) );
OAI221xp5_ASAP7_75t_L g400 ( .A1(n_395), .A2(n_353), .B1(n_320), .B2(n_296), .C(n_273), .Y(n_400) );
BUFx2_ASAP7_75t_SL g401 ( .A(n_363), .Y(n_401) );
AND2x2_ASAP7_75t_L g402 ( .A(n_387), .B(n_344), .Y(n_402) );
AOI22xp33_ASAP7_75t_L g403 ( .A1(n_379), .A2(n_315), .B1(n_316), .B2(n_348), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_362), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_379), .A2(n_316), .B1(n_325), .B2(n_331), .Y(n_405) );
BUFx3_ASAP7_75t_L g406 ( .A(n_364), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_375), .Y(n_407) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_387), .A2(n_83), .B1(n_288), .B2(n_350), .Y(n_408) );
BUFx2_ASAP7_75t_L g409 ( .A(n_364), .Y(n_409) );
BUFx12f_ASAP7_75t_L g410 ( .A(n_378), .Y(n_410) );
INVx2_ASAP7_75t_L g411 ( .A(n_376), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_373), .Y(n_412) );
AND2x2_ASAP7_75t_L g413 ( .A(n_390), .B(n_365), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_373), .Y(n_414) );
AOI22xp33_ASAP7_75t_SL g415 ( .A1(n_368), .A2(n_313), .B1(n_340), .B2(n_345), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_396), .A2(n_305), .B1(n_339), .B2(n_343), .Y(n_416) );
AOI22xp33_ASAP7_75t_L g417 ( .A1(n_377), .A2(n_83), .B1(n_342), .B2(n_321), .Y(n_417) );
BUFx2_ASAP7_75t_L g418 ( .A(n_364), .Y(n_418) );
AOI22xp33_ASAP7_75t_L g419 ( .A1(n_377), .A2(n_321), .B1(n_342), .B2(n_295), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_391), .A2(n_302), .B1(n_292), .B2(n_329), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_385), .B(n_311), .Y(n_421) );
BUFx2_ASAP7_75t_L g422 ( .A(n_389), .Y(n_422) );
OAI22xp5_ASAP7_75t_L g423 ( .A1(n_390), .A2(n_334), .B1(n_340), .B2(n_306), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_384), .A2(n_312), .B(n_308), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_385), .Y(n_426) );
HB1xp67_ASAP7_75t_L g427 ( .A(n_409), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_412), .B(n_386), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_404), .B(n_389), .Y(n_429) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_397), .A2(n_368), .B1(n_391), .B2(n_382), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g431 ( .A1(n_397), .A2(n_392), .B1(n_372), .B2(n_380), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_404), .B(n_389), .Y(n_432) );
AOI22xp5_ASAP7_75t_L g433 ( .A1(n_413), .A2(n_375), .B1(n_372), .B2(n_380), .Y(n_433) );
OAI21x1_ASAP7_75t_L g434 ( .A1(n_425), .A2(n_370), .B(n_308), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_404), .B(n_394), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_411), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_413), .B(n_388), .Y(n_437) );
OR2x2_ASAP7_75t_L g438 ( .A(n_413), .B(n_383), .Y(n_438) );
OAI211xp5_ASAP7_75t_L g439 ( .A1(n_415), .A2(n_378), .B(n_370), .C(n_363), .Y(n_439) );
AND2x4_ASAP7_75t_L g440 ( .A(n_412), .B(n_394), .Y(n_440) );
AOI33xp33_ASAP7_75t_L g441 ( .A1(n_403), .A2(n_345), .A3(n_372), .B1(n_380), .B2(n_381), .B3(n_196), .Y(n_441) );
AOI221xp5_ASAP7_75t_L g442 ( .A1(n_400), .A2(n_374), .B1(n_301), .B2(n_212), .C(n_369), .Y(n_442) );
INVxp67_ASAP7_75t_L g443 ( .A(n_409), .Y(n_443) );
AOI22xp33_ASAP7_75t_L g444 ( .A1(n_400), .A2(n_363), .B1(n_369), .B2(n_329), .Y(n_444) );
INVxp67_ASAP7_75t_SL g445 ( .A(n_411), .Y(n_445) );
AOI221xp5_ASAP7_75t_L g446 ( .A1(n_414), .A2(n_212), .B1(n_369), .B2(n_114), .C(n_82), .Y(n_446) );
INVx2_ASAP7_75t_L g447 ( .A(n_411), .Y(n_447) );
AO21x2_ASAP7_75t_L g448 ( .A1(n_414), .A2(n_383), .B(n_393), .Y(n_448) );
AND2x4_ASAP7_75t_L g449 ( .A(n_426), .B(n_394), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_424), .Y(n_450) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_418), .Y(n_451) );
NAND4xp25_ASAP7_75t_SL g452 ( .A(n_415), .B(n_317), .C(n_329), .D(n_16), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_398), .B(n_388), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_424), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_398), .B(n_383), .Y(n_455) );
HB1xp67_ASAP7_75t_L g456 ( .A(n_418), .Y(n_456) );
OAI221xp5_ASAP7_75t_L g457 ( .A1(n_417), .A2(n_393), .B1(n_346), .B2(n_366), .C(n_114), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_426), .B(n_317), .Y(n_458) );
INVx1_ASAP7_75t_L g459 ( .A(n_424), .Y(n_459) );
OAI31xp33_ASAP7_75t_L g460 ( .A1(n_399), .A2(n_346), .A3(n_356), .B(n_357), .Y(n_460) );
INVx1_ASAP7_75t_SL g461 ( .A(n_422), .Y(n_461) );
AND2x4_ASAP7_75t_L g462 ( .A(n_422), .B(n_332), .Y(n_462) );
NAND3xp33_ASAP7_75t_L g463 ( .A(n_446), .B(n_408), .C(n_405), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_455), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_436), .Y(n_465) );
AND2x2_ASAP7_75t_L g466 ( .A(n_438), .B(n_408), .Y(n_466) );
NOR2xp33_ASAP7_75t_L g467 ( .A(n_458), .B(n_410), .Y(n_467) );
OAI22xp33_ASAP7_75t_SL g468 ( .A1(n_443), .A2(n_406), .B1(n_423), .B2(n_407), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_455), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_448), .Y(n_470) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_452), .B(n_401), .Y(n_471) );
AND2x2_ASAP7_75t_L g472 ( .A(n_438), .B(n_401), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_437), .B(n_407), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_437), .B(n_419), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_436), .Y(n_475) );
INVx2_ASAP7_75t_L g476 ( .A(n_436), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g477 ( .A1(n_452), .A2(n_423), .B1(n_402), .B2(n_406), .Y(n_477) );
AOI33xp33_ASAP7_75t_L g478 ( .A1(n_430), .A2(n_402), .A3(n_417), .B1(n_419), .B2(n_416), .B3(n_420), .Y(n_478) );
BUFx3_ASAP7_75t_L g479 ( .A(n_462), .Y(n_479) );
INVx3_ASAP7_75t_L g480 ( .A(n_447), .Y(n_480) );
AND2x2_ASAP7_75t_L g481 ( .A(n_459), .B(n_425), .Y(n_481) );
INVx1_ASAP7_75t_L g482 ( .A(n_448), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_448), .Y(n_483) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_461), .B(n_406), .Y(n_484) );
AOI22xp5_ASAP7_75t_L g485 ( .A1(n_442), .A2(n_399), .B1(n_402), .B2(n_421), .Y(n_485) );
BUFx2_ASAP7_75t_L g486 ( .A(n_445), .Y(n_486) );
OAI222xp33_ASAP7_75t_L g487 ( .A1(n_433), .A2(n_421), .B1(n_13), .B2(n_14), .C1(n_410), .C2(n_357), .Y(n_487) );
INVxp67_ASAP7_75t_L g488 ( .A(n_427), .Y(n_488) );
OA332x1_ASAP7_75t_L g489 ( .A1(n_441), .A2(n_13), .A3(n_410), .B1(n_143), .B2(n_26), .B3(n_27), .C1(n_30), .C2(n_31), .Y(n_489) );
INVx1_ASAP7_75t_L g490 ( .A(n_448), .Y(n_490) );
INVxp67_ASAP7_75t_L g491 ( .A(n_451), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_459), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_447), .B(n_425), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_447), .Y(n_494) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_460), .A2(n_425), .B1(n_185), .B2(n_332), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_450), .Y(n_496) );
INVxp67_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_460), .A2(n_425), .B1(n_332), .B2(n_326), .Y(n_498) );
NAND3xp33_ASAP7_75t_L g499 ( .A(n_446), .B(n_212), .C(n_294), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_450), .B(n_212), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_450), .Y(n_501) );
OAI31xp33_ASAP7_75t_L g502 ( .A1(n_439), .A2(n_356), .A3(n_323), .B(n_319), .Y(n_502) );
AO21x2_ASAP7_75t_L g503 ( .A1(n_434), .A2(n_303), .B(n_238), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_454), .Y(n_504) );
INVx2_ASAP7_75t_SL g505 ( .A(n_461), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g506 ( .A1(n_442), .A2(n_212), .B1(n_323), .B2(n_294), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_453), .B(n_319), .Y(n_507) );
AOI22xp33_ASAP7_75t_SL g508 ( .A1(n_457), .A2(n_294), .B1(n_246), .B2(n_248), .Y(n_508) );
NAND3xp33_ASAP7_75t_L g509 ( .A(n_444), .B(n_294), .C(n_193), .Y(n_509) );
AND2x2_ASAP7_75t_L g510 ( .A(n_454), .B(n_20), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_454), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_453), .B(n_21), .Y(n_512) );
INVx2_ASAP7_75t_SL g513 ( .A(n_486), .Y(n_513) );
OR2x2_ASAP7_75t_L g514 ( .A(n_472), .B(n_429), .Y(n_514) );
NAND2xp5_ASAP7_75t_L g515 ( .A(n_473), .B(n_449), .Y(n_515) );
INVxp67_ASAP7_75t_L g516 ( .A(n_486), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_492), .Y(n_517) );
OR2x2_ASAP7_75t_L g518 ( .A(n_472), .B(n_429), .Y(n_518) );
AND2x2_ASAP7_75t_L g519 ( .A(n_474), .B(n_432), .Y(n_519) );
INVx2_ASAP7_75t_L g520 ( .A(n_480), .Y(n_520) );
INVx1_ASAP7_75t_L g521 ( .A(n_492), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_488), .Y(n_522) );
AND2x4_ASAP7_75t_SL g523 ( .A(n_477), .B(n_462), .Y(n_523) );
OR2x6_ASAP7_75t_L g524 ( .A(n_471), .B(n_462), .Y(n_524) );
NOR4xp75_ASAP7_75t_L g525 ( .A(n_484), .B(n_458), .C(n_457), .D(n_428), .Y(n_525) );
INVx1_ASAP7_75t_SL g526 ( .A(n_479), .Y(n_526) );
NOR3xp33_ASAP7_75t_SL g527 ( .A(n_487), .B(n_428), .C(n_431), .Y(n_527) );
NOR2x1_ASAP7_75t_L g528 ( .A(n_471), .B(n_462), .Y(n_528) );
AND2x2_ASAP7_75t_L g529 ( .A(n_464), .B(n_432), .Y(n_529) );
AND2x2_ASAP7_75t_L g530 ( .A(n_474), .B(n_449), .Y(n_530) );
BUFx3_ASAP7_75t_L g531 ( .A(n_505), .Y(n_531) );
NAND5xp2_ASAP7_75t_L g532 ( .A(n_502), .B(n_433), .C(n_434), .D(n_440), .E(n_449), .Y(n_532) );
NAND2xp5_ASAP7_75t_L g533 ( .A(n_491), .B(n_449), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_497), .B(n_440), .Y(n_534) );
NOR2xp33_ASAP7_75t_L g535 ( .A(n_467), .B(n_440), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_479), .B(n_440), .Y(n_536) );
AND2x2_ASAP7_75t_L g537 ( .A(n_512), .B(n_435), .Y(n_537) );
INVx1_ASAP7_75t_SL g538 ( .A(n_512), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_464), .Y(n_539) );
NAND4xp25_ASAP7_75t_L g540 ( .A(n_485), .B(n_435), .C(n_177), .D(n_184), .Y(n_540) );
INVx2_ASAP7_75t_L g541 ( .A(n_480), .Y(n_541) );
NOR3xp33_ASAP7_75t_L g542 ( .A(n_468), .B(n_435), .C(n_283), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_469), .Y(n_543) );
XNOR2xp5_ASAP7_75t_L g544 ( .A(n_485), .B(n_435), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_505), .B(n_32), .Y(n_545) );
OAI33xp33_ASAP7_75t_L g546 ( .A1(n_468), .A2(n_177), .A3(n_188), .B1(n_196), .B2(n_208), .B3(n_209), .Y(n_546) );
OAI31xp33_ASAP7_75t_L g547 ( .A1(n_489), .A2(n_282), .A3(n_283), .B(n_277), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_469), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_466), .B(n_33), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_466), .B(n_34), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_496), .B(n_294), .Y(n_551) );
NOR3xp33_ASAP7_75t_L g552 ( .A(n_463), .B(n_277), .C(n_271), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_496), .Y(n_553) );
NAND2xp5_ASAP7_75t_L g554 ( .A(n_501), .B(n_36), .Y(n_554) );
NOR2xp33_ASAP7_75t_L g555 ( .A(n_463), .B(n_38), .Y(n_555) );
OAI221xp5_ASAP7_75t_L g556 ( .A1(n_498), .A2(n_238), .B1(n_271), .B2(n_269), .C(n_248), .Y(n_556) );
HB1xp67_ASAP7_75t_L g557 ( .A(n_480), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_465), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_501), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_511), .B(n_46), .Y(n_560) );
NOR2xp33_ASAP7_75t_L g561 ( .A(n_507), .B(n_47), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_511), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_465), .B(n_52), .Y(n_563) );
OR2x2_ASAP7_75t_L g564 ( .A(n_475), .B(n_53), .Y(n_564) );
AND2x2_ASAP7_75t_L g565 ( .A(n_475), .B(n_55), .Y(n_565) );
INVx1_ASAP7_75t_L g566 ( .A(n_476), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_481), .B(n_56), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_510), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_476), .B(n_58), .Y(n_569) );
BUFx2_ASAP7_75t_L g570 ( .A(n_494), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_494), .Y(n_571) );
INVx3_ASAP7_75t_L g572 ( .A(n_504), .Y(n_572) );
NAND3xp33_ASAP7_75t_L g573 ( .A(n_542), .B(n_470), .C(n_490), .Y(n_573) );
XNOR2xp5_ASAP7_75t_L g574 ( .A(n_544), .B(n_481), .Y(n_574) );
INVx2_ASAP7_75t_L g575 ( .A(n_558), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_517), .Y(n_576) );
AND2x2_ASAP7_75t_L g577 ( .A(n_530), .B(n_519), .Y(n_577) );
AOI22xp33_ASAP7_75t_SL g578 ( .A1(n_523), .A2(n_509), .B1(n_499), .B2(n_510), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_521), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_514), .B(n_504), .Y(n_580) );
AND2x2_ASAP7_75t_L g581 ( .A(n_529), .B(n_493), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_522), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g583 ( .A(n_529), .B(n_493), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_513), .B(n_470), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g585 ( .A(n_539), .B(n_543), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_548), .Y(n_586) );
INVx2_ASAP7_75t_L g587 ( .A(n_558), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_553), .Y(n_588) );
INVx1_ASAP7_75t_L g589 ( .A(n_559), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_572), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_513), .B(n_490), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_516), .B(n_482), .Y(n_592) );
NAND4xp75_ASAP7_75t_L g593 ( .A(n_527), .B(n_482), .C(n_483), .D(n_500), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_572), .Y(n_594) );
AND2x2_ASAP7_75t_L g595 ( .A(n_572), .B(n_483), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_516), .B(n_478), .Y(n_596) );
NAND2xp33_ASAP7_75t_L g597 ( .A(n_538), .B(n_499), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_533), .B(n_495), .Y(n_598) );
AOI221x1_ASAP7_75t_L g599 ( .A1(n_542), .A2(n_509), .B1(n_500), .B2(n_503), .C(n_508), .Y(n_599) );
BUFx3_ASAP7_75t_L g600 ( .A(n_531), .Y(n_600) );
BUFx2_ASAP7_75t_L g601 ( .A(n_531), .Y(n_601) );
NAND2x1p5_ASAP7_75t_L g602 ( .A(n_528), .B(n_506), .Y(n_602) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_570), .B(n_503), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_518), .B(n_503), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_562), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_515), .B(n_534), .Y(n_606) );
AOI21xp5_ASAP7_75t_L g607 ( .A1(n_546), .A2(n_248), .B(n_246), .Y(n_607) );
AND2x4_ASAP7_75t_L g608 ( .A(n_524), .B(n_60), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_557), .B(n_62), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_566), .Y(n_610) );
NAND3xp33_ASAP7_75t_L g611 ( .A(n_555), .B(n_193), .C(n_192), .Y(n_611) );
AND2x2_ASAP7_75t_L g612 ( .A(n_557), .B(n_65), .Y(n_612) );
AND2x2_ASAP7_75t_L g613 ( .A(n_520), .B(n_71), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_526), .Y(n_614) );
INVx1_ASAP7_75t_SL g615 ( .A(n_536), .Y(n_615) );
INVx2_ASAP7_75t_SL g616 ( .A(n_524), .Y(n_616) );
AND2x2_ASAP7_75t_L g617 ( .A(n_520), .B(n_541), .Y(n_617) );
OAI21xp33_ASAP7_75t_L g618 ( .A1(n_532), .A2(n_192), .B(n_193), .Y(n_618) );
NOR2x1_ASAP7_75t_L g619 ( .A(n_540), .B(n_282), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_535), .B(n_72), .Y(n_620) );
NAND2xp5_ASAP7_75t_SL g621 ( .A(n_552), .B(n_248), .Y(n_621) );
AOI21xp5_ASAP7_75t_L g622 ( .A1(n_546), .A2(n_248), .B(n_246), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_541), .B(n_75), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_571), .Y(n_624) );
INVx2_ASAP7_75t_L g625 ( .A(n_551), .Y(n_625) );
AND2x2_ASAP7_75t_L g626 ( .A(n_537), .B(n_76), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_535), .B(n_80), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_596), .B(n_523), .Y(n_628) );
NAND2xp5_ASAP7_75t_L g629 ( .A(n_581), .B(n_568), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g630 ( .A1(n_621), .A2(n_524), .B(n_552), .Y(n_630) );
XNOR2x1_ASAP7_75t_L g631 ( .A(n_574), .B(n_525), .Y(n_631) );
AND2x2_ASAP7_75t_L g632 ( .A(n_577), .B(n_549), .Y(n_632) );
NAND2x1_ASAP7_75t_L g633 ( .A(n_601), .B(n_616), .Y(n_633) );
OAI21xp5_ASAP7_75t_SL g634 ( .A1(n_619), .A2(n_555), .B(n_561), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_580), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_584), .Y(n_636) );
AND2x2_ASAP7_75t_L g637 ( .A(n_577), .B(n_615), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_582), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_585), .Y(n_639) );
INVx1_ASAP7_75t_L g640 ( .A(n_586), .Y(n_640) );
XOR2x2_ASAP7_75t_L g641 ( .A(n_593), .B(n_550), .Y(n_641) );
OR2x2_ASAP7_75t_L g642 ( .A(n_583), .B(n_567), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_576), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_581), .B(n_527), .Y(n_644) );
NOR2xp67_ASAP7_75t_SL g645 ( .A(n_600), .B(n_564), .Y(n_645) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_588), .B(n_545), .Y(n_646) );
NAND3xp33_ASAP7_75t_L g647 ( .A(n_573), .B(n_599), .C(n_592), .Y(n_647) );
NOR2xp33_ASAP7_75t_L g648 ( .A(n_614), .B(n_561), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_579), .Y(n_649) );
XNOR2x2_ASAP7_75t_L g650 ( .A(n_620), .B(n_563), .Y(n_650) );
INVx1_ASAP7_75t_L g651 ( .A(n_589), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_605), .Y(n_652) );
INVx1_ASAP7_75t_SL g653 ( .A(n_600), .Y(n_653) );
INVxp67_ASAP7_75t_L g654 ( .A(n_614), .Y(n_654) );
OAI211xp5_ASAP7_75t_L g655 ( .A1(n_578), .A2(n_547), .B(n_560), .C(n_554), .Y(n_655) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_598), .A2(n_565), .B1(n_569), .B2(n_556), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_624), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_591), .Y(n_658) );
XNOR2xp5_ASAP7_75t_L g659 ( .A(n_606), .B(n_184), .Y(n_659) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_616), .B(n_193), .Y(n_660) );
OR2x2_ASAP7_75t_L g661 ( .A(n_604), .B(n_192), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_584), .Y(n_662) );
INVx1_ASAP7_75t_L g663 ( .A(n_610), .Y(n_663) );
INVx1_ASAP7_75t_L g664 ( .A(n_610), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_595), .B(n_193), .Y(n_665) );
INVx1_ASAP7_75t_L g666 ( .A(n_595), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_575), .Y(n_667) );
INVx2_ASAP7_75t_L g668 ( .A(n_575), .Y(n_668) );
INVx1_ASAP7_75t_L g669 ( .A(n_587), .Y(n_669) );
OAI32xp33_ASAP7_75t_L g670 ( .A1(n_602), .A2(n_269), .A3(n_188), .B1(n_208), .B2(n_209), .Y(n_670) );
A2O1A1Ixp33_ASAP7_75t_L g671 ( .A1(n_620), .A2(n_246), .B(n_192), .C(n_215), .Y(n_671) );
CKINVDCx5p33_ASAP7_75t_R g672 ( .A(n_626), .Y(n_672) );
INVx1_ASAP7_75t_L g673 ( .A(n_625), .Y(n_673) );
INVx1_ASAP7_75t_SL g674 ( .A(n_609), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_625), .B(n_192), .Y(n_675) );
HB1xp67_ASAP7_75t_L g676 ( .A(n_617), .Y(n_676) );
NAND2xp5_ASAP7_75t_SL g677 ( .A(n_608), .B(n_200), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_617), .Y(n_678) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_626), .A2(n_200), .B1(n_215), .B2(n_597), .Y(n_679) );
OAI21xp33_ASAP7_75t_L g680 ( .A1(n_603), .A2(n_215), .B(n_618), .Y(n_680) );
HB1xp67_ASAP7_75t_L g681 ( .A(n_590), .Y(n_681) );
OAI22xp5_ASAP7_75t_L g682 ( .A1(n_602), .A2(n_608), .B1(n_611), .B2(n_627), .Y(n_682) );
AOI22xp33_ASAP7_75t_L g683 ( .A1(n_597), .A2(n_609), .B1(n_612), .B2(n_621), .Y(n_683) );
O2A1O1Ixp5_ASAP7_75t_L g684 ( .A1(n_612), .A2(n_594), .B(n_613), .C(n_623), .Y(n_684) );
OR2x2_ASAP7_75t_L g685 ( .A(n_613), .B(n_623), .Y(n_685) );
CKINVDCx5p33_ASAP7_75t_R g686 ( .A(n_607), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_622), .Y(n_687) );
AOI22xp33_ASAP7_75t_L g688 ( .A1(n_574), .A2(n_532), .B1(n_452), .B2(n_523), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_582), .Y(n_689) );
O2A1O1Ixp33_ASAP7_75t_L g690 ( .A1(n_670), .A2(n_680), .B(n_671), .C(n_644), .Y(n_690) );
NOR2x1_ASAP7_75t_L g691 ( .A(n_633), .B(n_634), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_644), .B(n_658), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_672), .A2(n_653), .B1(n_688), .B2(n_683), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_662), .Y(n_694) );
INVx2_ASAP7_75t_L g695 ( .A(n_668), .Y(n_695) );
BUFx2_ASAP7_75t_L g696 ( .A(n_653), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g697 ( .A1(n_677), .A2(n_631), .B(n_630), .Y(n_697) );
OAI322xp33_ASAP7_75t_L g698 ( .A1(n_654), .A2(n_639), .A3(n_628), .B1(n_650), .B2(n_629), .C1(n_647), .C2(n_689), .Y(n_698) );
AOI211xp5_ASAP7_75t_L g699 ( .A1(n_634), .A2(n_682), .B(n_677), .C(n_655), .Y(n_699) );
AOI322xp5_ASAP7_75t_L g700 ( .A1(n_637), .A2(n_629), .A3(n_632), .B1(n_672), .B2(n_648), .C1(n_676), .C2(n_666), .Y(n_700) );
INVx1_ASAP7_75t_L g701 ( .A(n_643), .Y(n_701) );
XNOR2xp5_ASAP7_75t_L g702 ( .A(n_641), .B(n_659), .Y(n_702) );
CKINVDCx5p33_ASAP7_75t_R g703 ( .A(n_638), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_636), .B(n_649), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_699), .B(n_640), .Y(n_705) );
AOI222xp33_ASAP7_75t_L g706 ( .A1(n_693), .A2(n_651), .B1(n_652), .B2(n_657), .C1(n_646), .C2(n_674), .Y(n_706) );
OR2x2_ASAP7_75t_L g707 ( .A(n_692), .B(n_635), .Y(n_707) );
AOI22xp5_ASAP7_75t_L g708 ( .A1(n_697), .A2(n_679), .B1(n_686), .B2(n_646), .Y(n_708) );
OAI211xp5_ASAP7_75t_L g709 ( .A1(n_691), .A2(n_656), .B(n_671), .C(n_686), .Y(n_709) );
OAI22xp5_ASAP7_75t_L g710 ( .A1(n_696), .A2(n_642), .B1(n_678), .B2(n_685), .Y(n_710) );
AOI221xp5_ASAP7_75t_L g711 ( .A1(n_698), .A2(n_684), .B1(n_673), .B2(n_664), .C(n_663), .Y(n_711) );
INVx1_ASAP7_75t_L g712 ( .A(n_701), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_700), .B(n_681), .Y(n_713) );
OR4x1_ASAP7_75t_L g714 ( .A(n_712), .B(n_694), .C(n_702), .D(n_687), .Y(n_714) );
NOR2xp67_ASAP7_75t_SL g715 ( .A(n_709), .B(n_703), .Y(n_715) );
NAND3xp33_ASAP7_75t_SL g716 ( .A(n_708), .B(n_690), .C(n_661), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_705), .B(n_704), .Y(n_717) );
NAND3xp33_ASAP7_75t_L g718 ( .A(n_706), .B(n_690), .C(n_660), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_717), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
AOI22xp5_ASAP7_75t_L g721 ( .A1(n_715), .A2(n_713), .B1(n_711), .B2(n_710), .Y(n_721) );
AOI22xp5_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_716), .B1(n_714), .B2(n_707), .Y(n_722) );
NAND3xp33_ASAP7_75t_SL g723 ( .A(n_720), .B(n_665), .C(n_675), .Y(n_723) );
INVx1_ASAP7_75t_L g724 ( .A(n_723), .Y(n_724) );
OR2x6_ASAP7_75t_L g725 ( .A(n_722), .B(n_719), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_724), .Y(n_726) );
OAI22xp33_ASAP7_75t_L g727 ( .A1(n_726), .A2(n_725), .B1(n_695), .B2(n_665), .Y(n_727) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_727), .A2(n_695), .B1(n_645), .B2(n_669), .C(n_667), .Y(n_728) );
endmodule