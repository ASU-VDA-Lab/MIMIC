module real_jpeg_25483_n_14 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_2, n_13, n_6, n_7, n_3, n_10, n_9, n_14);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_2;
input n_13;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_14;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_146;
wire n_83;
wire n_78;
wire n_104;
wire n_153;
wire n_64;
wire n_131;
wire n_47;
wire n_22;
wire n_87;
wire n_105;
wire n_40;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_140;
wire n_126;
wire n_113;
wire n_155;
wire n_120;
wire n_93;
wire n_141;
wire n_95;
wire n_65;
wire n_33;
wire n_139;
wire n_142;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_156;
wire n_147;
wire n_66;
wire n_136;
wire n_44;
wire n_28;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_145;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_118;
wire n_17;
wire n_123;
wire n_116;
wire n_21;
wire n_50;
wire n_143;
wire n_69;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_134;
wire n_72;
wire n_151;
wire n_100;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_30;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_138;
wire n_25;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

AOI21xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_22),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_1),
.B(n_83),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g111 ( 
.A1(n_1),
.A2(n_26),
.B1(n_30),
.B2(n_32),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g115 ( 
.A1(n_1),
.A2(n_38),
.B(n_56),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_1),
.B(n_78),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g144 ( 
.A1(n_1),
.A2(n_35),
.B1(n_140),
.B2(n_145),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_2),
.A2(n_22),
.B1(n_23),
.B2(n_72),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_2),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_2),
.A2(n_26),
.B1(n_32),
.B2(n_72),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_2),
.A2(n_37),
.B1(n_38),
.B2(n_72),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g52 ( 
.A1(n_3),
.A2(n_26),
.B1(n_32),
.B2(n_53),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_3),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_3),
.A2(n_22),
.B1(n_23),
.B2(n_53),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_L g130 ( 
.A1(n_3),
.A2(n_37),
.B1(n_38),
.B2(n_53),
.Y(n_130)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_4),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

INVx8_ASAP7_75t_SL g87 ( 
.A(n_6),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_7),
.A2(n_37),
.B1(n_38),
.B2(n_44),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_7),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_7),
.A2(n_26),
.B1(n_32),
.B2(n_44),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_8),
.A2(n_37),
.B1(n_38),
.B2(n_50),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_8),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_11),
.A2(n_37),
.B1(n_38),
.B2(n_92),
.Y(n_91)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_11),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_12),
.A2(n_26),
.B1(n_32),
.B2(n_62),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_12),
.A2(n_37),
.B1(n_38),
.B2(n_62),
.Y(n_123)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_13),
.Y(n_41)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

INVx6_ASAP7_75t_L g133 ( 
.A(n_13),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g14 ( 
.A(n_15),
.B(n_105),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_104),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_17),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_73),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_18),
.B(n_73),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_51),
.C(n_63),
.Y(n_18)
);

AOI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_19),
.A2(n_20),
.B1(n_154),
.B2(n_156),
.Y(n_153)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_34),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_21),
.B(n_34),
.Y(n_96)
);

OAI32xp33_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_26),
.A3(n_28),
.B1(n_29),
.B2(n_31),
.Y(n_21)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_22),
.A2(n_23),
.B1(n_28),
.B2(n_33),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_22),
.A2(n_23),
.B1(n_85),
.B2(n_86),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_30),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp33_ASAP7_75t_L g55 ( 
.A1(n_26),
.A2(n_32),
.B1(n_56),
.B2(n_58),
.Y(n_55)
);

AOI22xp5_ASAP7_75t_L g69 ( 
.A1(n_26),
.A2(n_28),
.B1(n_32),
.B2(n_33),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_SL g114 ( 
.A1(n_26),
.A2(n_30),
.B(n_58),
.C(n_115),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_29),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g138 ( 
.A(n_30),
.B(n_59),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_30),
.B(n_41),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g34 ( 
.A1(n_35),
.A2(n_42),
.B(n_45),
.Y(n_34)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_35),
.A2(n_123),
.B(n_124),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_35),
.A2(n_130),
.B1(n_140),
.B2(n_141),
.Y(n_139)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_36),
.B(n_49),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_36),
.A2(n_129),
.B1(n_131),
.B2(n_132),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_37),
.B(n_40),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g59 ( 
.A1(n_37),
.A2(n_38),
.B1(n_56),
.B2(n_58),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_37),
.B(n_147),
.Y(n_146)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_40),
.Y(n_90)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_43),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_46),
.B(n_49),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_48),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_51),
.A2(n_63),
.B1(n_64),
.B2(n_155),
.Y(n_154)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_51),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_54),
.B1(n_60),
.B2(n_61),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_52),
.A2(n_54),
.B1(n_60),
.B2(n_113),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_54),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_59),
.Y(n_54)
);

INVx13_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

BUFx24_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_59),
.A2(n_98),
.B1(n_111),
.B2(n_112),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_60),
.B(n_101),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g99 ( 
.A(n_61),
.Y(n_99)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_68),
.A2(n_77),
.B1(n_78),
.B2(n_79),
.Y(n_76)
);

AND2x2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_70),
.Y(n_68)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_71),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_74),
.A2(n_75),
.B1(n_94),
.B2(n_95),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_80),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_88),
.B2(n_89),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx4_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g88 ( 
.A(n_89),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_91),
.B(n_93),
.Y(n_89)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_96),
.Y(n_102)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_97),
.Y(n_103)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_99),
.B(n_100),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_106),
.A2(n_151),
.B(n_157),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_107),
.A2(n_126),
.B(n_150),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_108),
.B(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g108 ( 
.A(n_109),
.B(n_114),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_109),
.A2(n_110),
.B1(n_114),
.B2(n_135),
.Y(n_134)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g135 ( 
.A(n_114),
.Y(n_135)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_122),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_118),
.A2(n_119),
.B1(n_120),
.B2(n_121),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_118),
.B(n_121),
.C(n_122),
.Y(n_152)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_120),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_123),
.Y(n_131)
);

AOI21xp5_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_136),
.B(n_149),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_128),
.B(n_134),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g149 ( 
.A(n_128),
.B(n_134),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g145 ( 
.A(n_132),
.Y(n_145)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_133),
.Y(n_142)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_143),
.B(n_148),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_138),
.B(n_139),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_138),
.B(n_139),
.Y(n_148)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_146),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_152),
.B(n_153),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_152),
.B(n_153),
.Y(n_157)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_154),
.Y(n_156)
);


endmodule