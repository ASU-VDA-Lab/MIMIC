module fake_aes_3636_n_23 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_23);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_23;
wire n_20;
wire n_22;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_19;
wire n_21;
NAND2xp5_ASAP7_75t_L g12 ( .A(n_4), .B(n_7), .Y(n_12) );
INVx1_ASAP7_75t_L g13 ( .A(n_8), .Y(n_13) );
CKINVDCx16_ASAP7_75t_R g14 ( .A(n_5), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_6), .B(n_3), .Y(n_15) );
NAND2xp5_ASAP7_75t_SL g16 ( .A(n_14), .B(n_0), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_17), .Y(n_18) );
INVx2_ASAP7_75t_SL g19 ( .A(n_18), .Y(n_19) );
AOI221xp5_ASAP7_75t_L g20 ( .A1(n_19), .A2(n_13), .B1(n_15), .B2(n_12), .C(n_10), .Y(n_20) );
BUFx2_ASAP7_75t_L g21 ( .A(n_20), .Y(n_21) );
NOR2xp67_ASAP7_75t_L g22 ( .A(n_21), .B(n_1), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_2), .B1(n_9), .B2(n_11), .Y(n_23) );
endmodule