module fake_jpeg_12567_n_43 (n_3, n_2, n_1, n_0, n_4, n_5, n_43);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_43;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_5),
.B(n_4),
.Y(n_6)
);

INVx2_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx8_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_3),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

AOI22xp33_ASAP7_75t_SL g11 ( 
.A1(n_0),
.A2(n_4),
.B1(n_1),
.B2(n_2),
.Y(n_11)
);

BUFx6f_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

INVx2_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_SL g14 ( 
.A(n_6),
.B(n_3),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_14),
.B(n_19),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g15 ( 
.A(n_6),
.B(n_9),
.Y(n_15)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_15),
.B(n_20),
.C(n_18),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_SL g16 ( 
.A1(n_8),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_16),
.A2(n_11),
.B1(n_13),
.B2(n_12),
.Y(n_27)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_7),
.A2(n_9),
.B1(n_10),
.B2(n_13),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g29 ( 
.A1(n_17),
.A2(n_0),
.B1(n_1),
.B2(n_5),
.Y(n_29)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_20),
.B(n_21),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

INVx4_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_22),
.Y(n_23)
);

AO22x1_ASAP7_75t_L g31 ( 
.A1(n_27),
.A2(n_28),
.B1(n_16),
.B2(n_22),
.Y(n_31)
);

AOI22xp5_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_14),
.B1(n_15),
.B2(n_21),
.Y(n_33)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

BUFx2_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_SL g36 ( 
.A1(n_31),
.A2(n_32),
.B1(n_33),
.B2(n_24),
.Y(n_36)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_33),
.A2(n_27),
.B1(n_29),
.B2(n_28),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_35),
.B(n_36),
.Y(n_39)
);

OAI21xp5_ASAP7_75t_SL g37 ( 
.A1(n_35),
.A2(n_31),
.B(n_30),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_37),
.B(n_22),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g38 ( 
.A1(n_34),
.A2(n_23),
.B(n_25),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_38),
.B(n_34),
.Y(n_40)
);

AOI221xp5_ASAP7_75t_L g42 ( 
.A1(n_40),
.A2(n_41),
.B1(n_39),
.B2(n_17),
.C(n_21),
.Y(n_42)
);

XNOR2xp5_ASAP7_75t_L g43 ( 
.A(n_42),
.B(n_1),
.Y(n_43)
);


endmodule