module fake_jpeg_29816_n_160 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_40, n_19, n_18, n_20, n_35, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_160);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_160;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx4_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_13),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

BUFx12f_ASAP7_75t_L g49 ( 
.A(n_2),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

BUFx10_ASAP7_75t_L g52 ( 
.A(n_44),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_23),
.Y(n_53)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_40),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g56 ( 
.A(n_11),
.Y(n_56)
);

BUFx10_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_18),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_42),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_4),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_31),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_28),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_27),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_15),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_1),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g67 ( 
.A(n_51),
.Y(n_67)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_67),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_46),
.B(n_0),
.Y(n_68)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_60),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g69 ( 
.A(n_51),
.Y(n_69)
);

BUFx8_ASAP7_75t_L g89 ( 
.A(n_69),
.Y(n_89)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_64),
.Y(n_70)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_70),
.Y(n_78)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_50),
.Y(n_71)
);

HB1xp67_ASAP7_75t_L g83 ( 
.A(n_71),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_48),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_72),
.Y(n_85)
);

INVx4_ASAP7_75t_SL g73 ( 
.A(n_56),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_74),
.Y(n_90)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_54),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_45),
.Y(n_75)
);

BUFx12_ASAP7_75t_L g87 ( 
.A(n_75),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_61),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_76),
.B(n_77),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_73),
.B(n_61),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_67),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_79),
.B(n_82),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_72),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_68),
.B(n_60),
.Y(n_82)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_84),
.B(n_88),
.Y(n_103)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_68),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_54),
.C(n_55),
.Y(n_88)
);

INVxp67_ASAP7_75t_L g91 ( 
.A(n_90),
.Y(n_91)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_91),
.B(n_8),
.Y(n_122)
);

OAI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_83),
.A2(n_59),
.B1(n_53),
.B2(n_63),
.Y(n_92)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_92),
.A2(n_100),
.B1(n_106),
.B2(n_108),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g94 ( 
.A1(n_84),
.A2(n_55),
.B(n_47),
.Y(n_94)
);

INVxp67_ASAP7_75t_L g126 ( 
.A(n_94),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_78),
.A2(n_49),
.B1(n_64),
.B2(n_57),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_95),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_62),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_96),
.B(n_3),
.Y(n_110)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_81),
.Y(n_97)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_97),
.Y(n_111)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_98),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_99),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_78),
.A2(n_65),
.B1(n_58),
.B2(n_3),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_89),
.B(n_49),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_101),
.B(n_107),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_87),
.A2(n_57),
.B(n_52),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_6),
.C(n_7),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_87),
.A2(n_52),
.B1(n_25),
.B2(n_26),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_89),
.B(n_0),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_80),
.A2(n_24),
.B1(n_43),
.B2(n_41),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g109 ( 
.A(n_84),
.B(n_1),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_109),
.B(n_8),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_110),
.B(n_120),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g113 ( 
.A1(n_92),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_113),
.A2(n_35),
.B1(n_37),
.B2(n_38),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_115),
.B(n_123),
.Y(n_137)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_99),
.Y(n_116)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_116),
.Y(n_130)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_117),
.Y(n_140)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_102),
.Y(n_119)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_119),
.Y(n_142)
);

OR2x2_ASAP7_75t_L g120 ( 
.A(n_109),
.B(n_104),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_122),
.B(n_125),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_103),
.B(n_9),
.Y(n_125)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_103),
.B(n_9),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_127),
.B(n_10),
.Y(n_131)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_95),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_128),
.B(n_129),
.Y(n_138)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_97),
.Y(n_129)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_136),
.C(n_126),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_121),
.A2(n_10),
.B1(n_12),
.B2(n_14),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_132),
.B(n_121),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g133 ( 
.A(n_111),
.Y(n_133)
);

OR2x2_ASAP7_75t_L g150 ( 
.A(n_133),
.B(n_127),
.Y(n_150)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_120),
.A2(n_17),
.B(n_20),
.C(n_21),
.D(n_22),
.Y(n_136)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_118),
.A2(n_29),
.B1(n_30),
.B2(n_32),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_139),
.B(n_143),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g141 ( 
.A(n_112),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_141),
.B(n_114),
.Y(n_145)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_130),
.Y(n_144)
);

NAND3xp33_ASAP7_75t_L g153 ( 
.A(n_144),
.B(n_146),
.C(n_149),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g151 ( 
.A(n_145),
.B(n_138),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_148),
.A2(n_150),
.B1(n_113),
.B2(n_135),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_124),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_151),
.B(n_140),
.C(n_137),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_152),
.A2(n_148),
.B(n_147),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_154),
.B(n_155),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_141),
.Y(n_157)
);

OAI221xp5_ASAP7_75t_L g158 ( 
.A1(n_157),
.A2(n_136),
.B1(n_134),
.B2(n_153),
.C(n_141),
.Y(n_158)
);

AOI21xp5_ASAP7_75t_L g159 ( 
.A1(n_158),
.A2(n_123),
.B(n_131),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_159),
.B(n_39),
.Y(n_160)
);


endmodule