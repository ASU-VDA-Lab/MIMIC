module fake_aes_10435_n_627 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_627);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_627;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_612;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_162;
wire n_387;
wire n_163;
wire n_476;
wire n_105;
wire n_227;
wire n_384;
wire n_434;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_586;
wire n_244;
wire n_540;
wire n_563;
wire n_73;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_554;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_610;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_621;
wire n_370;
wire n_589;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_363;
wire n_315;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_618;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_469;
wire n_585;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g73 ( .A(n_66), .Y(n_73) );
INVx1_ASAP7_75t_L g74 ( .A(n_0), .Y(n_74) );
CKINVDCx5p33_ASAP7_75t_R g75 ( .A(n_38), .Y(n_75) );
INVx1_ASAP7_75t_L g76 ( .A(n_44), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_34), .Y(n_77) );
NOR2xp67_ASAP7_75t_L g78 ( .A(n_72), .B(n_43), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_35), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_24), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_29), .Y(n_81) );
CKINVDCx16_ASAP7_75t_R g82 ( .A(n_59), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_32), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_13), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
BUFx6f_ASAP7_75t_L g86 ( .A(n_1), .Y(n_86) );
INVx1_ASAP7_75t_SL g87 ( .A(n_42), .Y(n_87) );
INVx1_ASAP7_75t_SL g88 ( .A(n_3), .Y(n_88) );
CKINVDCx5p33_ASAP7_75t_R g89 ( .A(n_4), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_33), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_50), .Y(n_91) );
INVx1_ASAP7_75t_L g92 ( .A(n_52), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_14), .Y(n_93) );
INVx2_ASAP7_75t_SL g94 ( .A(n_54), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_7), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_11), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_64), .Y(n_97) );
INVxp33_ASAP7_75t_L g98 ( .A(n_31), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_10), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_61), .Y(n_100) );
INVxp33_ASAP7_75t_SL g101 ( .A(n_20), .Y(n_101) );
NOR2xp67_ASAP7_75t_L g102 ( .A(n_7), .B(n_11), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_49), .Y(n_103) );
INVxp33_ASAP7_75t_L g104 ( .A(n_39), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_9), .Y(n_105) );
CKINVDCx5p33_ASAP7_75t_R g106 ( .A(n_30), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_13), .Y(n_107) );
INVxp67_ASAP7_75t_L g108 ( .A(n_2), .Y(n_108) );
BUFx6f_ASAP7_75t_L g109 ( .A(n_62), .Y(n_109) );
INVxp33_ASAP7_75t_L g110 ( .A(n_37), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_2), .Y(n_111) );
INVxp67_ASAP7_75t_SL g112 ( .A(n_22), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_3), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_4), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_6), .Y(n_115) );
BUFx2_ASAP7_75t_SL g116 ( .A(n_12), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_18), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_94), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_73), .Y(n_119) );
CKINVDCx20_ASAP7_75t_R g120 ( .A(n_89), .Y(n_120) );
NOR2xp67_ASAP7_75t_L g121 ( .A(n_94), .B(n_0), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_73), .Y(n_122) );
CKINVDCx5p33_ASAP7_75t_R g123 ( .A(n_82), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g124 ( .A(n_109), .B(n_1), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_83), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_83), .Y(n_126) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_89), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_127) );
CKINVDCx5p33_ASAP7_75t_R g128 ( .A(n_75), .Y(n_128) );
INVx2_ASAP7_75t_L g129 ( .A(n_90), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_76), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_77), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_86), .Y(n_132) );
BUFx3_ASAP7_75t_L g133 ( .A(n_90), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_79), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_80), .Y(n_135) );
NOR2xp33_ASAP7_75t_R g136 ( .A(n_75), .B(n_41), .Y(n_136) );
BUFx6f_ASAP7_75t_L g137 ( .A(n_109), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_106), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_81), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_91), .Y(n_140) );
BUFx6f_ASAP7_75t_L g141 ( .A(n_109), .Y(n_141) );
NAND2xp5_ASAP7_75t_L g142 ( .A(n_108), .B(n_5), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_106), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_109), .Y(n_144) );
INVx2_ASAP7_75t_L g145 ( .A(n_92), .Y(n_145) );
AND2x2_ASAP7_75t_L g146 ( .A(n_98), .B(n_8), .Y(n_146) );
BUFx6f_ASAP7_75t_L g147 ( .A(n_109), .Y(n_147) );
NOR2xp33_ASAP7_75t_L g148 ( .A(n_97), .B(n_9), .Y(n_148) );
NAND2xp5_ASAP7_75t_L g149 ( .A(n_99), .B(n_10), .Y(n_149) );
HB1xp67_ASAP7_75t_L g150 ( .A(n_99), .Y(n_150) );
INVx2_ASAP7_75t_SL g151 ( .A(n_100), .Y(n_151) );
INVx3_ASAP7_75t_L g152 ( .A(n_86), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_101), .Y(n_153) );
INVx1_ASAP7_75t_L g154 ( .A(n_103), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_117), .Y(n_155) );
INVxp67_ASAP7_75t_L g156 ( .A(n_116), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_132), .Y(n_157) );
CKINVDCx20_ASAP7_75t_R g158 ( .A(n_120), .Y(n_158) );
AND2x2_ASAP7_75t_L g159 ( .A(n_119), .B(n_104), .Y(n_159) );
INVx1_ASAP7_75t_L g160 ( .A(n_132), .Y(n_160) );
CKINVDCx5p33_ASAP7_75t_R g161 ( .A(n_128), .Y(n_161) );
NAND2xp5_ASAP7_75t_SL g162 ( .A(n_138), .B(n_110), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_137), .Y(n_163) );
INVx2_ASAP7_75t_L g164 ( .A(n_137), .Y(n_164) );
BUFx2_ASAP7_75t_L g165 ( .A(n_143), .Y(n_165) );
NAND2xp33_ASAP7_75t_L g166 ( .A(n_153), .B(n_130), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_137), .Y(n_167) );
NAND2xp5_ASAP7_75t_L g168 ( .A(n_119), .B(n_101), .Y(n_168) );
AND2x4_ASAP7_75t_L g169 ( .A(n_118), .B(n_115), .Y(n_169) );
INVx3_ASAP7_75t_L g170 ( .A(n_129), .Y(n_170) );
NAND2xp5_ASAP7_75t_SL g171 ( .A(n_156), .B(n_87), .Y(n_171) );
INVx1_ASAP7_75t_L g172 ( .A(n_132), .Y(n_172) );
INVx3_ASAP7_75t_L g173 ( .A(n_129), .Y(n_173) );
AOI22xp33_ASAP7_75t_L g174 ( .A1(n_122), .A2(n_85), .B1(n_115), .B2(n_84), .Y(n_174) );
HB1xp67_ASAP7_75t_L g175 ( .A(n_150), .Y(n_175) );
NOR2xp33_ASAP7_75t_L g176 ( .A(n_118), .B(n_112), .Y(n_176) );
INVx1_ASAP7_75t_L g177 ( .A(n_132), .Y(n_177) );
BUFx6f_ASAP7_75t_L g178 ( .A(n_137), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_152), .Y(n_179) );
INVx1_ASAP7_75t_SL g180 ( .A(n_146), .Y(n_180) );
INVx1_ASAP7_75t_L g181 ( .A(n_152), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_137), .Y(n_182) );
AND2x2_ASAP7_75t_L g183 ( .A(n_122), .B(n_84), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_137), .Y(n_184) );
BUFx3_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
AND2x2_ASAP7_75t_L g186 ( .A(n_125), .B(n_85), .Y(n_186) );
BUFx10_ASAP7_75t_L g187 ( .A(n_123), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_141), .Y(n_188) );
INVx2_ASAP7_75t_L g189 ( .A(n_141), .Y(n_189) );
NAND2x1p5_ASAP7_75t_L g190 ( .A(n_146), .B(n_78), .Y(n_190) );
NAND2xp5_ASAP7_75t_SL g191 ( .A(n_125), .B(n_114), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_126), .B(n_130), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_126), .B(n_74), .Y(n_193) );
INVx1_ASAP7_75t_L g194 ( .A(n_152), .Y(n_194) );
INVx4_ASAP7_75t_L g195 ( .A(n_133), .Y(n_195) );
NAND2xp5_ASAP7_75t_SL g196 ( .A(n_151), .B(n_114), .Y(n_196) );
AOI22xp33_ASAP7_75t_L g197 ( .A1(n_131), .A2(n_113), .B1(n_111), .B2(n_107), .Y(n_197) );
BUFx3_ASAP7_75t_L g198 ( .A(n_151), .Y(n_198) );
AND2x2_ASAP7_75t_L g199 ( .A(n_131), .B(n_95), .Y(n_199) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_134), .B(n_135), .Y(n_200) );
INVx3_ASAP7_75t_L g201 ( .A(n_152), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_141), .Y(n_202) );
INVx2_ASAP7_75t_L g203 ( .A(n_141), .Y(n_203) );
BUFx3_ASAP7_75t_L g204 ( .A(n_145), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_155), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_145), .Y(n_207) );
INVx1_ASAP7_75t_L g208 ( .A(n_204), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_180), .A2(n_149), .B1(n_142), .B2(n_121), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_201), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_204), .Y(n_211) );
BUFx3_ASAP7_75t_L g212 ( .A(n_185), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g213 ( .A(n_159), .B(n_154), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_204), .Y(n_214) );
INVx1_ASAP7_75t_L g215 ( .A(n_185), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g216 ( .A(n_159), .B(n_154), .Y(n_216) );
OAI22xp5_ASAP7_75t_L g217 ( .A1(n_180), .A2(n_139), .B1(n_134), .B2(n_135), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g218 ( .A(n_168), .B(n_140), .Y(n_218) );
CKINVDCx5p33_ASAP7_75t_R g219 ( .A(n_158), .Y(n_219) );
NOR2xp67_ASAP7_75t_SL g220 ( .A(n_159), .B(n_116), .Y(n_220) );
INVx4_ASAP7_75t_L g221 ( .A(n_195), .Y(n_221) );
AND2x2_ASAP7_75t_L g222 ( .A(n_175), .B(n_140), .Y(n_222) );
AOI22xp33_ASAP7_75t_L g223 ( .A1(n_183), .A2(n_139), .B1(n_148), .B2(n_105), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_168), .B(n_121), .Y(n_224) );
NOR3xp33_ASAP7_75t_SL g225 ( .A(n_161), .B(n_127), .C(n_96), .Y(n_225) );
AOI221xp5_ASAP7_75t_SL g226 ( .A1(n_174), .A2(n_124), .B1(n_93), .B2(n_86), .C(n_88), .Y(n_226) );
HB1xp67_ASAP7_75t_L g227 ( .A(n_175), .Y(n_227) );
INVx1_ASAP7_75t_L g228 ( .A(n_185), .Y(n_228) );
OAI22xp5_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_102), .B1(n_86), .B2(n_141), .Y(n_229) );
NOR2xp33_ASAP7_75t_SL g230 ( .A(n_165), .B(n_86), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_198), .B(n_136), .Y(n_231) );
OAI22xp5_ASAP7_75t_SL g232 ( .A1(n_165), .A2(n_12), .B1(n_14), .B2(n_15), .Y(n_232) );
NAND2xp5_ASAP7_75t_SL g233 ( .A(n_192), .B(n_147), .Y(n_233) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_198), .B(n_147), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_205), .Y(n_235) );
INVx1_ASAP7_75t_L g236 ( .A(n_205), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_206), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_192), .Y(n_238) );
AOI22xp5_ASAP7_75t_L g239 ( .A1(n_166), .A2(n_147), .B1(n_144), .B2(n_141), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g240 ( .A(n_171), .B(n_196), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_201), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_198), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_201), .Y(n_243) );
INVx3_ASAP7_75t_L g244 ( .A(n_195), .Y(n_244) );
O2A1O1Ixp33_ASAP7_75t_L g245 ( .A1(n_200), .A2(n_16), .B(n_17), .C(n_19), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_200), .B(n_147), .Y(n_246) );
NAND2xp5_ASAP7_75t_SL g247 ( .A(n_169), .B(n_147), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_169), .B(n_147), .Y(n_248) );
INVxp67_ASAP7_75t_L g249 ( .A(n_187), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_206), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_195), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_191), .A2(n_144), .B1(n_23), .B2(n_25), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_201), .Y(n_253) );
O2A1O1Ixp33_ASAP7_75t_L g254 ( .A1(n_193), .A2(n_21), .B(n_26), .C(n_27), .Y(n_254) );
AO22x1_ASAP7_75t_L g255 ( .A1(n_169), .A2(n_144), .B1(n_36), .B2(n_40), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_207), .Y(n_256) );
AND2x2_ASAP7_75t_L g257 ( .A(n_187), .B(n_144), .Y(n_257) );
AND2x4_ASAP7_75t_L g258 ( .A(n_183), .B(n_144), .Y(n_258) );
A2O1A1Ixp33_ASAP7_75t_L g259 ( .A1(n_183), .A2(n_144), .B(n_45), .C(n_46), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_169), .B(n_28), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g261 ( .A(n_195), .B(n_47), .Y(n_261) );
OR2x6_ASAP7_75t_L g262 ( .A(n_190), .B(n_48), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_238), .Y(n_263) );
NOR2xp33_ASAP7_75t_L g264 ( .A(n_213), .B(n_190), .Y(n_264) );
AOI21x1_ASAP7_75t_L g265 ( .A1(n_260), .A2(n_193), .B(n_186), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_210), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_221), .Y(n_267) );
AOI22xp33_ASAP7_75t_L g268 ( .A1(n_218), .A2(n_186), .B1(n_199), .B2(n_207), .Y(n_268) );
BUFx12f_ASAP7_75t_L g269 ( .A(n_219), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g270 ( .A(n_230), .B(n_190), .Y(n_270) );
A2O1A1Ixp33_ASAP7_75t_L g271 ( .A1(n_218), .A2(n_186), .B(n_199), .C(n_176), .Y(n_271) );
INVx3_ASAP7_75t_L g272 ( .A(n_221), .Y(n_272) );
INVx2_ASAP7_75t_L g273 ( .A(n_210), .Y(n_273) );
AOI21xp5_ASAP7_75t_L g274 ( .A1(n_233), .A2(n_162), .B(n_190), .Y(n_274) );
OR2x6_ASAP7_75t_SL g275 ( .A(n_219), .B(n_187), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_222), .B(n_199), .Y(n_276) );
AOI21xp5_ASAP7_75t_L g277 ( .A1(n_233), .A2(n_194), .B(n_181), .Y(n_277) );
AOI21xp5_ASAP7_75t_L g278 ( .A1(n_224), .A2(n_194), .B(n_181), .Y(n_278) );
O2A1O1Ixp33_ASAP7_75t_L g279 ( .A1(n_216), .A2(n_173), .B(n_170), .C(n_179), .Y(n_279) );
OAI22xp5_ASAP7_75t_SL g280 ( .A1(n_232), .A2(n_187), .B1(n_170), .B2(n_173), .Y(n_280) );
NAND2x1p5_ASAP7_75t_L g281 ( .A(n_242), .B(n_173), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_242), .Y(n_282) );
BUFx2_ASAP7_75t_L g283 ( .A(n_227), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_262), .B(n_173), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_212), .Y(n_285) );
AOI21xp33_ASAP7_75t_L g286 ( .A1(n_220), .A2(n_170), .B(n_179), .Y(n_286) );
AOI21xp5_ASAP7_75t_L g287 ( .A1(n_234), .A2(n_157), .B(n_177), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_217), .B(n_170), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_249), .Y(n_289) );
AOI21xp33_ASAP7_75t_L g290 ( .A1(n_240), .A2(n_157), .B(n_177), .Y(n_290) );
AOI22xp33_ASAP7_75t_SL g291 ( .A1(n_262), .A2(n_160), .B1(n_172), .B2(n_178), .Y(n_291) );
AND2x4_ASAP7_75t_L g292 ( .A(n_240), .B(n_172), .Y(n_292) );
AOI22x1_ASAP7_75t_L g293 ( .A1(n_257), .A2(n_203), .B1(n_202), .B2(n_189), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_241), .Y(n_294) );
INVx4_ASAP7_75t_L g295 ( .A(n_262), .Y(n_295) );
INVx4_ASAP7_75t_L g296 ( .A(n_212), .Y(n_296) );
BUFx3_ASAP7_75t_L g297 ( .A(n_251), .Y(n_297) );
INVx2_ASAP7_75t_L g298 ( .A(n_241), .Y(n_298) );
AOI221xp5_ASAP7_75t_L g299 ( .A1(n_223), .A2(n_160), .B1(n_202), .B2(n_189), .C(n_188), .Y(n_299) );
BUFx6f_ASAP7_75t_L g300 ( .A(n_251), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_235), .Y(n_301) );
BUFx6f_ASAP7_75t_L g302 ( .A(n_258), .Y(n_302) );
A2O1A1Ixp33_ASAP7_75t_L g303 ( .A1(n_236), .A2(n_203), .B(n_202), .C(n_189), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_237), .Y(n_304) );
BUFx6f_ASAP7_75t_L g305 ( .A(n_258), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_223), .B(n_51), .Y(n_306) );
O2A1O1Ixp5_ASAP7_75t_L g307 ( .A1(n_270), .A2(n_261), .B(n_255), .C(n_247), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_265), .A2(n_245), .B(n_254), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_263), .Y(n_309) );
OAI21xp5_ASAP7_75t_L g310 ( .A1(n_303), .A2(n_248), .B(n_247), .Y(n_310) );
INVx1_ASAP7_75t_SL g311 ( .A(n_283), .Y(n_311) );
AO31x2_ASAP7_75t_L g312 ( .A1(n_271), .A2(n_259), .A3(n_229), .B(n_246), .Y(n_312) );
AND2x2_ASAP7_75t_L g313 ( .A(n_268), .B(n_250), .Y(n_313) );
AOI221xp5_ASAP7_75t_L g314 ( .A1(n_276), .A2(n_225), .B1(n_209), .B2(n_226), .C(n_258), .Y(n_314) );
OAI21x1_ASAP7_75t_L g315 ( .A1(n_293), .A2(n_261), .B(n_252), .Y(n_315) );
OAI22xp33_ASAP7_75t_L g316 ( .A1(n_284), .A2(n_256), .B1(n_231), .B2(n_211), .Y(n_316) );
AND2x2_ASAP7_75t_L g317 ( .A(n_268), .B(n_208), .Y(n_317) );
AOI21x1_ASAP7_75t_L g318 ( .A1(n_270), .A2(n_164), .B(n_163), .Y(n_318) );
BUFx3_ASAP7_75t_L g319 ( .A(n_282), .Y(n_319) );
OAI21x1_ASAP7_75t_L g320 ( .A1(n_279), .A2(n_239), .B(n_228), .Y(n_320) );
NAND2x1p5_ASAP7_75t_L g321 ( .A(n_295), .B(n_244), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g322 ( .A(n_264), .B(n_214), .Y(n_322) );
CKINVDCx6p67_ASAP7_75t_R g323 ( .A(n_275), .Y(n_323) );
AOI22xp5_ASAP7_75t_L g324 ( .A1(n_284), .A2(n_215), .B1(n_244), .B2(n_253), .Y(n_324) );
BUFx3_ASAP7_75t_L g325 ( .A(n_282), .Y(n_325) );
BUFx6f_ASAP7_75t_L g326 ( .A(n_282), .Y(n_326) );
INVx6_ASAP7_75t_L g327 ( .A(n_302), .Y(n_327) );
OA21x2_ASAP7_75t_L g328 ( .A1(n_303), .A2(n_259), .B(n_184), .Y(n_328) );
AOI221xp5_ASAP7_75t_L g329 ( .A1(n_264), .A2(n_253), .B1(n_243), .B2(n_203), .C(n_188), .Y(n_329) );
AO21x2_ASAP7_75t_L g330 ( .A1(n_271), .A2(n_243), .B(n_188), .Y(n_330) );
NAND2xp5_ASAP7_75t_SL g331 ( .A(n_295), .B(n_178), .Y(n_331) );
AO21x1_ASAP7_75t_L g332 ( .A1(n_288), .A2(n_184), .B(n_182), .Y(n_332) );
NAND2xp5_ASAP7_75t_L g333 ( .A(n_301), .B(n_53), .Y(n_333) );
OAI21x1_ASAP7_75t_L g334 ( .A1(n_274), .A2(n_184), .B(n_182), .Y(n_334) );
AOI22xp33_ASAP7_75t_L g335 ( .A1(n_313), .A2(n_280), .B1(n_284), .B2(n_306), .Y(n_335) );
OAI21xp5_ASAP7_75t_L g336 ( .A1(n_314), .A2(n_291), .B(n_278), .Y(n_336) );
OAI21xp33_ASAP7_75t_L g337 ( .A1(n_311), .A2(n_291), .B(n_289), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_313), .B(n_309), .Y(n_339) );
AND2x4_ASAP7_75t_L g340 ( .A(n_317), .B(n_304), .Y(n_340) );
CKINVDCx12_ASAP7_75t_R g341 ( .A(n_323), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_317), .Y(n_342) );
OAI22xp33_ASAP7_75t_L g343 ( .A1(n_323), .A2(n_305), .B1(n_302), .B2(n_269), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_321), .B(n_302), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g345 ( .A1(n_322), .A2(n_290), .B1(n_302), .B2(n_305), .C(n_286), .Y(n_345) );
OAI21x1_ASAP7_75t_L g346 ( .A1(n_334), .A2(n_287), .B(n_277), .Y(n_346) );
AOI21xp5_ASAP7_75t_L g347 ( .A1(n_332), .A2(n_266), .B(n_273), .Y(n_347) );
INVx3_ASAP7_75t_L g348 ( .A(n_321), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g349 ( .A1(n_321), .A2(n_327), .B1(n_305), .B2(n_330), .Y(n_349) );
OAI22xp5_ASAP7_75t_L g350 ( .A1(n_316), .A2(n_281), .B1(n_305), .B2(n_296), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_334), .Y(n_351) );
A2O1A1Ixp33_ASAP7_75t_L g352 ( .A1(n_307), .A2(n_273), .B(n_298), .C(n_266), .Y(n_352) );
AOI221x1_ASAP7_75t_SL g353 ( .A1(n_333), .A2(n_292), .B1(n_298), .B2(n_294), .C(n_285), .Y(n_353) );
AOI22xp33_ASAP7_75t_L g354 ( .A1(n_330), .A2(n_327), .B1(n_310), .B2(n_292), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_327), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_327), .Y(n_356) );
AOI21xp5_ASAP7_75t_L g357 ( .A1(n_332), .A2(n_294), .B(n_299), .Y(n_357) );
OAI211xp5_ASAP7_75t_L g358 ( .A1(n_324), .A2(n_272), .B(n_267), .C(n_296), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_330), .B(n_272), .Y(n_359) );
OAI211xp5_ASAP7_75t_SL g360 ( .A1(n_337), .A2(n_331), .B(n_329), .C(n_267), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_338), .Y(n_361) );
INVx1_ASAP7_75t_L g362 ( .A(n_339), .Y(n_362) );
HB1xp67_ASAP7_75t_L g363 ( .A(n_344), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_347), .A2(n_318), .B(n_308), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_342), .B(n_312), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_339), .B(n_312), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_340), .Y(n_367) );
AND2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_312), .Y(n_368) );
INVx1_ASAP7_75t_SL g369 ( .A(n_348), .Y(n_369) );
BUFx2_ASAP7_75t_L g370 ( .A(n_359), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_340), .B(n_312), .Y(n_371) );
AND2x4_ASAP7_75t_L g372 ( .A(n_348), .B(n_326), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_335), .B(n_312), .Y(n_373) );
BUFx2_ASAP7_75t_L g374 ( .A(n_351), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_335), .B(n_325), .Y(n_375) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_354), .B(n_326), .Y(n_376) );
OR2x2_ASAP7_75t_L g377 ( .A(n_354), .B(n_325), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_352), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_352), .Y(n_379) );
HB1xp67_ASAP7_75t_L g380 ( .A(n_341), .Y(n_380) );
AND2x2_ASAP7_75t_L g381 ( .A(n_355), .B(n_319), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_356), .B(n_319), .Y(n_382) );
NAND2xp33_ASAP7_75t_R g383 ( .A(n_343), .B(n_328), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g384 ( .A(n_353), .B(n_326), .Y(n_384) );
BUFx2_ASAP7_75t_L g385 ( .A(n_351), .Y(n_385) );
INVxp67_ASAP7_75t_L g386 ( .A(n_343), .Y(n_386) );
HB1xp67_ASAP7_75t_L g387 ( .A(n_350), .Y(n_387) );
INVx2_ASAP7_75t_SL g388 ( .A(n_346), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
HB1xp67_ASAP7_75t_L g390 ( .A(n_358), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_349), .Y(n_391) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_363), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_368), .Y(n_393) );
INVx1_ASAP7_75t_L g394 ( .A(n_368), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_371), .B(n_336), .Y(n_395) );
INVx2_ASAP7_75t_L g396 ( .A(n_374), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_365), .B(n_357), .Y(n_397) );
AND2x2_ASAP7_75t_L g398 ( .A(n_371), .B(n_328), .Y(n_398) );
AND2x2_ASAP7_75t_L g399 ( .A(n_366), .B(n_328), .Y(n_399) );
INVxp67_ASAP7_75t_SL g400 ( .A(n_370), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_365), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_361), .B(n_326), .Y(n_402) );
NOR2xp33_ASAP7_75t_L g403 ( .A(n_380), .B(n_300), .Y(n_403) );
INVx1_ASAP7_75t_SL g404 ( .A(n_369), .Y(n_404) );
NOR2x1_ASAP7_75t_R g405 ( .A(n_370), .B(n_326), .Y(n_405) );
NOR3xp33_ASAP7_75t_SL g406 ( .A(n_383), .B(n_55), .C(n_56), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_366), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_361), .Y(n_408) );
AND2x2_ASAP7_75t_L g409 ( .A(n_373), .B(n_318), .Y(n_409) );
OR2x2_ASAP7_75t_SL g410 ( .A(n_384), .B(n_282), .Y(n_410) );
AND2x2_ASAP7_75t_L g411 ( .A(n_373), .B(n_308), .Y(n_411) );
INVx4_ASAP7_75t_L g412 ( .A(n_372), .Y(n_412) );
INVx5_ASAP7_75t_L g413 ( .A(n_372), .Y(n_413) );
AND2x2_ASAP7_75t_L g414 ( .A(n_367), .B(n_320), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_367), .B(n_320), .Y(n_415) );
BUFx2_ASAP7_75t_SL g416 ( .A(n_369), .Y(n_416) );
INVxp67_ASAP7_75t_SL g417 ( .A(n_374), .Y(n_417) );
OR2x2_ASAP7_75t_L g418 ( .A(n_391), .B(n_281), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_385), .Y(n_419) );
INVx2_ASAP7_75t_L g420 ( .A(n_385), .Y(n_420) );
AND2x2_ASAP7_75t_L g421 ( .A(n_375), .B(n_315), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_388), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_388), .Y(n_423) );
AO21x2_ASAP7_75t_L g424 ( .A1(n_384), .A2(n_315), .B(n_163), .Y(n_424) );
INVx2_ASAP7_75t_L g425 ( .A(n_364), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_375), .B(n_57), .Y(n_426) );
AOI22xp33_ASAP7_75t_L g427 ( .A1(n_386), .A2(n_300), .B1(n_297), .B2(n_178), .Y(n_427) );
OAI22xp5_ASAP7_75t_SL g428 ( .A1(n_390), .A2(n_300), .B1(n_297), .B2(n_63), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_362), .B(n_58), .Y(n_429) );
NAND3xp33_ASAP7_75t_L g430 ( .A(n_391), .B(n_300), .C(n_178), .Y(n_430) );
OAI21xp5_ASAP7_75t_L g431 ( .A1(n_389), .A2(n_182), .B(n_167), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_362), .B(n_60), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_377), .Y(n_433) );
INVx2_ASAP7_75t_SL g434 ( .A(n_372), .Y(n_434) );
AND2x4_ASAP7_75t_L g435 ( .A(n_377), .B(n_65), .Y(n_435) );
INVx2_ASAP7_75t_L g436 ( .A(n_364), .Y(n_436) );
INVxp67_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_376), .Y(n_438) );
HB1xp67_ASAP7_75t_L g439 ( .A(n_392), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_422), .Y(n_440) );
AND2x4_ASAP7_75t_L g441 ( .A(n_393), .B(n_376), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_422), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_408), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_394), .B(n_379), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_394), .B(n_379), .Y(n_445) );
OAI21xp33_ASAP7_75t_SL g446 ( .A1(n_400), .A2(n_389), .B(n_382), .Y(n_446) );
AND2x2_ASAP7_75t_L g447 ( .A(n_407), .B(n_378), .Y(n_447) );
AND2x2_ASAP7_75t_L g448 ( .A(n_407), .B(n_378), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_428), .B(n_389), .Y(n_449) );
INVx2_ASAP7_75t_SL g450 ( .A(n_413), .Y(n_450) );
NOR2xp33_ASAP7_75t_L g451 ( .A(n_403), .B(n_382), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_399), .B(n_381), .Y(n_452) );
INVx1_ASAP7_75t_L g453 ( .A(n_408), .Y(n_453) );
NAND2xp33_ASAP7_75t_L g454 ( .A(n_428), .B(n_381), .Y(n_454) );
OAI31xp33_ASAP7_75t_L g455 ( .A1(n_435), .A2(n_360), .A3(n_372), .B(n_69), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_399), .B(n_67), .Y(n_456) );
OR2x2_ASAP7_75t_L g457 ( .A(n_433), .B(n_68), .Y(n_457) );
OAI221xp5_ASAP7_75t_L g458 ( .A1(n_437), .A2(n_360), .B1(n_163), .B2(n_164), .C(n_167), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_401), .B(n_70), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_422), .Y(n_460) );
HB1xp67_ASAP7_75t_L g461 ( .A(n_404), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_401), .B(n_71), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_402), .Y(n_463) );
NOR2x1_ASAP7_75t_L g464 ( .A(n_430), .B(n_164), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_395), .B(n_167), .Y(n_465) );
INVx2_ASAP7_75t_SL g466 ( .A(n_413), .Y(n_466) );
BUFx2_ASAP7_75t_L g467 ( .A(n_405), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_395), .B(n_178), .Y(n_468) );
NAND2xp5_ASAP7_75t_L g469 ( .A(n_433), .B(n_178), .Y(n_469) );
AND2x2_ASAP7_75t_L g470 ( .A(n_398), .B(n_178), .Y(n_470) );
INVx2_ASAP7_75t_L g471 ( .A(n_423), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_402), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_437), .B(n_398), .Y(n_473) );
AND2x4_ASAP7_75t_L g474 ( .A(n_412), .B(n_421), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_421), .B(n_414), .Y(n_475) );
INVx1_ASAP7_75t_SL g476 ( .A(n_416), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_414), .B(n_411), .Y(n_477) );
INVxp67_ASAP7_75t_SL g478 ( .A(n_405), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_411), .B(n_396), .Y(n_479) );
BUFx3_ASAP7_75t_L g480 ( .A(n_413), .Y(n_480) );
INVx2_ASAP7_75t_L g481 ( .A(n_423), .Y(n_481) );
NAND2x1p5_ASAP7_75t_L g482 ( .A(n_435), .B(n_413), .Y(n_482) );
NOR2xp67_ASAP7_75t_L g483 ( .A(n_430), .B(n_413), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_423), .Y(n_484) );
INVx1_ASAP7_75t_L g485 ( .A(n_419), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_396), .B(n_420), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_396), .B(n_420), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_419), .Y(n_488) );
NAND2xp5_ASAP7_75t_L g489 ( .A(n_426), .B(n_404), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_426), .B(n_397), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_397), .B(n_418), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_463), .B(n_409), .Y(n_492) );
XOR2xp5_ASAP7_75t_L g493 ( .A(n_452), .B(n_435), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_473), .B(n_417), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_463), .B(n_409), .Y(n_495) );
AND2x2_ASAP7_75t_L g496 ( .A(n_452), .B(n_412), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_477), .B(n_475), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_439), .Y(n_498) );
INVx2_ASAP7_75t_L g499 ( .A(n_486), .Y(n_499) );
INVx1_ASAP7_75t_L g500 ( .A(n_443), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_443), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_453), .Y(n_502) );
AND2x2_ASAP7_75t_L g503 ( .A(n_477), .B(n_412), .Y(n_503) );
OR2x2_ASAP7_75t_L g504 ( .A(n_491), .B(n_420), .Y(n_504) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_472), .B(n_415), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_453), .Y(n_506) );
INVx2_ASAP7_75t_L g507 ( .A(n_486), .Y(n_507) );
NAND3xp33_ASAP7_75t_SL g508 ( .A(n_455), .B(n_406), .C(n_429), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_475), .B(n_412), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_472), .B(n_415), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_485), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_476), .Y(n_512) );
AND2x2_ASAP7_75t_L g513 ( .A(n_479), .B(n_434), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_485), .B(n_434), .Y(n_514) );
AO21x1_ASAP7_75t_L g515 ( .A1(n_454), .A2(n_435), .B(n_418), .Y(n_515) );
AND2x4_ASAP7_75t_L g516 ( .A(n_474), .B(n_413), .Y(n_516) );
INVx1_ASAP7_75t_L g517 ( .A(n_488), .Y(n_517) );
OR2x6_ASAP7_75t_L g518 ( .A(n_482), .B(n_416), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_488), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_479), .B(n_413), .Y(n_520) );
OR2x2_ASAP7_75t_L g521 ( .A(n_490), .B(n_410), .Y(n_521) );
INVx1_ASAP7_75t_L g522 ( .A(n_461), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_487), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_474), .B(n_424), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_487), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_444), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_444), .B(n_424), .Y(n_527) );
NAND2xp5_ASAP7_75t_L g528 ( .A(n_445), .B(n_424), .Y(n_528) );
INVx1_ASAP7_75t_L g529 ( .A(n_445), .Y(n_529) );
OR2x2_ASAP7_75t_L g530 ( .A(n_438), .B(n_410), .Y(n_530) );
OAI21xp33_ASAP7_75t_L g531 ( .A1(n_446), .A2(n_427), .B(n_429), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_474), .B(n_424), .Y(n_532) );
NOR2x1_ASAP7_75t_L g533 ( .A(n_467), .B(n_432), .Y(n_533) );
OR2x2_ASAP7_75t_L g534 ( .A(n_438), .B(n_425), .Y(n_534) );
INVx2_ASAP7_75t_L g535 ( .A(n_440), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_474), .B(n_432), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_447), .B(n_425), .Y(n_537) );
OR2x2_ASAP7_75t_L g538 ( .A(n_489), .B(n_425), .Y(n_538) );
NAND2xp5_ASAP7_75t_L g539 ( .A(n_447), .B(n_436), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g540 ( .A(n_449), .B(n_431), .Y(n_540) );
NOR3xp33_ASAP7_75t_SL g541 ( .A(n_508), .B(n_455), .C(n_446), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_526), .B(n_448), .Y(n_542) );
AOI32xp33_ASAP7_75t_L g543 ( .A1(n_533), .A2(n_467), .A3(n_476), .B1(n_478), .B2(n_456), .Y(n_543) );
AOI22xp5_ASAP7_75t_L g544 ( .A1(n_515), .A2(n_451), .B1(n_482), .B2(n_441), .Y(n_544) );
INVx2_ASAP7_75t_L g545 ( .A(n_535), .Y(n_545) );
INVx1_ASAP7_75t_SL g546 ( .A(n_512), .Y(n_546) );
OR2x6_ASAP7_75t_L g547 ( .A(n_518), .B(n_482), .Y(n_547) );
XNOR2x2_ASAP7_75t_L g548 ( .A(n_498), .B(n_457), .Y(n_548) );
AOI31xp33_ASAP7_75t_L g549 ( .A1(n_508), .A2(n_450), .A3(n_466), .B(n_457), .Y(n_549) );
OAI21xp33_ASAP7_75t_L g550 ( .A1(n_530), .A2(n_441), .B(n_448), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_529), .B(n_441), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_497), .B(n_441), .Y(n_552) );
AOI322xp5_ASAP7_75t_L g553 ( .A1(n_540), .A2(n_456), .A3(n_450), .B1(n_466), .B2(n_459), .C1(n_465), .C2(n_480), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_509), .B(n_480), .Y(n_554) );
OAI32xp33_ASAP7_75t_L g555 ( .A1(n_521), .A2(n_480), .A3(n_459), .B1(n_462), .B2(n_468), .Y(n_555) );
AO21x1_ASAP7_75t_L g556 ( .A1(n_540), .A2(n_484), .B(n_471), .Y(n_556) );
OAI22xp33_ASAP7_75t_L g557 ( .A1(n_518), .A2(n_483), .B1(n_464), .B2(n_440), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_516), .B(n_483), .Y(n_558) );
XNOR2xp5_ASAP7_75t_L g559 ( .A(n_493), .B(n_470), .Y(n_559) );
INVx1_ASAP7_75t_SL g560 ( .A(n_496), .Y(n_560) );
INVx2_ASAP7_75t_L g561 ( .A(n_535), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_518), .A2(n_464), .B(n_469), .Y(n_562) );
NAND2xp5_ASAP7_75t_L g563 ( .A(n_522), .B(n_460), .Y(n_563) );
OAI21xp5_ASAP7_75t_SL g564 ( .A1(n_531), .A2(n_470), .B(n_458), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g565 ( .A1(n_516), .A2(n_460), .B1(n_481), .B2(n_440), .Y(n_565) );
OAI22xp33_ASAP7_75t_L g566 ( .A1(n_494), .A2(n_442), .B1(n_460), .B2(n_471), .Y(n_566) );
AOI211xp5_ASAP7_75t_L g567 ( .A1(n_524), .A2(n_442), .B(n_471), .C(n_481), .Y(n_567) );
NOR2xp33_ASAP7_75t_L g568 ( .A(n_503), .B(n_442), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_511), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_517), .Y(n_570) );
NOR2xp33_ASAP7_75t_L g571 ( .A(n_523), .B(n_481), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_519), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_504), .B(n_484), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_538), .Y(n_574) );
INVxp67_ASAP7_75t_SL g575 ( .A(n_556), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_545), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_574), .B(n_525), .Y(n_577) );
INVx1_ASAP7_75t_L g578 ( .A(n_551), .Y(n_578) );
INVx1_ASAP7_75t_L g579 ( .A(n_569), .Y(n_579) );
AND2x2_ASAP7_75t_L g580 ( .A(n_560), .B(n_513), .Y(n_580) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_550), .A2(n_532), .B1(n_536), .B2(n_520), .Y(n_581) );
XNOR2xp5_ASAP7_75t_L g582 ( .A(n_559), .B(n_507), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_570), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_572), .Y(n_584) );
AOI21xp33_ASAP7_75t_SL g585 ( .A1(n_549), .A2(n_514), .B(n_492), .Y(n_585) );
A2O1A1Ixp33_ASAP7_75t_L g586 ( .A1(n_543), .A2(n_499), .B(n_514), .C(n_492), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_563), .Y(n_587) );
AND3x1_ASAP7_75t_L g588 ( .A(n_541), .B(n_495), .C(n_527), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_573), .B(n_542), .Y(n_589) );
NAND2xp5_ASAP7_75t_L g590 ( .A(n_571), .B(n_528), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_566), .B(n_528), .Y(n_591) );
AOI22xp5_ASAP7_75t_L g592 ( .A1(n_544), .A2(n_495), .B1(n_527), .B2(n_537), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_552), .Y(n_593) );
INVx2_ASAP7_75t_L g594 ( .A(n_561), .Y(n_594) );
INVx2_ASAP7_75t_L g595 ( .A(n_547), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g596 ( .A(n_587), .B(n_502), .Y(n_596) );
AOI221x1_ASAP7_75t_L g597 ( .A1(n_586), .A2(n_558), .B1(n_565), .B2(n_562), .C(n_568), .Y(n_597) );
AOI322xp5_ASAP7_75t_L g598 ( .A1(n_575), .A2(n_546), .A3(n_544), .B1(n_554), .B2(n_558), .C1(n_557), .C2(n_548), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_586), .A2(n_564), .B(n_553), .Y(n_599) );
OAI211xp5_ASAP7_75t_SL g600 ( .A1(n_575), .A2(n_567), .B(n_510), .C(n_505), .Y(n_600) );
INVxp67_ASAP7_75t_L g601 ( .A(n_588), .Y(n_601) );
INVx2_ASAP7_75t_L g602 ( .A(n_576), .Y(n_602) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_595), .A2(n_547), .B1(n_534), .B2(n_537), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_589), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_579), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_576), .Y(n_606) );
AOI222xp33_ASAP7_75t_L g607 ( .A1(n_591), .A2(n_582), .B1(n_595), .B2(n_578), .C1(n_577), .C2(n_590), .Y(n_607) );
INVx1_ASAP7_75t_L g608 ( .A(n_596), .Y(n_608) );
OAI21xp33_ASAP7_75t_L g609 ( .A1(n_598), .A2(n_592), .B(n_585), .Y(n_609) );
AOI21xp5_ASAP7_75t_L g610 ( .A1(n_599), .A2(n_597), .B(n_601), .Y(n_610) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_604), .B(n_584), .Y(n_611) );
AOI22xp5_ASAP7_75t_L g612 ( .A1(n_607), .A2(n_581), .B1(n_583), .B2(n_547), .Y(n_612) );
AOI211xp5_ASAP7_75t_L g613 ( .A1(n_600), .A2(n_555), .B(n_580), .C(n_593), .Y(n_613) );
AOI222xp33_ASAP7_75t_L g614 ( .A1(n_600), .A2(n_594), .B1(n_506), .B2(n_501), .C1(n_500), .C2(n_505), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_610), .B(n_605), .Y(n_615) );
OAI22xp5_ASAP7_75t_L g616 ( .A1(n_612), .A2(n_603), .B1(n_606), .B2(n_602), .Y(n_616) );
AOI221xp5_ASAP7_75t_L g617 ( .A1(n_609), .A2(n_596), .B1(n_594), .B2(n_510), .C(n_539), .Y(n_617) );
NOR2xp33_ASAP7_75t_R g618 ( .A(n_611), .B(n_539), .Y(n_618) );
NOR2x1p5_ASAP7_75t_L g619 ( .A(n_615), .B(n_608), .Y(n_619) );
AOI221xp5_ASAP7_75t_L g620 ( .A1(n_617), .A2(n_613), .B1(n_614), .B2(n_484), .C(n_431), .Y(n_620) );
BUFx2_ASAP7_75t_L g621 ( .A(n_619), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_620), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_621), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_623), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_624), .A2(n_622), .B1(n_621), .B2(n_616), .Y(n_625) );
XNOR2xp5_ASAP7_75t_L g626 ( .A(n_625), .B(n_618), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_626), .A2(n_436), .B(n_623), .Y(n_627) );
endmodule