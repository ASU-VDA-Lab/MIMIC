module fake_netlist_6_3342_n_1990 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_184, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_174, n_127, n_125, n_153, n_168, n_178, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_188, n_102, n_186, n_0, n_87, n_189, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_180, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_172, n_81, n_59, n_181, n_76, n_36, n_182, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_175, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_177, n_176, n_114, n_86, n_104, n_95, n_179, n_9, n_107, n_10, n_71, n_74, n_6, n_190, n_14, n_123, n_136, n_72, n_187, n_89, n_173, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_185, n_35, n_183, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_1990);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_184;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_174;
input n_127;
input n_125;
input n_153;
input n_168;
input n_178;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_188;
input n_102;
input n_186;
input n_0;
input n_87;
input n_189;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_180;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_172;
input n_81;
input n_59;
input n_181;
input n_76;
input n_36;
input n_182;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_175;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_177;
input n_176;
input n_114;
input n_86;
input n_104;
input n_95;
input n_179;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_190;
input n_14;
input n_123;
input n_136;
input n_72;
input n_187;
input n_89;
input n_173;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_185;
input n_35;
input n_183;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1990;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_1853;
wire n_783;
wire n_1738;
wire n_798;
wire n_1575;
wire n_1854;
wire n_1923;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_1708;
wire n_805;
wire n_1151;
wire n_396;
wire n_1739;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1691;
wire n_1688;
wire n_1975;
wire n_1009;
wire n_1743;
wire n_1930;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1724;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_1844;
wire n_424;
wire n_1700;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_1786;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_1985;
wire n_447;
wire n_1803;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1867;
wire n_1704;
wire n_1078;
wire n_544;
wire n_250;
wire n_1711;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1903;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1772;
wire n_1572;
wire n_616;
wire n_658;
wire n_1874;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1902;
wire n_1842;
wire n_1620;
wire n_1954;
wire n_1735;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1798;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_1781;
wire n_1971;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_1820;
wire n_494;
wire n_539;
wire n_493;
wire n_454;
wire n_1421;
wire n_1936;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1961;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1526;
wire n_1560;
wire n_734;
wire n_1088;
wire n_1894;
wire n_196;
wire n_1231;
wire n_1978;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_1815;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1967;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_1911;
wire n_1956;
wire n_1644;
wire n_1558;
wire n_1732;
wire n_281;
wire n_551;
wire n_699;
wire n_1986;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_1918;
wire n_577;
wire n_1843;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1909;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_1699;
wire n_916;
wire n_483;
wire n_1970;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_1957;
wire n_219;
wire n_1907;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1762;
wire n_1910;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_1876;
wire n_1895;
wire n_1697;
wire n_243;
wire n_979;
wire n_1873;
wire n_905;
wire n_1866;
wire n_1680;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1988;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1793;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_1703;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_1865;
wire n_1875;
wire n_1701;
wire n_318;
wire n_1111;
wire n_1713;
wire n_715;
wire n_1251;
wire n_1265;
wire n_1726;
wire n_1950;
wire n_530;
wire n_1563;
wire n_1912;
wire n_277;
wire n_1982;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_1760;
wire n_1927;
wire n_210;
wire n_1069;
wire n_1722;
wire n_1664;
wire n_612;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1926;
wire n_1175;
wire n_328;
wire n_1386;
wire n_1896;
wire n_429;
wire n_1747;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1977;
wire n_1802;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_835;
wire n_242;
wire n_928;
wire n_1214;
wire n_850;
wire n_690;
wire n_1801;
wire n_1886;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1750;
wire n_1462;
wire n_1188;
wire n_1752;
wire n_877;
wire n_1813;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_1965;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_697;
wire n_687;
wire n_890;
wire n_637;
wire n_701;
wire n_295;
wire n_950;
wire n_388;
wire n_484;
wire n_1709;
wire n_1825;
wire n_1796;
wire n_1757;
wire n_1792;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_1987;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_1033;
wire n_462;
wire n_1052;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_595;
wire n_297;
wire n_627;
wire n_1767;
wire n_1779;
wire n_524;
wire n_1465;
wire n_342;
wire n_1858;
wire n_1044;
wire n_1712;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1756;
wire n_1128;
wire n_382;
wire n_673;
wire n_1969;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_1968;
wire n_898;
wire n_255;
wire n_284;
wire n_1952;
wire n_865;
wire n_925;
wire n_1932;
wire n_1101;
wire n_1026;
wire n_1880;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_1839;
wire n_685;
wire n_1765;
wire n_353;
wire n_605;
wire n_1514;
wire n_1863;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_1714;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_1913;
wire n_510;
wire n_837;
wire n_1488;
wire n_1808;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_1947;
wire n_536;
wire n_1788;
wire n_622;
wire n_1469;
wire n_1838;
wire n_1835;
wire n_1776;
wire n_1766;
wire n_1959;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_1771;
wire n_631;
wire n_720;
wire n_842;
wire n_1707;
wire n_1432;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1723;
wire n_1246;
wire n_1878;
wire n_899;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1809;
wire n_1577;
wire n_1181;
wire n_1822;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_1717;
wire n_926;
wire n_1817;
wire n_927;
wire n_1849;
wire n_919;
wire n_1698;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_552;
wire n_1358;
wire n_1811;
wire n_1388;
wire n_216;
wire n_912;
wire n_1857;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1774;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_1955;
wire n_755;
wire n_1021;
wire n_931;
wire n_527;
wire n_474;
wire n_811;
wire n_683;
wire n_1207;
wire n_312;
wire n_1791;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_1897;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_1942;
wire n_1966;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_1837;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_1736;
wire n_211;
wire n_1483;
wire n_1834;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_1719;
wire n_319;
wire n_1339;
wire n_1787;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1919;
wire n_1080;
wire n_723;
wire n_1877;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1939;
wire n_1769;
wire n_1220;
wire n_1893;
wire n_556;
wire n_1755;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_1980;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_1951;
wire n_444;
wire n_1252;
wire n_1784;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1773;
wire n_1775;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1783;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_1745;
wire n_914;
wire n_759;
wire n_1831;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_1901;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1892;
wire n_1933;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1917;
wire n_1580;
wire n_1425;
wire n_1881;
wire n_1281;
wire n_1267;
wire n_1806;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1733;
wire n_1419;
wire n_351;
wire n_259;
wire n_1731;
wire n_1855;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_1832;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_736;
wire n_613;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1696;
wire n_1594;
wire n_664;
wire n_1869;
wire n_1764;
wire n_1429;
wire n_1610;
wire n_1889;
wire n_435;
wire n_1905;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_1937;
wire n_465;
wire n_1790;
wire n_1778;
wire n_1635;
wire n_1079;
wire n_341;
wire n_1744;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1934;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_1728;
wire n_557;
wire n_1871;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_1859;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1718;
wire n_1749;
wire n_1683;
wire n_1916;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1852;
wire n_1024;
wire n_1768;
wire n_198;
wire n_1847;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1841;
wire n_1639;
wire n_1623;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1818;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1960;
wire n_1686;
wire n_1356;
wire n_1589;
wire n_1740;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1943;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_1694;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_1734;
wire n_397;
wire n_1983;
wire n_1938;
wire n_1262;
wire n_218;
wire n_1891;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_1715;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1797;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_1870;
wire n_352;
wire n_1692;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1827;
wire n_1361;
wire n_1864;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_1840;
wire n_1705;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_1695;
wire n_1828;
wire n_650;
wire n_1046;
wire n_1940;
wire n_1979;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_1963;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1883;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_1823;
wire n_227;
wire n_1974;
wire n_1720;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_1795;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1845;
wire n_1489;
wire n_942;
wire n_1524;
wire n_543;
wire n_1964;
wire n_1920;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1946;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_1846;
wire n_533;
wire n_806;
wire n_959;
wire n_879;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_1782;
wire n_282;
wire n_1676;
wire n_833;
wire n_1830;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_1900;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_1086;
wire n_1066;
wire n_1948;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1906;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_1758;
wire n_1925;
wire n_737;
wire n_1318;
wire n_1914;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1706;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1984;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_1931;
wire n_502;
wire n_672;
wire n_1257;
wire n_1751;
wire n_285;
wire n_1375;
wire n_1941;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1794;
wire n_1236;
wire n_1962;
wire n_1559;
wire n_1725;
wire n_1928;
wire n_1872;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1746;
wire n_1325;
wire n_1002;
wire n_1741;
wire n_1949;
wire n_545;
wire n_489;
wire n_1804;
wire n_1727;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1860;
wire n_1904;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1777;
wire n_1908;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1800;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1742;
wire n_1562;
wire n_1690;
wire n_398;
wire n_1191;
wire n_1826;
wire n_566;
wire n_1023;
wire n_1882;
wire n_1076;
wire n_1118;
wire n_194;
wire n_1007;
wire n_1807;
wire n_1929;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1759;
wire n_1814;
wire n_1631;
wire n_591;
wire n_1377;
wire n_1879;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_680;
wire n_367;
wire n_1678;
wire n_661;
wire n_1716;
wire n_278;
wire n_1256;
wire n_671;
wire n_1953;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1976;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_1824;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_1810;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_1730;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_1729;
wire n_669;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_1785;
wire n_763;
wire n_1147;
wire n_1848;
wire n_360;
wire n_1754;
wire n_1506;
wire n_1652;
wire n_1812;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_1173;
wire n_1924;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1702;
wire n_1219;
wire n_1780;
wire n_1689;
wire n_1174;
wire n_1944;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_1945;
wire n_910;
wire n_1656;
wire n_1721;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1737;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_1922;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_1973;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1821;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1693;
wire n_1109;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1989;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1972;
wire n_1525;
wire n_455;
wire n_1585;
wire n_1851;
wire n_363;
wire n_1799;
wire n_1090;
wire n_592;
wire n_1816;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_1829;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_1789;
wire n_1770;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1710;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1763;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1981;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_1753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1921;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_404;
wire n_271;
wire n_1884;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1819;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_1761;
wire n_534;
wire n_1578;
wire n_1006;
wire n_1861;
wire n_373;
wire n_1632;
wire n_1890;
wire n_1805;
wire n_257;
wire n_1557;
wire n_1888;
wire n_1833;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_1850;
wire n_1898;
wire n_1868;
wire n_207;
wire n_1089;
wire n_1887;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_1836;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1899;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_1862;
wire n_1856;
wire n_1958;
wire n_339;
wire n_784;
wire n_434;
wire n_315;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_540;
wire n_1423;
wire n_1935;
wire n_457;
wire n_364;
wire n_1915;
wire n_629;
wire n_1621;
wire n_1748;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1885;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_43),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_135),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_78),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_141),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_27),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_162),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_109),
.Y(n_198)
);

CKINVDCx5p33_ASAP7_75t_R g199 ( 
.A(n_41),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_174),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_163),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_85),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_56),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_63),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_29),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_175),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_149),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_43),
.Y(n_208)
);

INVx2_ASAP7_75t_SL g209 ( 
.A(n_144),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_123),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g211 ( 
.A(n_10),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_24),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_131),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_8),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_36),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_103),
.Y(n_216)
);

BUFx2_ASAP7_75t_SL g217 ( 
.A(n_1),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_158),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_190),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_26),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_186),
.Y(n_221)
);

INVx2_ASAP7_75t_SL g222 ( 
.A(n_56),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_112),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_22),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_5),
.Y(n_225)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_117),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_127),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_148),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_164),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_36),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_42),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_73),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_81),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_53),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_65),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_21),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_24),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_6),
.Y(n_239)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_47),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_132),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_53),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_178),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_166),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_108),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_44),
.Y(n_246)
);

INVx1_ASAP7_75t_SL g247 ( 
.A(n_45),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_70),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_84),
.Y(n_249)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_62),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_114),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_69),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_40),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_104),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_59),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_179),
.Y(n_256)
);

INVx3_ASAP7_75t_L g257 ( 
.A(n_68),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_87),
.Y(n_258)
);

BUFx3_ASAP7_75t_L g259 ( 
.A(n_20),
.Y(n_259)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_75),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_136),
.Y(n_261)
);

INVx1_ASAP7_75t_SL g262 ( 
.A(n_67),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_159),
.Y(n_263)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_110),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_33),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_169),
.Y(n_266)
);

CKINVDCx20_ASAP7_75t_R g267 ( 
.A(n_101),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_57),
.Y(n_268)
);

CKINVDCx14_ASAP7_75t_R g269 ( 
.A(n_26),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_115),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_95),
.Y(n_271)
);

INVx2_ASAP7_75t_SL g272 ( 
.A(n_122),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_142),
.Y(n_273)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_155),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_35),
.Y(n_275)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_146),
.Y(n_276)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_137),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_88),
.Y(n_278)
);

BUFx5_ASAP7_75t_L g279 ( 
.A(n_98),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_40),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_29),
.Y(n_281)
);

BUFx3_ASAP7_75t_L g282 ( 
.A(n_106),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_167),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_57),
.Y(n_284)
);

BUFx3_ASAP7_75t_L g285 ( 
.A(n_89),
.Y(n_285)
);

BUFx2_ASAP7_75t_L g286 ( 
.A(n_156),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_42),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_187),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_44),
.Y(n_289)
);

CKINVDCx5p33_ASAP7_75t_R g290 ( 
.A(n_27),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_143),
.Y(n_291)
);

HB1xp67_ASAP7_75t_L g292 ( 
.A(n_49),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_176),
.Y(n_293)
);

INVx2_ASAP7_75t_SL g294 ( 
.A(n_37),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_22),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_41),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_71),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_10),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g299 ( 
.A(n_5),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g300 ( 
.A(n_82),
.Y(n_300)
);

CKINVDCx5p33_ASAP7_75t_R g301 ( 
.A(n_76),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_184),
.Y(n_302)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_86),
.Y(n_303)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_66),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_180),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_3),
.Y(n_306)
);

BUFx3_ASAP7_75t_L g307 ( 
.A(n_151),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_74),
.Y(n_308)
);

CKINVDCx5p33_ASAP7_75t_R g309 ( 
.A(n_128),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_116),
.Y(n_310)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_147),
.Y(n_311)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_102),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_12),
.Y(n_313)
);

BUFx3_ASAP7_75t_L g314 ( 
.A(n_34),
.Y(n_314)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_182),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_7),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_17),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_14),
.Y(n_318)
);

BUFx6f_ASAP7_75t_L g319 ( 
.A(n_52),
.Y(n_319)
);

INVx3_ASAP7_75t_L g320 ( 
.A(n_48),
.Y(n_320)
);

INVx1_ASAP7_75t_L g321 ( 
.A(n_47),
.Y(n_321)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_97),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_50),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_12),
.Y(n_324)
);

CKINVDCx5p33_ASAP7_75t_R g325 ( 
.A(n_55),
.Y(n_325)
);

INVx2_ASAP7_75t_SL g326 ( 
.A(n_119),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_34),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_99),
.Y(n_328)
);

CKINVDCx5p33_ASAP7_75t_R g329 ( 
.A(n_124),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_48),
.Y(n_330)
);

CKINVDCx20_ASAP7_75t_R g331 ( 
.A(n_90),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_130),
.Y(n_332)
);

INVxp67_ASAP7_75t_SL g333 ( 
.A(n_125),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_31),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g335 ( 
.A(n_173),
.Y(n_335)
);

BUFx3_ASAP7_75t_L g336 ( 
.A(n_18),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_96),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_37),
.Y(n_338)
);

CKINVDCx5p33_ASAP7_75t_R g339 ( 
.A(n_80),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_31),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_79),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_9),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_54),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_55),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_171),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_8),
.Y(n_346)
);

INVx1_ASAP7_75t_SL g347 ( 
.A(n_35),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_172),
.Y(n_348)
);

INVx2_ASAP7_75t_L g349 ( 
.A(n_64),
.Y(n_349)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_185),
.Y(n_350)
);

CKINVDCx5p33_ASAP7_75t_R g351 ( 
.A(n_39),
.Y(n_351)
);

CKINVDCx5p33_ASAP7_75t_R g352 ( 
.A(n_107),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_181),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_168),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_72),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_18),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_33),
.Y(n_357)
);

CKINVDCx20_ASAP7_75t_R g358 ( 
.A(n_11),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_45),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_54),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_7),
.Y(n_361)
);

BUFx3_ASAP7_75t_L g362 ( 
.A(n_61),
.Y(n_362)
);

CKINVDCx5p33_ASAP7_75t_R g363 ( 
.A(n_152),
.Y(n_363)
);

INVx2_ASAP7_75t_SL g364 ( 
.A(n_25),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_58),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_16),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_145),
.Y(n_367)
);

BUFx8_ASAP7_75t_SL g368 ( 
.A(n_9),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_189),
.Y(n_369)
);

CKINVDCx20_ASAP7_75t_R g370 ( 
.A(n_51),
.Y(n_370)
);

INVx1_ASAP7_75t_SL g371 ( 
.A(n_120),
.Y(n_371)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_17),
.Y(n_372)
);

INVx1_ASAP7_75t_SL g373 ( 
.A(n_111),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_1),
.Y(n_374)
);

CKINVDCx20_ASAP7_75t_R g375 ( 
.A(n_92),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_93),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_49),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_118),
.Y(n_378)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_183),
.Y(n_379)
);

CKINVDCx5p33_ASAP7_75t_R g380 ( 
.A(n_38),
.Y(n_380)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_280),
.Y(n_381)
);

INVx3_ASAP7_75t_L g382 ( 
.A(n_280),
.Y(n_382)
);

CKINVDCx5p33_ASAP7_75t_R g383 ( 
.A(n_368),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_280),
.Y(n_384)
);

INVx1_ASAP7_75t_SL g385 ( 
.A(n_211),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_286),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_280),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_280),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_319),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_319),
.Y(n_390)
);

INVxp67_ASAP7_75t_L g391 ( 
.A(n_292),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_319),
.Y(n_392)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_319),
.Y(n_393)
);

CKINVDCx16_ASAP7_75t_R g394 ( 
.A(n_240),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_269),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g396 ( 
.A(n_198),
.Y(n_396)
);

INVxp67_ASAP7_75t_L g397 ( 
.A(n_217),
.Y(n_397)
);

INVxp67_ASAP7_75t_SL g398 ( 
.A(n_320),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_319),
.Y(n_399)
);

CKINVDCx20_ASAP7_75t_R g400 ( 
.A(n_221),
.Y(n_400)
);

INVxp67_ASAP7_75t_L g401 ( 
.A(n_205),
.Y(n_401)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_320),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_226),
.Y(n_403)
);

INVxp67_ASAP7_75t_SL g404 ( 
.A(n_320),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_215),
.Y(n_405)
);

CKINVDCx5p33_ASAP7_75t_R g406 ( 
.A(n_243),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_215),
.Y(n_407)
);

HB1xp67_ASAP7_75t_L g408 ( 
.A(n_192),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_267),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_237),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_237),
.Y(n_411)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_279),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_259),
.Y(n_413)
);

INVxp33_ASAP7_75t_L g414 ( 
.A(n_208),
.Y(n_414)
);

INVxp67_ASAP7_75t_SL g415 ( 
.A(n_282),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_245),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_276),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_259),
.Y(n_418)
);

INVx3_ASAP7_75t_L g419 ( 
.A(n_282),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_299),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_300),
.Y(n_421)
);

INVxp67_ASAP7_75t_SL g422 ( 
.A(n_285),
.Y(n_422)
);

INVx2_ASAP7_75t_L g423 ( 
.A(n_279),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_299),
.Y(n_424)
);

CKINVDCx5p33_ASAP7_75t_R g425 ( 
.A(n_248),
.Y(n_425)
);

INVxp33_ASAP7_75t_L g426 ( 
.A(n_220),
.Y(n_426)
);

INVxp67_ASAP7_75t_L g427 ( 
.A(n_230),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_314),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_314),
.Y(n_429)
);

INVx2_ASAP7_75t_SL g430 ( 
.A(n_336),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_336),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_246),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_255),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_249),
.Y(n_434)
);

INVxp67_ASAP7_75t_SL g435 ( 
.A(n_285),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_265),
.Y(n_436)
);

CKINVDCx5p33_ASAP7_75t_R g437 ( 
.A(n_251),
.Y(n_437)
);

CKINVDCx20_ASAP7_75t_R g438 ( 
.A(n_331),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_192),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_287),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_296),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_353),
.Y(n_442)
);

CKINVDCx5p33_ASAP7_75t_R g443 ( 
.A(n_252),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_313),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_279),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g446 ( 
.A(n_375),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_318),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_321),
.Y(n_448)
);

CKINVDCx5p33_ASAP7_75t_R g449 ( 
.A(n_254),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_327),
.Y(n_450)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_330),
.Y(n_451)
);

CKINVDCx20_ASAP7_75t_R g452 ( 
.A(n_256),
.Y(n_452)
);

CKINVDCx5p33_ASAP7_75t_R g453 ( 
.A(n_261),
.Y(n_453)
);

HB1xp67_ASAP7_75t_L g454 ( 
.A(n_199),
.Y(n_454)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_334),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_263),
.Y(n_456)
);

BUFx2_ASAP7_75t_L g457 ( 
.A(n_199),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_279),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_360),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_366),
.Y(n_460)
);

CKINVDCx16_ASAP7_75t_R g461 ( 
.A(n_346),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_266),
.Y(n_462)
);

CKINVDCx5p33_ASAP7_75t_R g463 ( 
.A(n_270),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_273),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_372),
.Y(n_465)
);

INVx2_ASAP7_75t_L g466 ( 
.A(n_279),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_222),
.Y(n_467)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_222),
.Y(n_468)
);

INVx1_ASAP7_75t_L g469 ( 
.A(n_294),
.Y(n_469)
);

CKINVDCx5p33_ASAP7_75t_R g470 ( 
.A(n_288),
.Y(n_470)
);

BUFx3_ASAP7_75t_L g471 ( 
.A(n_304),
.Y(n_471)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_294),
.Y(n_472)
);

CKINVDCx20_ASAP7_75t_R g473 ( 
.A(n_291),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_364),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_364),
.Y(n_475)
);

NOR2xp67_ASAP7_75t_L g476 ( 
.A(n_419),
.B(n_257),
.Y(n_476)
);

BUFx6f_ASAP7_75t_L g477 ( 
.A(n_382),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_SL g478 ( 
.A(n_395),
.B(n_394),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_381),
.Y(n_479)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_385),
.A2(n_358),
.B1(n_370),
.B2(n_374),
.Y(n_480)
);

INVx3_ASAP7_75t_L g481 ( 
.A(n_382),
.Y(n_481)
);

CKINVDCx16_ASAP7_75t_R g482 ( 
.A(n_461),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_381),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_406),
.B(n_304),
.Y(n_484)
);

INVx2_ASAP7_75t_L g485 ( 
.A(n_382),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_416),
.Y(n_487)
);

INVx2_ASAP7_75t_L g488 ( 
.A(n_384),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_425),
.Y(n_489)
);

INVx3_ASAP7_75t_L g490 ( 
.A(n_412),
.Y(n_490)
);

INVx2_ASAP7_75t_L g491 ( 
.A(n_387),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_387),
.Y(n_492)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_388),
.Y(n_493)
);

AND2x6_ASAP7_75t_L g494 ( 
.A(n_412),
.B(n_257),
.Y(n_494)
);

AND2x4_ASAP7_75t_L g495 ( 
.A(n_398),
.B(n_307),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_434),
.B(n_307),
.Y(n_496)
);

BUFx6f_ASAP7_75t_L g497 ( 
.A(n_388),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_437),
.B(n_362),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_389),
.Y(n_499)
);

HB1xp67_ASAP7_75t_L g500 ( 
.A(n_408),
.Y(n_500)
);

INVx2_ASAP7_75t_L g501 ( 
.A(n_389),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_SL g502 ( 
.A(n_443),
.B(n_209),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_449),
.Y(n_503)
);

CKINVDCx20_ASAP7_75t_R g504 ( 
.A(n_396),
.Y(n_504)
);

AND2x2_ASAP7_75t_L g505 ( 
.A(n_415),
.B(n_422),
.Y(n_505)
);

INVx1_ASAP7_75t_L g506 ( 
.A(n_390),
.Y(n_506)
);

INVxp67_ASAP7_75t_SL g507 ( 
.A(n_419),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_R g508 ( 
.A(n_452),
.B(n_301),
.Y(n_508)
);

BUFx6f_ASAP7_75t_L g509 ( 
.A(n_390),
.Y(n_509)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_392),
.Y(n_510)
);

AOI22xp5_ASAP7_75t_L g511 ( 
.A1(n_386),
.A2(n_380),
.B1(n_377),
.B2(n_374),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_392),
.Y(n_512)
);

INVx1_ASAP7_75t_L g513 ( 
.A(n_393),
.Y(n_513)
);

AND2x6_ASAP7_75t_L g514 ( 
.A(n_423),
.B(n_257),
.Y(n_514)
);

INVx2_ASAP7_75t_L g515 ( 
.A(n_393),
.Y(n_515)
);

INVx2_ASAP7_75t_L g516 ( 
.A(n_399),
.Y(n_516)
);

INVx2_ASAP7_75t_L g517 ( 
.A(n_399),
.Y(n_517)
);

AND2x2_ASAP7_75t_L g518 ( 
.A(n_435),
.B(n_362),
.Y(n_518)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_432),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_432),
.Y(n_520)
);

AND2x2_ASAP7_75t_L g521 ( 
.A(n_404),
.B(n_196),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_453),
.Y(n_522)
);

BUFx2_ASAP7_75t_L g523 ( 
.A(n_457),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_402),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_423),
.Y(n_525)
);

CKINVDCx5p33_ASAP7_75t_R g526 ( 
.A(n_456),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_433),
.Y(n_527)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_391),
.A2(n_380),
.B1(n_377),
.B2(n_365),
.Y(n_528)
);

INVx1_ASAP7_75t_L g529 ( 
.A(n_433),
.Y(n_529)
);

INVx3_ASAP7_75t_L g530 ( 
.A(n_445),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_436),
.Y(n_531)
);

INVx2_ASAP7_75t_L g532 ( 
.A(n_402),
.Y(n_532)
);

INVx1_ASAP7_75t_L g533 ( 
.A(n_436),
.Y(n_533)
);

INVx3_ASAP7_75t_L g534 ( 
.A(n_445),
.Y(n_534)
);

CKINVDCx20_ASAP7_75t_R g535 ( 
.A(n_400),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_419),
.Y(n_536)
);

NAND2xp5_ASAP7_75t_L g537 ( 
.A(n_462),
.B(n_209),
.Y(n_537)
);

AND2x2_ASAP7_75t_SL g538 ( 
.A(n_458),
.B(n_195),
.Y(n_538)
);

INVx1_ASAP7_75t_L g539 ( 
.A(n_440),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_440),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_471),
.Y(n_541)
);

INVx1_ASAP7_75t_L g542 ( 
.A(n_441),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_458),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_441),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_444),
.Y(n_545)
);

INVx1_ASAP7_75t_L g546 ( 
.A(n_444),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_447),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_447),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_457),
.A2(n_325),
.B1(n_203),
.B2(n_212),
.Y(n_549)
);

BUFx6f_ASAP7_75t_L g550 ( 
.A(n_466),
.Y(n_550)
);

INVx1_ASAP7_75t_L g551 ( 
.A(n_448),
.Y(n_551)
);

AND2x4_ASAP7_75t_L g552 ( 
.A(n_471),
.B(n_272),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_463),
.B(n_272),
.Y(n_553)
);

CKINVDCx5p33_ASAP7_75t_R g554 ( 
.A(n_464),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_519),
.Y(n_555)
);

NAND2xp5_ASAP7_75t_SL g556 ( 
.A(n_554),
.B(n_470),
.Y(n_556)
);

BUFx6f_ASAP7_75t_L g557 ( 
.A(n_477),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_505),
.B(n_430),
.Y(n_558)
);

INVx2_ASAP7_75t_SL g559 ( 
.A(n_541),
.Y(n_559)
);

CKINVDCx16_ASAP7_75t_R g560 ( 
.A(n_482),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_505),
.B(n_430),
.Y(n_561)
);

INVx2_ASAP7_75t_L g562 ( 
.A(n_488),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g563 ( 
.A(n_507),
.B(n_326),
.Y(n_563)
);

INVx2_ASAP7_75t_L g564 ( 
.A(n_488),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_543),
.Y(n_565)
);

INVx2_ASAP7_75t_L g566 ( 
.A(n_491),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_525),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_519),
.Y(n_568)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_487),
.B(n_473),
.Y(n_569)
);

INVxp67_ASAP7_75t_L g570 ( 
.A(n_523),
.Y(n_570)
);

BUFx2_ASAP7_75t_L g571 ( 
.A(n_541),
.Y(n_571)
);

NAND2xp5_ASAP7_75t_SL g572 ( 
.A(n_489),
.B(n_397),
.Y(n_572)
);

INVx2_ASAP7_75t_L g573 ( 
.A(n_491),
.Y(n_573)
);

INVx3_ASAP7_75t_L g574 ( 
.A(n_525),
.Y(n_574)
);

INVx1_ASAP7_75t_L g575 ( 
.A(n_543),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g576 ( 
.A(n_503),
.B(n_383),
.Y(n_576)
);

INVxp33_ASAP7_75t_L g577 ( 
.A(n_480),
.Y(n_577)
);

AND2x2_ASAP7_75t_L g578 ( 
.A(n_518),
.B(n_413),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_518),
.B(n_413),
.Y(n_579)
);

INVx3_ASAP7_75t_L g580 ( 
.A(n_525),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_523),
.B(n_439),
.Y(n_581)
);

AND2x6_ASAP7_75t_L g582 ( 
.A(n_552),
.B(n_195),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_501),
.Y(n_583)
);

BUFx3_ASAP7_75t_L g584 ( 
.A(n_541),
.Y(n_584)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_536),
.B(n_326),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_479),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_479),
.Y(n_587)
);

NOR2xp33_ASAP7_75t_L g588 ( 
.A(n_537),
.B(n_454),
.Y(n_588)
);

INVx2_ASAP7_75t_L g589 ( 
.A(n_501),
.Y(n_589)
);

NOR2xp33_ASAP7_75t_L g590 ( 
.A(n_553),
.B(n_414),
.Y(n_590)
);

BUFx4f_ASAP7_75t_L g591 ( 
.A(n_538),
.Y(n_591)
);

INVx1_ASAP7_75t_SL g592 ( 
.A(n_504),
.Y(n_592)
);

NAND2xp33_ASAP7_75t_R g593 ( 
.A(n_508),
.B(n_200),
.Y(n_593)
);

INVx2_ASAP7_75t_L g594 ( 
.A(n_516),
.Y(n_594)
);

INVx1_ASAP7_75t_L g595 ( 
.A(n_483),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_483),
.Y(n_596)
);

NAND2xp5_ASAP7_75t_SL g597 ( 
.A(n_522),
.B(n_200),
.Y(n_597)
);

INVx1_ASAP7_75t_L g598 ( 
.A(n_486),
.Y(n_598)
);

AND2x4_ASAP7_75t_L g599 ( 
.A(n_495),
.B(n_448),
.Y(n_599)
);

INVx5_ASAP7_75t_L g600 ( 
.A(n_494),
.Y(n_600)
);

INVx2_ASAP7_75t_L g601 ( 
.A(n_516),
.Y(n_601)
);

INVx1_ASAP7_75t_SL g602 ( 
.A(n_535),
.Y(n_602)
);

INVx2_ASAP7_75t_L g603 ( 
.A(n_517),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_536),
.B(n_262),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_536),
.B(n_303),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_SL g606 ( 
.A(n_526),
.B(n_201),
.Y(n_606)
);

OAI22xp33_ASAP7_75t_SL g607 ( 
.A1(n_502),
.A2(n_401),
.B1(n_427),
.B2(n_315),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_SL g608 ( 
.A(n_484),
.B(n_201),
.Y(n_608)
);

INVx1_ASAP7_75t_L g609 ( 
.A(n_520),
.Y(n_609)
);

INVx1_ASAP7_75t_L g610 ( 
.A(n_520),
.Y(n_610)
);

BUFx6f_ASAP7_75t_L g611 ( 
.A(n_477),
.Y(n_611)
);

AND2x4_ASAP7_75t_L g612 ( 
.A(n_495),
.B(n_450),
.Y(n_612)
);

INVx2_ASAP7_75t_L g613 ( 
.A(n_517),
.Y(n_613)
);

INVx2_ASAP7_75t_SL g614 ( 
.A(n_495),
.Y(n_614)
);

NOR2xp33_ASAP7_75t_L g615 ( 
.A(n_496),
.B(n_426),
.Y(n_615)
);

INVx1_ASAP7_75t_L g616 ( 
.A(n_527),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_527),
.Y(n_617)
);

NOR3xp33_ASAP7_75t_L g618 ( 
.A(n_549),
.B(n_347),
.C(n_247),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_529),
.Y(n_619)
);

INVx2_ASAP7_75t_L g620 ( 
.A(n_485),
.Y(n_620)
);

INVxp67_ASAP7_75t_SL g621 ( 
.A(n_525),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_529),
.Y(n_622)
);

INVx2_ASAP7_75t_L g623 ( 
.A(n_485),
.Y(n_623)
);

INVx1_ASAP7_75t_SL g624 ( 
.A(n_482),
.Y(n_624)
);

INVx3_ASAP7_75t_L g625 ( 
.A(n_525),
.Y(n_625)
);

INVx2_ASAP7_75t_SL g626 ( 
.A(n_495),
.Y(n_626)
);

AOI22xp5_ASAP7_75t_L g627 ( 
.A1(n_521),
.A2(n_403),
.B1(n_446),
.B2(n_442),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_486),
.Y(n_628)
);

INVx2_ASAP7_75t_L g629 ( 
.A(n_515),
.Y(n_629)
);

NAND2xp5_ASAP7_75t_SL g630 ( 
.A(n_498),
.B(n_206),
.Y(n_630)
);

OR2x6_ASAP7_75t_L g631 ( 
.A(n_478),
.B(n_418),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_515),
.Y(n_632)
);

INVx2_ASAP7_75t_L g633 ( 
.A(n_515),
.Y(n_633)
);

INVx1_ASAP7_75t_L g634 ( 
.A(n_492),
.Y(n_634)
);

INVx2_ASAP7_75t_L g635 ( 
.A(n_492),
.Y(n_635)
);

INVx1_ASAP7_75t_L g636 ( 
.A(n_493),
.Y(n_636)
);

CKINVDCx16_ASAP7_75t_R g637 ( 
.A(n_480),
.Y(n_637)
);

INVxp33_ASAP7_75t_L g638 ( 
.A(n_500),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_531),
.Y(n_639)
);

NAND2xp5_ASAP7_75t_SL g640 ( 
.A(n_511),
.B(n_206),
.Y(n_640)
);

CKINVDCx12_ASAP7_75t_R g641 ( 
.A(n_521),
.Y(n_641)
);

BUFx10_ASAP7_75t_L g642 ( 
.A(n_552),
.Y(n_642)
);

BUFx6f_ASAP7_75t_L g643 ( 
.A(n_477),
.Y(n_643)
);

AOI22xp33_ASAP7_75t_L g644 ( 
.A1(n_538),
.A2(n_202),
.B1(n_274),
.B2(n_277),
.Y(n_644)
);

INVx2_ASAP7_75t_L g645 ( 
.A(n_493),
.Y(n_645)
);

INVx1_ASAP7_75t_L g646 ( 
.A(n_499),
.Y(n_646)
);

NAND2xp5_ASAP7_75t_L g647 ( 
.A(n_536),
.B(n_335),
.Y(n_647)
);

OA22x2_ASAP7_75t_L g648 ( 
.A1(n_511),
.A2(n_475),
.B1(n_474),
.B2(n_472),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_499),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_506),
.Y(n_650)
);

INVx3_ASAP7_75t_L g651 ( 
.A(n_525),
.Y(n_651)
);

INVx1_ASAP7_75t_L g652 ( 
.A(n_531),
.Y(n_652)
);

NAND2xp33_ASAP7_75t_L g653 ( 
.A(n_494),
.B(n_204),
.Y(n_653)
);

CKINVDCx5p33_ASAP7_75t_R g654 ( 
.A(n_528),
.Y(n_654)
);

AOI22xp33_ASAP7_75t_L g655 ( 
.A1(n_538),
.A2(n_202),
.B1(n_274),
.B2(n_277),
.Y(n_655)
);

AOI22xp5_ASAP7_75t_L g656 ( 
.A1(n_552),
.A2(n_409),
.B1(n_438),
.B2(n_417),
.Y(n_656)
);

INVx2_ASAP7_75t_L g657 ( 
.A(n_506),
.Y(n_657)
);

INVx1_ASAP7_75t_L g658 ( 
.A(n_533),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_510),
.Y(n_659)
);

INVx1_ASAP7_75t_SL g660 ( 
.A(n_552),
.Y(n_660)
);

CKINVDCx14_ASAP7_75t_R g661 ( 
.A(n_528),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_481),
.B(n_371),
.Y(n_662)
);

OR2x6_ASAP7_75t_L g663 ( 
.A(n_533),
.B(n_418),
.Y(n_663)
);

INVx1_ASAP7_75t_L g664 ( 
.A(n_510),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_512),
.Y(n_665)
);

NAND2xp33_ASAP7_75t_L g666 ( 
.A(n_494),
.B(n_204),
.Y(n_666)
);

INVx2_ASAP7_75t_L g667 ( 
.A(n_512),
.Y(n_667)
);

INVx2_ASAP7_75t_L g668 ( 
.A(n_513),
.Y(n_668)
);

INVx4_ASAP7_75t_L g669 ( 
.A(n_550),
.Y(n_669)
);

AOI22xp33_ASAP7_75t_L g670 ( 
.A1(n_494),
.A2(n_349),
.B1(n_283),
.B2(n_379),
.Y(n_670)
);

AO21x2_ASAP7_75t_L g671 ( 
.A1(n_476),
.A2(n_193),
.B(n_191),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_513),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_490),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_490),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_539),
.Y(n_675)
);

INVx2_ASAP7_75t_L g676 ( 
.A(n_490),
.Y(n_676)
);

INVx2_ASAP7_75t_L g677 ( 
.A(n_490),
.Y(n_677)
);

INVx2_ASAP7_75t_L g678 ( 
.A(n_530),
.Y(n_678)
);

AOI22xp33_ASAP7_75t_L g679 ( 
.A1(n_494),
.A2(n_349),
.B1(n_283),
.B2(n_379),
.Y(n_679)
);

AOI22xp5_ASAP7_75t_L g680 ( 
.A1(n_476),
.A2(n_421),
.B1(n_216),
.B2(n_223),
.Y(n_680)
);

INVx2_ASAP7_75t_L g681 ( 
.A(n_530),
.Y(n_681)
);

INVx1_ASAP7_75t_L g682 ( 
.A(n_530),
.Y(n_682)
);

INVx2_ASAP7_75t_L g683 ( 
.A(n_530),
.Y(n_683)
);

INVx2_ASAP7_75t_L g684 ( 
.A(n_534),
.Y(n_684)
);

OAI22xp33_ASAP7_75t_SL g685 ( 
.A1(n_539),
.A2(n_271),
.B1(n_325),
.B2(n_203),
.Y(n_685)
);

INVx5_ASAP7_75t_L g686 ( 
.A(n_494),
.Y(n_686)
);

INVx1_ASAP7_75t_L g687 ( 
.A(n_534),
.Y(n_687)
);

INVx2_ASAP7_75t_L g688 ( 
.A(n_534),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_534),
.Y(n_689)
);

BUFx6f_ASAP7_75t_L g690 ( 
.A(n_477),
.Y(n_690)
);

OR2x6_ASAP7_75t_L g691 ( 
.A(n_540),
.B(n_420),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_540),
.B(n_207),
.Y(n_692)
);

NAND2xp5_ASAP7_75t_L g693 ( 
.A(n_481),
.B(n_373),
.Y(n_693)
);

INVx1_ASAP7_75t_L g694 ( 
.A(n_481),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_481),
.Y(n_695)
);

HB1xp67_ASAP7_75t_L g696 ( 
.A(n_542),
.Y(n_696)
);

NOR2xp33_ASAP7_75t_L g697 ( 
.A(n_542),
.B(n_420),
.Y(n_697)
);

INVx2_ASAP7_75t_SL g698 ( 
.A(n_544),
.Y(n_698)
);

BUFx6f_ASAP7_75t_SL g699 ( 
.A(n_544),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_545),
.B(n_207),
.Y(n_700)
);

NAND2xp5_ASAP7_75t_SL g701 ( 
.A(n_545),
.B(n_210),
.Y(n_701)
);

INVx1_ASAP7_75t_L g702 ( 
.A(n_524),
.Y(n_702)
);

INVx2_ASAP7_75t_L g703 ( 
.A(n_477),
.Y(n_703)
);

INVx2_ASAP7_75t_L g704 ( 
.A(n_477),
.Y(n_704)
);

INVx1_ASAP7_75t_L g705 ( 
.A(n_524),
.Y(n_705)
);

NOR2xp33_ASAP7_75t_L g706 ( 
.A(n_546),
.B(n_424),
.Y(n_706)
);

NAND2xp5_ASAP7_75t_L g707 ( 
.A(n_614),
.B(n_550),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_L g708 ( 
.A(n_614),
.B(n_550),
.Y(n_708)
);

INVx1_ASAP7_75t_L g709 ( 
.A(n_696),
.Y(n_709)
);

NAND3xp33_ASAP7_75t_L g710 ( 
.A(n_590),
.B(n_239),
.C(n_238),
.Y(n_710)
);

INVx2_ASAP7_75t_L g711 ( 
.A(n_635),
.Y(n_711)
);

AOI22xp33_ASAP7_75t_L g712 ( 
.A1(n_591),
.A2(n_514),
.B1(n_494),
.B2(n_204),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_582),
.B(n_279),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_591),
.B(n_204),
.Y(n_714)
);

INVx2_ASAP7_75t_L g715 ( 
.A(n_635),
.Y(n_715)
);

INVx2_ASAP7_75t_SL g716 ( 
.A(n_578),
.Y(n_716)
);

OR2x2_ASAP7_75t_L g717 ( 
.A(n_581),
.B(n_424),
.Y(n_717)
);

INVx2_ASAP7_75t_L g718 ( 
.A(n_674),
.Y(n_718)
);

NOR2xp33_ASAP7_75t_L g719 ( 
.A(n_615),
.B(n_210),
.Y(n_719)
);

CKINVDCx5p33_ASAP7_75t_R g720 ( 
.A(n_593),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_L g721 ( 
.A(n_626),
.B(n_550),
.Y(n_721)
);

INVx2_ASAP7_75t_L g722 ( 
.A(n_674),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_676),
.Y(n_723)
);

AOI22xp33_ASAP7_75t_L g724 ( 
.A1(n_591),
.A2(n_514),
.B1(n_494),
.B2(n_204),
.Y(n_724)
);

NOR2xp33_ASAP7_75t_L g725 ( 
.A(n_588),
.B(n_216),
.Y(n_725)
);

INVx1_ASAP7_75t_L g726 ( 
.A(n_555),
.Y(n_726)
);

HB1xp67_ASAP7_75t_L g727 ( 
.A(n_641),
.Y(n_727)
);

NAND2xp5_ASAP7_75t_L g728 ( 
.A(n_626),
.B(n_660),
.Y(n_728)
);

AOI22xp33_ASAP7_75t_L g729 ( 
.A1(n_644),
.A2(n_514),
.B1(n_233),
.B2(n_322),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_568),
.Y(n_730)
);

BUFx6f_ASAP7_75t_L g731 ( 
.A(n_584),
.Y(n_731)
);

NAND2xp5_ASAP7_75t_L g732 ( 
.A(n_698),
.B(n_550),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_609),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_L g734 ( 
.A(n_698),
.B(n_532),
.Y(n_734)
);

AND2x2_ASAP7_75t_L g735 ( 
.A(n_558),
.B(n_428),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_610),
.Y(n_736)
);

NAND2xp5_ASAP7_75t_SL g737 ( 
.A(n_599),
.B(n_233),
.Y(n_737)
);

INVx1_ASAP7_75t_L g738 ( 
.A(n_616),
.Y(n_738)
);

HB1xp67_ASAP7_75t_L g739 ( 
.A(n_641),
.Y(n_739)
);

AND2x2_ASAP7_75t_L g740 ( 
.A(n_558),
.B(n_428),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_599),
.B(n_532),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_645),
.Y(n_742)
);

NAND2xp5_ASAP7_75t_L g743 ( 
.A(n_599),
.B(n_497),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_612),
.B(n_497),
.Y(n_744)
);

OAI221xp5_ASAP7_75t_L g745 ( 
.A1(n_655),
.A2(n_551),
.B1(n_548),
.B2(n_547),
.C(n_546),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_617),
.Y(n_746)
);

AND2x4_ASAP7_75t_L g747 ( 
.A(n_584),
.B(n_547),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_612),
.B(n_497),
.Y(n_748)
);

OR2x2_ASAP7_75t_L g749 ( 
.A(n_581),
.B(n_429),
.Y(n_749)
);

NAND2xp5_ASAP7_75t_L g750 ( 
.A(n_612),
.B(n_497),
.Y(n_750)
);

NOR2xp33_ASAP7_75t_L g751 ( 
.A(n_561),
.B(n_218),
.Y(n_751)
);

NAND2xp5_ASAP7_75t_L g752 ( 
.A(n_604),
.B(n_497),
.Y(n_752)
);

AND2x4_ASAP7_75t_L g753 ( 
.A(n_559),
.B(n_571),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_619),
.Y(n_754)
);

NOR2xp67_ASAP7_75t_L g755 ( 
.A(n_656),
.B(n_548),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_561),
.B(n_640),
.Y(n_756)
);

BUFx3_ASAP7_75t_L g757 ( 
.A(n_571),
.Y(n_757)
);

NAND2xp33_ASAP7_75t_L g758 ( 
.A(n_582),
.B(n_279),
.Y(n_758)
);

INVx1_ASAP7_75t_L g759 ( 
.A(n_622),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_L g760 ( 
.A(n_608),
.B(n_218),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_605),
.B(n_647),
.Y(n_761)
);

OAI22xp33_ASAP7_75t_L g762 ( 
.A1(n_577),
.A2(n_342),
.B1(n_365),
.B2(n_361),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_648),
.A2(n_514),
.B1(n_233),
.B2(n_322),
.Y(n_763)
);

INVx2_ASAP7_75t_L g764 ( 
.A(n_645),
.Y(n_764)
);

AND2x2_ASAP7_75t_L g765 ( 
.A(n_578),
.B(n_429),
.Y(n_765)
);

NAND2xp5_ASAP7_75t_L g766 ( 
.A(n_639),
.B(n_497),
.Y(n_766)
);

NAND2xp5_ASAP7_75t_L g767 ( 
.A(n_652),
.B(n_658),
.Y(n_767)
);

NOR2xp33_ASAP7_75t_L g768 ( 
.A(n_630),
.B(n_223),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_675),
.B(n_509),
.Y(n_769)
);

BUFx6f_ASAP7_75t_L g770 ( 
.A(n_642),
.Y(n_770)
);

NOR2xp33_ASAP7_75t_L g771 ( 
.A(n_579),
.B(n_228),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_L g772 ( 
.A(n_579),
.B(n_662),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_L g773 ( 
.A(n_693),
.B(n_509),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_559),
.B(n_509),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_586),
.B(n_509),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_694),
.Y(n_776)
);

AND2x4_ASAP7_75t_L g777 ( 
.A(n_663),
.B(n_551),
.Y(n_777)
);

CKINVDCx20_ASAP7_75t_R g778 ( 
.A(n_560),
.Y(n_778)
);

OAI22xp5_ASAP7_75t_L g779 ( 
.A1(n_631),
.A2(n_333),
.B1(n_312),
.B2(n_311),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_586),
.B(n_509),
.Y(n_780)
);

AOI221xp5_ASAP7_75t_L g781 ( 
.A1(n_654),
.A2(n_231),
.B1(n_338),
.B2(n_340),
.C(n_342),
.Y(n_781)
);

NAND2xp33_ASAP7_75t_L g782 ( 
.A(n_582),
.B(n_585),
.Y(n_782)
);

NAND2xp33_ASAP7_75t_L g783 ( 
.A(n_582),
.B(n_563),
.Y(n_783)
);

NOR2xp33_ASAP7_75t_L g784 ( 
.A(n_597),
.B(n_228),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_638),
.B(n_431),
.Y(n_785)
);

NAND2xp33_ASAP7_75t_L g786 ( 
.A(n_582),
.B(n_279),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_570),
.B(n_431),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_676),
.Y(n_788)
);

INVx2_ASAP7_75t_L g789 ( 
.A(n_677),
.Y(n_789)
);

OAI22xp5_ASAP7_75t_SL g790 ( 
.A1(n_661),
.A2(n_235),
.B1(n_232),
.B2(n_231),
.Y(n_790)
);

INVx1_ASAP7_75t_L g791 ( 
.A(n_694),
.Y(n_791)
);

AND2x2_ASAP7_75t_L g792 ( 
.A(n_624),
.B(n_467),
.Y(n_792)
);

AOI221xp5_ASAP7_75t_L g793 ( 
.A1(n_654),
.A2(n_212),
.B1(n_338),
.B2(n_214),
.C(n_340),
.Y(n_793)
);

NAND2xp5_ASAP7_75t_L g794 ( 
.A(n_587),
.B(n_509),
.Y(n_794)
);

NAND2xp33_ASAP7_75t_SL g795 ( 
.A(n_699),
.B(n_214),
.Y(n_795)
);

INVx1_ASAP7_75t_L g796 ( 
.A(n_695),
.Y(n_796)
);

NOR2xp33_ASAP7_75t_L g797 ( 
.A(n_606),
.B(n_229),
.Y(n_797)
);

NOR3xp33_ASAP7_75t_L g798 ( 
.A(n_637),
.B(n_468),
.C(n_467),
.Y(n_798)
);

INVx4_ASAP7_75t_L g799 ( 
.A(n_557),
.Y(n_799)
);

INVx1_ASAP7_75t_L g800 ( 
.A(n_695),
.Y(n_800)
);

INVx2_ASAP7_75t_L g801 ( 
.A(n_657),
.Y(n_801)
);

BUFx6f_ASAP7_75t_L g802 ( 
.A(n_642),
.Y(n_802)
);

NAND2xp5_ASAP7_75t_L g803 ( 
.A(n_587),
.B(n_514),
.Y(n_803)
);

INVx2_ASAP7_75t_L g804 ( 
.A(n_677),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_657),
.Y(n_805)
);

NAND2xp5_ASAP7_75t_L g806 ( 
.A(n_595),
.B(n_514),
.Y(n_806)
);

NAND2xp5_ASAP7_75t_SL g807 ( 
.A(n_642),
.B(n_233),
.Y(n_807)
);

NAND2xp5_ASAP7_75t_L g808 ( 
.A(n_595),
.B(n_514),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_SL g809 ( 
.A(n_600),
.B(n_686),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_596),
.Y(n_810)
);

BUFx6f_ASAP7_75t_L g811 ( 
.A(n_557),
.Y(n_811)
);

OAI22xp5_ASAP7_75t_L g812 ( 
.A1(n_631),
.A2(n_250),
.B1(n_297),
.B2(n_293),
.Y(n_812)
);

BUFx3_ASAP7_75t_L g813 ( 
.A(n_663),
.Y(n_813)
);

NAND2xp5_ASAP7_75t_L g814 ( 
.A(n_596),
.B(n_514),
.Y(n_814)
);

NAND2xp5_ASAP7_75t_L g815 ( 
.A(n_598),
.B(n_194),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_598),
.Y(n_816)
);

NOR2xp33_ASAP7_75t_L g817 ( 
.A(n_572),
.B(n_229),
.Y(n_817)
);

INVx2_ASAP7_75t_SL g818 ( 
.A(n_631),
.Y(n_818)
);

AND2x2_ASAP7_75t_L g819 ( 
.A(n_627),
.B(n_468),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_628),
.Y(n_820)
);

NAND2xp5_ASAP7_75t_L g821 ( 
.A(n_628),
.B(n_197),
.Y(n_821)
);

OAI22xp5_ASAP7_75t_L g822 ( 
.A1(n_631),
.A2(n_680),
.B1(n_691),
.B2(n_663),
.Y(n_822)
);

INVx2_ASAP7_75t_L g823 ( 
.A(n_659),
.Y(n_823)
);

NAND2xp5_ASAP7_75t_L g824 ( 
.A(n_634),
.B(n_213),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_634),
.B(n_219),
.Y(n_825)
);

NOR2xp33_ASAP7_75t_R g826 ( 
.A(n_592),
.B(n_234),
.Y(n_826)
);

INVx2_ASAP7_75t_L g827 ( 
.A(n_659),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_636),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_636),
.B(n_227),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_667),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_646),
.B(n_236),
.Y(n_831)
);

NOR2xp67_ASAP7_75t_L g832 ( 
.A(n_576),
.B(n_469),
.Y(n_832)
);

AO221x1_ASAP7_75t_L g833 ( 
.A1(n_567),
.A2(n_322),
.B1(n_233),
.B2(n_376),
.C(n_354),
.Y(n_833)
);

NAND2xp5_ASAP7_75t_L g834 ( 
.A(n_646),
.B(n_241),
.Y(n_834)
);

BUFx4_ASAP7_75t_L g835 ( 
.A(n_602),
.Y(n_835)
);

BUFx3_ASAP7_75t_L g836 ( 
.A(n_663),
.Y(n_836)
);

AOI22xp5_ASAP7_75t_L g837 ( 
.A1(n_582),
.A2(n_310),
.B1(n_305),
.B2(n_309),
.Y(n_837)
);

INVx1_ASAP7_75t_L g838 ( 
.A(n_649),
.Y(n_838)
);

INVx1_ASAP7_75t_L g839 ( 
.A(n_649),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_648),
.A2(n_322),
.B1(n_264),
.B2(n_260),
.Y(n_840)
);

OR2x6_ASAP7_75t_L g841 ( 
.A(n_569),
.B(n_469),
.Y(n_841)
);

NOR3xp33_ASAP7_75t_L g842 ( 
.A(n_685),
.B(n_475),
.C(n_474),
.Y(n_842)
);

NAND2xp5_ASAP7_75t_L g843 ( 
.A(n_650),
.B(n_664),
.Y(n_843)
);

AOI22xp5_ASAP7_75t_L g844 ( 
.A1(n_699),
.A2(n_328),
.B1(n_234),
.B2(n_329),
.Y(n_844)
);

AOI22xp5_ASAP7_75t_L g845 ( 
.A1(n_699),
.A2(n_691),
.B1(n_648),
.B2(n_618),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_SL g846 ( 
.A(n_600),
.B(n_322),
.Y(n_846)
);

NAND2xp5_ASAP7_75t_L g847 ( 
.A(n_650),
.B(n_244),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_L g848 ( 
.A(n_664),
.B(n_258),
.Y(n_848)
);

NAND2xp5_ASAP7_75t_L g849 ( 
.A(n_665),
.B(n_278),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_665),
.Y(n_850)
);

OAI221xp5_ASAP7_75t_L g851 ( 
.A1(n_697),
.A2(n_378),
.B1(n_302),
.B2(n_332),
.C(n_341),
.Y(n_851)
);

OAI21xp5_ASAP7_75t_L g852 ( 
.A1(n_621),
.A2(n_345),
.B(n_350),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_667),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_672),
.B(n_308),
.Y(n_854)
);

BUFx6f_ASAP7_75t_SL g855 ( 
.A(n_691),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_672),
.Y(n_856)
);

NOR2xp33_ASAP7_75t_SL g857 ( 
.A(n_607),
.B(n_328),
.Y(n_857)
);

AOI22xp5_ASAP7_75t_L g858 ( 
.A1(n_691),
.A2(n_556),
.B1(n_692),
.B2(n_700),
.Y(n_858)
);

NOR2xp33_ASAP7_75t_L g859 ( 
.A(n_701),
.B(n_329),
.Y(n_859)
);

NAND2xp5_ASAP7_75t_SL g860 ( 
.A(n_600),
.B(n_337),
.Y(n_860)
);

OAI22xp5_ASAP7_75t_L g861 ( 
.A1(n_670),
.A2(n_367),
.B1(n_337),
.B2(n_348),
.Y(n_861)
);

A2O1A1Ixp33_ASAP7_75t_L g862 ( 
.A1(n_706),
.A2(n_465),
.B(n_460),
.C(n_459),
.Y(n_862)
);

NAND2xp5_ASAP7_75t_SL g863 ( 
.A(n_600),
.B(n_339),
.Y(n_863)
);

NOR2xp33_ASAP7_75t_L g864 ( 
.A(n_668),
.B(n_339),
.Y(n_864)
);

NOR2xp33_ASAP7_75t_L g865 ( 
.A(n_668),
.B(n_348),
.Y(n_865)
);

INVx2_ASAP7_75t_L g866 ( 
.A(n_678),
.Y(n_866)
);

NAND2xp5_ASAP7_75t_L g867 ( 
.A(n_702),
.B(n_352),
.Y(n_867)
);

AND2x2_ASAP7_75t_L g868 ( 
.A(n_702),
.B(n_472),
.Y(n_868)
);

NAND2xp5_ASAP7_75t_L g869 ( 
.A(n_705),
.B(n_352),
.Y(n_869)
);

NAND2xp5_ASAP7_75t_L g870 ( 
.A(n_567),
.B(n_355),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_673),
.B(n_355),
.Y(n_871)
);

NOR3xp33_ASAP7_75t_L g872 ( 
.A(n_653),
.B(n_465),
.C(n_460),
.Y(n_872)
);

BUFx3_ASAP7_75t_L g873 ( 
.A(n_703),
.Y(n_873)
);

NAND2xp33_ASAP7_75t_L g874 ( 
.A(n_703),
.B(n_363),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_567),
.B(n_363),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_SL g876 ( 
.A(n_600),
.B(n_367),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_SL g877 ( 
.A(n_761),
.B(n_686),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_776),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_770),
.B(n_686),
.Y(n_879)
);

INVx1_ASAP7_75t_SL g880 ( 
.A(n_835),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_772),
.B(n_673),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_711),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_SL g883 ( 
.A(n_770),
.B(n_686),
.Y(n_883)
);

NOR2xp33_ASAP7_75t_L g884 ( 
.A(n_725),
.B(n_574),
.Y(n_884)
);

OR2x2_ASAP7_75t_L g885 ( 
.A(n_717),
.B(n_451),
.Y(n_885)
);

NAND2xp5_ASAP7_75t_L g886 ( 
.A(n_719),
.B(n_682),
.Y(n_886)
);

NOR2x1p5_ASAP7_75t_L g887 ( 
.A(n_720),
.B(n_224),
.Y(n_887)
);

INVx1_ASAP7_75t_SL g888 ( 
.A(n_785),
.Y(n_888)
);

INVxp67_ASAP7_75t_L g889 ( 
.A(n_792),
.Y(n_889)
);

AO22x1_ASAP7_75t_L g890 ( 
.A1(n_725),
.A2(n_719),
.B1(n_817),
.B2(n_797),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_791),
.Y(n_891)
);

OR2x6_ASAP7_75t_L g892 ( 
.A(n_757),
.B(n_451),
.Y(n_892)
);

INVx3_ASAP7_75t_L g893 ( 
.A(n_873),
.Y(n_893)
);

INVx1_ASAP7_75t_L g894 ( 
.A(n_796),
.Y(n_894)
);

BUFx8_ASAP7_75t_L g895 ( 
.A(n_855),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_L g896 ( 
.A(n_810),
.B(n_682),
.Y(n_896)
);

NOR2x2_ASAP7_75t_L g897 ( 
.A(n_841),
.B(n_704),
.Y(n_897)
);

BUFx6f_ASAP7_75t_L g898 ( 
.A(n_770),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_L g899 ( 
.A(n_816),
.B(n_687),
.Y(n_899)
);

AOI22xp33_ASAP7_75t_L g900 ( 
.A1(n_840),
.A2(n_671),
.B1(n_679),
.B2(n_565),
.Y(n_900)
);

INVx1_ASAP7_75t_L g901 ( 
.A(n_800),
.Y(n_901)
);

OR2x2_ASAP7_75t_SL g902 ( 
.A(n_727),
.B(n_455),
.Y(n_902)
);

NAND2xp5_ASAP7_75t_L g903 ( 
.A(n_820),
.B(n_687),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_L g904 ( 
.A(n_828),
.B(n_689),
.Y(n_904)
);

AND2x6_ASAP7_75t_L g905 ( 
.A(n_770),
.B(n_704),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_711),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_838),
.B(n_689),
.Y(n_907)
);

HB1xp67_ASAP7_75t_L g908 ( 
.A(n_757),
.Y(n_908)
);

BUFx6f_ASAP7_75t_L g909 ( 
.A(n_802),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_839),
.B(n_574),
.Y(n_910)
);

HB1xp67_ASAP7_75t_L g911 ( 
.A(n_753),
.Y(n_911)
);

NAND2xp5_ASAP7_75t_L g912 ( 
.A(n_850),
.B(n_856),
.Y(n_912)
);

INVx2_ASAP7_75t_L g913 ( 
.A(n_715),
.Y(n_913)
);

INVxp67_ASAP7_75t_SL g914 ( 
.A(n_811),
.Y(n_914)
);

INVx2_ASAP7_75t_L g915 ( 
.A(n_715),
.Y(n_915)
);

INVx2_ASAP7_75t_L g916 ( 
.A(n_742),
.Y(n_916)
);

INVx2_ASAP7_75t_L g917 ( 
.A(n_742),
.Y(n_917)
);

INVx2_ASAP7_75t_L g918 ( 
.A(n_764),
.Y(n_918)
);

INVx2_ASAP7_75t_L g919 ( 
.A(n_764),
.Y(n_919)
);

INVx2_ASAP7_75t_L g920 ( 
.A(n_801),
.Y(n_920)
);

INVx3_ASAP7_75t_L g921 ( 
.A(n_873),
.Y(n_921)
);

NAND2xp5_ASAP7_75t_L g922 ( 
.A(n_751),
.B(n_574),
.Y(n_922)
);

AND2x2_ASAP7_75t_L g923 ( 
.A(n_787),
.B(n_455),
.Y(n_923)
);

NAND2xp33_ASAP7_75t_R g924 ( 
.A(n_826),
.B(n_224),
.Y(n_924)
);

NAND2xp5_ASAP7_75t_SL g925 ( 
.A(n_802),
.B(n_686),
.Y(n_925)
);

AOI22xp5_ASAP7_75t_L g926 ( 
.A1(n_756),
.A2(n_580),
.B1(n_625),
.B2(n_651),
.Y(n_926)
);

OAI22xp5_ASAP7_75t_L g927 ( 
.A1(n_756),
.A2(n_625),
.B1(n_580),
.B2(n_651),
.Y(n_927)
);

OR2x6_ASAP7_75t_L g928 ( 
.A(n_818),
.B(n_459),
.Y(n_928)
);

INVx5_ASAP7_75t_L g929 ( 
.A(n_802),
.Y(n_929)
);

INVx2_ASAP7_75t_L g930 ( 
.A(n_801),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_747),
.B(n_620),
.Y(n_931)
);

INVx5_ASAP7_75t_L g932 ( 
.A(n_802),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_805),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_L g934 ( 
.A(n_751),
.B(n_580),
.Y(n_934)
);

INVx3_ASAP7_75t_L g935 ( 
.A(n_731),
.Y(n_935)
);

NAND2xp5_ASAP7_75t_SL g936 ( 
.A(n_753),
.B(n_625),
.Y(n_936)
);

AOI22xp33_ASAP7_75t_L g937 ( 
.A1(n_840),
.A2(n_671),
.B1(n_575),
.B2(n_565),
.Y(n_937)
);

NAND2xp5_ASAP7_75t_L g938 ( 
.A(n_735),
.B(n_651),
.Y(n_938)
);

NOR2xp33_ASAP7_75t_L g939 ( 
.A(n_709),
.B(n_669),
.Y(n_939)
);

AND2x6_ASAP7_75t_SL g940 ( 
.A(n_841),
.B(n_405),
.Y(n_940)
);

NAND2xp5_ASAP7_75t_L g941 ( 
.A(n_740),
.B(n_575),
.Y(n_941)
);

INVx5_ASAP7_75t_L g942 ( 
.A(n_811),
.Y(n_942)
);

NOR2xp33_ASAP7_75t_SL g943 ( 
.A(n_778),
.B(n_369),
.Y(n_943)
);

INVx3_ASAP7_75t_L g944 ( 
.A(n_731),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_731),
.Y(n_945)
);

INVx2_ASAP7_75t_L g946 ( 
.A(n_805),
.Y(n_946)
);

NOR2xp33_ASAP7_75t_L g947 ( 
.A(n_728),
.B(n_669),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_823),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_843),
.B(n_678),
.Y(n_949)
);

BUFx3_ASAP7_75t_L g950 ( 
.A(n_731),
.Y(n_950)
);

AND2x2_ASAP7_75t_L g951 ( 
.A(n_716),
.B(n_671),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_823),
.Y(n_952)
);

OAI22xp5_ASAP7_75t_L g953 ( 
.A1(n_714),
.A2(n_669),
.B1(n_620),
.B2(n_623),
.Y(n_953)
);

INVx5_ASAP7_75t_L g954 ( 
.A(n_811),
.Y(n_954)
);

NAND2xp5_ASAP7_75t_SL g955 ( 
.A(n_858),
.B(n_557),
.Y(n_955)
);

AOI22xp5_ASAP7_75t_L g956 ( 
.A1(n_822),
.A2(n_688),
.B1(n_684),
.B2(n_683),
.Y(n_956)
);

NAND2xp5_ASAP7_75t_L g957 ( 
.A(n_771),
.B(n_681),
.Y(n_957)
);

BUFx2_ASAP7_75t_L g958 ( 
.A(n_739),
.Y(n_958)
);

NAND2xp5_ASAP7_75t_SL g959 ( 
.A(n_845),
.B(n_557),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_827),
.Y(n_960)
);

INVx1_ASAP7_75t_L g961 ( 
.A(n_827),
.Y(n_961)
);

NAND2xp5_ASAP7_75t_SL g962 ( 
.A(n_777),
.B(n_557),
.Y(n_962)
);

INVx2_ASAP7_75t_L g963 ( 
.A(n_830),
.Y(n_963)
);

OAI22xp5_ASAP7_75t_L g964 ( 
.A1(n_714),
.A2(n_623),
.B1(n_369),
.B2(n_566),
.Y(n_964)
);

NAND3xp33_ASAP7_75t_SL g965 ( 
.A(n_781),
.B(n_225),
.C(n_232),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_765),
.B(n_681),
.Y(n_966)
);

INVx1_ASAP7_75t_L g967 ( 
.A(n_830),
.Y(n_967)
);

INVx2_ASAP7_75t_L g968 ( 
.A(n_853),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_853),
.Y(n_969)
);

BUFx6f_ASAP7_75t_L g970 ( 
.A(n_811),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_749),
.B(n_683),
.Y(n_971)
);

NAND2xp5_ASAP7_75t_L g972 ( 
.A(n_734),
.B(n_684),
.Y(n_972)
);

INVx2_ASAP7_75t_SL g973 ( 
.A(n_841),
.Y(n_973)
);

NAND2xp5_ASAP7_75t_L g974 ( 
.A(n_726),
.B(n_688),
.Y(n_974)
);

NAND2x1p5_ASAP7_75t_L g975 ( 
.A(n_813),
.B(n_611),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_777),
.B(n_611),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_730),
.B(n_562),
.Y(n_977)
);

OAI22xp5_ASAP7_75t_L g978 ( 
.A1(n_741),
.A2(n_566),
.B1(n_562),
.B2(n_564),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_733),
.B(n_564),
.Y(n_979)
);

INVx1_ASAP7_75t_SL g980 ( 
.A(n_826),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_736),
.Y(n_981)
);

NAND2xp5_ASAP7_75t_L g982 ( 
.A(n_738),
.B(n_573),
.Y(n_982)
);

AND2x2_ASAP7_75t_L g983 ( 
.A(n_819),
.B(n_405),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_855),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_SL g985 ( 
.A(n_803),
.B(n_611),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_806),
.B(n_808),
.Y(n_986)
);

AOI22xp33_ASAP7_75t_L g987 ( 
.A1(n_729),
.A2(n_573),
.B1(n_601),
.B2(n_603),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_817),
.B(n_407),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_746),
.B(n_583),
.Y(n_989)
);

BUFx3_ASAP7_75t_L g990 ( 
.A(n_813),
.Y(n_990)
);

INVx1_ASAP7_75t_L g991 ( 
.A(n_754),
.Y(n_991)
);

BUFx8_ASAP7_75t_L g992 ( 
.A(n_836),
.Y(n_992)
);

AOI21xp5_ASAP7_75t_L g993 ( 
.A1(n_707),
.A2(n_690),
.B(n_643),
.Y(n_993)
);

NAND2xp5_ASAP7_75t_L g994 ( 
.A(n_759),
.B(n_583),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_868),
.Y(n_995)
);

INVx2_ASAP7_75t_L g996 ( 
.A(n_718),
.Y(n_996)
);

O2A1O1Ixp33_ASAP7_75t_L g997 ( 
.A1(n_862),
.A2(n_666),
.B(n_653),
.C(n_613),
.Y(n_997)
);

AOI22xp33_ASAP7_75t_L g998 ( 
.A1(n_729),
.A2(n_589),
.B1(n_601),
.B2(n_594),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_795),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_L g1000 ( 
.A(n_767),
.B(n_589),
.Y(n_1000)
);

NAND2xp5_ASAP7_75t_L g1001 ( 
.A(n_864),
.B(n_594),
.Y(n_1001)
);

NOR2xp33_ASAP7_75t_L g1002 ( 
.A(n_784),
.B(n_242),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_755),
.Y(n_1003)
);

HB1xp67_ASAP7_75t_L g1004 ( 
.A(n_747),
.Y(n_1004)
);

INVx4_ASAP7_75t_L g1005 ( 
.A(n_799),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_708),
.A2(n_690),
.B(n_643),
.Y(n_1006)
);

AOI22xp33_ASAP7_75t_L g1007 ( 
.A1(n_763),
.A2(n_603),
.B1(n_613),
.B2(n_666),
.Y(n_1007)
);

INVx1_ASAP7_75t_L g1008 ( 
.A(n_722),
.Y(n_1008)
);

INVx3_ASAP7_75t_L g1009 ( 
.A(n_799),
.Y(n_1009)
);

INVx1_ASAP7_75t_L g1010 ( 
.A(n_723),
.Y(n_1010)
);

INVx2_ASAP7_75t_L g1011 ( 
.A(n_788),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_789),
.Y(n_1012)
);

BUFx3_ASAP7_75t_L g1013 ( 
.A(n_836),
.Y(n_1013)
);

BUFx2_ASAP7_75t_L g1014 ( 
.A(n_867),
.Y(n_1014)
);

NAND2x1p5_ASAP7_75t_L g1015 ( 
.A(n_809),
.B(n_737),
.Y(n_1015)
);

O2A1O1Ixp33_ASAP7_75t_L g1016 ( 
.A1(n_862),
.A2(n_632),
.B(n_629),
.C(n_633),
.Y(n_1016)
);

INVx2_ASAP7_75t_L g1017 ( 
.A(n_804),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_866),
.Y(n_1018)
);

INVx1_ASAP7_75t_L g1019 ( 
.A(n_775),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_780),
.Y(n_1020)
);

HB1xp67_ASAP7_75t_L g1021 ( 
.A(n_743),
.Y(n_1021)
);

INVx3_ASAP7_75t_L g1022 ( 
.A(n_744),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_864),
.B(n_611),
.Y(n_1023)
);

BUFx6f_ASAP7_75t_L g1024 ( 
.A(n_748),
.Y(n_1024)
);

BUFx3_ASAP7_75t_L g1025 ( 
.A(n_750),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_865),
.B(n_611),
.Y(n_1026)
);

BUFx6f_ASAP7_75t_L g1027 ( 
.A(n_721),
.Y(n_1027)
);

INVx1_ASAP7_75t_L g1028 ( 
.A(n_794),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_766),
.Y(n_1029)
);

OAI21xp33_ASAP7_75t_L g1030 ( 
.A1(n_793),
.A2(n_225),
.B(n_235),
.Y(n_1030)
);

NOR2xp33_ASAP7_75t_L g1031 ( 
.A(n_784),
.B(n_253),
.Y(n_1031)
);

INVx2_ASAP7_75t_L g1032 ( 
.A(n_732),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_865),
.B(n_852),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_769),
.Y(n_1034)
);

INVx2_ASAP7_75t_L g1035 ( 
.A(n_814),
.Y(n_1035)
);

NAND2xp5_ASAP7_75t_L g1036 ( 
.A(n_871),
.B(n_643),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_774),
.Y(n_1037)
);

INVx2_ASAP7_75t_SL g1038 ( 
.A(n_869),
.Y(n_1038)
);

INVx1_ASAP7_75t_SL g1039 ( 
.A(n_790),
.Y(n_1039)
);

OR2x6_ASAP7_75t_L g1040 ( 
.A(n_832),
.B(n_407),
.Y(n_1040)
);

INVx2_ASAP7_75t_SL g1041 ( 
.A(n_815),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_821),
.Y(n_1042)
);

NAND2xp5_ASAP7_75t_SL g1043 ( 
.A(n_712),
.B(n_643),
.Y(n_1043)
);

INVx2_ASAP7_75t_L g1044 ( 
.A(n_773),
.Y(n_1044)
);

INVx1_ASAP7_75t_L g1045 ( 
.A(n_824),
.Y(n_1045)
);

INVx1_ASAP7_75t_L g1046 ( 
.A(n_825),
.Y(n_1046)
);

AND2x2_ASAP7_75t_L g1047 ( 
.A(n_797),
.B(n_410),
.Y(n_1047)
);

BUFx6f_ASAP7_75t_L g1048 ( 
.A(n_809),
.Y(n_1048)
);

INVx1_ASAP7_75t_L g1049 ( 
.A(n_829),
.Y(n_1049)
);

INVx4_ASAP7_75t_L g1050 ( 
.A(n_783),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_831),
.Y(n_1051)
);

BUFx2_ASAP7_75t_L g1052 ( 
.A(n_870),
.Y(n_1052)
);

INVx2_ASAP7_75t_L g1053 ( 
.A(n_834),
.Y(n_1053)
);

INVx4_ASAP7_75t_L g1054 ( 
.A(n_874),
.Y(n_1054)
);

NAND2xp5_ASAP7_75t_SL g1055 ( 
.A(n_712),
.B(n_643),
.Y(n_1055)
);

INVx1_ASAP7_75t_L g1056 ( 
.A(n_847),
.Y(n_1056)
);

BUFx8_ASAP7_75t_L g1057 ( 
.A(n_798),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_848),
.Y(n_1058)
);

NOR2xp33_ASAP7_75t_L g1059 ( 
.A(n_710),
.B(n_857),
.Y(n_1059)
);

NAND2xp5_ASAP7_75t_SL g1060 ( 
.A(n_724),
.B(n_763),
.Y(n_1060)
);

INVx1_ASAP7_75t_L g1061 ( 
.A(n_849),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_871),
.B(n_690),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_760),
.B(n_768),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_737),
.Y(n_1064)
);

NAND2xp5_ASAP7_75t_SL g1065 ( 
.A(n_724),
.B(n_690),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_SL g1066 ( 
.A(n_752),
.B(n_690),
.Y(n_1066)
);

A2O1A1Ixp33_ASAP7_75t_L g1067 ( 
.A1(n_760),
.A2(n_343),
.B(n_344),
.C(n_351),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_844),
.Y(n_1068)
);

INVx3_ASAP7_75t_L g1069 ( 
.A(n_854),
.Y(n_1069)
);

NAND2xp5_ASAP7_75t_SL g1070 ( 
.A(n_1063),
.B(n_768),
.Y(n_1070)
);

A2O1A1Ixp33_ASAP7_75t_L g1071 ( 
.A1(n_1002),
.A2(n_859),
.B(n_779),
.C(n_812),
.Y(n_1071)
);

NOR3xp33_ASAP7_75t_L g1072 ( 
.A(n_890),
.B(n_859),
.C(n_762),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_981),
.Y(n_1073)
);

BUFx12f_ASAP7_75t_L g1074 ( 
.A(n_895),
.Y(n_1074)
);

OA21x2_ASAP7_75t_L g1075 ( 
.A1(n_955),
.A2(n_1062),
.B(n_1036),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_991),
.Y(n_1076)
);

O2A1O1Ixp5_ASAP7_75t_L g1077 ( 
.A1(n_1033),
.A2(n_807),
.B(n_876),
.C(n_863),
.Y(n_1077)
);

NAND3xp33_ASAP7_75t_SL g1078 ( 
.A(n_1002),
.B(n_851),
.C(n_842),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_1031),
.A2(n_745),
.B(n_807),
.C(n_875),
.Y(n_1079)
);

INVx2_ASAP7_75t_L g1080 ( 
.A(n_882),
.Y(n_1080)
);

NOR2xp33_ASAP7_75t_SL g1081 ( 
.A(n_980),
.B(n_762),
.Y(n_1081)
);

OAI22x1_ASAP7_75t_L g1082 ( 
.A1(n_1068),
.A2(n_343),
.B1(n_344),
.B2(n_351),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_908),
.Y(n_1083)
);

O2A1O1Ixp5_ASAP7_75t_L g1084 ( 
.A1(n_1031),
.A2(n_876),
.B(n_863),
.C(n_860),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_L g1085 ( 
.A1(n_1060),
.A2(n_837),
.B1(n_860),
.B2(n_861),
.Y(n_1085)
);

NOR2xp33_ASAP7_75t_L g1086 ( 
.A(n_888),
.B(n_268),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_906),
.Y(n_1087)
);

AND2x2_ASAP7_75t_L g1088 ( 
.A(n_889),
.B(n_872),
.Y(n_1088)
);

AND2x2_ASAP7_75t_L g1089 ( 
.A(n_983),
.B(n_410),
.Y(n_1089)
);

NAND2xp5_ASAP7_75t_L g1090 ( 
.A(n_1047),
.B(n_833),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_988),
.B(n_629),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_933),
.Y(n_1092)
);

INVx2_ASAP7_75t_L g1093 ( 
.A(n_882),
.Y(n_1093)
);

NOR2xp67_ASAP7_75t_L g1094 ( 
.A(n_1003),
.B(n_846),
.Y(n_1094)
);

OAI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_1060),
.A2(n_846),
.B1(n_782),
.B2(n_632),
.Y(n_1095)
);

A2O1A1Ixp33_ASAP7_75t_L g1096 ( 
.A1(n_1059),
.A2(n_786),
.B(n_758),
.C(n_713),
.Y(n_1096)
);

AOI22xp33_ASAP7_75t_L g1097 ( 
.A1(n_965),
.A2(n_356),
.B1(n_357),
.B2(n_361),
.Y(n_1097)
);

OAI22xp5_ASAP7_75t_L g1098 ( 
.A1(n_884),
.A2(n_633),
.B1(n_316),
.B2(n_306),
.Y(n_1098)
);

AO21x2_ASAP7_75t_L g1099 ( 
.A1(n_955),
.A2(n_411),
.B(n_105),
.Y(n_1099)
);

INVx2_ASAP7_75t_L g1100 ( 
.A(n_915),
.Y(n_1100)
);

OAI22xp5_ASAP7_75t_L g1101 ( 
.A1(n_884),
.A2(n_298),
.B1(n_281),
.B2(n_284),
.Y(n_1101)
);

AOI21xp5_ASAP7_75t_L g1102 ( 
.A1(n_1023),
.A2(n_411),
.B(n_323),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_948),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1026),
.A2(n_317),
.B(n_289),
.Y(n_1104)
);

AOI221xp5_ASAP7_75t_L g1105 ( 
.A1(n_1030),
.A2(n_359),
.B1(n_357),
.B2(n_356),
.C(n_324),
.Y(n_1105)
);

NAND2x1p5_ASAP7_75t_L g1106 ( 
.A(n_929),
.B(n_77),
.Y(n_1106)
);

AOI22xp5_ASAP7_75t_L g1107 ( 
.A1(n_1059),
.A2(n_295),
.B1(n_290),
.B2(n_275),
.Y(n_1107)
);

INVx2_ASAP7_75t_SL g1108 ( 
.A(n_958),
.Y(n_1108)
);

OAI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_886),
.A2(n_359),
.B1(n_188),
.B2(n_177),
.Y(n_1109)
);

BUFx12f_ASAP7_75t_L g1110 ( 
.A(n_895),
.Y(n_1110)
);

INVx1_ASAP7_75t_L g1111 ( 
.A(n_952),
.Y(n_1111)
);

A2O1A1Ixp33_ASAP7_75t_L g1112 ( 
.A1(n_1042),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_1112)
);

OR2x6_ASAP7_75t_L g1113 ( 
.A(n_892),
.B(n_170),
.Y(n_1113)
);

INVx2_ASAP7_75t_L g1114 ( 
.A(n_915),
.Y(n_1114)
);

INVx2_ASAP7_75t_L g1115 ( 
.A(n_916),
.Y(n_1115)
);

A2O1A1Ixp33_ASAP7_75t_L g1116 ( 
.A1(n_1045),
.A2(n_1046),
.B(n_1051),
.C(n_1049),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_1056),
.B(n_0),
.Y(n_1117)
);

NAND2xp5_ASAP7_75t_L g1118 ( 
.A(n_1058),
.B(n_2),
.Y(n_1118)
);

NAND2xp5_ASAP7_75t_L g1119 ( 
.A(n_1061),
.B(n_4),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_922),
.A2(n_134),
.B(n_161),
.Y(n_1120)
);

INVx2_ASAP7_75t_L g1121 ( 
.A(n_916),
.Y(n_1121)
);

A2O1A1Ixp33_ASAP7_75t_L g1122 ( 
.A1(n_1038),
.A2(n_4),
.B(n_6),
.C(n_11),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_SL g1123 ( 
.A(n_1014),
.B(n_929),
.Y(n_1123)
);

INVx1_ASAP7_75t_L g1124 ( 
.A(n_960),
.Y(n_1124)
);

BUFx3_ASAP7_75t_L g1125 ( 
.A(n_992),
.Y(n_1125)
);

INVx1_ASAP7_75t_L g1126 ( 
.A(n_961),
.Y(n_1126)
);

AOI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1052),
.A2(n_165),
.B1(n_160),
.B2(n_157),
.Y(n_1127)
);

INVx3_ASAP7_75t_L g1128 ( 
.A(n_898),
.Y(n_1128)
);

BUFx2_ASAP7_75t_L g1129 ( 
.A(n_908),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_967),
.Y(n_1130)
);

NAND2xp5_ASAP7_75t_SL g1131 ( 
.A(n_929),
.B(n_154),
.Y(n_1131)
);

O2A1O1Ixp33_ASAP7_75t_L g1132 ( 
.A1(n_1067),
.A2(n_13),
.B(n_14),
.C(n_15),
.Y(n_1132)
);

AND2x2_ASAP7_75t_L g1133 ( 
.A(n_923),
.B(n_13),
.Y(n_1133)
);

NOR2xp33_ASAP7_75t_L g1134 ( 
.A(n_1041),
.B(n_16),
.Y(n_1134)
);

NOR2xp33_ASAP7_75t_R g1135 ( 
.A(n_999),
.B(n_924),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_917),
.Y(n_1136)
);

INVx2_ASAP7_75t_L g1137 ( 
.A(n_917),
.Y(n_1137)
);

BUFx2_ASAP7_75t_L g1138 ( 
.A(n_892),
.Y(n_1138)
);

NAND2xp5_ASAP7_75t_L g1139 ( 
.A(n_1053),
.B(n_19),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_934),
.A2(n_150),
.B(n_140),
.Y(n_1140)
);

OAI22xp5_ASAP7_75t_L g1141 ( 
.A1(n_1050),
.A2(n_139),
.B1(n_138),
.B2(n_133),
.Y(n_1141)
);

NOR2xp33_ASAP7_75t_L g1142 ( 
.A(n_911),
.B(n_19),
.Y(n_1142)
);

INVx4_ASAP7_75t_L g1143 ( 
.A(n_898),
.Y(n_1143)
);

XOR2xp5_ASAP7_75t_L g1144 ( 
.A(n_984),
.B(n_129),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_878),
.Y(n_1145)
);

A2O1A1Ixp33_ASAP7_75t_L g1146 ( 
.A1(n_1069),
.A2(n_20),
.B(n_21),
.C(n_23),
.Y(n_1146)
);

NOR2xp33_ASAP7_75t_SL g1147 ( 
.A(n_880),
.B(n_126),
.Y(n_1147)
);

AO32x1_ASAP7_75t_L g1148 ( 
.A1(n_964),
.A2(n_23),
.A3(n_25),
.B1(n_28),
.B2(n_30),
.Y(n_1148)
);

INVx2_ASAP7_75t_L g1149 ( 
.A(n_918),
.Y(n_1149)
);

OAI21x1_ASAP7_75t_L g1150 ( 
.A1(n_993),
.A2(n_121),
.B(n_113),
.Y(n_1150)
);

INVx2_ASAP7_75t_L g1151 ( 
.A(n_918),
.Y(n_1151)
);

OR2x6_ASAP7_75t_SL g1152 ( 
.A(n_885),
.B(n_28),
.Y(n_1152)
);

INVx3_ASAP7_75t_L g1153 ( 
.A(n_898),
.Y(n_1153)
);

AND2x2_ASAP7_75t_L g1154 ( 
.A(n_995),
.B(n_911),
.Y(n_1154)
);

AOI21xp5_ASAP7_75t_L g1155 ( 
.A1(n_947),
.A2(n_94),
.B(n_91),
.Y(n_1155)
);

NAND3xp33_ASAP7_75t_SL g1156 ( 
.A(n_1067),
.B(n_943),
.C(n_941),
.Y(n_1156)
);

INVx1_ASAP7_75t_L g1157 ( 
.A(n_891),
.Y(n_1157)
);

HB1xp67_ASAP7_75t_L g1158 ( 
.A(n_1004),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_894),
.Y(n_1159)
);

NAND2xp5_ASAP7_75t_L g1160 ( 
.A(n_971),
.B(n_30),
.Y(n_1160)
);

NAND2xp5_ASAP7_75t_L g1161 ( 
.A(n_971),
.B(n_32),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_901),
.Y(n_1162)
);

INVx2_ASAP7_75t_L g1163 ( 
.A(n_919),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_898),
.Y(n_1164)
);

INVx2_ASAP7_75t_L g1165 ( 
.A(n_919),
.Y(n_1165)
);

A2O1A1Ixp33_ASAP7_75t_L g1166 ( 
.A1(n_1069),
.A2(n_32),
.B(n_38),
.C(n_39),
.Y(n_1166)
);

OAI22x1_ASAP7_75t_L g1167 ( 
.A1(n_1039),
.A2(n_46),
.B1(n_50),
.B2(n_51),
.Y(n_1167)
);

NOR3xp33_ASAP7_75t_L g1168 ( 
.A(n_973),
.B(n_46),
.C(n_52),
.Y(n_1168)
);

NAND2xp5_ASAP7_75t_L g1169 ( 
.A(n_1021),
.B(n_58),
.Y(n_1169)
);

O2A1O1Ixp33_ASAP7_75t_L g1170 ( 
.A1(n_881),
.A2(n_59),
.B(n_60),
.C(n_83),
.Y(n_1170)
);

AOI21xp5_ASAP7_75t_L g1171 ( 
.A1(n_947),
.A2(n_100),
.B(n_60),
.Y(n_1171)
);

O2A1O1Ixp33_ASAP7_75t_L g1172 ( 
.A1(n_959),
.A2(n_957),
.B(n_912),
.C(n_1000),
.Y(n_1172)
);

BUFx8_ASAP7_75t_L g1173 ( 
.A(n_990),
.Y(n_1173)
);

A2O1A1Ixp33_ASAP7_75t_L g1174 ( 
.A1(n_939),
.A2(n_959),
.B(n_1028),
.C(n_1020),
.Y(n_1174)
);

INVx3_ASAP7_75t_L g1175 ( 
.A(n_909),
.Y(n_1175)
);

OR2x6_ASAP7_75t_SL g1176 ( 
.A(n_977),
.B(n_979),
.Y(n_1176)
);

NAND2xp5_ASAP7_75t_L g1177 ( 
.A(n_1021),
.B(n_1044),
.Y(n_1177)
);

INVx1_ASAP7_75t_L g1178 ( 
.A(n_920),
.Y(n_1178)
);

O2A1O1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_1001),
.A2(n_966),
.B(n_994),
.C(n_989),
.Y(n_1179)
);

NAND2xp5_ASAP7_75t_SL g1180 ( 
.A(n_932),
.B(n_909),
.Y(n_1180)
);

NAND3xp33_ASAP7_75t_L g1181 ( 
.A(n_924),
.B(n_1004),
.C(n_892),
.Y(n_1181)
);

BUFx2_ASAP7_75t_L g1182 ( 
.A(n_902),
.Y(n_1182)
);

NAND2xp5_ASAP7_75t_L g1183 ( 
.A(n_1019),
.B(n_1029),
.Y(n_1183)
);

INVx1_ASAP7_75t_SL g1184 ( 
.A(n_897),
.Y(n_1184)
);

NAND2xp5_ASAP7_75t_L g1185 ( 
.A(n_1034),
.B(n_1032),
.Y(n_1185)
);

O2A1O1Ixp33_ASAP7_75t_L g1186 ( 
.A1(n_982),
.A2(n_938),
.B(n_896),
.C(n_899),
.Y(n_1186)
);

AOI22xp5_ASAP7_75t_L g1187 ( 
.A1(n_939),
.A2(n_931),
.B1(n_951),
.B2(n_936),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_R g1188 ( 
.A(n_909),
.B(n_935),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_920),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_913),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_930),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_986),
.A2(n_1065),
.B(n_1055),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_986),
.A2(n_1065),
.B(n_1055),
.Y(n_1193)
);

AND2x2_ASAP7_75t_L g1194 ( 
.A(n_887),
.B(n_990),
.Y(n_1194)
);

OAI22xp5_ASAP7_75t_L g1195 ( 
.A1(n_1050),
.A2(n_937),
.B1(n_1054),
.B2(n_1064),
.Y(n_1195)
);

AOI21xp5_ASAP7_75t_L g1196 ( 
.A1(n_1043),
.A2(n_1066),
.B(n_877),
.Y(n_1196)
);

AOI22xp5_ASAP7_75t_L g1197 ( 
.A1(n_931),
.A2(n_936),
.B1(n_1024),
.B2(n_962),
.Y(n_1197)
);

AND2x2_ASAP7_75t_L g1198 ( 
.A(n_1013),
.B(n_928),
.Y(n_1198)
);

AOI22xp5_ASAP7_75t_L g1199 ( 
.A1(n_1024),
.A2(n_962),
.B1(n_976),
.B2(n_1064),
.Y(n_1199)
);

AND2x2_ASAP7_75t_L g1200 ( 
.A(n_1013),
.B(n_928),
.Y(n_1200)
);

NAND2xp5_ASAP7_75t_L g1201 ( 
.A(n_1025),
.B(n_1037),
.Y(n_1201)
);

AOI21xp5_ASAP7_75t_L g1202 ( 
.A1(n_1043),
.A2(n_1066),
.B(n_877),
.Y(n_1202)
);

AOI21xp5_ASAP7_75t_L g1203 ( 
.A1(n_949),
.A2(n_985),
.B(n_1006),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_928),
.B(n_1040),
.Y(n_1204)
);

INVx1_ASAP7_75t_L g1205 ( 
.A(n_946),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_SL g1206 ( 
.A(n_932),
.B(n_909),
.Y(n_1206)
);

INVx2_ASAP7_75t_L g1207 ( 
.A(n_963),
.Y(n_1207)
);

BUFx3_ASAP7_75t_L g1208 ( 
.A(n_992),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_968),
.Y(n_1209)
);

BUFx3_ASAP7_75t_L g1210 ( 
.A(n_1057),
.Y(n_1210)
);

AOI21xp5_ASAP7_75t_L g1211 ( 
.A1(n_985),
.A2(n_972),
.B(n_1009),
.Y(n_1211)
);

NAND2xp5_ASAP7_75t_L g1212 ( 
.A(n_1025),
.B(n_1022),
.Y(n_1212)
);

INVxp67_ASAP7_75t_SL g1213 ( 
.A(n_914),
.Y(n_1213)
);

NOR2xp33_ASAP7_75t_L g1214 ( 
.A(n_940),
.B(n_1024),
.Y(n_1214)
);

A2O1A1Ixp33_ASAP7_75t_L g1215 ( 
.A1(n_1022),
.A2(n_1035),
.B(n_956),
.C(n_1016),
.Y(n_1215)
);

OAI21x1_ASAP7_75t_L g1216 ( 
.A1(n_978),
.A2(n_953),
.B(n_927),
.Y(n_1216)
);

BUFx6f_ASAP7_75t_L g1217 ( 
.A(n_970),
.Y(n_1217)
);

AOI21xp5_ASAP7_75t_L g1218 ( 
.A1(n_1009),
.A2(n_914),
.B(n_954),
.Y(n_1218)
);

AOI22xp5_ASAP7_75t_L g1219 ( 
.A1(n_1024),
.A2(n_976),
.B1(n_1064),
.B2(n_1040),
.Y(n_1219)
);

BUFx3_ASAP7_75t_L g1220 ( 
.A(n_1057),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_942),
.A2(n_954),
.B(n_932),
.Y(n_1221)
);

NOR3xp33_ASAP7_75t_SL g1222 ( 
.A(n_903),
.B(n_907),
.C(n_904),
.Y(n_1222)
);

AOI21xp5_ASAP7_75t_L g1223 ( 
.A1(n_942),
.A2(n_954),
.B(n_937),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_969),
.Y(n_1224)
);

O2A1O1Ixp33_ASAP7_75t_L g1225 ( 
.A1(n_974),
.A2(n_997),
.B(n_910),
.C(n_1012),
.Y(n_1225)
);

BUFx2_ASAP7_75t_R g1226 ( 
.A(n_945),
.Y(n_1226)
);

NAND2xp5_ASAP7_75t_L g1227 ( 
.A(n_1027),
.B(n_893),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_893),
.B(n_921),
.Y(n_1228)
);

NOR2xp33_ASAP7_75t_L g1229 ( 
.A(n_921),
.B(n_1027),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_996),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1027),
.B(n_944),
.Y(n_1231)
);

AOI21xp5_ASAP7_75t_L g1232 ( 
.A1(n_942),
.A2(n_954),
.B(n_900),
.Y(n_1232)
);

BUFx3_ASAP7_75t_L g1233 ( 
.A(n_1173),
.Y(n_1233)
);

BUFx2_ASAP7_75t_L g1234 ( 
.A(n_1108),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1203),
.A2(n_926),
.B(n_1018),
.Y(n_1235)
);

AO32x2_ASAP7_75t_L g1236 ( 
.A1(n_1195),
.A2(n_1054),
.A3(n_1005),
.B1(n_900),
.B2(n_1007),
.Y(n_1236)
);

INVx1_ASAP7_75t_L g1237 ( 
.A(n_1073),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1080),
.Y(n_1238)
);

INVx1_ASAP7_75t_SL g1239 ( 
.A(n_1226),
.Y(n_1239)
);

CKINVDCx8_ASAP7_75t_R g1240 ( 
.A(n_1182),
.Y(n_1240)
);

CKINVDCx11_ASAP7_75t_R g1241 ( 
.A(n_1074),
.Y(n_1241)
);

OA21x2_ASAP7_75t_L g1242 ( 
.A1(n_1216),
.A2(n_998),
.B(n_987),
.Y(n_1242)
);

NAND3x1_ASAP7_75t_L g1243 ( 
.A(n_1072),
.B(n_935),
.C(n_1010),
.Y(n_1243)
);

OAI21x1_ASAP7_75t_L g1244 ( 
.A1(n_1203),
.A2(n_996),
.B(n_1018),
.Y(n_1244)
);

OAI21x1_ASAP7_75t_L g1245 ( 
.A1(n_1196),
.A2(n_1017),
.B(n_975),
.Y(n_1245)
);

OAI21xp5_ASAP7_75t_L g1246 ( 
.A1(n_1192),
.A2(n_998),
.B(n_987),
.Y(n_1246)
);

AOI21xp5_ASAP7_75t_L g1247 ( 
.A1(n_1096),
.A2(n_942),
.B(n_1007),
.Y(n_1247)
);

OAI21x1_ASAP7_75t_L g1248 ( 
.A1(n_1196),
.A2(n_1017),
.B(n_975),
.Y(n_1248)
);

NOR2xp33_ASAP7_75t_L g1249 ( 
.A(n_1081),
.B(n_1040),
.Y(n_1249)
);

INVx1_ASAP7_75t_L g1250 ( 
.A(n_1076),
.Y(n_1250)
);

INVx4_ASAP7_75t_L g1251 ( 
.A(n_1217),
.Y(n_1251)
);

OR2x2_ASAP7_75t_L g1252 ( 
.A(n_1070),
.B(n_1008),
.Y(n_1252)
);

AOI221xp5_ASAP7_75t_L g1253 ( 
.A1(n_1072),
.A2(n_1064),
.B1(n_1011),
.B2(n_950),
.C(n_945),
.Y(n_1253)
);

NAND2xp5_ASAP7_75t_L g1254 ( 
.A(n_1183),
.B(n_1116),
.Y(n_1254)
);

A2O1A1Ixp33_ASAP7_75t_L g1255 ( 
.A1(n_1071),
.A2(n_1079),
.B(n_1078),
.C(n_1084),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1145),
.Y(n_1256)
);

O2A1O1Ixp5_ASAP7_75t_L g1257 ( 
.A1(n_1084),
.A2(n_879),
.B(n_883),
.C(n_925),
.Y(n_1257)
);

NAND2xp5_ASAP7_75t_L g1258 ( 
.A(n_1185),
.B(n_1048),
.Y(n_1258)
);

INVx2_ASAP7_75t_L g1259 ( 
.A(n_1093),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1157),
.Y(n_1260)
);

OAI21x1_ASAP7_75t_L g1261 ( 
.A1(n_1202),
.A2(n_1015),
.B(n_883),
.Y(n_1261)
);

INVx3_ASAP7_75t_L g1262 ( 
.A(n_1143),
.Y(n_1262)
);

OA21x2_ASAP7_75t_L g1263 ( 
.A1(n_1077),
.A2(n_879),
.B(n_925),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_SL g1264 ( 
.A1(n_1097),
.A2(n_950),
.B1(n_1015),
.B2(n_1048),
.Y(n_1264)
);

NAND2xp5_ASAP7_75t_SL g1265 ( 
.A(n_1135),
.B(n_1005),
.Y(n_1265)
);

NAND2xp5_ASAP7_75t_SL g1266 ( 
.A(n_1214),
.B(n_1048),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1100),
.Y(n_1267)
);

OA21x2_ASAP7_75t_L g1268 ( 
.A1(n_1077),
.A2(n_905),
.B(n_970),
.Y(n_1268)
);

AO31x2_ASAP7_75t_L g1269 ( 
.A1(n_1174),
.A2(n_905),
.A3(n_970),
.B(n_1048),
.Y(n_1269)
);

O2A1O1Ixp33_ASAP7_75t_L g1270 ( 
.A1(n_1078),
.A2(n_905),
.B(n_970),
.C(n_1156),
.Y(n_1270)
);

NAND2xp5_ASAP7_75t_L g1271 ( 
.A(n_1213),
.B(n_905),
.Y(n_1271)
);

NAND2xp5_ASAP7_75t_L g1272 ( 
.A(n_1213),
.B(n_905),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1159),
.Y(n_1273)
);

AND2x2_ASAP7_75t_L g1274 ( 
.A(n_1154),
.B(n_1133),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_L g1275 ( 
.A(n_1177),
.B(n_1089),
.Y(n_1275)
);

O2A1O1Ixp5_ASAP7_75t_SL g1276 ( 
.A1(n_1109),
.A2(n_1161),
.B(n_1160),
.C(n_1098),
.Y(n_1276)
);

OAI22xp5_ASAP7_75t_L g1277 ( 
.A1(n_1232),
.A2(n_1223),
.B1(n_1187),
.B2(n_1219),
.Y(n_1277)
);

AOI21xp5_ASAP7_75t_L g1278 ( 
.A1(n_1223),
.A2(n_1172),
.B(n_1186),
.Y(n_1278)
);

BUFx4_ASAP7_75t_SL g1279 ( 
.A(n_1125),
.Y(n_1279)
);

AO31x2_ASAP7_75t_L g1280 ( 
.A1(n_1095),
.A2(n_1215),
.A3(n_1085),
.B(n_1171),
.Y(n_1280)
);

OAI21x1_ASAP7_75t_L g1281 ( 
.A1(n_1150),
.A2(n_1218),
.B(n_1225),
.Y(n_1281)
);

NAND2xp5_ASAP7_75t_L g1282 ( 
.A(n_1201),
.B(n_1091),
.Y(n_1282)
);

INVx2_ASAP7_75t_L g1283 ( 
.A(n_1114),
.Y(n_1283)
);

OR2x2_ASAP7_75t_L g1284 ( 
.A(n_1083),
.B(n_1129),
.Y(n_1284)
);

BUFx10_ASAP7_75t_L g1285 ( 
.A(n_1142),
.Y(n_1285)
);

BUFx12f_ASAP7_75t_L g1286 ( 
.A(n_1110),
.Y(n_1286)
);

AOI21xp5_ASAP7_75t_L g1287 ( 
.A1(n_1186),
.A2(n_1179),
.B(n_1079),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_1173),
.Y(n_1288)
);

AOI221xp5_ASAP7_75t_L g1289 ( 
.A1(n_1097),
.A2(n_1132),
.B1(n_1167),
.B2(n_1105),
.C(n_1082),
.Y(n_1289)
);

AO21x2_ASAP7_75t_L g1290 ( 
.A1(n_1102),
.A2(n_1222),
.B(n_1099),
.Y(n_1290)
);

INVx3_ASAP7_75t_L g1291 ( 
.A(n_1143),
.Y(n_1291)
);

NAND2xp5_ASAP7_75t_SL g1292 ( 
.A(n_1181),
.B(n_1086),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_1221),
.A2(n_1179),
.B(n_1140),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1184),
.B(n_1158),
.Y(n_1294)
);

OAI21x1_ASAP7_75t_L g1295 ( 
.A1(n_1120),
.A2(n_1212),
.B(n_1155),
.Y(n_1295)
);

NAND2xp5_ASAP7_75t_L g1296 ( 
.A(n_1229),
.B(n_1227),
.Y(n_1296)
);

BUFx2_ASAP7_75t_R g1297 ( 
.A(n_1208),
.Y(n_1297)
);

BUFx2_ASAP7_75t_L g1298 ( 
.A(n_1138),
.Y(n_1298)
);

OAI21xp5_ASAP7_75t_L g1299 ( 
.A1(n_1090),
.A2(n_1102),
.B(n_1171),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1162),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_SL g1301 ( 
.A(n_1198),
.B(n_1200),
.Y(n_1301)
);

INVx1_ASAP7_75t_L g1302 ( 
.A(n_1087),
.Y(n_1302)
);

NOR2xp33_ASAP7_75t_L g1303 ( 
.A(n_1176),
.B(n_1158),
.Y(n_1303)
);

AND2x2_ASAP7_75t_L g1304 ( 
.A(n_1088),
.B(n_1204),
.Y(n_1304)
);

AOI21xp5_ASAP7_75t_L g1305 ( 
.A1(n_1075),
.A2(n_1228),
.B(n_1231),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_1092),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1103),
.Y(n_1307)
);

NOR2xp33_ASAP7_75t_L g1308 ( 
.A(n_1156),
.B(n_1117),
.Y(n_1308)
);

OA21x2_ASAP7_75t_L g1309 ( 
.A1(n_1222),
.A2(n_1104),
.B(n_1178),
.Y(n_1309)
);

AND2x6_ASAP7_75t_L g1310 ( 
.A(n_1199),
.B(n_1197),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1194),
.B(n_1107),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1111),
.Y(n_1312)
);

O2A1O1Ixp33_ASAP7_75t_L g1313 ( 
.A1(n_1132),
.A2(n_1118),
.B(n_1119),
.C(n_1122),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1134),
.B(n_1152),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1101),
.B(n_1169),
.Y(n_1315)
);

NAND3xp33_ASAP7_75t_L g1316 ( 
.A(n_1168),
.B(n_1170),
.C(n_1112),
.Y(n_1316)
);

NAND2xp5_ASAP7_75t_SL g1317 ( 
.A(n_1139),
.B(n_1094),
.Y(n_1317)
);

NAND2xp5_ASAP7_75t_SL g1318 ( 
.A(n_1123),
.B(n_1147),
.Y(n_1318)
);

A2O1A1Ixp33_ASAP7_75t_L g1319 ( 
.A1(n_1104),
.A2(n_1170),
.B(n_1127),
.C(n_1146),
.Y(n_1319)
);

NAND2xp33_ASAP7_75t_L g1320 ( 
.A(n_1188),
.B(n_1217),
.Y(n_1320)
);

OAI21x1_ASAP7_75t_L g1321 ( 
.A1(n_1115),
.A2(n_1165),
.B(n_1151),
.Y(n_1321)
);

NOR2xp33_ASAP7_75t_L g1322 ( 
.A(n_1190),
.B(n_1224),
.Y(n_1322)
);

INVx1_ASAP7_75t_SL g1323 ( 
.A(n_1217),
.Y(n_1323)
);

AO31x2_ASAP7_75t_L g1324 ( 
.A1(n_1166),
.A2(n_1130),
.A3(n_1126),
.B(n_1124),
.Y(n_1324)
);

OAI21x1_ASAP7_75t_L g1325 ( 
.A1(n_1121),
.A2(n_1189),
.B(n_1163),
.Y(n_1325)
);

O2A1O1Ixp5_ASAP7_75t_L g1326 ( 
.A1(n_1131),
.A2(n_1206),
.B(n_1180),
.C(n_1141),
.Y(n_1326)
);

OA21x2_ASAP7_75t_L g1327 ( 
.A1(n_1230),
.A2(n_1137),
.B(n_1136),
.Y(n_1327)
);

NOR2xp33_ASAP7_75t_L g1328 ( 
.A(n_1205),
.B(n_1209),
.Y(n_1328)
);

AOI21xp5_ASAP7_75t_L g1329 ( 
.A1(n_1099),
.A2(n_1149),
.B(n_1207),
.Y(n_1329)
);

OAI21x1_ASAP7_75t_L g1330 ( 
.A1(n_1106),
.A2(n_1191),
.B(n_1128),
.Y(n_1330)
);

OAI22x1_ASAP7_75t_L g1331 ( 
.A1(n_1144),
.A2(n_1106),
.B1(n_1164),
.B2(n_1128),
.Y(n_1331)
);

AOI21xp5_ASAP7_75t_L g1332 ( 
.A1(n_1148),
.A2(n_1113),
.B(n_1164),
.Y(n_1332)
);

BUFx2_ASAP7_75t_R g1333 ( 
.A(n_1210),
.Y(n_1333)
);

BUFx2_ASAP7_75t_L g1334 ( 
.A(n_1113),
.Y(n_1334)
);

AOI22xp5_ASAP7_75t_L g1335 ( 
.A1(n_1113),
.A2(n_1168),
.B1(n_1220),
.B2(n_1175),
.Y(n_1335)
);

INVx2_ASAP7_75t_L g1336 ( 
.A(n_1153),
.Y(n_1336)
);

INVx1_ASAP7_75t_SL g1337 ( 
.A(n_1148),
.Y(n_1337)
);

AOI21xp5_ASAP7_75t_L g1338 ( 
.A1(n_1148),
.A2(n_591),
.B(n_1033),
.Y(n_1338)
);

AOI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1072),
.A2(n_1031),
.B1(n_1002),
.B2(n_890),
.Y(n_1339)
);

BUFx3_ASAP7_75t_L g1340 ( 
.A(n_1173),
.Y(n_1340)
);

BUFx2_ASAP7_75t_L g1341 ( 
.A(n_1108),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1192),
.A2(n_1193),
.B(n_1077),
.Y(n_1342)
);

OAI21xp5_ASAP7_75t_SL g1343 ( 
.A1(n_1072),
.A2(n_1031),
.B(n_1002),
.Y(n_1343)
);

BUFx12f_ASAP7_75t_L g1344 ( 
.A(n_1074),
.Y(n_1344)
);

AOI21xp5_ASAP7_75t_L g1345 ( 
.A1(n_1096),
.A2(n_591),
.B(n_1033),
.Y(n_1345)
);

AOI21x1_ASAP7_75t_L g1346 ( 
.A1(n_1203),
.A2(n_1211),
.B(n_1202),
.Y(n_1346)
);

AO31x2_ASAP7_75t_L g1347 ( 
.A1(n_1174),
.A2(n_1196),
.A3(n_1202),
.B(n_1095),
.Y(n_1347)
);

BUFx2_ASAP7_75t_L g1348 ( 
.A(n_1108),
.Y(n_1348)
);

AND2x4_ASAP7_75t_L g1349 ( 
.A(n_1198),
.B(n_990),
.Y(n_1349)
);

AOI21xp5_ASAP7_75t_L g1350 ( 
.A1(n_1096),
.A2(n_591),
.B(n_1033),
.Y(n_1350)
);

AND2x4_ASAP7_75t_L g1351 ( 
.A(n_1198),
.B(n_990),
.Y(n_1351)
);

OAI21x1_ASAP7_75t_L g1352 ( 
.A1(n_1203),
.A2(n_1202),
.B(n_1196),
.Y(n_1352)
);

NAND3x1_ASAP7_75t_L g1353 ( 
.A(n_1072),
.B(n_1031),
.C(n_1002),
.Y(n_1353)
);

NAND2xp5_ASAP7_75t_L g1354 ( 
.A(n_1183),
.B(n_890),
.Y(n_1354)
);

OAI21xp5_ASAP7_75t_L g1355 ( 
.A1(n_1192),
.A2(n_1193),
.B(n_1077),
.Y(n_1355)
);

NAND2xp5_ASAP7_75t_L g1356 ( 
.A(n_1183),
.B(n_890),
.Y(n_1356)
);

AOI21xp5_ASAP7_75t_L g1357 ( 
.A1(n_1096),
.A2(n_591),
.B(n_1033),
.Y(n_1357)
);

NAND2xp5_ASAP7_75t_L g1358 ( 
.A(n_1183),
.B(n_890),
.Y(n_1358)
);

BUFx2_ASAP7_75t_L g1359 ( 
.A(n_1108),
.Y(n_1359)
);

BUFx12f_ASAP7_75t_L g1360 ( 
.A(n_1074),
.Y(n_1360)
);

NAND2xp5_ASAP7_75t_L g1361 ( 
.A(n_1183),
.B(n_890),
.Y(n_1361)
);

AOI22xp5_ASAP7_75t_L g1362 ( 
.A1(n_1072),
.A2(n_1031),
.B1(n_1002),
.B2(n_890),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1154),
.B(n_888),
.Y(n_1363)
);

NAND2xp5_ASAP7_75t_L g1364 ( 
.A(n_1183),
.B(n_890),
.Y(n_1364)
);

AOI21xp5_ASAP7_75t_L g1365 ( 
.A1(n_1096),
.A2(n_591),
.B(n_1033),
.Y(n_1365)
);

AOI21xp5_ASAP7_75t_L g1366 ( 
.A1(n_1096),
.A2(n_591),
.B(n_1033),
.Y(n_1366)
);

INVx2_ASAP7_75t_L g1367 ( 
.A(n_1080),
.Y(n_1367)
);

AND2x4_ASAP7_75t_L g1368 ( 
.A(n_1198),
.B(n_990),
.Y(n_1368)
);

INVx5_ASAP7_75t_L g1369 ( 
.A(n_1217),
.Y(n_1369)
);

INVxp67_ASAP7_75t_SL g1370 ( 
.A(n_1213),
.Y(n_1370)
);

AO32x2_ASAP7_75t_L g1371 ( 
.A1(n_1195),
.A2(n_1085),
.A3(n_1095),
.B1(n_1098),
.B2(n_1109),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_L g1372 ( 
.A(n_1183),
.B(n_890),
.Y(n_1372)
);

INVx2_ASAP7_75t_SL g1373 ( 
.A(n_1173),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1080),
.Y(n_1374)
);

AOI21x1_ASAP7_75t_L g1375 ( 
.A1(n_1203),
.A2(n_1211),
.B(n_1202),
.Y(n_1375)
);

AO32x2_ASAP7_75t_L g1376 ( 
.A1(n_1195),
.A2(n_1085),
.A3(n_1095),
.B1(n_1098),
.B2(n_1109),
.Y(n_1376)
);

AOI21xp5_ASAP7_75t_SL g1377 ( 
.A1(n_1195),
.A2(n_1096),
.B(n_1232),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1203),
.A2(n_1202),
.B(n_1196),
.Y(n_1378)
);

BUFx2_ASAP7_75t_L g1379 ( 
.A(n_1108),
.Y(n_1379)
);

AND2x4_ASAP7_75t_L g1380 ( 
.A(n_1198),
.B(n_990),
.Y(n_1380)
);

AND2x4_ASAP7_75t_L g1381 ( 
.A(n_1198),
.B(n_990),
.Y(n_1381)
);

AOI21xp5_ASAP7_75t_L g1382 ( 
.A1(n_1096),
.A2(n_591),
.B(n_1033),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1154),
.B(n_888),
.Y(n_1383)
);

NAND2x1p5_ASAP7_75t_L g1384 ( 
.A(n_1143),
.B(n_929),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1183),
.B(n_890),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_L g1386 ( 
.A(n_1183),
.B(n_890),
.Y(n_1386)
);

BUFx2_ASAP7_75t_L g1387 ( 
.A(n_1108),
.Y(n_1387)
);

NAND2xp5_ASAP7_75t_L g1388 ( 
.A(n_1183),
.B(n_890),
.Y(n_1388)
);

INVx3_ASAP7_75t_L g1389 ( 
.A(n_1143),
.Y(n_1389)
);

OA21x2_ASAP7_75t_L g1390 ( 
.A1(n_1278),
.A2(n_1287),
.B(n_1299),
.Y(n_1390)
);

BUFx8_ASAP7_75t_L g1391 ( 
.A(n_1286),
.Y(n_1391)
);

AOI22xp5_ASAP7_75t_L g1392 ( 
.A1(n_1343),
.A2(n_1353),
.B1(n_1362),
.B2(n_1339),
.Y(n_1392)
);

O2A1O1Ixp33_ASAP7_75t_L g1393 ( 
.A1(n_1343),
.A2(n_1319),
.B(n_1292),
.C(n_1255),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1237),
.Y(n_1394)
);

OAI21x1_ASAP7_75t_L g1395 ( 
.A1(n_1281),
.A2(n_1375),
.B(n_1346),
.Y(n_1395)
);

INVx2_ASAP7_75t_SL g1396 ( 
.A(n_1284),
.Y(n_1396)
);

INVxp67_ASAP7_75t_L g1397 ( 
.A(n_1294),
.Y(n_1397)
);

CKINVDCx11_ASAP7_75t_R g1398 ( 
.A(n_1241),
.Y(n_1398)
);

INVx2_ASAP7_75t_L g1399 ( 
.A(n_1327),
.Y(n_1399)
);

INVx1_ASAP7_75t_SL g1400 ( 
.A(n_1234),
.Y(n_1400)
);

INVx3_ASAP7_75t_L g1401 ( 
.A(n_1262),
.Y(n_1401)
);

INVx1_ASAP7_75t_L g1402 ( 
.A(n_1250),
.Y(n_1402)
);

AOI22xp33_ASAP7_75t_L g1403 ( 
.A1(n_1289),
.A2(n_1315),
.B1(n_1316),
.B2(n_1308),
.Y(n_1403)
);

NAND2xp5_ASAP7_75t_L g1404 ( 
.A(n_1275),
.B(n_1363),
.Y(n_1404)
);

O2A1O1Ixp33_ASAP7_75t_SL g1405 ( 
.A1(n_1254),
.A2(n_1289),
.B(n_1317),
.C(n_1313),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1370),
.Y(n_1406)
);

OAI22xp5_ASAP7_75t_L g1407 ( 
.A1(n_1354),
.A2(n_1364),
.B1(n_1388),
.B2(n_1356),
.Y(n_1407)
);

NAND2xp5_ASAP7_75t_L g1408 ( 
.A(n_1275),
.B(n_1383),
.Y(n_1408)
);

O2A1O1Ixp5_ASAP7_75t_L g1409 ( 
.A1(n_1278),
.A2(n_1299),
.B(n_1338),
.C(n_1332),
.Y(n_1409)
);

OAI21x1_ASAP7_75t_L g1410 ( 
.A1(n_1235),
.A2(n_1244),
.B(n_1352),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1341),
.Y(n_1412)
);

AO31x2_ASAP7_75t_L g1413 ( 
.A1(n_1277),
.A2(n_1329),
.A3(n_1305),
.B(n_1382),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1256),
.Y(n_1414)
);

OR2x6_ASAP7_75t_L g1415 ( 
.A(n_1377),
.B(n_1264),
.Y(n_1415)
);

INVx2_ASAP7_75t_SL g1416 ( 
.A(n_1348),
.Y(n_1416)
);

BUFx3_ASAP7_75t_L g1417 ( 
.A(n_1359),
.Y(n_1417)
);

OAI21x1_ASAP7_75t_L g1418 ( 
.A1(n_1378),
.A2(n_1329),
.B(n_1248),
.Y(n_1418)
);

NOR2xp33_ASAP7_75t_L g1419 ( 
.A(n_1354),
.B(n_1356),
.Y(n_1419)
);

HB1xp67_ASAP7_75t_L g1420 ( 
.A(n_1327),
.Y(n_1420)
);

OAI22xp5_ASAP7_75t_L g1421 ( 
.A1(n_1358),
.A2(n_1385),
.B1(n_1388),
.B2(n_1372),
.Y(n_1421)
);

AO31x2_ASAP7_75t_L g1422 ( 
.A1(n_1277),
.A2(n_1305),
.A3(n_1365),
.B(n_1345),
.Y(n_1422)
);

CKINVDCx20_ASAP7_75t_R g1423 ( 
.A(n_1288),
.Y(n_1423)
);

OAI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1358),
.A2(n_1372),
.B1(n_1364),
.B2(n_1361),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1276),
.A2(n_1357),
.B(n_1366),
.Y(n_1425)
);

INVx2_ASAP7_75t_SL g1426 ( 
.A(n_1379),
.Y(n_1426)
);

OAI21x1_ASAP7_75t_L g1427 ( 
.A1(n_1245),
.A2(n_1261),
.B(n_1295),
.Y(n_1427)
);

INVx1_ASAP7_75t_L g1428 ( 
.A(n_1260),
.Y(n_1428)
);

AOI22xp5_ASAP7_75t_L g1429 ( 
.A1(n_1249),
.A2(n_1314),
.B1(n_1311),
.B2(n_1318),
.Y(n_1429)
);

OAI21x1_ASAP7_75t_L g1430 ( 
.A1(n_1293),
.A2(n_1247),
.B(n_1342),
.Y(n_1430)
);

INVx1_ASAP7_75t_L g1431 ( 
.A(n_1273),
.Y(n_1431)
);

BUFx6f_ASAP7_75t_L g1432 ( 
.A(n_1369),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1300),
.Y(n_1433)
);

AOI222xp33_ASAP7_75t_L g1434 ( 
.A1(n_1361),
.A2(n_1385),
.B1(n_1386),
.B2(n_1301),
.C1(n_1334),
.C2(n_1310),
.Y(n_1434)
);

OAI21x1_ASAP7_75t_L g1435 ( 
.A1(n_1355),
.A2(n_1350),
.B(n_1366),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1302),
.Y(n_1436)
);

AND2x4_ASAP7_75t_L g1437 ( 
.A(n_1349),
.B(n_1351),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1279),
.Y(n_1438)
);

AOI22xp5_ASAP7_75t_L g1439 ( 
.A1(n_1335),
.A2(n_1303),
.B1(n_1386),
.B2(n_1310),
.Y(n_1439)
);

OA21x2_ASAP7_75t_L g1440 ( 
.A1(n_1246),
.A2(n_1332),
.B(n_1257),
.Y(n_1440)
);

OA21x2_ASAP7_75t_L g1441 ( 
.A1(n_1337),
.A2(n_1254),
.B(n_1253),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1321),
.Y(n_1442)
);

BUFx3_ASAP7_75t_L g1443 ( 
.A(n_1387),
.Y(n_1443)
);

OAI21x1_ASAP7_75t_L g1444 ( 
.A1(n_1270),
.A2(n_1268),
.B(n_1330),
.Y(n_1444)
);

NAND2x1p5_ASAP7_75t_L g1445 ( 
.A(n_1369),
.B(n_1266),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_1306),
.Y(n_1446)
);

INVx2_ASAP7_75t_L g1447 ( 
.A(n_1325),
.Y(n_1447)
);

INVx2_ASAP7_75t_L g1448 ( 
.A(n_1238),
.Y(n_1448)
);

OA21x2_ASAP7_75t_L g1449 ( 
.A1(n_1337),
.A2(n_1272),
.B(n_1271),
.Y(n_1449)
);

OAI21x1_ASAP7_75t_L g1450 ( 
.A1(n_1268),
.A2(n_1243),
.B(n_1263),
.Y(n_1450)
);

INVx1_ASAP7_75t_L g1451 ( 
.A(n_1307),
.Y(n_1451)
);

OA21x2_ASAP7_75t_L g1452 ( 
.A1(n_1326),
.A2(n_1282),
.B(n_1296),
.Y(n_1452)
);

HB1xp67_ASAP7_75t_L g1453 ( 
.A(n_1269),
.Y(n_1453)
);

OAI21x1_ASAP7_75t_L g1454 ( 
.A1(n_1263),
.A2(n_1242),
.B(n_1309),
.Y(n_1454)
);

BUFx3_ASAP7_75t_L g1455 ( 
.A(n_1368),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1368),
.B(n_1381),
.Y(n_1456)
);

OAI21x1_ASAP7_75t_L g1457 ( 
.A1(n_1309),
.A2(n_1296),
.B(n_1258),
.Y(n_1457)
);

OAI21x1_ASAP7_75t_L g1458 ( 
.A1(n_1384),
.A2(n_1312),
.B(n_1267),
.Y(n_1458)
);

BUFx2_ASAP7_75t_L g1459 ( 
.A(n_1298),
.Y(n_1459)
);

AND2x4_ASAP7_75t_L g1460 ( 
.A(n_1380),
.B(n_1381),
.Y(n_1460)
);

INVx1_ASAP7_75t_L g1461 ( 
.A(n_1259),
.Y(n_1461)
);

OAI21x1_ASAP7_75t_L g1462 ( 
.A1(n_1384),
.A2(n_1283),
.B(n_1374),
.Y(n_1462)
);

CKINVDCx5p33_ASAP7_75t_R g1463 ( 
.A(n_1344),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1367),
.A2(n_1252),
.B(n_1336),
.Y(n_1464)
);

BUFx12f_ASAP7_75t_L g1465 ( 
.A(n_1360),
.Y(n_1465)
);

OAI221xp5_ASAP7_75t_SL g1466 ( 
.A1(n_1239),
.A2(n_1373),
.B1(n_1233),
.B2(n_1340),
.C(n_1376),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1322),
.Y(n_1467)
);

NAND2xp5_ASAP7_75t_SL g1468 ( 
.A(n_1285),
.B(n_1331),
.Y(n_1468)
);

OAI21x1_ASAP7_75t_L g1469 ( 
.A1(n_1262),
.A2(n_1389),
.B(n_1291),
.Y(n_1469)
);

BUFx12f_ASAP7_75t_L g1470 ( 
.A(n_1251),
.Y(n_1470)
);

OAI22xp5_ASAP7_75t_L g1471 ( 
.A1(n_1265),
.A2(n_1240),
.B1(n_1328),
.B2(n_1239),
.Y(n_1471)
);

AOI22xp33_ASAP7_75t_L g1472 ( 
.A1(n_1310),
.A2(n_1290),
.B1(n_1371),
.B2(n_1376),
.Y(n_1472)
);

INVx2_ASAP7_75t_L g1473 ( 
.A(n_1324),
.Y(n_1473)
);

INVx6_ASAP7_75t_L g1474 ( 
.A(n_1369),
.Y(n_1474)
);

BUFx2_ASAP7_75t_L g1475 ( 
.A(n_1323),
.Y(n_1475)
);

INVx2_ASAP7_75t_L g1476 ( 
.A(n_1324),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1310),
.B(n_1323),
.Y(n_1477)
);

OAI22xp33_ASAP7_75t_SL g1478 ( 
.A1(n_1371),
.A2(n_1376),
.B1(n_1369),
.B2(n_1251),
.Y(n_1478)
);

AO21x2_ASAP7_75t_L g1479 ( 
.A1(n_1290),
.A2(n_1371),
.B(n_1280),
.Y(n_1479)
);

OAI221xp5_ASAP7_75t_SL g1480 ( 
.A1(n_1280),
.A2(n_1297),
.B1(n_1333),
.B2(n_1236),
.C(n_1347),
.Y(n_1480)
);

AO21x2_ASAP7_75t_L g1481 ( 
.A1(n_1280),
.A2(n_1347),
.B(n_1236),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1269),
.Y(n_1482)
);

OAI21x1_ASAP7_75t_L g1483 ( 
.A1(n_1347),
.A2(n_1269),
.B(n_1236),
.Y(n_1483)
);

NAND2xp5_ASAP7_75t_L g1484 ( 
.A(n_1320),
.B(n_1297),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1333),
.Y(n_1485)
);

AO31x2_ASAP7_75t_L g1486 ( 
.A1(n_1255),
.A2(n_1287),
.A3(n_1278),
.B(n_1277),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1237),
.Y(n_1487)
);

AOI22xp5_ASAP7_75t_L g1488 ( 
.A1(n_1343),
.A2(n_1031),
.B1(n_1002),
.B2(n_1353),
.Y(n_1488)
);

NOR2xp33_ASAP7_75t_L g1489 ( 
.A(n_1343),
.B(n_1063),
.Y(n_1489)
);

AND2x2_ASAP7_75t_L g1490 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1237),
.Y(n_1491)
);

INVx1_ASAP7_75t_L g1492 ( 
.A(n_1237),
.Y(n_1492)
);

OAI21x1_ASAP7_75t_L g1493 ( 
.A1(n_1281),
.A2(n_1375),
.B(n_1346),
.Y(n_1493)
);

NAND2xp5_ASAP7_75t_L g1494 ( 
.A(n_1275),
.B(n_1363),
.Y(n_1494)
);

OR2x6_ASAP7_75t_L g1495 ( 
.A(n_1377),
.B(n_1232),
.Y(n_1495)
);

BUFx2_ASAP7_75t_L g1496 ( 
.A(n_1234),
.Y(n_1496)
);

OR2x2_ASAP7_75t_L g1497 ( 
.A(n_1275),
.B(n_1284),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1327),
.Y(n_1498)
);

NOR2xp33_ASAP7_75t_L g1499 ( 
.A(n_1343),
.B(n_1063),
.Y(n_1499)
);

INVx3_ASAP7_75t_L g1500 ( 
.A(n_1262),
.Y(n_1500)
);

AO21x1_ASAP7_75t_L g1501 ( 
.A1(n_1343),
.A2(n_1063),
.B(n_1339),
.Y(n_1501)
);

AOI22xp33_ASAP7_75t_L g1502 ( 
.A1(n_1289),
.A2(n_1072),
.B1(n_1063),
.B2(n_1002),
.Y(n_1502)
);

AO31x2_ASAP7_75t_L g1503 ( 
.A1(n_1255),
.A2(n_1287),
.A3(n_1278),
.B(n_1277),
.Y(n_1503)
);

AO221x2_ASAP7_75t_L g1504 ( 
.A1(n_1343),
.A2(n_890),
.B1(n_1167),
.B2(n_1316),
.C(n_1063),
.Y(n_1504)
);

INVx3_ASAP7_75t_L g1505 ( 
.A(n_1262),
.Y(n_1505)
);

BUFx12f_ASAP7_75t_L g1506 ( 
.A(n_1241),
.Y(n_1506)
);

AOI22xp5_ASAP7_75t_L g1507 ( 
.A1(n_1343),
.A2(n_1031),
.B1(n_1002),
.B2(n_1353),
.Y(n_1507)
);

OAI22xp33_ASAP7_75t_L g1508 ( 
.A1(n_1339),
.A2(n_1362),
.B1(n_1063),
.B2(n_1343),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1237),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_1237),
.Y(n_1510)
);

HB1xp67_ASAP7_75t_L g1511 ( 
.A(n_1370),
.Y(n_1511)
);

OA21x2_ASAP7_75t_L g1512 ( 
.A1(n_1278),
.A2(n_1287),
.B(n_1299),
.Y(n_1512)
);

BUFx8_ASAP7_75t_L g1513 ( 
.A(n_1286),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1275),
.B(n_1363),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1237),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1237),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1237),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1275),
.B(n_1363),
.Y(n_1520)
);

A2O1A1Ixp33_ASAP7_75t_L g1521 ( 
.A1(n_1343),
.A2(n_1063),
.B(n_1362),
.C(n_1339),
.Y(n_1521)
);

NOR2xp33_ASAP7_75t_SL g1522 ( 
.A(n_1333),
.B(n_504),
.Y(n_1522)
);

INVx1_ASAP7_75t_L g1523 ( 
.A(n_1237),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1327),
.Y(n_1524)
);

AOI22xp33_ASAP7_75t_L g1525 ( 
.A1(n_1289),
.A2(n_1072),
.B1(n_1063),
.B2(n_1002),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1237),
.Y(n_1526)
);

INVx2_ASAP7_75t_L g1527 ( 
.A(n_1327),
.Y(n_1527)
);

BUFx2_ASAP7_75t_L g1528 ( 
.A(n_1234),
.Y(n_1528)
);

NOR2xp33_ASAP7_75t_SL g1529 ( 
.A(n_1333),
.B(n_504),
.Y(n_1529)
);

AND2x2_ASAP7_75t_L g1530 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1237),
.Y(n_1531)
);

AND2x2_ASAP7_75t_L g1532 ( 
.A(n_1274),
.B(n_1304),
.Y(n_1532)
);

NOR2xp33_ASAP7_75t_L g1533 ( 
.A(n_1343),
.B(n_1063),
.Y(n_1533)
);

NAND2xp5_ASAP7_75t_L g1534 ( 
.A(n_1404),
.B(n_1408),
.Y(n_1534)
);

NOR2xp33_ASAP7_75t_R g1535 ( 
.A(n_1522),
.B(n_1529),
.Y(n_1535)
);

OAI22xp5_ASAP7_75t_L g1536 ( 
.A1(n_1403),
.A2(n_1507),
.B1(n_1488),
.B2(n_1525),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1406),
.Y(n_1537)
);

AOI21x1_ASAP7_75t_SL g1538 ( 
.A1(n_1477),
.A2(n_1453),
.B(n_1484),
.Y(n_1538)
);

AND2x2_ASAP7_75t_L g1539 ( 
.A(n_1411),
.B(n_1490),
.Y(n_1539)
);

INVx1_ASAP7_75t_L g1540 ( 
.A(n_1511),
.Y(n_1540)
);

OAI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1403),
.A2(n_1502),
.B1(n_1525),
.B2(n_1429),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1497),
.B(n_1494),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1515),
.B(n_1518),
.Y(n_1543)
);

AOI21x1_ASAP7_75t_SL g1544 ( 
.A1(n_1453),
.A2(n_1520),
.B(n_1514),
.Y(n_1544)
);

AND2x2_ASAP7_75t_L g1545 ( 
.A(n_1530),
.B(n_1532),
.Y(n_1545)
);

INVx2_ASAP7_75t_L g1546 ( 
.A(n_1399),
.Y(n_1546)
);

OAI22xp5_ASAP7_75t_L g1547 ( 
.A1(n_1502),
.A2(n_1415),
.B1(n_1439),
.B2(n_1392),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1415),
.A2(n_1467),
.B1(n_1419),
.B2(n_1471),
.Y(n_1548)
);

O2A1O1Ixp33_ASAP7_75t_L g1549 ( 
.A1(n_1521),
.A2(n_1508),
.B(n_1405),
.C(n_1533),
.Y(n_1549)
);

O2A1O1Ixp5_ASAP7_75t_L g1550 ( 
.A1(n_1425),
.A2(n_1409),
.B(n_1501),
.C(n_1508),
.Y(n_1550)
);

AOI21xp5_ASAP7_75t_L g1551 ( 
.A1(n_1495),
.A2(n_1415),
.B(n_1390),
.Y(n_1551)
);

OA21x2_ASAP7_75t_L g1552 ( 
.A1(n_1430),
.A2(n_1435),
.B(n_1395),
.Y(n_1552)
);

NAND2xp5_ASAP7_75t_L g1553 ( 
.A(n_1419),
.B(n_1407),
.Y(n_1553)
);

AND2x4_ASAP7_75t_L g1554 ( 
.A(n_1455),
.B(n_1437),
.Y(n_1554)
);

NAND2xp5_ASAP7_75t_L g1555 ( 
.A(n_1421),
.B(n_1424),
.Y(n_1555)
);

HB1xp67_ASAP7_75t_L g1556 ( 
.A(n_1420),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1498),
.Y(n_1557)
);

INVx1_ASAP7_75t_L g1558 ( 
.A(n_1511),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1489),
.B(n_1499),
.Y(n_1559)
);

BUFx6f_ASAP7_75t_SL g1560 ( 
.A(n_1412),
.Y(n_1560)
);

O2A1O1Ixp5_ASAP7_75t_L g1561 ( 
.A1(n_1521),
.A2(n_1533),
.B(n_1489),
.C(n_1499),
.Y(n_1561)
);

NOR2x1_ASAP7_75t_SL g1562 ( 
.A(n_1495),
.B(n_1468),
.Y(n_1562)
);

AND2x2_ASAP7_75t_L g1563 ( 
.A(n_1460),
.B(n_1456),
.Y(n_1563)
);

AOI21xp5_ASAP7_75t_L g1564 ( 
.A1(n_1495),
.A2(n_1390),
.B(n_1512),
.Y(n_1564)
);

BUFx12f_ASAP7_75t_L g1565 ( 
.A(n_1398),
.Y(n_1565)
);

OA21x2_ASAP7_75t_L g1566 ( 
.A1(n_1430),
.A2(n_1435),
.B(n_1493),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1393),
.A2(n_1432),
.B(n_1441),
.Y(n_1567)
);

NAND2xp5_ASAP7_75t_L g1568 ( 
.A(n_1396),
.B(n_1397),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1504),
.B(n_1434),
.Y(n_1569)
);

AOI21x1_ASAP7_75t_SL g1570 ( 
.A1(n_1420),
.A2(n_1504),
.B(n_1405),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1394),
.Y(n_1571)
);

OR2x2_ASAP7_75t_L g1572 ( 
.A(n_1459),
.B(n_1402),
.Y(n_1572)
);

AND2x2_ASAP7_75t_L g1573 ( 
.A(n_1504),
.B(n_1475),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1524),
.Y(n_1574)
);

CKINVDCx5p33_ASAP7_75t_R g1575 ( 
.A(n_1438),
.Y(n_1575)
);

AOI21x1_ASAP7_75t_SL g1576 ( 
.A1(n_1466),
.A2(n_1480),
.B(n_1478),
.Y(n_1576)
);

NAND2xp5_ASAP7_75t_L g1577 ( 
.A(n_1461),
.B(n_1448),
.Y(n_1577)
);

O2A1O1Ixp33_ASAP7_75t_L g1578 ( 
.A1(n_1468),
.A2(n_1426),
.B(n_1416),
.C(n_1400),
.Y(n_1578)
);

OR2x2_ASAP7_75t_L g1579 ( 
.A(n_1414),
.B(n_1428),
.Y(n_1579)
);

NAND2xp5_ASAP7_75t_L g1580 ( 
.A(n_1448),
.B(n_1496),
.Y(n_1580)
);

AND2x2_ASAP7_75t_L g1581 ( 
.A(n_1464),
.B(n_1431),
.Y(n_1581)
);

AND2x2_ASAP7_75t_L g1582 ( 
.A(n_1531),
.B(n_1433),
.Y(n_1582)
);

OR2x2_ASAP7_75t_L g1583 ( 
.A(n_1436),
.B(n_1446),
.Y(n_1583)
);

AND2x4_ASAP7_75t_L g1584 ( 
.A(n_1417),
.B(n_1443),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1451),
.B(n_1487),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1491),
.Y(n_1586)
);

CKINVDCx14_ASAP7_75t_R g1587 ( 
.A(n_1438),
.Y(n_1587)
);

NAND2xp5_ASAP7_75t_L g1588 ( 
.A(n_1528),
.B(n_1492),
.Y(n_1588)
);

AND2x2_ASAP7_75t_L g1589 ( 
.A(n_1509),
.B(n_1510),
.Y(n_1589)
);

INVx1_ASAP7_75t_L g1590 ( 
.A(n_1516),
.Y(n_1590)
);

HB1xp67_ASAP7_75t_L g1591 ( 
.A(n_1527),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1517),
.B(n_1519),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1523),
.B(n_1526),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1485),
.B(n_1500),
.Y(n_1594)
);

NOR2xp33_ASAP7_75t_L g1595 ( 
.A(n_1445),
.B(n_1485),
.Y(n_1595)
);

AND2x4_ASAP7_75t_L g1596 ( 
.A(n_1401),
.B(n_1505),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1527),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1470),
.Y(n_1598)
);

BUFx3_ASAP7_75t_L g1599 ( 
.A(n_1474),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_L g1600 ( 
.A(n_1452),
.B(n_1503),
.Y(n_1600)
);

OAI22xp5_ASAP7_75t_L g1601 ( 
.A1(n_1472),
.A2(n_1445),
.B1(n_1474),
.B2(n_1452),
.Y(n_1601)
);

OAI22xp5_ASAP7_75t_L g1602 ( 
.A1(n_1474),
.A2(n_1441),
.B1(n_1505),
.B2(n_1401),
.Y(n_1602)
);

OR2x2_ASAP7_75t_L g1603 ( 
.A(n_1486),
.B(n_1503),
.Y(n_1603)
);

HB1xp67_ASAP7_75t_L g1604 ( 
.A(n_1473),
.Y(n_1604)
);

AOI21x1_ASAP7_75t_SL g1605 ( 
.A1(n_1486),
.A2(n_1503),
.B(n_1457),
.Y(n_1605)
);

OR2x2_ASAP7_75t_L g1606 ( 
.A(n_1486),
.B(n_1449),
.Y(n_1606)
);

OAI22xp5_ASAP7_75t_L g1607 ( 
.A1(n_1432),
.A2(n_1423),
.B1(n_1463),
.B2(n_1482),
.Y(n_1607)
);

OAI22xp5_ASAP7_75t_L g1608 ( 
.A1(n_1432),
.A2(n_1423),
.B1(n_1463),
.B2(n_1476),
.Y(n_1608)
);

AND2x2_ASAP7_75t_L g1609 ( 
.A(n_1458),
.B(n_1486),
.Y(n_1609)
);

AND2x4_ASAP7_75t_L g1610 ( 
.A(n_1458),
.B(n_1469),
.Y(n_1610)
);

BUFx2_ASAP7_75t_L g1611 ( 
.A(n_1469),
.Y(n_1611)
);

HB1xp67_ASAP7_75t_L g1612 ( 
.A(n_1473),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1398),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1449),
.B(n_1422),
.Y(n_1614)
);

AND2x2_ASAP7_75t_L g1615 ( 
.A(n_1462),
.B(n_1422),
.Y(n_1615)
);

AND2x2_ASAP7_75t_L g1616 ( 
.A(n_1422),
.B(n_1481),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_L g1617 ( 
.A(n_1413),
.B(n_1479),
.Y(n_1617)
);

O2A1O1Ixp5_ASAP7_75t_L g1618 ( 
.A1(n_1442),
.A2(n_1447),
.B(n_1440),
.C(n_1413),
.Y(n_1618)
);

OAI22xp5_ASAP7_75t_L g1619 ( 
.A1(n_1465),
.A2(n_1506),
.B1(n_1447),
.B2(n_1513),
.Y(n_1619)
);

AOI21xp5_ASAP7_75t_SL g1620 ( 
.A1(n_1479),
.A2(n_1391),
.B(n_1513),
.Y(n_1620)
);

OAI22xp5_ASAP7_75t_L g1621 ( 
.A1(n_1465),
.A2(n_1506),
.B1(n_1513),
.B2(n_1391),
.Y(n_1621)
);

AND2x2_ASAP7_75t_L g1622 ( 
.A(n_1483),
.B(n_1413),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1391),
.A2(n_1444),
.B1(n_1450),
.B2(n_1454),
.Y(n_1623)
);

OAI22xp5_ASAP7_75t_L g1624 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1507),
.B2(n_1488),
.Y(n_1624)
);

OR2x2_ASAP7_75t_L g1625 ( 
.A(n_1410),
.B(n_1427),
.Y(n_1625)
);

CKINVDCx6p67_ASAP7_75t_R g1626 ( 
.A(n_1427),
.Y(n_1626)
);

OAI22xp5_ASAP7_75t_L g1627 ( 
.A1(n_1418),
.A2(n_1403),
.B1(n_1507),
.B2(n_1488),
.Y(n_1627)
);

OA22x2_ASAP7_75t_L g1628 ( 
.A1(n_1488),
.A2(n_1507),
.B1(n_1362),
.B2(n_1339),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1404),
.B(n_1408),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1497),
.B(n_1404),
.Y(n_1630)
);

AND2x2_ASAP7_75t_L g1631 ( 
.A(n_1411),
.B(n_1490),
.Y(n_1631)
);

OAI22xp5_ASAP7_75t_L g1632 ( 
.A1(n_1403),
.A2(n_1507),
.B1(n_1488),
.B2(n_1339),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1404),
.B(n_1408),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1411),
.B(n_1490),
.Y(n_1634)
);

AOI21x1_ASAP7_75t_SL g1635 ( 
.A1(n_1477),
.A2(n_1063),
.B(n_1354),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1404),
.B(n_1408),
.Y(n_1636)
);

AND2x4_ASAP7_75t_L g1637 ( 
.A(n_1455),
.B(n_1437),
.Y(n_1637)
);

AOI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1495),
.A2(n_890),
.B(n_1033),
.Y(n_1638)
);

OAI22xp5_ASAP7_75t_L g1639 ( 
.A1(n_1403),
.A2(n_1507),
.B1(n_1488),
.B2(n_1339),
.Y(n_1639)
);

BUFx10_ASAP7_75t_L g1640 ( 
.A(n_1438),
.Y(n_1640)
);

HB1xp67_ASAP7_75t_L g1641 ( 
.A(n_1420),
.Y(n_1641)
);

CKINVDCx5p33_ASAP7_75t_R g1642 ( 
.A(n_1438),
.Y(n_1642)
);

BUFx2_ASAP7_75t_L g1643 ( 
.A(n_1437),
.Y(n_1643)
);

OR2x2_ASAP7_75t_L g1644 ( 
.A(n_1497),
.B(n_1404),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1411),
.B(n_1490),
.Y(n_1645)
);

O2A1O1Ixp33_ASAP7_75t_L g1646 ( 
.A1(n_1521),
.A2(n_1343),
.B(n_1063),
.C(n_1031),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1574),
.Y(n_1647)
);

OAI21xp5_ASAP7_75t_L g1648 ( 
.A1(n_1646),
.A2(n_1549),
.B(n_1561),
.Y(n_1648)
);

INVx1_ASAP7_75t_L g1649 ( 
.A(n_1574),
.Y(n_1649)
);

AND2x2_ASAP7_75t_L g1650 ( 
.A(n_1573),
.B(n_1622),
.Y(n_1650)
);

INVx1_ASAP7_75t_L g1651 ( 
.A(n_1591),
.Y(n_1651)
);

OR2x6_ASAP7_75t_L g1652 ( 
.A(n_1551),
.B(n_1564),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1591),
.Y(n_1653)
);

INVx1_ASAP7_75t_SL g1654 ( 
.A(n_1572),
.Y(n_1654)
);

BUFx3_ASAP7_75t_L g1655 ( 
.A(n_1611),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1616),
.B(n_1559),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1604),
.Y(n_1657)
);

OR2x2_ASAP7_75t_L g1658 ( 
.A(n_1603),
.B(n_1606),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1604),
.Y(n_1659)
);

INVx1_ASAP7_75t_L g1660 ( 
.A(n_1612),
.Y(n_1660)
);

BUFx4f_ASAP7_75t_SL g1661 ( 
.A(n_1565),
.Y(n_1661)
);

INVx2_ASAP7_75t_L g1662 ( 
.A(n_1546),
.Y(n_1662)
);

AND2x2_ASAP7_75t_L g1663 ( 
.A(n_1609),
.B(n_1581),
.Y(n_1663)
);

BUFx4f_ASAP7_75t_SL g1664 ( 
.A(n_1565),
.Y(n_1664)
);

BUFx2_ASAP7_75t_L g1665 ( 
.A(n_1556),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_L g1666 ( 
.A(n_1553),
.B(n_1555),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1641),
.B(n_1614),
.Y(n_1667)
);

AOI22xp33_ASAP7_75t_L g1668 ( 
.A1(n_1536),
.A2(n_1628),
.B1(n_1541),
.B2(n_1632),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1597),
.Y(n_1669)
);

BUFx2_ASAP7_75t_SL g1670 ( 
.A(n_1560),
.Y(n_1670)
);

OR2x2_ASAP7_75t_L g1671 ( 
.A(n_1641),
.B(n_1600),
.Y(n_1671)
);

BUFx3_ASAP7_75t_L g1672 ( 
.A(n_1599),
.Y(n_1672)
);

BUFx12f_ASAP7_75t_L g1673 ( 
.A(n_1575),
.Y(n_1673)
);

OR2x2_ASAP7_75t_L g1674 ( 
.A(n_1617),
.B(n_1537),
.Y(n_1674)
);

INVx2_ASAP7_75t_L g1675 ( 
.A(n_1557),
.Y(n_1675)
);

AND2x2_ASAP7_75t_L g1676 ( 
.A(n_1571),
.B(n_1586),
.Y(n_1676)
);

BUFx2_ASAP7_75t_L g1677 ( 
.A(n_1610),
.Y(n_1677)
);

AO222x2_ASAP7_75t_L g1678 ( 
.A1(n_1569),
.A2(n_1645),
.B1(n_1631),
.B2(n_1545),
.C1(n_1539),
.C2(n_1543),
.Y(n_1678)
);

AND2x2_ASAP7_75t_L g1679 ( 
.A(n_1590),
.B(n_1615),
.Y(n_1679)
);

INVxp67_ASAP7_75t_L g1680 ( 
.A(n_1579),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1540),
.B(n_1558),
.Y(n_1681)
);

AO21x2_ASAP7_75t_L g1682 ( 
.A1(n_1624),
.A2(n_1627),
.B(n_1623),
.Y(n_1682)
);

BUFx2_ASAP7_75t_L g1683 ( 
.A(n_1626),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1542),
.B(n_1644),
.Y(n_1684)
);

OA21x2_ASAP7_75t_L g1685 ( 
.A1(n_1618),
.A2(n_1550),
.B(n_1561),
.Y(n_1685)
);

NOR2xp33_ASAP7_75t_L g1686 ( 
.A(n_1534),
.B(n_1629),
.Y(n_1686)
);

AO21x2_ASAP7_75t_L g1687 ( 
.A1(n_1601),
.A2(n_1638),
.B(n_1602),
.Y(n_1687)
);

OR2x6_ASAP7_75t_L g1688 ( 
.A(n_1567),
.B(n_1620),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1592),
.Y(n_1689)
);

AND2x2_ASAP7_75t_L g1690 ( 
.A(n_1582),
.B(n_1589),
.Y(n_1690)
);

INVxp67_ASAP7_75t_SL g1691 ( 
.A(n_1593),
.Y(n_1691)
);

AND2x4_ASAP7_75t_L g1692 ( 
.A(n_1562),
.B(n_1625),
.Y(n_1692)
);

AND2x2_ASAP7_75t_L g1693 ( 
.A(n_1585),
.B(n_1634),
.Y(n_1693)
);

AO21x2_ASAP7_75t_L g1694 ( 
.A1(n_1639),
.A2(n_1547),
.B(n_1548),
.Y(n_1694)
);

AO21x2_ASAP7_75t_L g1695 ( 
.A1(n_1577),
.A2(n_1605),
.B(n_1566),
.Y(n_1695)
);

INVx1_ASAP7_75t_L g1696 ( 
.A(n_1583),
.Y(n_1696)
);

AO21x2_ASAP7_75t_L g1697 ( 
.A1(n_1552),
.A2(n_1566),
.B(n_1580),
.Y(n_1697)
);

INVx1_ASAP7_75t_L g1698 ( 
.A(n_1552),
.Y(n_1698)
);

AOI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1628),
.A2(n_1578),
.B(n_1636),
.Y(n_1699)
);

OR2x2_ASAP7_75t_L g1700 ( 
.A(n_1630),
.B(n_1588),
.Y(n_1700)
);

AOI22xp33_ASAP7_75t_L g1701 ( 
.A1(n_1535),
.A2(n_1643),
.B1(n_1595),
.B2(n_1619),
.Y(n_1701)
);

OA21x2_ASAP7_75t_L g1702 ( 
.A1(n_1635),
.A2(n_1570),
.B(n_1595),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1596),
.Y(n_1703)
);

INVx1_ASAP7_75t_L g1704 ( 
.A(n_1594),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1663),
.B(n_1584),
.Y(n_1705)
);

AND2x2_ASAP7_75t_L g1706 ( 
.A(n_1663),
.B(n_1584),
.Y(n_1706)
);

AND2x2_ASAP7_75t_SL g1707 ( 
.A(n_1668),
.B(n_1576),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1647),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1691),
.B(n_1633),
.Y(n_1709)
);

NAND2x1_ASAP7_75t_L g1710 ( 
.A(n_1688),
.B(n_1637),
.Y(n_1710)
);

NAND2xp5_ASAP7_75t_L g1711 ( 
.A(n_1691),
.B(n_1568),
.Y(n_1711)
);

OR2x2_ASAP7_75t_L g1712 ( 
.A(n_1667),
.B(n_1658),
.Y(n_1712)
);

AOI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1694),
.A2(n_1608),
.B1(n_1607),
.B2(n_1554),
.Y(n_1713)
);

BUFx3_ASAP7_75t_L g1714 ( 
.A(n_1683),
.Y(n_1714)
);

NAND2xp5_ASAP7_75t_L g1715 ( 
.A(n_1656),
.B(n_1563),
.Y(n_1715)
);

INVx1_ASAP7_75t_L g1716 ( 
.A(n_1647),
.Y(n_1716)
);

HB1xp67_ASAP7_75t_L g1717 ( 
.A(n_1665),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1649),
.Y(n_1718)
);

AND2x4_ASAP7_75t_L g1719 ( 
.A(n_1677),
.B(n_1598),
.Y(n_1719)
);

AOI22xp33_ASAP7_75t_L g1720 ( 
.A1(n_1694),
.A2(n_1535),
.B1(n_1613),
.B2(n_1560),
.Y(n_1720)
);

AND2x4_ASAP7_75t_L g1721 ( 
.A(n_1652),
.B(n_1570),
.Y(n_1721)
);

AND2x2_ASAP7_75t_L g1722 ( 
.A(n_1679),
.B(n_1544),
.Y(n_1722)
);

OR2x6_ASAP7_75t_L g1723 ( 
.A(n_1652),
.B(n_1538),
.Y(n_1723)
);

AND2x2_ASAP7_75t_L g1724 ( 
.A(n_1679),
.B(n_1656),
.Y(n_1724)
);

AND2x2_ASAP7_75t_L g1725 ( 
.A(n_1697),
.B(n_1698),
.Y(n_1725)
);

HB1xp67_ASAP7_75t_L g1726 ( 
.A(n_1671),
.Y(n_1726)
);

HB1xp67_ASAP7_75t_L g1727 ( 
.A(n_1671),
.Y(n_1727)
);

AND2x2_ASAP7_75t_L g1728 ( 
.A(n_1697),
.B(n_1544),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1689),
.B(n_1538),
.Y(n_1729)
);

AND2x2_ASAP7_75t_L g1730 ( 
.A(n_1697),
.B(n_1576),
.Y(n_1730)
);

AND2x4_ASAP7_75t_L g1731 ( 
.A(n_1662),
.B(n_1675),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1689),
.B(n_1666),
.Y(n_1732)
);

NOR2xp33_ASAP7_75t_L g1733 ( 
.A(n_1699),
.B(n_1621),
.Y(n_1733)
);

AND2x2_ASAP7_75t_L g1734 ( 
.A(n_1697),
.B(n_1695),
.Y(n_1734)
);

OR2x2_ASAP7_75t_L g1735 ( 
.A(n_1712),
.B(n_1726),
.Y(n_1735)
);

OR2x2_ASAP7_75t_L g1736 ( 
.A(n_1712),
.B(n_1654),
.Y(n_1736)
);

INVx3_ASAP7_75t_L g1737 ( 
.A(n_1731),
.Y(n_1737)
);

AND2x4_ASAP7_75t_L g1738 ( 
.A(n_1714),
.B(n_1692),
.Y(n_1738)
);

AOI22xp33_ASAP7_75t_L g1739 ( 
.A1(n_1707),
.A2(n_1694),
.B1(n_1648),
.B2(n_1733),
.Y(n_1739)
);

OAI22xp33_ASAP7_75t_L g1740 ( 
.A1(n_1713),
.A2(n_1648),
.B1(n_1666),
.B2(n_1699),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1705),
.B(n_1650),
.Y(n_1741)
);

OR2x6_ASAP7_75t_L g1742 ( 
.A(n_1723),
.B(n_1688),
.Y(n_1742)
);

NAND4xp25_ASAP7_75t_L g1743 ( 
.A(n_1733),
.B(n_1686),
.C(n_1701),
.D(n_1654),
.Y(n_1743)
);

OAI22xp5_ASAP7_75t_L g1744 ( 
.A1(n_1707),
.A2(n_1688),
.B1(n_1670),
.B2(n_1700),
.Y(n_1744)
);

OAI211xp5_ASAP7_75t_L g1745 ( 
.A1(n_1720),
.A2(n_1678),
.B(n_1685),
.C(n_1702),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1712),
.B(n_1684),
.Y(n_1746)
);

CKINVDCx20_ASAP7_75t_R g1747 ( 
.A(n_1715),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1708),
.Y(n_1748)
);

INVx1_ASAP7_75t_L g1749 ( 
.A(n_1708),
.Y(n_1749)
);

INVx5_ASAP7_75t_L g1750 ( 
.A(n_1723),
.Y(n_1750)
);

AOI221xp5_ASAP7_75t_L g1751 ( 
.A1(n_1730),
.A2(n_1694),
.B1(n_1682),
.B2(n_1680),
.C(n_1684),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1709),
.B(n_1700),
.Y(n_1752)
);

INVx3_ASAP7_75t_L g1753 ( 
.A(n_1731),
.Y(n_1753)
);

NAND2xp33_ASAP7_75t_R g1754 ( 
.A(n_1730),
.B(n_1688),
.Y(n_1754)
);

BUFx2_ASAP7_75t_L g1755 ( 
.A(n_1714),
.Y(n_1755)
);

INVxp67_ASAP7_75t_L g1756 ( 
.A(n_1722),
.Y(n_1756)
);

AOI221xp5_ASAP7_75t_L g1757 ( 
.A1(n_1730),
.A2(n_1682),
.B1(n_1680),
.B2(n_1696),
.C(n_1704),
.Y(n_1757)
);

AOI22xp33_ASAP7_75t_SL g1758 ( 
.A1(n_1707),
.A2(n_1682),
.B1(n_1688),
.B2(n_1702),
.Y(n_1758)
);

AOI33xp33_ASAP7_75t_L g1759 ( 
.A1(n_1720),
.A2(n_1696),
.A3(n_1704),
.B1(n_1676),
.B2(n_1693),
.B3(n_1690),
.Y(n_1759)
);

NAND2xp33_ASAP7_75t_R g1760 ( 
.A(n_1732),
.B(n_1575),
.Y(n_1760)
);

INVx1_ASAP7_75t_L g1761 ( 
.A(n_1716),
.Y(n_1761)
);

BUFx2_ASAP7_75t_L g1762 ( 
.A(n_1714),
.Y(n_1762)
);

INVxp67_ASAP7_75t_L g1763 ( 
.A(n_1722),
.Y(n_1763)
);

AND2x2_ASAP7_75t_L g1764 ( 
.A(n_1706),
.B(n_1693),
.Y(n_1764)
);

AOI33xp33_ASAP7_75t_L g1765 ( 
.A1(n_1722),
.A2(n_1676),
.A3(n_1690),
.B1(n_1653),
.B2(n_1651),
.B3(n_1669),
.Y(n_1765)
);

AOI22xp5_ASAP7_75t_L g1766 ( 
.A1(n_1707),
.A2(n_1682),
.B1(n_1687),
.B2(n_1692),
.Y(n_1766)
);

BUFx10_ASAP7_75t_L g1767 ( 
.A(n_1719),
.Y(n_1767)
);

OAI22xp5_ASAP7_75t_SL g1768 ( 
.A1(n_1713),
.A2(n_1664),
.B1(n_1661),
.B2(n_1673),
.Y(n_1768)
);

AND2x2_ASAP7_75t_L g1769 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1769)
);

OAI33xp33_ASAP7_75t_L g1770 ( 
.A1(n_1729),
.A2(n_1674),
.A3(n_1681),
.B1(n_1659),
.B2(n_1660),
.B3(n_1657),
.Y(n_1770)
);

NOR4xp25_ASAP7_75t_L g1771 ( 
.A(n_1729),
.B(n_1681),
.C(n_1674),
.D(n_1703),
.Y(n_1771)
);

AND2x6_ASAP7_75t_SL g1772 ( 
.A(n_1719),
.B(n_1664),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1716),
.Y(n_1773)
);

NAND3xp33_ASAP7_75t_L g1774 ( 
.A(n_1711),
.B(n_1702),
.C(n_1652),
.Y(n_1774)
);

AND2x2_ASAP7_75t_L g1775 ( 
.A(n_1706),
.B(n_1692),
.Y(n_1775)
);

INVx1_ASAP7_75t_L g1776 ( 
.A(n_1718),
.Y(n_1776)
);

HB1xp67_ASAP7_75t_L g1777 ( 
.A(n_1717),
.Y(n_1777)
);

OAI31xp33_ASAP7_75t_L g1778 ( 
.A1(n_1721),
.A2(n_1655),
.A3(n_1703),
.B(n_1672),
.Y(n_1778)
);

AND2x2_ASAP7_75t_L g1779 ( 
.A(n_1756),
.B(n_1763),
.Y(n_1779)
);

OA21x2_ASAP7_75t_L g1780 ( 
.A1(n_1751),
.A2(n_1734),
.B(n_1725),
.Y(n_1780)
);

HB1xp67_ASAP7_75t_L g1781 ( 
.A(n_1777),
.Y(n_1781)
);

INVx2_ASAP7_75t_L g1782 ( 
.A(n_1737),
.Y(n_1782)
);

INVx4_ASAP7_75t_SL g1783 ( 
.A(n_1768),
.Y(n_1783)
);

INVx2_ASAP7_75t_SL g1784 ( 
.A(n_1767),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1767),
.Y(n_1785)
);

OR2x2_ASAP7_75t_L g1786 ( 
.A(n_1771),
.B(n_1763),
.Y(n_1786)
);

OR2x6_ASAP7_75t_L g1787 ( 
.A(n_1742),
.B(n_1710),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1748),
.Y(n_1788)
);

INVx1_ASAP7_75t_SL g1789 ( 
.A(n_1755),
.Y(n_1789)
);

BUFx12f_ASAP7_75t_L g1790 ( 
.A(n_1772),
.Y(n_1790)
);

NAND3xp33_ASAP7_75t_SL g1791 ( 
.A(n_1739),
.B(n_1751),
.C(n_1745),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1749),
.Y(n_1792)
);

INVx2_ASAP7_75t_L g1793 ( 
.A(n_1753),
.Y(n_1793)
);

INVx1_ASAP7_75t_L g1794 ( 
.A(n_1761),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1773),
.B(n_1726),
.Y(n_1795)
);

INVx2_ASAP7_75t_L g1796 ( 
.A(n_1776),
.Y(n_1796)
);

HB1xp67_ASAP7_75t_L g1797 ( 
.A(n_1777),
.Y(n_1797)
);

NOR2x1p5_ASAP7_75t_L g1798 ( 
.A(n_1743),
.B(n_1710),
.Y(n_1798)
);

INVx1_ASAP7_75t_L g1799 ( 
.A(n_1735),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1736),
.Y(n_1800)
);

AO21x1_ASAP7_75t_L g1801 ( 
.A1(n_1740),
.A2(n_1734),
.B(n_1728),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1746),
.Y(n_1802)
);

AND2x2_ASAP7_75t_L g1803 ( 
.A(n_1762),
.B(n_1724),
.Y(n_1803)
);

HB1xp67_ASAP7_75t_L g1804 ( 
.A(n_1752),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1738),
.Y(n_1805)
);

AOI21xp33_ASAP7_75t_L g1806 ( 
.A1(n_1740),
.A2(n_1711),
.B(n_1723),
.Y(n_1806)
);

OA21x2_ASAP7_75t_L g1807 ( 
.A1(n_1774),
.A2(n_1734),
.B(n_1725),
.Y(n_1807)
);

AOI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1745),
.A2(n_1723),
.B(n_1685),
.Y(n_1808)
);

AND2x2_ASAP7_75t_L g1809 ( 
.A(n_1758),
.B(n_1724),
.Y(n_1809)
);

INVx5_ASAP7_75t_L g1810 ( 
.A(n_1742),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1765),
.Y(n_1811)
);

INVx1_ASAP7_75t_L g1812 ( 
.A(n_1738),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1788),
.Y(n_1813)
);

AND2x2_ASAP7_75t_L g1814 ( 
.A(n_1809),
.B(n_1769),
.Y(n_1814)
);

INVx1_ASAP7_75t_SL g1815 ( 
.A(n_1789),
.Y(n_1815)
);

AND2x2_ASAP7_75t_L g1816 ( 
.A(n_1809),
.B(n_1775),
.Y(n_1816)
);

BUFx2_ASAP7_75t_L g1817 ( 
.A(n_1790),
.Y(n_1817)
);

OR2x2_ASAP7_75t_L g1818 ( 
.A(n_1786),
.B(n_1727),
.Y(n_1818)
);

INVx1_ASAP7_75t_L g1819 ( 
.A(n_1788),
.Y(n_1819)
);

NOR2x1_ASAP7_75t_L g1820 ( 
.A(n_1791),
.B(n_1670),
.Y(n_1820)
);

INVx5_ASAP7_75t_SL g1821 ( 
.A(n_1787),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_L g1822 ( 
.A(n_1811),
.B(n_1739),
.Y(n_1822)
);

NAND3xp33_ASAP7_75t_L g1823 ( 
.A(n_1786),
.B(n_1806),
.C(n_1808),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1792),
.Y(n_1824)
);

INVx2_ASAP7_75t_L g1825 ( 
.A(n_1796),
.Y(n_1825)
);

NAND2xp5_ASAP7_75t_L g1826 ( 
.A(n_1811),
.B(n_1764),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1804),
.B(n_1759),
.Y(n_1827)
);

AND3x1_ASAP7_75t_L g1828 ( 
.A(n_1783),
.B(n_1766),
.C(n_1757),
.Y(n_1828)
);

A2O1A1Ixp33_ASAP7_75t_L g1829 ( 
.A1(n_1791),
.A2(n_1757),
.B(n_1758),
.C(n_1778),
.Y(n_1829)
);

BUFx3_ASAP7_75t_L g1830 ( 
.A(n_1790),
.Y(n_1830)
);

INVx1_ASAP7_75t_L g1831 ( 
.A(n_1792),
.Y(n_1831)
);

OR2x2_ASAP7_75t_L g1832 ( 
.A(n_1786),
.B(n_1727),
.Y(n_1832)
);

CKINVDCx5p33_ASAP7_75t_R g1833 ( 
.A(n_1790),
.Y(n_1833)
);

INVx1_ASAP7_75t_L g1834 ( 
.A(n_1794),
.Y(n_1834)
);

BUFx3_ASAP7_75t_L g1835 ( 
.A(n_1810),
.Y(n_1835)
);

NAND2xp33_ASAP7_75t_SL g1836 ( 
.A(n_1798),
.B(n_1760),
.Y(n_1836)
);

INVx1_ASAP7_75t_SL g1837 ( 
.A(n_1783),
.Y(n_1837)
);

OR2x6_ASAP7_75t_L g1838 ( 
.A(n_1801),
.B(n_1723),
.Y(n_1838)
);

NAND3xp33_ASAP7_75t_SL g1839 ( 
.A(n_1801),
.B(n_1808),
.C(n_1789),
.Y(n_1839)
);

INVx1_ASAP7_75t_L g1840 ( 
.A(n_1794),
.Y(n_1840)
);

INVx2_ASAP7_75t_L g1841 ( 
.A(n_1796),
.Y(n_1841)
);

NAND3xp33_ASAP7_75t_SL g1842 ( 
.A(n_1801),
.B(n_1744),
.C(n_1747),
.Y(n_1842)
);

AND2x2_ASAP7_75t_L g1843 ( 
.A(n_1805),
.B(n_1750),
.Y(n_1843)
);

AND2x2_ASAP7_75t_L g1844 ( 
.A(n_1805),
.B(n_1750),
.Y(n_1844)
);

AND2x2_ASAP7_75t_L g1845 ( 
.A(n_1812),
.B(n_1741),
.Y(n_1845)
);

INVxp67_ASAP7_75t_SL g1846 ( 
.A(n_1798),
.Y(n_1846)
);

INVx1_ASAP7_75t_SL g1847 ( 
.A(n_1817),
.Y(n_1847)
);

INVx1_ASAP7_75t_SL g1848 ( 
.A(n_1817),
.Y(n_1848)
);

NAND2xp5_ASAP7_75t_L g1849 ( 
.A(n_1822),
.B(n_1800),
.Y(n_1849)
);

OR2x6_ASAP7_75t_L g1850 ( 
.A(n_1820),
.B(n_1830),
.Y(n_1850)
);

OA21x2_ASAP7_75t_L g1851 ( 
.A1(n_1823),
.A2(n_1782),
.B(n_1793),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1815),
.B(n_1800),
.Y(n_1852)
);

NAND2xp5_ASAP7_75t_L g1853 ( 
.A(n_1815),
.B(n_1802),
.Y(n_1853)
);

NOR2xp67_ASAP7_75t_L g1854 ( 
.A(n_1839),
.B(n_1823),
.Y(n_1854)
);

AND2x2_ASAP7_75t_L g1855 ( 
.A(n_1814),
.B(n_1783),
.Y(n_1855)
);

NAND2xp5_ASAP7_75t_L g1856 ( 
.A(n_1826),
.B(n_1802),
.Y(n_1856)
);

AND2x2_ASAP7_75t_L g1857 ( 
.A(n_1814),
.B(n_1783),
.Y(n_1857)
);

INVx1_ASAP7_75t_L g1858 ( 
.A(n_1813),
.Y(n_1858)
);

INVx2_ASAP7_75t_L g1859 ( 
.A(n_1825),
.Y(n_1859)
);

OR2x2_ASAP7_75t_L g1860 ( 
.A(n_1827),
.B(n_1799),
.Y(n_1860)
);

OAI22xp33_ASAP7_75t_L g1861 ( 
.A1(n_1842),
.A2(n_1754),
.B1(n_1780),
.B2(n_1810),
.Y(n_1861)
);

AND2x4_ASAP7_75t_L g1862 ( 
.A(n_1835),
.B(n_1783),
.Y(n_1862)
);

INVxp67_ASAP7_75t_L g1863 ( 
.A(n_1820),
.Y(n_1863)
);

INVxp67_ASAP7_75t_L g1864 ( 
.A(n_1830),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1813),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1819),
.Y(n_1866)
);

NAND2xp5_ASAP7_75t_L g1867 ( 
.A(n_1845),
.B(n_1799),
.Y(n_1867)
);

AND2x2_ASAP7_75t_L g1868 ( 
.A(n_1816),
.B(n_1783),
.Y(n_1868)
);

INVx3_ASAP7_75t_L g1869 ( 
.A(n_1835),
.Y(n_1869)
);

OR2x2_ASAP7_75t_L g1870 ( 
.A(n_1818),
.B(n_1780),
.Y(n_1870)
);

OAI21xp33_ASAP7_75t_L g1871 ( 
.A1(n_1829),
.A2(n_1806),
.B(n_1779),
.Y(n_1871)
);

INVx1_ASAP7_75t_L g1872 ( 
.A(n_1819),
.Y(n_1872)
);

A2O1A1Ixp33_ASAP7_75t_L g1873 ( 
.A1(n_1830),
.A2(n_1810),
.B(n_1721),
.C(n_1797),
.Y(n_1873)
);

INVxp67_ASAP7_75t_SL g1874 ( 
.A(n_1818),
.Y(n_1874)
);

AND2x2_ASAP7_75t_L g1875 ( 
.A(n_1816),
.B(n_1779),
.Y(n_1875)
);

INVx1_ASAP7_75t_L g1876 ( 
.A(n_1824),
.Y(n_1876)
);

NAND2xp5_ASAP7_75t_L g1877 ( 
.A(n_1845),
.B(n_1803),
.Y(n_1877)
);

INVx2_ASAP7_75t_L g1878 ( 
.A(n_1825),
.Y(n_1878)
);

OAI211xp5_ASAP7_75t_L g1879 ( 
.A1(n_1837),
.A2(n_1780),
.B(n_1807),
.C(n_1810),
.Y(n_1879)
);

OR2x6_ASAP7_75t_L g1880 ( 
.A(n_1835),
.B(n_1673),
.Y(n_1880)
);

AND2x2_ASAP7_75t_L g1881 ( 
.A(n_1821),
.B(n_1779),
.Y(n_1881)
);

INVx1_ASAP7_75t_L g1882 ( 
.A(n_1824),
.Y(n_1882)
);

NOR4xp25_ASAP7_75t_L g1883 ( 
.A(n_1832),
.B(n_1795),
.C(n_1784),
.D(n_1785),
.Y(n_1883)
);

AND2x4_ASAP7_75t_L g1884 ( 
.A(n_1854),
.B(n_1828),
.Y(n_1884)
);

AND2x2_ASAP7_75t_L g1885 ( 
.A(n_1850),
.B(n_1821),
.Y(n_1885)
);

AOI22xp33_ASAP7_75t_L g1886 ( 
.A1(n_1871),
.A2(n_1836),
.B1(n_1780),
.B2(n_1838),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1850),
.B(n_1855),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1850),
.B(n_1821),
.Y(n_1888)
);

NAND2xp5_ASAP7_75t_SL g1889 ( 
.A(n_1861),
.B(n_1828),
.Y(n_1889)
);

AND2x2_ASAP7_75t_L g1890 ( 
.A(n_1850),
.B(n_1821),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1874),
.Y(n_1891)
);

BUFx3_ASAP7_75t_L g1892 ( 
.A(n_1869),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1851),
.Y(n_1893)
);

INVx3_ASAP7_75t_SL g1894 ( 
.A(n_1847),
.Y(n_1894)
);

OAI21x1_ASAP7_75t_L g1895 ( 
.A1(n_1851),
.A2(n_1832),
.B(n_1825),
.Y(n_1895)
);

AND2x2_ASAP7_75t_L g1896 ( 
.A(n_1855),
.B(n_1857),
.Y(n_1896)
);

NOR2xp33_ASAP7_75t_R g1897 ( 
.A(n_1848),
.B(n_1833),
.Y(n_1897)
);

AOI22xp33_ASAP7_75t_L g1898 ( 
.A1(n_1863),
.A2(n_1780),
.B1(n_1838),
.B2(n_1846),
.Y(n_1898)
);

INVx2_ASAP7_75t_L g1899 ( 
.A(n_1851),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1849),
.B(n_1831),
.Y(n_1900)
);

AOI222xp33_ASAP7_75t_L g1901 ( 
.A1(n_1864),
.A2(n_1770),
.B1(n_1797),
.B2(n_1781),
.C1(n_1831),
.C2(n_1834),
.Y(n_1901)
);

INVx1_ASAP7_75t_L g1902 ( 
.A(n_1858),
.Y(n_1902)
);

INVx1_ASAP7_75t_L g1903 ( 
.A(n_1865),
.Y(n_1903)
);

AND2x2_ASAP7_75t_L g1904 ( 
.A(n_1857),
.B(n_1821),
.Y(n_1904)
);

INVx2_ASAP7_75t_L g1905 ( 
.A(n_1875),
.Y(n_1905)
);

INVx1_ASAP7_75t_L g1906 ( 
.A(n_1866),
.Y(n_1906)
);

INVx1_ASAP7_75t_SL g1907 ( 
.A(n_1862),
.Y(n_1907)
);

INVxp67_ASAP7_75t_L g1908 ( 
.A(n_1852),
.Y(n_1908)
);

OR2x2_ASAP7_75t_L g1909 ( 
.A(n_1870),
.B(n_1841),
.Y(n_1909)
);

OAI211xp5_ASAP7_75t_L g1910 ( 
.A1(n_1889),
.A2(n_1883),
.B(n_1879),
.C(n_1873),
.Y(n_1910)
);

BUFx2_ASAP7_75t_L g1911 ( 
.A(n_1897),
.Y(n_1911)
);

BUFx12f_ASAP7_75t_L g1912 ( 
.A(n_1884),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1892),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1894),
.B(n_1880),
.Y(n_1914)
);

AOI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1884),
.A2(n_1868),
.B1(n_1862),
.B2(n_1838),
.Y(n_1915)
);

INVx2_ASAP7_75t_SL g1916 ( 
.A(n_1892),
.Y(n_1916)
);

OAI21xp5_ASAP7_75t_SL g1917 ( 
.A1(n_1884),
.A2(n_1868),
.B(n_1862),
.Y(n_1917)
);

OAI22xp33_ASAP7_75t_SL g1918 ( 
.A1(n_1884),
.A2(n_1838),
.B1(n_1894),
.B2(n_1870),
.Y(n_1918)
);

OR2x2_ASAP7_75t_L g1919 ( 
.A(n_1894),
.B(n_1853),
.Y(n_1919)
);

OAI221xp5_ASAP7_75t_SL g1920 ( 
.A1(n_1886),
.A2(n_1838),
.B1(n_1860),
.B2(n_1873),
.C(n_1880),
.Y(n_1920)
);

INVx1_ASAP7_75t_L g1921 ( 
.A(n_1905),
.Y(n_1921)
);

INVx1_ASAP7_75t_SL g1922 ( 
.A(n_1897),
.Y(n_1922)
);

AOI33xp33_ASAP7_75t_L g1923 ( 
.A1(n_1884),
.A2(n_1881),
.A3(n_1875),
.B1(n_1872),
.B2(n_1882),
.B3(n_1876),
.Y(n_1923)
);

AOI221xp5_ASAP7_75t_L g1924 ( 
.A1(n_1886),
.A2(n_1881),
.B1(n_1856),
.B2(n_1869),
.C(n_1867),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1894),
.B(n_1896),
.Y(n_1925)
);

AOI22xp33_ASAP7_75t_L g1926 ( 
.A1(n_1898),
.A2(n_1780),
.B1(n_1880),
.B2(n_1810),
.Y(n_1926)
);

INVxp67_ASAP7_75t_SL g1927 ( 
.A(n_1893),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1905),
.Y(n_1928)
);

AOI21xp33_ASAP7_75t_L g1929 ( 
.A1(n_1885),
.A2(n_1880),
.B(n_1869),
.Y(n_1929)
);

NAND2x1_ASAP7_75t_SL g1930 ( 
.A(n_1915),
.B(n_1885),
.Y(n_1930)
);

INVx1_ASAP7_75t_L g1931 ( 
.A(n_1927),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1910),
.A2(n_1899),
.B(n_1893),
.Y(n_1932)
);

NOR2xp67_ASAP7_75t_SL g1933 ( 
.A(n_1912),
.B(n_1642),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_SL g1934 ( 
.A(n_1918),
.B(n_1885),
.Y(n_1934)
);

INVx1_ASAP7_75t_L g1935 ( 
.A(n_1927),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_L g1936 ( 
.A(n_1916),
.B(n_1896),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1921),
.Y(n_1937)
);

NAND2xp5_ASAP7_75t_L g1938 ( 
.A(n_1925),
.B(n_1896),
.Y(n_1938)
);

OAI22xp33_ASAP7_75t_L g1939 ( 
.A1(n_1919),
.A2(n_1899),
.B1(n_1893),
.B2(n_1810),
.Y(n_1939)
);

INVx1_ASAP7_75t_L g1940 ( 
.A(n_1928),
.Y(n_1940)
);

OAI22xp5_ASAP7_75t_SL g1941 ( 
.A1(n_1911),
.A2(n_1587),
.B1(n_1898),
.B2(n_1907),
.Y(n_1941)
);

INVx1_ASAP7_75t_SL g1942 ( 
.A(n_1930),
.Y(n_1942)
);

NAND3xp33_ASAP7_75t_L g1943 ( 
.A(n_1932),
.B(n_1910),
.C(n_1920),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_L g1944 ( 
.A(n_1936),
.B(n_1907),
.Y(n_1944)
);

OAI211xp5_ASAP7_75t_SL g1945 ( 
.A1(n_1934),
.A2(n_1923),
.B(n_1922),
.C(n_1924),
.Y(n_1945)
);

OAI221xp5_ASAP7_75t_L g1946 ( 
.A1(n_1941),
.A2(n_1920),
.B1(n_1926),
.B2(n_1917),
.C(n_1914),
.Y(n_1946)
);

NOR3xp33_ASAP7_75t_L g1947 ( 
.A(n_1938),
.B(n_1929),
.C(n_1913),
.Y(n_1947)
);

INVxp67_ASAP7_75t_SL g1948 ( 
.A(n_1933),
.Y(n_1948)
);

AOI211xp5_ASAP7_75t_L g1949 ( 
.A1(n_1932),
.A2(n_1887),
.B(n_1888),
.C(n_1890),
.Y(n_1949)
);

OR2x2_ASAP7_75t_L g1950 ( 
.A(n_1931),
.B(n_1891),
.Y(n_1950)
);

AOI221xp5_ASAP7_75t_L g1951 ( 
.A1(n_1935),
.A2(n_1908),
.B1(n_1891),
.B2(n_1887),
.C(n_1900),
.Y(n_1951)
);

O2A1O1Ixp5_ASAP7_75t_L g1952 ( 
.A1(n_1939),
.A2(n_1899),
.B(n_1888),
.C(n_1890),
.Y(n_1952)
);

AOI21xp33_ASAP7_75t_L g1953 ( 
.A1(n_1937),
.A2(n_1890),
.B(n_1888),
.Y(n_1953)
);

AOI22xp5_ASAP7_75t_L g1954 ( 
.A1(n_1943),
.A2(n_1904),
.B1(n_1887),
.B2(n_1905),
.Y(n_1954)
);

OAI22xp5_ASAP7_75t_L g1955 ( 
.A1(n_1942),
.A2(n_1908),
.B1(n_1904),
.B2(n_1892),
.Y(n_1955)
);

XNOR2x1_ASAP7_75t_L g1956 ( 
.A(n_1944),
.B(n_1642),
.Y(n_1956)
);

AOI22xp33_ASAP7_75t_L g1957 ( 
.A1(n_1945),
.A2(n_1904),
.B1(n_1901),
.B2(n_1940),
.Y(n_1957)
);

INVx1_ASAP7_75t_L g1958 ( 
.A(n_1950),
.Y(n_1958)
);

OAI22xp5_ASAP7_75t_L g1959 ( 
.A1(n_1948),
.A2(n_1900),
.B1(n_1877),
.B2(n_1810),
.Y(n_1959)
);

A2O1A1Ixp33_ASAP7_75t_L g1960 ( 
.A1(n_1952),
.A2(n_1895),
.B(n_1902),
.C(n_1906),
.Y(n_1960)
);

NOR2x1_ASAP7_75t_L g1961 ( 
.A(n_1958),
.B(n_1946),
.Y(n_1961)
);

NAND2xp5_ASAP7_75t_SL g1962 ( 
.A(n_1955),
.B(n_1949),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1954),
.Y(n_1963)
);

INVx2_ASAP7_75t_L g1964 ( 
.A(n_1956),
.Y(n_1964)
);

INVxp67_ASAP7_75t_L g1965 ( 
.A(n_1959),
.Y(n_1965)
);

OR2x2_ASAP7_75t_L g1966 ( 
.A(n_1957),
.B(n_1947),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1960),
.B(n_1951),
.Y(n_1967)
);

AOI22xp33_ASAP7_75t_L g1968 ( 
.A1(n_1961),
.A2(n_1966),
.B1(n_1967),
.B2(n_1963),
.Y(n_1968)
);

INVx2_ASAP7_75t_SL g1969 ( 
.A(n_1964),
.Y(n_1969)
);

NAND2x1p5_ASAP7_75t_L g1970 ( 
.A(n_1962),
.B(n_1902),
.Y(n_1970)
);

OAI22xp33_ASAP7_75t_L g1971 ( 
.A1(n_1965),
.A2(n_1953),
.B1(n_1903),
.B2(n_1906),
.Y(n_1971)
);

BUFx8_ASAP7_75t_SL g1972 ( 
.A(n_1964),
.Y(n_1972)
);

INVx1_ASAP7_75t_SL g1973 ( 
.A(n_1961),
.Y(n_1973)
);

INVx2_ASAP7_75t_L g1974 ( 
.A(n_1970),
.Y(n_1974)
);

OAI21xp33_ASAP7_75t_L g1975 ( 
.A1(n_1968),
.A2(n_1903),
.B(n_1901),
.Y(n_1975)
);

INVx1_ASAP7_75t_L g1976 ( 
.A(n_1973),
.Y(n_1976)
);

NOR3xp33_ASAP7_75t_L g1977 ( 
.A(n_1976),
.B(n_1969),
.C(n_1971),
.Y(n_1977)
);

NAND3xp33_ASAP7_75t_SL g1978 ( 
.A(n_1977),
.B(n_1974),
.C(n_1975),
.Y(n_1978)
);

INVx3_ASAP7_75t_L g1979 ( 
.A(n_1978),
.Y(n_1979)
);

OR3x2_ASAP7_75t_L g1980 ( 
.A(n_1978),
.B(n_1972),
.C(n_1909),
.Y(n_1980)
);

NAND2x1p5_ASAP7_75t_L g1981 ( 
.A(n_1979),
.B(n_1640),
.Y(n_1981)
);

INVx1_ASAP7_75t_L g1982 ( 
.A(n_1980),
.Y(n_1982)
);

NAND2xp5_ASAP7_75t_L g1983 ( 
.A(n_1982),
.B(n_1587),
.Y(n_1983)
);

OAI22xp5_ASAP7_75t_SL g1984 ( 
.A1(n_1981),
.A2(n_1673),
.B1(n_1640),
.B2(n_1909),
.Y(n_1984)
);

AOI22xp5_ASAP7_75t_L g1985 ( 
.A1(n_1984),
.A2(n_1895),
.B1(n_1878),
.B2(n_1859),
.Y(n_1985)
);

NOR2xp33_ASAP7_75t_SL g1986 ( 
.A(n_1985),
.B(n_1983),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1986),
.A2(n_1909),
.B(n_1859),
.Y(n_1987)
);

AOI22x1_ASAP7_75t_L g1988 ( 
.A1(n_1987),
.A2(n_1878),
.B1(n_1895),
.B2(n_1841),
.Y(n_1988)
);

OAI22xp33_ASAP7_75t_L g1989 ( 
.A1(n_1988),
.A2(n_1841),
.B1(n_1834),
.B2(n_1840),
.Y(n_1989)
);

AOI211xp5_ASAP7_75t_L g1990 ( 
.A1(n_1989),
.A2(n_1840),
.B(n_1843),
.C(n_1844),
.Y(n_1990)
);


endmodule