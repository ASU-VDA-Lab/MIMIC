module fake_jpeg_20522_n_278 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_278);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_278;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_212;
wire n_131;
wire n_56;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx3_ASAP7_75t_L g16 ( 
.A(n_15),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_2),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_13),
.Y(n_23)
);

BUFx10_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx8_ASAP7_75t_L g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx4f_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx3_ASAP7_75t_L g30 ( 
.A(n_9),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_6),
.Y(n_31)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_28),
.Y(n_33)
);

INVx11_ASAP7_75t_L g51 ( 
.A(n_33),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_18),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_34),
.B(n_35),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_19),
.Y(n_36)
);

INVx5_ASAP7_75t_SL g54 ( 
.A(n_36),
.Y(n_54)
);

INVx4_ASAP7_75t_SL g37 ( 
.A(n_30),
.Y(n_37)
);

INVx6_ASAP7_75t_SL g53 ( 
.A(n_37),
.Y(n_53)
);

NAND2xp33_ASAP7_75t_SL g38 ( 
.A(n_29),
.B(n_0),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_20),
.Y(n_39)
);

INVx2_ASAP7_75t_SL g40 ( 
.A(n_19),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_40),
.Y(n_43)
);

INVx6_ASAP7_75t_L g41 ( 
.A(n_33),
.Y(n_41)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_41),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_42),
.B(n_48),
.Y(n_69)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_33),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_45),
.B(n_24),
.Y(n_71)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_30),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g66 ( 
.A1(n_46),
.A2(n_40),
.B1(n_36),
.B2(n_37),
.Y(n_66)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_37),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_24),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_33),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_49),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_52),
.B(n_39),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_36),
.A2(n_30),
.B1(n_32),
.B2(n_31),
.Y(n_55)
);

OA22x2_ASAP7_75t_L g83 ( 
.A1(n_55),
.A2(n_28),
.B1(n_26),
.B2(n_20),
.Y(n_83)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_33),
.Y(n_57)
);

BUFx6f_ASAP7_75t_SL g59 ( 
.A(n_57),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g58 ( 
.A1(n_36),
.A2(n_32),
.B1(n_31),
.B2(n_19),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_L g67 ( 
.A1(n_58),
.A2(n_40),
.B1(n_54),
.B2(n_37),
.Y(n_67)
);

INVxp67_ASAP7_75t_L g97 ( 
.A(n_60),
.Y(n_97)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_42),
.Y(n_61)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_61),
.Y(n_113)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_51),
.Y(n_63)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_63),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_50),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_65),
.B(n_72),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_66),
.A2(n_77),
.B1(n_79),
.B2(n_87),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_67),
.A2(n_73),
.B1(n_57),
.B2(n_44),
.Y(n_107)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_52),
.Y(n_70)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_70),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g110 ( 
.A(n_71),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_50),
.B(n_35),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_L g73 ( 
.A1(n_56),
.A2(n_40),
.B1(n_37),
.B2(n_39),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_55),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_74),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_75),
.B(n_76),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_27),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_51),
.A2(n_40),
.B1(n_21),
.B2(n_25),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g78 ( 
.A(n_55),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_78),
.B(n_82),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_51),
.A2(n_40),
.B1(n_21),
.B2(n_25),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_81),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_53),
.B(n_27),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g90 ( 
.A1(n_83),
.A2(n_54),
.B1(n_53),
.B2(n_57),
.Y(n_90)
);

OR2x2_ASAP7_75t_L g84 ( 
.A(n_43),
.B(n_28),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_85),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_53),
.B(n_26),
.Y(n_85)
);

AND2x2_ASAP7_75t_SL g86 ( 
.A(n_43),
.B(n_29),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_86),
.B(n_47),
.C(n_24),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_54),
.A2(n_28),
.B1(n_29),
.B2(n_16),
.Y(n_87)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_80),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_89),
.B(n_100),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_90),
.A2(n_86),
.B1(n_60),
.B2(n_41),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_80),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

CKINVDCx12_ASAP7_75t_R g92 ( 
.A(n_65),
.Y(n_92)
);

CKINVDCx14_ASAP7_75t_R g121 ( 
.A(n_92),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_69),
.B(n_70),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_108),
.Y(n_122)
);

AND2x6_ASAP7_75t_L g96 ( 
.A(n_61),
.B(n_58),
.Y(n_96)
);

NAND3xp33_ASAP7_75t_L g138 ( 
.A(n_96),
.B(n_109),
.C(n_68),
.Y(n_138)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_68),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_69),
.B(n_45),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_101),
.B(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_49),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g126 ( 
.A1(n_107),
.A2(n_103),
.B1(n_84),
.B2(n_113),
.Y(n_126)
);

NOR2x1_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_28),
.Y(n_109)
);

INVx13_ASAP7_75t_L g111 ( 
.A(n_63),
.Y(n_111)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_86),
.B(n_47),
.C(n_29),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_112),
.B(n_41),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g115 ( 
.A1(n_96),
.A2(n_78),
.B1(n_74),
.B2(n_61),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_115),
.A2(n_125),
.B1(n_126),
.B2(n_139),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_117),
.A2(n_127),
.B1(n_137),
.B2(n_112),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g118 ( 
.A(n_101),
.B(n_72),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_118),
.B(n_119),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g119 ( 
.A(n_93),
.B(n_86),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g123 ( 
.A(n_98),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_123),
.B(n_129),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_106),
.A2(n_84),
.B1(n_83),
.B2(n_71),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_90),
.A2(n_83),
.B1(n_85),
.B2(n_82),
.Y(n_127)
);

XOR2xp5_ASAP7_75t_L g155 ( 
.A(n_128),
.B(n_100),
.Y(n_155)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_98),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_93),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_130),
.B(n_135),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_95),
.B(n_83),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_131),
.B(n_132),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_105),
.B(n_83),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_102),
.B(n_80),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_133),
.B(n_141),
.Y(n_163)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_91),
.Y(n_134)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_134),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_94),
.B(n_16),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_110),
.A2(n_44),
.B(n_59),
.Y(n_136)
);

OAI21xp5_ASAP7_75t_SL g159 ( 
.A1(n_136),
.A2(n_89),
.B(n_104),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g137 ( 
.A1(n_102),
.A2(n_68),
.B1(n_64),
.B2(n_59),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_138),
.A2(n_23),
.B(n_22),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_107),
.A2(n_64),
.B1(n_19),
.B2(n_22),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_94),
.B(n_64),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g142 ( 
.A(n_99),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_142),
.B(n_129),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_121),
.B(n_114),
.Y(n_143)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_143),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g144 ( 
.A1(n_136),
.A2(n_97),
.B(n_110),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_144),
.A2(n_159),
.B(n_162),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_145),
.A2(n_160),
.B1(n_0),
.B2(n_1),
.Y(n_183)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_140),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_147),
.B(n_150),
.Y(n_193)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_124),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_148),
.B(n_134),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_141),
.B(n_99),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_123),
.A2(n_108),
.B1(n_109),
.B2(n_88),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g178 ( 
.A1(n_151),
.A2(n_165),
.B(n_124),
.Y(n_178)
);

NOR4xp25_ASAP7_75t_L g154 ( 
.A(n_115),
.B(n_97),
.C(n_88),
.D(n_16),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_154),
.B(n_166),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_155),
.B(n_156),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g156 ( 
.A(n_137),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_111),
.Y(n_158)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_158),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_132),
.A2(n_104),
.B1(n_22),
.B2(n_17),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_161),
.B(n_167),
.Y(n_175)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_125),
.B(n_23),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g166 ( 
.A(n_122),
.B(n_23),
.Y(n_166)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_117),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_131),
.A2(n_17),
.B(n_1),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g196 ( 
.A1(n_168),
.A2(n_169),
.B(n_8),
.Y(n_196)
);

OAI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_128),
.A2(n_119),
.B(n_127),
.Y(n_169)
);

OAI22x1_ASAP7_75t_SL g170 ( 
.A1(n_126),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g174 ( 
.A1(n_170),
.A2(n_118),
.B1(n_116),
.B2(n_120),
.Y(n_174)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_133),
.Y(n_171)
);

INVx1_ASAP7_75t_SL g186 ( 
.A(n_171),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_152),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_172),
.B(n_177),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_174),
.A2(n_181),
.B1(n_184),
.B2(n_188),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g177 ( 
.A(n_146),
.B(n_116),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_178),
.A2(n_162),
.B1(n_159),
.B2(n_164),
.Y(n_210)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_180),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_167),
.A2(n_139),
.B1(n_122),
.B2(n_120),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_183),
.A2(n_195),
.B1(n_149),
.B2(n_156),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_170),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_166),
.B(n_14),
.C(n_4),
.Y(n_185)
);

XNOR2xp5_ASAP7_75t_L g211 ( 
.A(n_185),
.B(n_190),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_171),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g189 ( 
.A(n_148),
.Y(n_189)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_155),
.B(n_3),
.C(n_5),
.Y(n_190)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_169),
.B(n_14),
.C(n_6),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_191),
.B(n_196),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_153),
.B(n_5),
.Y(n_192)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_146),
.B(n_7),
.Y(n_194)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_194),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g195 ( 
.A1(n_163),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_195)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_182),
.B(n_144),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_197),
.B(n_207),
.Y(n_217)
);

BUFx4f_ASAP7_75t_SL g198 ( 
.A(n_186),
.Y(n_198)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_198),
.Y(n_223)
);

MAJx2_ASAP7_75t_L g199 ( 
.A(n_182),
.B(n_168),
.C(n_165),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_210),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g200 ( 
.A(n_193),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_200),
.B(n_201),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g201 ( 
.A(n_179),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_187),
.B(n_157),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_202),
.B(n_205),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_188),
.B(n_149),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_173),
.B(n_145),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g209 ( 
.A(n_192),
.B(n_151),
.Y(n_209)
);

AOI31xp33_ASAP7_75t_L g228 ( 
.A1(n_209),
.A2(n_215),
.A3(n_213),
.B(n_203),
.Y(n_228)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_189),
.Y(n_215)
);

OAI322xp33_ASAP7_75t_L g218 ( 
.A1(n_208),
.A2(n_191),
.A3(n_196),
.B1(n_185),
.B2(n_178),
.C1(n_190),
.C2(n_177),
.Y(n_218)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_218),
.B(n_220),
.Y(n_240)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_212),
.A2(n_183),
.B1(n_175),
.B2(n_186),
.Y(n_219)
);

AOI22xp5_ASAP7_75t_L g241 ( 
.A1(n_219),
.A2(n_198),
.B1(n_12),
.B2(n_13),
.Y(n_241)
);

MAJx2_ASAP7_75t_L g220 ( 
.A(n_197),
.B(n_176),
.C(n_173),
.Y(n_220)
);

INVx13_ASAP7_75t_L g224 ( 
.A(n_204),
.Y(n_224)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_224),
.Y(n_242)
);

A2O1A1Ixp33_ASAP7_75t_SL g225 ( 
.A1(n_210),
.A2(n_176),
.B(n_175),
.C(n_181),
.Y(n_225)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_225),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_195),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g234 ( 
.A(n_226),
.B(n_214),
.Y(n_234)
);

AOI21x1_ASAP7_75t_L g227 ( 
.A1(n_199),
.A2(n_163),
.B(n_162),
.Y(n_227)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_227),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_228),
.B(n_230),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_211),
.B(n_152),
.C(n_160),
.Y(n_230)
);

MAJx2_ASAP7_75t_L g231 ( 
.A(n_207),
.B(n_184),
.C(n_12),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_231),
.B(n_198),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_229),
.B(n_214),
.C(n_212),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_233),
.B(n_237),
.Y(n_254)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_234),
.B(n_239),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_232),
.B(n_205),
.C(n_216),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_217),
.B(n_222),
.C(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_238),
.B(n_244),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_241),
.B(n_224),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g244 ( 
.A(n_217),
.B(n_225),
.C(n_231),
.Y(n_244)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_246),
.Y(n_256)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_242),
.Y(n_248)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_248),
.Y(n_258)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

XNOR2xp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_220),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g257 ( 
.A(n_250),
.B(n_221),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_236),
.B(n_223),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_251),
.B(n_252),
.Y(n_259)
);

INVx6_ASAP7_75t_L g252 ( 
.A(n_235),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_234),
.B(n_225),
.C(n_223),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_253),
.B(n_11),
.Y(n_260)
);

AOI21xp33_ASAP7_75t_L g255 ( 
.A1(n_243),
.A2(n_240),
.B(n_221),
.Y(n_255)
);

OAI21x1_ASAP7_75t_L g263 ( 
.A1(n_255),
.A2(n_11),
.B(n_247),
.Y(n_263)
);

XNOR2xp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_250),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g265 ( 
.A1(n_260),
.A2(n_11),
.B(n_254),
.Y(n_265)
);

INVxp67_ASAP7_75t_L g262 ( 
.A(n_253),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_262),
.B(n_256),
.Y(n_269)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_263),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_264),
.B(n_269),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_265),
.B(n_266),
.Y(n_272)
);

AOI21xp5_ASAP7_75t_L g266 ( 
.A1(n_262),
.A2(n_252),
.B(n_245),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_261),
.B(n_245),
.C(n_259),
.Y(n_268)
);

AND2x2_ASAP7_75t_L g271 ( 
.A(n_268),
.B(n_258),
.Y(n_271)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_271),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g273 ( 
.A(n_268),
.B(n_267),
.Y(n_273)
);

AO21x1_ASAP7_75t_L g275 ( 
.A1(n_273),
.A2(n_272),
.B(n_270),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_275),
.Y(n_276)
);

AOI21xp5_ASAP7_75t_L g277 ( 
.A1(n_276),
.A2(n_274),
.B(n_272),
.Y(n_277)
);

HB1xp67_ASAP7_75t_L g278 ( 
.A(n_277),
.Y(n_278)
);


endmodule