module fake_jpeg_18926_n_377 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_377);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_377;

wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

BUFx5_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_8),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_15),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_14),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx12_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_0),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_15),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_2),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_29),
.Y(n_46)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx4_ASAP7_75t_L g47 ( 
.A(n_19),
.Y(n_47)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_47),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_48),
.Y(n_109)
);

INVx4_ASAP7_75t_L g49 ( 
.A(n_19),
.Y(n_49)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_50),
.Y(n_119)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_51),
.Y(n_122)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_34),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g89 ( 
.A(n_52),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_31),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_31),
.Y(n_54)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_54),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_38),
.B(n_16),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g88 ( 
.A(n_55),
.B(n_59),
.Y(n_88)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_56),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_17),
.Y(n_57)
);

INVx5_ASAP7_75t_SL g116 ( 
.A(n_57),
.Y(n_116)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_38),
.B(n_16),
.Y(n_59)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_17),
.Y(n_60)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_60),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_61),
.Y(n_87)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_41),
.Y(n_62)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_62),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_23),
.Y(n_63)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_63),
.Y(n_117)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_29),
.Y(n_64)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_64),
.Y(n_104)
);

INVx6_ASAP7_75t_L g65 ( 
.A(n_41),
.Y(n_65)
);

NAND2xp33_ASAP7_75t_SL g99 ( 
.A(n_65),
.B(n_77),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_23),
.Y(n_66)
);

INVx2_ASAP7_75t_L g125 ( 
.A(n_66),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_67),
.B(n_68),
.Y(n_106)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_26),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_35),
.Y(n_69)
);

INVx2_ASAP7_75t_L g130 ( 
.A(n_69),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_35),
.Y(n_70)
);

INVx5_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_20),
.B(n_27),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_71),
.B(n_74),
.Y(n_94)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_34),
.Y(n_72)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_72),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_35),
.Y(n_73)
);

INVx5_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_20),
.B(n_1),
.Y(n_74)
);

INVx5_ASAP7_75t_L g75 ( 
.A(n_26),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_75),
.B(n_79),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g76 ( 
.A(n_41),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g84 ( 
.A(n_76),
.Y(n_84)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_41),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g78 ( 
.A(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_78),
.B(n_37),
.Y(n_107)
);

INVx8_ASAP7_75t_L g79 ( 
.A(n_39),
.Y(n_79)
);

INVx4_ASAP7_75t_L g80 ( 
.A(n_28),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_80),
.B(n_81),
.Y(n_113)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx6_ASAP7_75t_L g82 ( 
.A(n_36),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g97 ( 
.A1(n_82),
.A2(n_26),
.B1(n_39),
.B2(n_32),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_SL g90 ( 
.A(n_74),
.B(n_43),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_90),
.B(n_95),
.Y(n_160)
);

NAND2x1_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_32),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g136 ( 
.A(n_93),
.B(n_121),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_43),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_97),
.A2(n_30),
.B1(n_38),
.B2(n_32),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_82),
.A2(n_79),
.B1(n_51),
.B2(n_42),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_103),
.A2(n_105),
.B1(n_112),
.B2(n_123),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g105 ( 
.A1(n_59),
.A2(n_27),
.B1(n_25),
.B2(n_42),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g148 ( 
.A(n_107),
.Y(n_148)
);

AND2x2_ASAP7_75t_L g108 ( 
.A(n_76),
.B(n_37),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_108),
.B(n_115),
.Y(n_139)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_61),
.A2(n_21),
.B1(n_25),
.B2(n_33),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_48),
.B(n_44),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_126),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_63),
.B(n_21),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_50),
.B(n_44),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_118),
.B(n_124),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_53),
.B(n_37),
.C(n_36),
.Y(n_121)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_73),
.A2(n_18),
.B1(n_22),
.B2(n_24),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_54),
.B(n_24),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_70),
.B(n_18),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_66),
.A2(n_40),
.B1(n_33),
.B2(n_30),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_127),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_69),
.B(n_22),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_128),
.B(n_129),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_74),
.B(n_40),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_71),
.B(n_38),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_131),
.B(n_133),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_55),
.B(n_28),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g199 ( 
.A(n_134),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_84),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_135),
.B(n_142),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_112),
.A2(n_32),
.B1(n_28),
.B2(n_3),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_137),
.A2(n_138),
.B1(n_155),
.B2(n_171),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_L g138 ( 
.A1(n_87),
.A2(n_8),
.B1(n_14),
.B2(n_13),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_94),
.B(n_88),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_140),
.B(n_89),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_84),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_88),
.B(n_1),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_143),
.B(n_144),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_85),
.B(n_1),
.Y(n_144)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_100),
.Y(n_146)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_146),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_104),
.B(n_2),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_147),
.B(n_170),
.Y(n_186)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_100),
.Y(n_149)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_149),
.Y(n_191)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_151),
.Y(n_192)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_96),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_156),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_109),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_154),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_127),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_155)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_110),
.Y(n_156)
);

INVx3_ASAP7_75t_L g157 ( 
.A(n_96),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_157),
.B(n_168),
.Y(n_188)
);

BUFx2_ASAP7_75t_L g159 ( 
.A(n_109),
.Y(n_159)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_159),
.Y(n_202)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_93),
.B(n_133),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_161),
.B(n_172),
.C(n_175),
.Y(n_180)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_111),
.Y(n_162)
);

BUFx12f_ASAP7_75t_L g198 ( 
.A(n_162),
.Y(n_198)
);

INVx11_ASAP7_75t_L g164 ( 
.A(n_89),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_164),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g165 ( 
.A(n_86),
.Y(n_165)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_165),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_4),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g204 ( 
.A(n_166),
.B(n_174),
.Y(n_204)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_120),
.Y(n_167)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_167),
.Y(n_212)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_120),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_91),
.Y(n_169)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_169),
.Y(n_213)
);

A2O1A1Ixp33_ASAP7_75t_L g170 ( 
.A1(n_99),
.A2(n_5),
.B(n_6),
.C(n_8),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_L g171 ( 
.A1(n_87),
.A2(n_5),
.B1(n_6),
.B2(n_10),
.Y(n_171)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_99),
.B(n_6),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_121),
.B(n_10),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_173),
.B(n_89),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_106),
.B(n_11),
.Y(n_174)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_102),
.B(n_11),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_176),
.A2(n_125),
.B1(n_117),
.B2(n_91),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_148),
.B(n_130),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g228 ( 
.A1(n_178),
.A2(n_195),
.B(n_205),
.Y(n_228)
);

INVxp33_ASAP7_75t_L g179 ( 
.A(n_165),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_179),
.B(n_184),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_136),
.B(n_161),
.C(n_145),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_183),
.B(n_187),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_149),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_185),
.B(n_189),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_136),
.B(n_108),
.C(n_132),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_141),
.B(n_86),
.Y(n_189)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_98),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_193),
.B(n_196),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_194),
.B(n_144),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g195 ( 
.A(n_139),
.B(n_130),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_160),
.B(n_98),
.Y(n_196)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_197),
.B(n_203),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_150),
.B(n_101),
.Y(n_203)
);

NAND2x1_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_172),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_140),
.B(n_83),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_206),
.B(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g224 ( 
.A1(n_209),
.A2(n_103),
.B1(n_92),
.B2(n_117),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_163),
.B(n_83),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_214),
.B(n_172),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_223),
.Y(n_251)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_186),
.A2(n_205),
.B(n_199),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_219),
.A2(n_233),
.B(n_180),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_187),
.A2(n_161),
.B1(n_175),
.B2(n_170),
.Y(n_220)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_220),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_186),
.B(n_143),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_SL g247 ( 
.A(n_221),
.B(n_245),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g222 ( 
.A(n_205),
.B(n_173),
.Y(n_222)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_222),
.B(n_180),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_224),
.A2(n_232),
.B1(n_234),
.B2(n_244),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_194),
.B(n_147),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_225),
.B(n_240),
.Y(n_255)
);

INVxp33_ASAP7_75t_SL g227 ( 
.A(n_182),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g269 ( 
.A(n_227),
.Y(n_269)
);

CKINVDCx16_ASAP7_75t_R g229 ( 
.A(n_177),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_192),
.B(n_165),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_190),
.Y(n_231)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_231),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_208),
.A2(n_158),
.B1(n_137),
.B2(n_97),
.Y(n_232)
);

OAI21xp5_ASAP7_75t_SL g233 ( 
.A1(n_199),
.A2(n_175),
.B(n_155),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_SL g234 ( 
.A1(n_208),
.A2(n_125),
.B1(n_92),
.B2(n_119),
.Y(n_234)
);

NOR2x1_ASAP7_75t_L g235 ( 
.A(n_178),
.B(n_171),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_L g270 ( 
.A1(n_235),
.A2(n_207),
.B(n_202),
.Y(n_270)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_190),
.Y(n_236)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_236),
.Y(n_253)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_211),
.Y(n_238)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_238),
.Y(n_258)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_191),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_239),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g240 ( 
.A(n_181),
.B(n_167),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_181),
.B(n_214),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_241),
.B(n_242),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_178),
.B(n_159),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_209),
.A2(n_119),
.B1(n_157),
.B2(n_152),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g245 ( 
.A(n_195),
.B(n_162),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_195),
.B(n_168),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g260 ( 
.A(n_246),
.B(n_197),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_248),
.A2(n_221),
.B(n_242),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_231),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_256),
.B(n_259),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g259 ( 
.A(n_216),
.Y(n_259)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_241),
.B(n_183),
.Y(n_261)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_261),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_SL g282 ( 
.A(n_262),
.B(n_271),
.Y(n_282)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_236),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_263),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_223),
.B(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_264),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_232),
.A2(n_191),
.B1(n_184),
.B2(n_185),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_268),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_234),
.A2(n_200),
.B1(n_212),
.B2(n_213),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_219),
.A2(n_192),
.B1(n_212),
.B2(n_200),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_L g268 ( 
.A1(n_235),
.A2(n_213),
.B1(n_188),
.B2(n_207),
.Y(n_268)
);

AO21x1_ASAP7_75t_L g281 ( 
.A1(n_270),
.A2(n_228),
.B(n_245),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_222),
.B(n_204),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_252),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_275),
.B(n_279),
.Y(n_310)
);

OAI22xp33_ASAP7_75t_SL g278 ( 
.A1(n_250),
.A2(n_235),
.B1(n_233),
.B2(n_216),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g304 ( 
.A1(n_278),
.A2(n_267),
.B1(n_268),
.B2(n_270),
.Y(n_304)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_252),
.Y(n_279)
);

AOI322xp5_ASAP7_75t_SL g280 ( 
.A1(n_249),
.A2(n_217),
.A3(n_220),
.B1(n_229),
.B2(n_237),
.C1(n_243),
.C2(n_218),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_280),
.B(n_291),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_281),
.B(n_285),
.Y(n_299)
);

AOI22xp33_ASAP7_75t_SL g284 ( 
.A1(n_250),
.A2(n_238),
.B1(n_224),
.B2(n_164),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_284),
.A2(n_238),
.B1(n_258),
.B2(n_265),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g285 ( 
.A(n_253),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_262),
.B(n_237),
.C(n_228),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_286),
.B(n_292),
.C(n_271),
.Y(n_303)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_253),
.Y(n_288)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_288),
.Y(n_302)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_260),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_272),
.Y(n_290)
);

INVx1_ASAP7_75t_L g312 ( 
.A(n_290),
.Y(n_312)
);

NOR3xp33_ASAP7_75t_SL g291 ( 
.A(n_272),
.B(n_217),
.C(n_243),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_262),
.B(n_240),
.C(n_246),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g293 ( 
.A(n_270),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g300 ( 
.A(n_293),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_251),
.Y(n_306)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_265),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_295),
.B(n_257),
.Y(n_309)
);

XOR2x1_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_248),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g324 ( 
.A(n_296),
.B(n_305),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g297 ( 
.A(n_286),
.B(n_271),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_297),
.B(n_303),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_298),
.A2(n_311),
.B1(n_313),
.B2(n_287),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_304),
.B(n_306),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_SL g305 ( 
.A(n_292),
.B(n_261),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_282),
.B(n_264),
.C(n_255),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g320 ( 
.A(n_308),
.B(n_314),
.C(n_294),
.Y(n_320)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_309),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_295),
.A2(n_254),
.B1(n_257),
.B2(n_255),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_L g313 ( 
.A1(n_290),
.A2(n_254),
.B1(n_269),
.B2(n_226),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_282),
.B(n_251),
.C(n_247),
.Y(n_314)
);

HB1xp67_ASAP7_75t_L g315 ( 
.A(n_299),
.Y(n_315)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_315),
.Y(n_333)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_310),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_317),
.B(n_319),
.Y(n_341)
);

INVx2_ASAP7_75t_L g319 ( 
.A(n_296),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_320),
.B(n_321),
.C(n_325),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_303),
.B(n_274),
.C(n_283),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_L g332 ( 
.A1(n_322),
.A2(n_326),
.B1(n_254),
.B2(n_304),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_SL g323 ( 
.A(n_301),
.B(n_312),
.Y(n_323)
);

NOR2xp33_ASAP7_75t_SL g335 ( 
.A(n_323),
.B(n_247),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_297),
.B(n_274),
.C(n_283),
.Y(n_325)
);

OA21x2_ASAP7_75t_L g326 ( 
.A1(n_299),
.A2(n_277),
.B(n_289),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g327 ( 
.A(n_306),
.B(n_291),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g331 ( 
.A(n_327),
.B(n_329),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_305),
.B(n_277),
.C(n_287),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g338 ( 
.A(n_328),
.B(n_308),
.C(n_314),
.Y(n_338)
);

INVx1_ASAP7_75t_SL g329 ( 
.A(n_302),
.Y(n_329)
);

AOI22xp5_ASAP7_75t_L g346 ( 
.A1(n_332),
.A2(n_273),
.B1(n_285),
.B2(n_326),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_328),
.B(n_269),
.Y(n_334)
);

OAI221xp5_ASAP7_75t_L g354 ( 
.A1(n_334),
.A2(n_340),
.B1(n_266),
.B2(n_239),
.C(n_215),
.Y(n_354)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_335),
.B(n_339),
.Y(n_348)
);

AO21x1_ASAP7_75t_L g336 ( 
.A1(n_318),
.A2(n_309),
.B(n_300),
.Y(n_336)
);

AOI21xp5_ASAP7_75t_L g349 ( 
.A1(n_336),
.A2(n_331),
.B(n_342),
.Y(n_349)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_266),
.Y(n_353)
);

HB1xp67_ASAP7_75t_L g339 ( 
.A(n_321),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_320),
.B(n_226),
.Y(n_340)
);

OAI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_316),
.A2(n_307),
.B1(n_273),
.B2(n_276),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_342),
.A2(n_263),
.B1(n_256),
.B2(n_288),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_325),
.B(n_330),
.C(n_324),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_343),
.B(n_330),
.C(n_326),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_SL g344 ( 
.A1(n_341),
.A2(n_276),
.B(n_329),
.Y(n_344)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_344),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g363 ( 
.A(n_345),
.B(n_350),
.Y(n_363)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_346),
.A2(n_122),
.B1(n_116),
.B2(n_211),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_347),
.B(n_351),
.Y(n_359)
);

OAI21xp5_ASAP7_75t_L g355 ( 
.A1(n_349),
.A2(n_352),
.B(n_244),
.Y(n_355)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_338),
.B(n_337),
.Y(n_350)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_333),
.A2(n_311),
.B(n_215),
.Y(n_351)
);

OAI21xp5_ASAP7_75t_L g352 ( 
.A1(n_336),
.A2(n_337),
.B(n_343),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_353),
.B(n_169),
.C(n_198),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g361 ( 
.A(n_354),
.B(n_198),
.Y(n_361)
);

CKINVDCx16_ASAP7_75t_R g366 ( 
.A(n_355),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_348),
.A2(n_202),
.B1(n_201),
.B2(n_211),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_356),
.B(n_357),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_358),
.B(n_360),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_353),
.B(n_198),
.C(n_154),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g369 ( 
.A1(n_361),
.A2(n_352),
.B(n_345),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_359),
.B(n_347),
.Y(n_367)
);

NAND2xp5_ASAP7_75t_SL g372 ( 
.A(n_367),
.B(n_368),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g368 ( 
.A(n_362),
.B(n_350),
.Y(n_368)
);

XOR2xp5_ASAP7_75t_L g371 ( 
.A(n_369),
.B(n_358),
.Y(n_371)
);

OAI21x1_ASAP7_75t_L g370 ( 
.A1(n_369),
.A2(n_363),
.B(n_355),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g375 ( 
.A(n_370),
.B(n_371),
.Y(n_375)
);

OAI21xp5_ASAP7_75t_L g373 ( 
.A1(n_365),
.A2(n_360),
.B(n_356),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_373),
.A2(n_366),
.B(n_364),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_L g376 ( 
.A(n_374),
.B(n_372),
.Y(n_376)
);

XOR2xp5_ASAP7_75t_L g377 ( 
.A(n_376),
.B(n_375),
.Y(n_377)
);


endmodule