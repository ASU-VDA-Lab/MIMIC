module fake_aes_3305_n_15 (n_1, n_2, n_4, n_3, n_5, n_0, n_15);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_15;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_9;
wire n_14;
wire n_7;
wire n_10;
wire n_8;
AND2x2_ASAP7_75t_L g6 ( .A(n_2), .B(n_5), .Y(n_6) );
INVx1_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
NAND3xp33_ASAP7_75t_L g8 ( .A(n_2), .B(n_3), .C(n_0), .Y(n_8) );
NAND2xp5_ASAP7_75t_SL g9 ( .A(n_0), .B(n_1), .Y(n_9) );
INVx2_ASAP7_75t_L g10 ( .A(n_7), .Y(n_10) );
HB1xp67_ASAP7_75t_L g11 ( .A(n_9), .Y(n_11) );
NOR2x1_ASAP7_75t_L g12 ( .A(n_10), .B(n_8), .Y(n_12) );
NAND2xp5_ASAP7_75t_SL g13 ( .A(n_12), .B(n_11), .Y(n_13) );
XOR2xp5_ASAP7_75t_L g14 ( .A(n_13), .B(n_9), .Y(n_14) );
OAI21x1_ASAP7_75t_SL g15 ( .A1(n_14), .A2(n_1), .B(n_6), .Y(n_15) );
endmodule