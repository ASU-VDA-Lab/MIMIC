module fake_netlist_6_4785_n_1689 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_68, n_28, n_50, n_49, n_7, n_83, n_5, n_101, n_144, n_127, n_125, n_153, n_77, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_31, n_57, n_53, n_51, n_44, n_56, n_1689);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_68;
input n_28;
input n_50;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_144;
input n_127;
input n_125;
input n_153;
input n_77;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_31;
input n_57;
input n_53;
input n_51;
input n_44;
input n_56;

output n_1689;

wire n_992;
wire n_1671;
wire n_801;
wire n_1613;
wire n_1234;
wire n_1458;
wire n_1199;
wire n_1674;
wire n_741;
wire n_1027;
wire n_1351;
wire n_625;
wire n_1189;
wire n_223;
wire n_1212;
wire n_226;
wire n_208;
wire n_726;
wire n_212;
wire n_700;
wire n_1307;
wire n_1038;
wire n_578;
wire n_1581;
wire n_1003;
wire n_365;
wire n_168;
wire n_1237;
wire n_1061;
wire n_1357;
wire n_783;
wire n_798;
wire n_188;
wire n_1575;
wire n_509;
wire n_1342;
wire n_245;
wire n_1209;
wire n_1348;
wire n_1387;
wire n_677;
wire n_805;
wire n_1151;
wire n_396;
wire n_350;
wire n_1380;
wire n_442;
wire n_480;
wire n_1402;
wire n_1688;
wire n_1009;
wire n_1160;
wire n_883;
wire n_1238;
wire n_1032;
wire n_1247;
wire n_1547;
wire n_1553;
wire n_893;
wire n_1099;
wire n_1264;
wire n_1192;
wire n_471;
wire n_424;
wire n_1555;
wire n_1415;
wire n_1370;
wire n_369;
wire n_287;
wire n_415;
wire n_830;
wire n_230;
wire n_461;
wire n_873;
wire n_383;
wire n_1285;
wire n_1371;
wire n_200;
wire n_447;
wire n_1172;
wire n_852;
wire n_229;
wire n_1590;
wire n_1532;
wire n_1393;
wire n_1517;
wire n_1078;
wire n_544;
wire n_250;
wire n_1140;
wire n_1444;
wire n_1670;
wire n_1603;
wire n_1579;
wire n_1263;
wire n_836;
wire n_375;
wire n_522;
wire n_1261;
wire n_945;
wire n_1649;
wire n_1511;
wire n_1143;
wire n_1422;
wire n_1232;
wire n_1572;
wire n_616;
wire n_658;
wire n_1119;
wire n_428;
wire n_1433;
wire n_1620;
wire n_1541;
wire n_1300;
wire n_641;
wire n_822;
wire n_693;
wire n_1313;
wire n_1056;
wire n_758;
wire n_516;
wire n_1455;
wire n_1163;
wire n_1180;
wire n_943;
wire n_1550;
wire n_491;
wire n_1591;
wire n_772;
wire n_1344;
wire n_666;
wire n_371;
wire n_940;
wire n_770;
wire n_567;
wire n_405;
wire n_213;
wire n_538;
wire n_1106;
wire n_886;
wire n_1471;
wire n_343;
wire n_953;
wire n_1094;
wire n_1345;
wire n_494;
wire n_539;
wire n_493;
wire n_155;
wire n_454;
wire n_1421;
wire n_638;
wire n_1404;
wire n_1211;
wire n_381;
wire n_887;
wire n_1660;
wire n_1280;
wire n_713;
wire n_1400;
wire n_1467;
wire n_976;
wire n_224;
wire n_1445;
wire n_1560;
wire n_1526;
wire n_734;
wire n_1088;
wire n_196;
wire n_1231;
wire n_917;
wire n_574;
wire n_907;
wire n_1446;
wire n_659;
wire n_407;
wire n_913;
wire n_1658;
wire n_808;
wire n_867;
wire n_1230;
wire n_473;
wire n_1193;
wire n_1054;
wire n_559;
wire n_1333;
wire n_1648;
wire n_163;
wire n_1644;
wire n_1558;
wire n_281;
wire n_551;
wire n_699;
wire n_564;
wire n_451;
wire n_824;
wire n_279;
wire n_686;
wire n_757;
wire n_594;
wire n_1641;
wire n_577;
wire n_166;
wire n_619;
wire n_1367;
wire n_1336;
wire n_521;
wire n_572;
wire n_395;
wire n_813;
wire n_1481;
wire n_323;
wire n_606;
wire n_1441;
wire n_818;
wire n_1123;
wire n_1309;
wire n_513;
wire n_645;
wire n_1381;
wire n_331;
wire n_916;
wire n_483;
wire n_608;
wire n_261;
wire n_630;
wire n_541;
wire n_512;
wire n_433;
wire n_792;
wire n_476;
wire n_1328;
wire n_219;
wire n_264;
wire n_263;
wire n_1162;
wire n_860;
wire n_1530;
wire n_788;
wire n_939;
wire n_1543;
wire n_821;
wire n_938;
wire n_1302;
wire n_1068;
wire n_1599;
wire n_329;
wire n_982;
wire n_549;
wire n_1075;
wire n_408;
wire n_932;
wire n_237;
wire n_243;
wire n_979;
wire n_905;
wire n_1680;
wire n_175;
wire n_322;
wire n_993;
wire n_689;
wire n_354;
wire n_1330;
wire n_1413;
wire n_1605;
wire n_1278;
wire n_547;
wire n_558;
wire n_1064;
wire n_1396;
wire n_634;
wire n_966;
wire n_764;
wire n_1663;
wire n_692;
wire n_733;
wire n_1233;
wire n_1289;
wire n_487;
wire n_241;
wire n_1107;
wire n_1014;
wire n_1290;
wire n_882;
wire n_1354;
wire n_586;
wire n_423;
wire n_318;
wire n_1111;
wire n_715;
wire n_1251;
wire n_1265;
wire n_530;
wire n_1563;
wire n_277;
wire n_618;
wire n_1297;
wire n_1662;
wire n_1312;
wire n_199;
wire n_1167;
wire n_1359;
wire n_674;
wire n_871;
wire n_922;
wire n_268;
wire n_1335;
wire n_210;
wire n_1069;
wire n_1664;
wire n_612;
wire n_178;
wire n_247;
wire n_1165;
wire n_355;
wire n_702;
wire n_347;
wire n_1175;
wire n_328;
wire n_1386;
wire n_429;
wire n_1012;
wire n_195;
wire n_780;
wire n_675;
wire n_903;
wire n_1540;
wire n_1504;
wire n_286;
wire n_254;
wire n_1655;
wire n_242;
wire n_835;
wire n_928;
wire n_1214;
wire n_690;
wire n_850;
wire n_1654;
wire n_816;
wire n_1157;
wire n_1462;
wire n_1188;
wire n_877;
wire n_604;
wire n_825;
wire n_728;
wire n_1063;
wire n_1588;
wire n_267;
wire n_1124;
wire n_1624;
wire n_515;
wire n_598;
wire n_696;
wire n_1515;
wire n_961;
wire n_437;
wire n_1082;
wire n_1317;
wire n_593;
wire n_514;
wire n_687;
wire n_697;
wire n_890;
wire n_637;
wire n_295;
wire n_701;
wire n_950;
wire n_388;
wire n_190;
wire n_484;
wire n_170;
wire n_891;
wire n_1412;
wire n_949;
wire n_1630;
wire n_678;
wire n_283;
wire n_507;
wire n_968;
wire n_909;
wire n_1369;
wire n_881;
wire n_1008;
wire n_760;
wire n_1546;
wire n_590;
wire n_362;
wire n_161;
wire n_462;
wire n_1052;
wire n_1033;
wire n_1296;
wire n_304;
wire n_694;
wire n_1294;
wire n_1420;
wire n_1634;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_1465;
wire n_342;
wire n_1044;
wire n_1391;
wire n_449;
wire n_1523;
wire n_1208;
wire n_1164;
wire n_1295;
wire n_1627;
wire n_1072;
wire n_1527;
wire n_1495;
wire n_1438;
wire n_495;
wire n_815;
wire n_1100;
wire n_585;
wire n_1487;
wire n_840;
wire n_874;
wire n_1128;
wire n_382;
wire n_673;
wire n_1071;
wire n_1067;
wire n_1565;
wire n_1493;
wire n_898;
wire n_255;
wire n_284;
wire n_865;
wire n_925;
wire n_1101;
wire n_1026;
wire n_289;
wire n_1364;
wire n_615;
wire n_1249;
wire n_1293;
wire n_1127;
wire n_1512;
wire n_1451;
wire n_320;
wire n_639;
wire n_963;
wire n_794;
wire n_727;
wire n_894;
wire n_685;
wire n_353;
wire n_605;
wire n_1514;
wire n_826;
wire n_1646;
wire n_872;
wire n_1139;
wire n_718;
wire n_1018;
wire n_1521;
wire n_1366;
wire n_542;
wire n_847;
wire n_644;
wire n_682;
wire n_851;
wire n_305;
wire n_996;
wire n_532;
wire n_173;
wire n_1308;
wire n_1376;
wire n_1513;
wire n_413;
wire n_791;
wire n_510;
wire n_837;
wire n_1488;
wire n_948;
wire n_704;
wire n_977;
wire n_1005;
wire n_536;
wire n_622;
wire n_1469;
wire n_581;
wire n_765;
wire n_432;
wire n_987;
wire n_1492;
wire n_1340;
wire n_631;
wire n_720;
wire n_842;
wire n_1432;
wire n_156;
wire n_843;
wire n_656;
wire n_989;
wire n_1277;
wire n_797;
wire n_1473;
wire n_1246;
wire n_899;
wire n_189;
wire n_738;
wire n_1304;
wire n_1035;
wire n_294;
wire n_499;
wire n_1426;
wire n_705;
wire n_1004;
wire n_1176;
wire n_1529;
wire n_1022;
wire n_614;
wire n_529;
wire n_425;
wire n_684;
wire n_1431;
wire n_1615;
wire n_1474;
wire n_1571;
wire n_1577;
wire n_1181;
wire n_486;
wire n_947;
wire n_1117;
wire n_1087;
wire n_1448;
wire n_648;
wire n_657;
wire n_1049;
wire n_1666;
wire n_1505;
wire n_803;
wire n_290;
wire n_926;
wire n_927;
wire n_919;
wire n_478;
wire n_929;
wire n_1228;
wire n_417;
wire n_446;
wire n_1568;
wire n_1490;
wire n_777;
wire n_1299;
wire n_272;
wire n_526;
wire n_1183;
wire n_1436;
wire n_1384;
wire n_293;
wire n_458;
wire n_1070;
wire n_998;
wire n_717;
wire n_1665;
wire n_1383;
wire n_1178;
wire n_1424;
wire n_1073;
wire n_1000;
wire n_796;
wire n_252;
wire n_1195;
wire n_1626;
wire n_1507;
wire n_184;
wire n_552;
wire n_1358;
wire n_1388;
wire n_216;
wire n_912;
wire n_1519;
wire n_745;
wire n_1284;
wire n_1604;
wire n_1142;
wire n_716;
wire n_1475;
wire n_623;
wire n_1048;
wire n_1201;
wire n_1398;
wire n_884;
wire n_1395;
wire n_731;
wire n_1502;
wire n_1659;
wire n_755;
wire n_931;
wire n_1021;
wire n_474;
wire n_527;
wire n_683;
wire n_811;
wire n_1207;
wire n_312;
wire n_1368;
wire n_1418;
wire n_958;
wire n_292;
wire n_1250;
wire n_1137;
wire n_880;
wire n_889;
wire n_1478;
wire n_589;
wire n_1310;
wire n_819;
wire n_1363;
wire n_1334;
wire n_767;
wire n_1314;
wire n_600;
wire n_964;
wire n_831;
wire n_477;
wire n_954;
wire n_864;
wire n_1110;
wire n_1410;
wire n_399;
wire n_1440;
wire n_1382;
wire n_1534;
wire n_1564;
wire n_211;
wire n_1483;
wire n_1372;
wire n_231;
wire n_1457;
wire n_505;
wire n_319;
wire n_1339;
wire n_537;
wire n_1427;
wire n_311;
wire n_1466;
wire n_403;
wire n_1080;
wire n_723;
wire n_596;
wire n_546;
wire n_562;
wire n_1141;
wire n_1268;
wire n_386;
wire n_1220;
wire n_556;
wire n_162;
wire n_1602;
wire n_1136;
wire n_1125;
wire n_970;
wire n_642;
wire n_995;
wire n_276;
wire n_1159;
wire n_1092;
wire n_441;
wire n_221;
wire n_1060;
wire n_444;
wire n_1252;
wire n_1223;
wire n_303;
wire n_511;
wire n_193;
wire n_1286;
wire n_1053;
wire n_416;
wire n_1681;
wire n_520;
wire n_418;
wire n_1093;
wire n_1533;
wire n_1597;
wire n_266;
wire n_296;
wire n_775;
wire n_651;
wire n_1153;
wire n_439;
wire n_1618;
wire n_217;
wire n_518;
wire n_1531;
wire n_1185;
wire n_453;
wire n_215;
wire n_914;
wire n_759;
wire n_426;
wire n_317;
wire n_1653;
wire n_1679;
wire n_1625;
wire n_1453;
wire n_488;
wire n_497;
wire n_773;
wire n_920;
wire n_1374;
wire n_1315;
wire n_1647;
wire n_1224;
wire n_1614;
wire n_1459;
wire n_1135;
wire n_1169;
wire n_1179;
wire n_401;
wire n_324;
wire n_1617;
wire n_335;
wire n_1470;
wire n_463;
wire n_1243;
wire n_848;
wire n_301;
wire n_274;
wire n_1096;
wire n_1091;
wire n_1580;
wire n_1425;
wire n_1281;
wire n_1267;
wire n_983;
wire n_427;
wire n_1520;
wire n_496;
wire n_906;
wire n_1390;
wire n_688;
wire n_1077;
wire n_1419;
wire n_351;
wire n_259;
wire n_177;
wire n_1636;
wire n_1437;
wire n_1645;
wire n_385;
wire n_1687;
wire n_1439;
wire n_1323;
wire n_858;
wire n_1331;
wire n_613;
wire n_736;
wire n_501;
wire n_956;
wire n_960;
wire n_663;
wire n_856;
wire n_379;
wire n_778;
wire n_1668;
wire n_1134;
wire n_410;
wire n_1129;
wire n_554;
wire n_602;
wire n_1594;
wire n_664;
wire n_171;
wire n_169;
wire n_1429;
wire n_1610;
wire n_435;
wire n_793;
wire n_326;
wire n_587;
wire n_1593;
wire n_580;
wire n_762;
wire n_1030;
wire n_1202;
wire n_465;
wire n_1635;
wire n_1079;
wire n_341;
wire n_828;
wire n_607;
wire n_316;
wire n_419;
wire n_1551;
wire n_1103;
wire n_1203;
wire n_820;
wire n_951;
wire n_725;
wire n_952;
wire n_999;
wire n_358;
wire n_1254;
wire n_160;
wire n_186;
wire n_368;
wire n_575;
wire n_994;
wire n_1508;
wire n_732;
wire n_974;
wire n_392;
wire n_724;
wire n_1020;
wire n_1042;
wire n_628;
wire n_1273;
wire n_1434;
wire n_1573;
wire n_557;
wire n_349;
wire n_617;
wire n_845;
wire n_807;
wire n_1036;
wire n_1138;
wire n_1661;
wire n_1275;
wire n_485;
wire n_1549;
wire n_443;
wire n_1510;
wire n_892;
wire n_768;
wire n_421;
wire n_1468;
wire n_238;
wire n_1095;
wire n_1595;
wire n_202;
wire n_1683;
wire n_597;
wire n_280;
wire n_1270;
wire n_1187;
wire n_610;
wire n_1403;
wire n_1669;
wire n_1024;
wire n_198;
wire n_179;
wire n_248;
wire n_517;
wire n_1667;
wire n_667;
wire n_1206;
wire n_621;
wire n_1037;
wire n_1397;
wire n_1279;
wire n_1115;
wire n_750;
wire n_901;
wire n_1499;
wire n_468;
wire n_923;
wire n_504;
wire n_1409;
wire n_1639;
wire n_1623;
wire n_183;
wire n_1015;
wire n_1503;
wire n_466;
wire n_1057;
wire n_603;
wire n_991;
wire n_1657;
wire n_235;
wire n_1126;
wire n_340;
wire n_710;
wire n_1108;
wire n_1182;
wire n_1298;
wire n_1611;
wire n_785;
wire n_746;
wire n_609;
wire n_1601;
wire n_1686;
wire n_167;
wire n_1356;
wire n_1589;
wire n_1497;
wire n_1168;
wire n_1216;
wire n_1320;
wire n_1430;
wire n_1316;
wire n_1287;
wire n_1452;
wire n_1622;
wire n_1586;
wire n_302;
wire n_380;
wire n_1535;
wire n_1596;
wire n_1190;
wire n_397;
wire n_1262;
wire n_218;
wire n_1213;
wire n_1350;
wire n_1673;
wire n_172;
wire n_1443;
wire n_1272;
wire n_239;
wire n_782;
wire n_1539;
wire n_490;
wire n_220;
wire n_809;
wire n_1043;
wire n_1608;
wire n_986;
wire n_1472;
wire n_1081;
wire n_402;
wire n_352;
wire n_800;
wire n_1084;
wire n_1171;
wire n_460;
wire n_1361;
wire n_1491;
wire n_662;
wire n_374;
wire n_1152;
wire n_450;
wire n_1684;
wire n_921;
wire n_1346;
wire n_711;
wire n_1642;
wire n_579;
wire n_1352;
wire n_937;
wire n_1682;
wire n_370;
wire n_650;
wire n_1046;
wire n_1145;
wire n_330;
wire n_1121;
wire n_1102;
wire n_972;
wire n_1405;
wire n_258;
wire n_1406;
wire n_456;
wire n_1332;
wire n_260;
wire n_313;
wire n_624;
wire n_962;
wire n_1041;
wire n_565;
wire n_356;
wire n_1569;
wire n_936;
wire n_1288;
wire n_1186;
wire n_1062;
wire n_885;
wire n_896;
wire n_654;
wire n_411;
wire n_1222;
wire n_599;
wire n_776;
wire n_321;
wire n_227;
wire n_204;
wire n_482;
wire n_934;
wire n_1637;
wire n_1407;
wire n_420;
wire n_1341;
wire n_394;
wire n_1456;
wire n_1489;
wire n_164;
wire n_942;
wire n_1524;
wire n_543;
wire n_1496;
wire n_1271;
wire n_1545;
wire n_1355;
wire n_1225;
wire n_1544;
wire n_1485;
wire n_325;
wire n_1640;
wire n_804;
wire n_464;
wire n_533;
wire n_806;
wire n_879;
wire n_959;
wire n_584;
wire n_244;
wire n_1343;
wire n_1522;
wire n_548;
wire n_282;
wire n_1676;
wire n_833;
wire n_1567;
wire n_523;
wire n_1319;
wire n_707;
wire n_345;
wire n_799;
wire n_1548;
wire n_1155;
wire n_273;
wire n_1633;
wire n_787;
wire n_1416;
wire n_1528;
wire n_1146;
wire n_159;
wire n_1086;
wire n_1066;
wire n_157;
wire n_1282;
wire n_550;
wire n_275;
wire n_652;
wire n_560;
wire n_1484;
wire n_1241;
wire n_1321;
wire n_1672;
wire n_569;
wire n_737;
wire n_1318;
wire n_1235;
wire n_1229;
wire n_306;
wire n_1292;
wire n_1373;
wire n_346;
wire n_1029;
wire n_1447;
wire n_790;
wire n_1498;
wire n_1210;
wire n_299;
wire n_1248;
wire n_1556;
wire n_902;
wire n_333;
wire n_1047;
wire n_1385;
wire n_431;
wire n_459;
wire n_1269;
wire n_502;
wire n_672;
wire n_1257;
wire n_285;
wire n_1375;
wire n_655;
wire n_706;
wire n_1045;
wire n_1650;
wire n_786;
wire n_1236;
wire n_1559;
wire n_834;
wire n_743;
wire n_766;
wire n_430;
wire n_1325;
wire n_1002;
wire n_545;
wire n_489;
wire n_251;
wire n_1019;
wire n_636;
wire n_729;
wire n_876;
wire n_774;
wire n_1337;
wire n_660;
wire n_438;
wire n_1477;
wire n_1360;
wire n_1200;
wire n_479;
wire n_1607;
wire n_1353;
wire n_1454;
wire n_869;
wire n_1154;
wire n_1113;
wire n_1600;
wire n_646;
wire n_528;
wire n_391;
wire n_1098;
wire n_1329;
wire n_817;
wire n_262;
wire n_187;
wire n_897;
wire n_846;
wire n_841;
wire n_1476;
wire n_1001;
wire n_508;
wire n_1050;
wire n_1411;
wire n_1463;
wire n_1177;
wire n_332;
wire n_1150;
wire n_1562;
wire n_398;
wire n_1191;
wire n_566;
wire n_1023;
wire n_1118;
wire n_1076;
wire n_194;
wire n_1007;
wire n_1378;
wire n_855;
wire n_1592;
wire n_1631;
wire n_591;
wire n_1377;
wire n_256;
wire n_853;
wire n_440;
wire n_695;
wire n_1542;
wire n_875;
wire n_209;
wire n_367;
wire n_680;
wire n_1678;
wire n_661;
wire n_278;
wire n_1256;
wire n_671;
wire n_933;
wire n_740;
wire n_703;
wire n_978;
wire n_384;
wire n_1291;
wire n_1217;
wire n_751;
wire n_749;
wire n_310;
wire n_1628;
wire n_1324;
wire n_1399;
wire n_1435;
wire n_969;
wire n_988;
wire n_1065;
wire n_1401;
wire n_1255;
wire n_568;
wire n_1516;
wire n_1536;
wire n_180;
wire n_1204;
wire n_823;
wire n_1132;
wire n_643;
wire n_233;
wire n_698;
wire n_1074;
wire n_1394;
wire n_1327;
wire n_1326;
wire n_739;
wire n_400;
wire n_955;
wire n_337;
wire n_1379;
wire n_214;
wire n_246;
wire n_1338;
wire n_1097;
wire n_935;
wire n_781;
wire n_789;
wire n_1554;
wire n_1130;
wire n_181;
wire n_182;
wire n_573;
wire n_769;
wire n_676;
wire n_327;
wire n_1120;
wire n_832;
wire n_1583;
wire n_555;
wire n_389;
wire n_814;
wire n_1643;
wire n_669;
wire n_176;
wire n_300;
wire n_222;
wire n_747;
wire n_1389;
wire n_1105;
wire n_721;
wire n_1461;
wire n_742;
wire n_535;
wire n_691;
wire n_372;
wire n_314;
wire n_1408;
wire n_378;
wire n_1196;
wire n_377;
wire n_1598;
wire n_863;
wire n_601;
wire n_338;
wire n_1283;
wire n_918;
wire n_748;
wire n_506;
wire n_1114;
wire n_763;
wire n_1147;
wire n_360;
wire n_1506;
wire n_1652;
wire n_957;
wire n_895;
wire n_866;
wire n_1227;
wire n_191;
wire n_387;
wire n_452;
wire n_744;
wire n_971;
wire n_946;
wire n_344;
wire n_761;
wire n_1303;
wire n_1205;
wire n_1258;
wire n_1392;
wire n_174;
wire n_1173;
wire n_525;
wire n_1677;
wire n_1116;
wire n_611;
wire n_1570;
wire n_1219;
wire n_1174;
wire n_1016;
wire n_1347;
wire n_795;
wire n_1501;
wire n_1221;
wire n_1245;
wire n_838;
wire n_647;
wire n_197;
wire n_844;
wire n_448;
wire n_1017;
wire n_1083;
wire n_445;
wire n_1561;
wire n_930;
wire n_888;
wire n_1112;
wire n_234;
wire n_910;
wire n_1656;
wire n_1460;
wire n_911;
wire n_1464;
wire n_236;
wire n_653;
wire n_1414;
wire n_752;
wire n_908;
wire n_944;
wire n_576;
wire n_1028;
wire n_472;
wire n_270;
wire n_414;
wire n_563;
wire n_1011;
wire n_1566;
wire n_1215;
wire n_839;
wire n_708;
wire n_668;
wire n_626;
wire n_990;
wire n_1500;
wire n_779;
wire n_1537;
wire n_1104;
wire n_854;
wire n_1058;
wire n_498;
wire n_1122;
wire n_870;
wire n_904;
wire n_1253;
wire n_709;
wire n_1266;
wire n_366;
wire n_1509;
wire n_1109;
wire n_185;
wire n_712;
wire n_348;
wire n_1276;
wire n_376;
wire n_390;
wire n_1148;
wire n_334;
wire n_1161;
wire n_1085;
wire n_232;
wire n_1239;
wire n_771;
wire n_1584;
wire n_470;
wire n_475;
wire n_924;
wire n_298;
wire n_1582;
wire n_492;
wire n_1149;
wire n_265;
wire n_1184;
wire n_228;
wire n_719;
wire n_1525;
wire n_455;
wire n_1585;
wire n_363;
wire n_1090;
wire n_592;
wire n_1518;
wire n_829;
wire n_1156;
wire n_1362;
wire n_393;
wire n_984;
wire n_503;
wire n_1450;
wire n_1638;
wire n_868;
wire n_570;
wire n_859;
wire n_406;
wire n_735;
wire n_878;
wire n_620;
wire n_519;
wire n_307;
wire n_469;
wire n_1218;
wire n_500;
wire n_1482;
wire n_981;
wire n_714;
wire n_1349;
wire n_291;
wire n_1144;
wire n_357;
wire n_985;
wire n_481;
wire n_997;
wire n_1301;
wire n_802;
wire n_561;
wire n_980;
wire n_1306;
wire n_1651;
wire n_1198;
wire n_1609;
wire n_436;
wire n_409;
wire n_1244;
wire n_1685;
wire n_1574;
wire n_240;
wire n_756;
wire n_1619;
wire n_1606;
wire n_810;
wire n_1133;
wire n_635;
wire n_1194;
wire n_1051;
wire n_253;
wire n_1552;
wire n_583;
wire n_249;
wire n_201;
wire n_1039;
wire n_1442;
wire n_1034;
wire n_1480;
wire n_1158;
wire n_754;
wire n_941;
wire n_975;
wire n_1031;
wire n_1305;
wire n_553;
wire n_849;
wire n_753;
wire n_467;
wire n_269;
wire n_359;
wire n_973;
wire n_1479;
wire n_1055;
wire n_1675;
wire n_582;
wire n_861;
wire n_857;
wire n_967;
wire n_571;
wire n_271;
wire n_404;
wire n_158;
wire n_206;
wire n_679;
wire n_633;
wire n_1170;
wire n_665;
wire n_1629;
wire n_588;
wire n_225;
wire n_1260;
wire n_308;
wire n_309;
wire n_1010;
wire n_1040;
wire n_915;
wire n_632;
wire n_1166;
wire n_812;
wire n_1131;
wire n_534;
wire n_1578;
wire n_1006;
wire n_373;
wire n_1632;
wire n_257;
wire n_1557;
wire n_730;
wire n_1311;
wire n_1494;
wire n_670;
wire n_203;
wire n_207;
wire n_1089;
wire n_1587;
wire n_1365;
wire n_1417;
wire n_205;
wire n_1242;
wire n_681;
wire n_1226;
wire n_1274;
wire n_1486;
wire n_412;
wire n_640;
wire n_1322;
wire n_965;
wire n_1428;
wire n_1616;
wire n_1576;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_288;
wire n_1059;
wire n_1197;
wire n_422;
wire n_722;
wire n_862;
wire n_165;
wire n_540;
wire n_1423;
wire n_457;
wire n_364;
wire n_629;
wire n_1621;
wire n_900;
wire n_1449;
wire n_531;
wire n_827;
wire n_361;
wire n_1025;
wire n_336;
wire n_1013;
wire n_1259;
wire n_192;
wire n_1538;
wire n_649;
wire n_1612;
wire n_1240;

INVx1_ASAP7_75t_L g155 ( 
.A(n_149),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_1),
.Y(n_156)
);

CKINVDCx5p33_ASAP7_75t_R g157 ( 
.A(n_14),
.Y(n_157)
);

CKINVDCx5p33_ASAP7_75t_R g158 ( 
.A(n_23),
.Y(n_158)
);

CKINVDCx5p33_ASAP7_75t_R g159 ( 
.A(n_131),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_145),
.Y(n_160)
);

CKINVDCx5p33_ASAP7_75t_R g161 ( 
.A(n_115),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_86),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_64),
.Y(n_164)
);

CKINVDCx5p33_ASAP7_75t_R g165 ( 
.A(n_24),
.Y(n_165)
);

CKINVDCx5p33_ASAP7_75t_R g166 ( 
.A(n_154),
.Y(n_166)
);

CKINVDCx5p33_ASAP7_75t_R g167 ( 
.A(n_30),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_151),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_18),
.Y(n_169)
);

CKINVDCx5p33_ASAP7_75t_R g170 ( 
.A(n_62),
.Y(n_170)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_93),
.Y(n_172)
);

CKINVDCx5p33_ASAP7_75t_R g173 ( 
.A(n_130),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_80),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_37),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_138),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_21),
.Y(n_177)
);

CKINVDCx5p33_ASAP7_75t_R g178 ( 
.A(n_32),
.Y(n_178)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_153),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_59),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_27),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_118),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_29),
.Y(n_183)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_103),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g185 ( 
.A(n_150),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_28),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_123),
.Y(n_187)
);

BUFx10_ASAP7_75t_L g188 ( 
.A(n_39),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_141),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_143),
.Y(n_190)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_6),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_55),
.Y(n_192)
);

INVx1_ASAP7_75t_SL g193 ( 
.A(n_0),
.Y(n_193)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_107),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_134),
.Y(n_195)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_137),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_23),
.Y(n_197)
);

BUFx3_ASAP7_75t_L g198 ( 
.A(n_39),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_3),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_12),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_152),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_24),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_112),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_42),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_33),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_102),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g207 ( 
.A(n_5),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_108),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_144),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_25),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_36),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_96),
.Y(n_212)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_146),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_27),
.Y(n_214)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_116),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_33),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_106),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_113),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_110),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_124),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g221 ( 
.A(n_42),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_126),
.Y(n_222)
);

INVx2_ASAP7_75t_SL g223 ( 
.A(n_117),
.Y(n_223)
);

INVx2_ASAP7_75t_SL g224 ( 
.A(n_97),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_66),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_101),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_65),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_47),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_140),
.Y(n_229)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_57),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_36),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_81),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_21),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_135),
.Y(n_234)
);

INVx2_ASAP7_75t_L g235 ( 
.A(n_90),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_20),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_92),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_73),
.Y(n_238)
);

BUFx3_ASAP7_75t_L g239 ( 
.A(n_54),
.Y(n_239)
);

CKINVDCx5p33_ASAP7_75t_R g240 ( 
.A(n_30),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_147),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_68),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_48),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_14),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_45),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_129),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_77),
.Y(n_247)
);

BUFx2_ASAP7_75t_R g248 ( 
.A(n_52),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_69),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_8),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_34),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_95),
.Y(n_252)
);

INVx3_ASAP7_75t_L g253 ( 
.A(n_0),
.Y(n_253)
);

INVx1_ASAP7_75t_SL g254 ( 
.A(n_44),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_4),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_63),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_85),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_83),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_43),
.Y(n_259)
);

BUFx3_ASAP7_75t_L g260 ( 
.A(n_26),
.Y(n_260)
);

CKINVDCx5p33_ASAP7_75t_R g261 ( 
.A(n_142),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g262 ( 
.A(n_40),
.Y(n_262)
);

CKINVDCx5p33_ASAP7_75t_R g263 ( 
.A(n_104),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_4),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_3),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_99),
.Y(n_266)
);

BUFx6f_ASAP7_75t_L g267 ( 
.A(n_17),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_31),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_37),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g270 ( 
.A(n_26),
.Y(n_270)
);

HB1xp67_ASAP7_75t_L g271 ( 
.A(n_119),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_114),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_74),
.Y(n_273)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_79),
.Y(n_274)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_139),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_17),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_18),
.Y(n_277)
);

INVx1_ASAP7_75t_SL g278 ( 
.A(n_122),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_88),
.Y(n_279)
);

CKINVDCx5p33_ASAP7_75t_R g280 ( 
.A(n_35),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_56),
.Y(n_281)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_25),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_44),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_11),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_75),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_6),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_72),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_12),
.Y(n_288)
);

CKINVDCx5p33_ASAP7_75t_R g289 ( 
.A(n_132),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_46),
.Y(n_290)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_109),
.Y(n_291)
);

CKINVDCx14_ASAP7_75t_R g292 ( 
.A(n_82),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_22),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_38),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_29),
.Y(n_295)
);

INVx1_ASAP7_75t_SL g296 ( 
.A(n_13),
.Y(n_296)
);

INVx1_ASAP7_75t_SL g297 ( 
.A(n_1),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_71),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_5),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_111),
.Y(n_300)
);

INVx1_ASAP7_75t_SL g301 ( 
.A(n_32),
.Y(n_301)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_8),
.Y(n_302)
);

BUFx10_ASAP7_75t_L g303 ( 
.A(n_22),
.Y(n_303)
);

BUFx8_ASAP7_75t_SL g304 ( 
.A(n_133),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_2),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_43),
.Y(n_306)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_10),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_51),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_267),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_267),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_304),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_189),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_267),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_172),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_267),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_267),
.Y(n_316)
);

CKINVDCx5p33_ASAP7_75t_R g317 ( 
.A(n_190),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_307),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_307),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_271),
.B(n_2),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_223),
.B(n_7),
.Y(n_321)
);

BUFx3_ASAP7_75t_L g322 ( 
.A(n_239),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g323 ( 
.A(n_176),
.Y(n_323)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_307),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_262),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_307),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g327 ( 
.A(n_222),
.Y(n_327)
);

CKINVDCx5p33_ASAP7_75t_R g328 ( 
.A(n_192),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_253),
.Y(n_330)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_198),
.B(n_7),
.Y(n_331)
);

CKINVDCx5p33_ASAP7_75t_R g332 ( 
.A(n_195),
.Y(n_332)
);

BUFx3_ASAP7_75t_L g333 ( 
.A(n_239),
.Y(n_333)
);

INVxp67_ASAP7_75t_SL g334 ( 
.A(n_253),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_253),
.Y(n_335)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_245),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_210),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g338 ( 
.A(n_230),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_210),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_282),
.Y(n_340)
);

BUFx6f_ASAP7_75t_SL g341 ( 
.A(n_186),
.Y(n_341)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_282),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_198),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_201),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_223),
.B(n_9),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_203),
.Y(n_346)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_260),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_206),
.Y(n_348)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_260),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_208),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_156),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_175),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_209),
.Y(n_353)
);

INVxp33_ASAP7_75t_L g354 ( 
.A(n_191),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_212),
.Y(n_355)
);

NOR2xp67_ASAP7_75t_L g356 ( 
.A(n_199),
.B(n_9),
.Y(n_356)
);

CKINVDCx5p33_ASAP7_75t_R g357 ( 
.A(n_219),
.Y(n_357)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_214),
.Y(n_358)
);

OR2x2_ASAP7_75t_L g359 ( 
.A(n_216),
.B(n_10),
.Y(n_359)
);

HB1xp67_ASAP7_75t_L g360 ( 
.A(n_207),
.Y(n_360)
);

CKINVDCx20_ASAP7_75t_R g361 ( 
.A(n_274),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_236),
.Y(n_362)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_251),
.Y(n_363)
);

NOR2xp67_ASAP7_75t_L g364 ( 
.A(n_276),
.B(n_11),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_220),
.Y(n_365)
);

NAND2xp33_ASAP7_75t_R g366 ( 
.A(n_159),
.B(n_13),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_292),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_226),
.Y(n_368)
);

CKINVDCx20_ASAP7_75t_R g369 ( 
.A(n_232),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_234),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_284),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_237),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_290),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_238),
.Y(n_374)
);

HB1xp67_ASAP7_75t_L g375 ( 
.A(n_221),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_241),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_295),
.Y(n_377)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_302),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_242),
.Y(n_379)
);

BUFx6f_ASAP7_75t_L g380 ( 
.A(n_309),
.Y(n_380)
);

AND2x2_ASAP7_75t_SL g381 ( 
.A(n_331),
.B(n_160),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_334),
.B(n_224),
.Y(n_382)
);

INVx1_ASAP7_75t_L g383 ( 
.A(n_309),
.Y(n_383)
);

BUFx6f_ASAP7_75t_L g384 ( 
.A(n_310),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g385 ( 
.A(n_321),
.B(n_224),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_345),
.B(n_300),
.Y(n_386)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_310),
.Y(n_387)
);

INVx2_ASAP7_75t_L g388 ( 
.A(n_313),
.Y(n_388)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_313),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_315),
.Y(n_390)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_315),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_316),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g393 ( 
.A(n_316),
.B(n_300),
.Y(n_393)
);

AND2x4_ASAP7_75t_L g394 ( 
.A(n_330),
.B(n_160),
.Y(n_394)
);

BUFx6f_ASAP7_75t_L g395 ( 
.A(n_318),
.Y(n_395)
);

INVx3_ASAP7_75t_L g396 ( 
.A(n_318),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_319),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_319),
.Y(n_398)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_331),
.B(n_179),
.Y(n_399)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_324),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_324),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g402 ( 
.A1(n_314),
.A2(n_269),
.B1(n_183),
.B2(n_202),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_326),
.Y(n_403)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_326),
.Y(n_404)
);

CKINVDCx5p33_ASAP7_75t_R g405 ( 
.A(n_368),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_329),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_329),
.Y(n_407)
);

AND2x2_ASAP7_75t_L g408 ( 
.A(n_330),
.B(n_179),
.Y(n_408)
);

OA21x2_ASAP7_75t_L g409 ( 
.A1(n_335),
.A2(n_305),
.B(n_235),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_335),
.Y(n_410)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_322),
.Y(n_411)
);

INVx1_ASAP7_75t_L g412 ( 
.A(n_351),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_351),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_337),
.Y(n_414)
);

AND2x4_ASAP7_75t_L g415 ( 
.A(n_356),
.B(n_235),
.Y(n_415)
);

BUFx6f_ASAP7_75t_L g416 ( 
.A(n_337),
.Y(n_416)
);

INVx2_ASAP7_75t_L g417 ( 
.A(n_339),
.Y(n_417)
);

NAND2xp5_ASAP7_75t_L g418 ( 
.A(n_322),
.B(n_159),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_333),
.B(n_161),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_352),
.Y(n_420)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_352),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_339),
.Y(n_422)
);

BUFx6f_ASAP7_75t_L g423 ( 
.A(n_340),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_340),
.Y(n_424)
);

NAND2xp33_ASAP7_75t_SL g425 ( 
.A(n_359),
.B(n_157),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_358),
.Y(n_426)
);

BUFx6f_ASAP7_75t_L g427 ( 
.A(n_342),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_342),
.Y(n_428)
);

NAND2xp33_ASAP7_75t_R g429 ( 
.A(n_311),
.B(n_157),
.Y(n_429)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_358),
.Y(n_430)
);

INVx3_ASAP7_75t_L g431 ( 
.A(n_362),
.Y(n_431)
);

BUFx3_ASAP7_75t_L g432 ( 
.A(n_333),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_362),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_363),
.Y(n_434)
);

HB1xp67_ASAP7_75t_L g435 ( 
.A(n_360),
.Y(n_435)
);

INVx2_ASAP7_75t_L g436 ( 
.A(n_363),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_371),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_364),
.B(n_162),
.Y(n_438)
);

BUFx6f_ASAP7_75t_L g439 ( 
.A(n_371),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_373),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_373),
.Y(n_441)
);

INVx2_ASAP7_75t_L g442 ( 
.A(n_377),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_343),
.B(n_161),
.Y(n_443)
);

INVx3_ASAP7_75t_L g444 ( 
.A(n_377),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_SL g445 ( 
.A(n_381),
.B(n_312),
.Y(n_445)
);

OAI22xp33_ASAP7_75t_L g446 ( 
.A1(n_385),
.A2(n_366),
.B1(n_254),
.B2(n_296),
.Y(n_446)
);

INVx2_ASAP7_75t_L g447 ( 
.A(n_388),
.Y(n_447)
);

BUFx3_ASAP7_75t_L g448 ( 
.A(n_432),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_408),
.B(n_343),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_409),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_381),
.B(n_317),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_409),
.Y(n_452)
);

AOI22xp33_ASAP7_75t_L g453 ( 
.A1(n_381),
.A2(n_320),
.B1(n_325),
.B2(n_359),
.Y(n_453)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_409),
.Y(n_454)
);

NAND2xp5_ASAP7_75t_L g455 ( 
.A(n_399),
.B(n_328),
.Y(n_455)
);

NAND2xp5_ASAP7_75t_SL g456 ( 
.A(n_418),
.B(n_332),
.Y(n_456)
);

NAND2xp33_ASAP7_75t_R g457 ( 
.A(n_405),
.B(n_385),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_409),
.Y(n_458)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_408),
.B(n_347),
.Y(n_459)
);

AND2x2_ASAP7_75t_L g460 ( 
.A(n_408),
.B(n_347),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_409),
.Y(n_461)
);

AOI22xp5_ASAP7_75t_L g462 ( 
.A1(n_425),
.A2(n_297),
.B1(n_301),
.B2(n_193),
.Y(n_462)
);

NOR3xp33_ASAP7_75t_L g463 ( 
.A(n_402),
.B(n_336),
.C(n_375),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_388),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g465 ( 
.A(n_432),
.Y(n_465)
);

NOR2x1p5_ASAP7_75t_L g466 ( 
.A(n_386),
.B(n_158),
.Y(n_466)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_409),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_405),
.B(n_248),
.Y(n_468)
);

INVx4_ASAP7_75t_L g469 ( 
.A(n_380),
.Y(n_469)
);

AOI22xp33_ASAP7_75t_L g470 ( 
.A1(n_386),
.A2(n_354),
.B1(n_162),
.B2(n_349),
.Y(n_470)
);

AO21x2_ASAP7_75t_L g471 ( 
.A1(n_382),
.A2(n_164),
.B(n_155),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_418),
.B(n_344),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g473 ( 
.A(n_419),
.B(n_346),
.Y(n_473)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_411),
.B(n_348),
.Y(n_474)
);

INVxp67_ASAP7_75t_SL g475 ( 
.A(n_432),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_388),
.Y(n_476)
);

AOI22xp33_ASAP7_75t_L g477 ( 
.A1(n_399),
.A2(n_162),
.B1(n_349),
.B2(n_378),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_389),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_388),
.Y(n_479)
);

OR2x2_ASAP7_75t_L g480 ( 
.A(n_419),
.B(n_350),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_398),
.Y(n_481)
);

INVx4_ASAP7_75t_L g482 ( 
.A(n_380),
.Y(n_482)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_389),
.Y(n_483)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_380),
.Y(n_484)
);

INVx3_ASAP7_75t_L g485 ( 
.A(n_380),
.Y(n_485)
);

NOR2xp33_ASAP7_75t_L g486 ( 
.A(n_411),
.B(n_353),
.Y(n_486)
);

CKINVDCx5p33_ASAP7_75t_R g487 ( 
.A(n_429),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_399),
.B(n_378),
.Y(n_488)
);

CKINVDCx5p33_ASAP7_75t_R g489 ( 
.A(n_429),
.Y(n_489)
);

INVx2_ASAP7_75t_L g490 ( 
.A(n_398),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_L g491 ( 
.A(n_411),
.B(n_355),
.Y(n_491)
);

BUFx10_ASAP7_75t_L g492 ( 
.A(n_435),
.Y(n_492)
);

AOI22xp33_ASAP7_75t_L g493 ( 
.A1(n_415),
.A2(n_425),
.B1(n_382),
.B2(n_438),
.Y(n_493)
);

BUFx4f_ASAP7_75t_L g494 ( 
.A(n_380),
.Y(n_494)
);

NAND2xp33_ASAP7_75t_L g495 ( 
.A(n_443),
.B(n_357),
.Y(n_495)
);

INVx1_ASAP7_75t_L g496 ( 
.A(n_389),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_L g497 ( 
.A(n_411),
.B(n_365),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_383),
.Y(n_498)
);

INVx2_ASAP7_75t_L g499 ( 
.A(n_398),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_383),
.Y(n_500)
);

INVx3_ASAP7_75t_L g501 ( 
.A(n_380),
.Y(n_501)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_439),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_411),
.B(n_370),
.Y(n_503)
);

INVx2_ASAP7_75t_L g504 ( 
.A(n_398),
.Y(n_504)
);

INVx2_ASAP7_75t_L g505 ( 
.A(n_404),
.Y(n_505)
);

INVx4_ASAP7_75t_L g506 ( 
.A(n_380),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_432),
.B(n_372),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_387),
.Y(n_508)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_387),
.Y(n_509)
);

OR2x2_ASAP7_75t_L g510 ( 
.A(n_435),
.B(n_374),
.Y(n_510)
);

INVx2_ASAP7_75t_L g511 ( 
.A(n_404),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_404),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_415),
.A2(n_165),
.B1(n_158),
.B2(n_167),
.Y(n_513)
);

AND2x2_ASAP7_75t_L g514 ( 
.A(n_410),
.B(n_376),
.Y(n_514)
);

BUFx4f_ASAP7_75t_L g515 ( 
.A(n_380),
.Y(n_515)
);

OR2x6_ASAP7_75t_L g516 ( 
.A(n_443),
.B(n_171),
.Y(n_516)
);

NAND2xp33_ASAP7_75t_L g517 ( 
.A(n_439),
.B(n_379),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_431),
.B(n_369),
.Y(n_518)
);

INVx3_ASAP7_75t_L g519 ( 
.A(n_384),
.Y(n_519)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_431),
.Y(n_520)
);

NOR2x1p5_ASAP7_75t_L g521 ( 
.A(n_412),
.B(n_165),
.Y(n_521)
);

INVx1_ASAP7_75t_L g522 ( 
.A(n_431),
.Y(n_522)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_431),
.B(n_367),
.Y(n_523)
);

INVx5_ASAP7_75t_L g524 ( 
.A(n_384),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_431),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_438),
.B(n_217),
.Y(n_526)
);

AND2x4_ASAP7_75t_L g527 ( 
.A(n_394),
.B(n_184),
.Y(n_527)
);

NAND2xp33_ASAP7_75t_L g528 ( 
.A(n_439),
.B(n_162),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_404),
.Y(n_529)
);

INVx2_ASAP7_75t_L g530 ( 
.A(n_406),
.Y(n_530)
);

NAND2xp5_ASAP7_75t_L g531 ( 
.A(n_438),
.B(n_278),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_SL g532 ( 
.A(n_415),
.B(n_338),
.Y(n_532)
);

AOI22x1_ASAP7_75t_L g533 ( 
.A1(n_415),
.A2(n_167),
.B1(n_169),
.B2(n_177),
.Y(n_533)
);

AOI22xp33_ASAP7_75t_L g534 ( 
.A1(n_415),
.A2(n_162),
.B1(n_227),
.B2(n_247),
.Y(n_534)
);

INVx4_ASAP7_75t_L g535 ( 
.A(n_384),
.Y(n_535)
);

INVx4_ASAP7_75t_L g536 ( 
.A(n_384),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_444),
.Y(n_537)
);

AOI22xp33_ASAP7_75t_L g538 ( 
.A1(n_415),
.A2(n_196),
.B1(n_258),
.B2(n_273),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g539 ( 
.A(n_438),
.B(n_361),
.Y(n_539)
);

BUFx6f_ASAP7_75t_L g540 ( 
.A(n_439),
.Y(n_540)
);

BUFx3_ASAP7_75t_L g541 ( 
.A(n_438),
.Y(n_541)
);

INVx3_ASAP7_75t_L g542 ( 
.A(n_384),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_406),
.Y(n_543)
);

AND2x2_ASAP7_75t_SL g544 ( 
.A(n_438),
.B(n_194),
.Y(n_544)
);

CKINVDCx20_ASAP7_75t_R g545 ( 
.A(n_402),
.Y(n_545)
);

INVx3_ASAP7_75t_L g546 ( 
.A(n_384),
.Y(n_546)
);

BUFx10_ASAP7_75t_L g547 ( 
.A(n_394),
.Y(n_547)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_410),
.B(n_213),
.Y(n_548)
);

AND2x2_ASAP7_75t_L g549 ( 
.A(n_410),
.B(n_215),
.Y(n_549)
);

BUFx8_ASAP7_75t_SL g550 ( 
.A(n_394),
.Y(n_550)
);

INVxp67_ASAP7_75t_SL g551 ( 
.A(n_393),
.Y(n_551)
);

INVx3_ASAP7_75t_L g552 ( 
.A(n_384),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_L g553 ( 
.A(n_390),
.B(n_246),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g554 ( 
.A(n_412),
.B(n_323),
.Y(n_554)
);

BUFx3_ASAP7_75t_L g555 ( 
.A(n_444),
.Y(n_555)
);

AND2x2_ASAP7_75t_L g556 ( 
.A(n_422),
.B(n_218),
.Y(n_556)
);

INVx3_ASAP7_75t_L g557 ( 
.A(n_384),
.Y(n_557)
);

BUFx6f_ASAP7_75t_L g558 ( 
.A(n_439),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_406),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_390),
.B(n_249),
.Y(n_560)
);

AOI22xp33_ASAP7_75t_L g561 ( 
.A1(n_394),
.A2(n_291),
.B1(n_281),
.B2(n_257),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_390),
.B(n_391),
.Y(n_562)
);

INVx1_ASAP7_75t_L g563 ( 
.A(n_444),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_444),
.Y(n_564)
);

INVx1_ASAP7_75t_L g565 ( 
.A(n_444),
.Y(n_565)
);

INVx2_ASAP7_75t_SL g566 ( 
.A(n_394),
.Y(n_566)
);

INVx3_ASAP7_75t_L g567 ( 
.A(n_395),
.Y(n_567)
);

INVx1_ASAP7_75t_L g568 ( 
.A(n_391),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_406),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_394),
.A2(n_433),
.B1(n_434),
.B2(n_442),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_SL g571 ( 
.A(n_439),
.B(n_163),
.Y(n_571)
);

BUFx3_ASAP7_75t_L g572 ( 
.A(n_391),
.Y(n_572)
);

INVx3_ASAP7_75t_L g573 ( 
.A(n_395),
.Y(n_573)
);

AOI22xp33_ASAP7_75t_L g574 ( 
.A1(n_433),
.A2(n_229),
.B1(n_225),
.B2(n_185),
.Y(n_574)
);

BUFx3_ASAP7_75t_L g575 ( 
.A(n_392),
.Y(n_575)
);

AOI22xp33_ASAP7_75t_L g576 ( 
.A1(n_433),
.A2(n_185),
.B1(n_341),
.B2(n_186),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_SL g577 ( 
.A(n_439),
.B(n_163),
.Y(n_577)
);

NOR2xp33_ASAP7_75t_L g578 ( 
.A(n_413),
.B(n_341),
.Y(n_578)
);

NAND2xp5_ASAP7_75t_L g579 ( 
.A(n_392),
.B(n_252),
.Y(n_579)
);

AO22x2_ASAP7_75t_L g580 ( 
.A1(n_393),
.A2(n_186),
.B1(n_188),
.B2(n_303),
.Y(n_580)
);

HB1xp67_ASAP7_75t_L g581 ( 
.A(n_413),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_420),
.Y(n_582)
);

AOI22xp33_ASAP7_75t_L g583 ( 
.A1(n_434),
.A2(n_185),
.B1(n_341),
.B2(n_188),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_392),
.Y(n_584)
);

INVx2_ASAP7_75t_L g585 ( 
.A(n_396),
.Y(n_585)
);

AND2x4_ASAP7_75t_L g586 ( 
.A(n_434),
.B(n_420),
.Y(n_586)
);

INVx3_ASAP7_75t_L g587 ( 
.A(n_395),
.Y(n_587)
);

INVx2_ASAP7_75t_L g588 ( 
.A(n_397),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_397),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_439),
.B(n_166),
.Y(n_590)
);

NOR2xp33_ASAP7_75t_SL g591 ( 
.A(n_487),
.B(n_327),
.Y(n_591)
);

INVx1_ASAP7_75t_L g592 ( 
.A(n_581),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_551),
.B(n_397),
.Y(n_593)
);

NAND2xp5_ASAP7_75t_SL g594 ( 
.A(n_518),
.B(n_166),
.Y(n_594)
);

AND2x6_ASAP7_75t_SL g595 ( 
.A(n_523),
.B(n_421),
.Y(n_595)
);

INVx1_ASAP7_75t_L g596 ( 
.A(n_586),
.Y(n_596)
);

NOR2xp33_ASAP7_75t_L g597 ( 
.A(n_455),
.B(n_168),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_493),
.B(n_400),
.Y(n_598)
);

INVx2_ASAP7_75t_L g599 ( 
.A(n_588),
.Y(n_599)
);

OAI22xp5_ASAP7_75t_L g600 ( 
.A1(n_544),
.A2(n_285),
.B1(n_170),
.B2(n_173),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_480),
.B(n_168),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_582),
.B(n_400),
.Y(n_602)
);

NAND2xp5_ASAP7_75t_L g603 ( 
.A(n_582),
.B(n_400),
.Y(n_603)
);

NAND2xp5_ASAP7_75t_L g604 ( 
.A(n_544),
.B(n_401),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_588),
.Y(n_605)
);

AOI22xp33_ASAP7_75t_L g606 ( 
.A1(n_544),
.A2(n_185),
.B1(n_441),
.B2(n_440),
.Y(n_606)
);

NOR3xp33_ASAP7_75t_L g607 ( 
.A(n_532),
.B(n_421),
.C(n_441),
.Y(n_607)
);

NAND2xp5_ASAP7_75t_L g608 ( 
.A(n_586),
.B(n_401),
.Y(n_608)
);

INVxp67_ASAP7_75t_L g609 ( 
.A(n_457),
.Y(n_609)
);

NAND3xp33_ASAP7_75t_L g610 ( 
.A(n_453),
.B(n_205),
.C(n_197),
.Y(n_610)
);

NAND2xp5_ASAP7_75t_L g611 ( 
.A(n_586),
.B(n_401),
.Y(n_611)
);

NAND2xp5_ASAP7_75t_L g612 ( 
.A(n_586),
.B(n_403),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_526),
.B(n_403),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_SL g614 ( 
.A(n_480),
.B(n_514),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_531),
.B(n_514),
.Y(n_615)
);

NOR2xp67_ASAP7_75t_L g616 ( 
.A(n_489),
.B(n_510),
.Y(n_616)
);

NAND2xp5_ASAP7_75t_L g617 ( 
.A(n_566),
.B(n_465),
.Y(n_617)
);

INVx1_ASAP7_75t_L g618 ( 
.A(n_478),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_L g619 ( 
.A(n_566),
.B(n_403),
.Y(n_619)
);

NAND2xp5_ASAP7_75t_L g620 ( 
.A(n_465),
.B(n_407),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_SL g621 ( 
.A(n_445),
.B(n_451),
.Y(n_621)
);

NOR2xp33_ASAP7_75t_L g622 ( 
.A(n_446),
.B(n_170),
.Y(n_622)
);

NAND2xp5_ASAP7_75t_L g623 ( 
.A(n_488),
.B(n_407),
.Y(n_623)
);

INVx2_ASAP7_75t_L g624 ( 
.A(n_568),
.Y(n_624)
);

INVx2_ASAP7_75t_L g625 ( 
.A(n_568),
.Y(n_625)
);

AND2x4_ASAP7_75t_L g626 ( 
.A(n_448),
.B(n_426),
.Y(n_626)
);

BUFx3_ASAP7_75t_L g627 ( 
.A(n_448),
.Y(n_627)
);

INVx2_ASAP7_75t_L g628 ( 
.A(n_584),
.Y(n_628)
);

NAND2xp5_ASAP7_75t_L g629 ( 
.A(n_488),
.B(n_396),
.Y(n_629)
);

NOR2xp67_ASAP7_75t_L g630 ( 
.A(n_510),
.B(n_426),
.Y(n_630)
);

NAND2xp5_ASAP7_75t_SL g631 ( 
.A(n_554),
.B(n_173),
.Y(n_631)
);

NAND2xp5_ASAP7_75t_L g632 ( 
.A(n_572),
.B(n_575),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_L g633 ( 
.A(n_572),
.B(n_396),
.Y(n_633)
);

OAI221xp5_ASAP7_75t_L g634 ( 
.A1(n_470),
.A2(n_513),
.B1(n_462),
.B2(n_533),
.C(n_538),
.Y(n_634)
);

AOI221xp5_ASAP7_75t_L g635 ( 
.A1(n_462),
.A2(n_181),
.B1(n_178),
.B2(n_177),
.C(n_169),
.Y(n_635)
);

BUFx6f_ASAP7_75t_L g636 ( 
.A(n_541),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_483),
.Y(n_637)
);

INVx1_ASAP7_75t_L g638 ( 
.A(n_483),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_L g639 ( 
.A(n_572),
.B(n_396),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_496),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_SL g641 ( 
.A(n_507),
.B(n_174),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_575),
.B(n_396),
.Y(n_642)
);

AO221x1_ASAP7_75t_L g643 ( 
.A1(n_580),
.A2(n_440),
.B1(n_422),
.B2(n_428),
.C(n_303),
.Y(n_643)
);

INVx1_ASAP7_75t_L g644 ( 
.A(n_496),
.Y(n_644)
);

INVx2_ASAP7_75t_SL g645 ( 
.A(n_492),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_L g646 ( 
.A(n_575),
.B(n_430),
.Y(n_646)
);

NOR2x1p5_ASAP7_75t_L g647 ( 
.A(n_491),
.B(n_178),
.Y(n_647)
);

AND2x2_ASAP7_75t_L g648 ( 
.A(n_449),
.B(n_188),
.Y(n_648)
);

NOR2xp33_ASAP7_75t_L g649 ( 
.A(n_456),
.B(n_174),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_SL g650 ( 
.A(n_474),
.B(n_180),
.Y(n_650)
);

INVx2_ASAP7_75t_L g651 ( 
.A(n_584),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_L g652 ( 
.A(n_450),
.B(n_430),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_449),
.B(n_303),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_498),
.Y(n_654)
);

NOR2xp33_ASAP7_75t_L g655 ( 
.A(n_472),
.B(n_180),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_450),
.B(n_436),
.Y(n_656)
);

AOI22xp33_ASAP7_75t_L g657 ( 
.A1(n_452),
.A2(n_185),
.B1(n_422),
.B2(n_428),
.Y(n_657)
);

NAND2xp5_ASAP7_75t_SL g658 ( 
.A(n_486),
.B(n_182),
.Y(n_658)
);

AOI22xp33_ASAP7_75t_L g659 ( 
.A1(n_452),
.A2(n_185),
.B1(n_428),
.B2(n_181),
.Y(n_659)
);

NOR2xp33_ASAP7_75t_L g660 ( 
.A(n_473),
.B(n_182),
.Y(n_660)
);

NOR2xp33_ASAP7_75t_L g661 ( 
.A(n_516),
.B(n_187),
.Y(n_661)
);

INVx2_ASAP7_75t_L g662 ( 
.A(n_589),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_498),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_454),
.B(n_436),
.Y(n_664)
);

NAND2xp5_ASAP7_75t_L g665 ( 
.A(n_454),
.B(n_458),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_L g666 ( 
.A(n_458),
.B(n_436),
.Y(n_666)
);

NAND2xp5_ASAP7_75t_L g667 ( 
.A(n_461),
.B(n_436),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_516),
.B(n_187),
.Y(n_668)
);

INVx2_ASAP7_75t_L g669 ( 
.A(n_589),
.Y(n_669)
);

NOR2xp33_ASAP7_75t_L g670 ( 
.A(n_516),
.B(n_279),
.Y(n_670)
);

NOR2xp33_ASAP7_75t_L g671 ( 
.A(n_516),
.B(n_279),
.Y(n_671)
);

INVx1_ASAP7_75t_L g672 ( 
.A(n_500),
.Y(n_672)
);

INVx1_ASAP7_75t_L g673 ( 
.A(n_500),
.Y(n_673)
);

BUFx6f_ASAP7_75t_SL g674 ( 
.A(n_492),
.Y(n_674)
);

A2O1A1Ixp33_ASAP7_75t_L g675 ( 
.A1(n_461),
.A2(n_442),
.B(n_437),
.C(n_424),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_508),
.Y(n_676)
);

OR2x6_ASAP7_75t_L g677 ( 
.A(n_539),
.B(n_437),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_467),
.B(n_437),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_467),
.B(n_437),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_L g680 ( 
.A(n_541),
.B(n_442),
.Y(n_680)
);

INVx1_ASAP7_75t_L g681 ( 
.A(n_508),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_541),
.B(n_442),
.Y(n_682)
);

INVx8_ASAP7_75t_L g683 ( 
.A(n_550),
.Y(n_683)
);

NAND2xp5_ASAP7_75t_SL g684 ( 
.A(n_503),
.B(n_285),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_492),
.Y(n_685)
);

NAND2xp5_ASAP7_75t_SL g686 ( 
.A(n_576),
.B(n_287),
.Y(n_686)
);

INVx2_ASAP7_75t_L g687 ( 
.A(n_509),
.Y(n_687)
);

INVx1_ASAP7_75t_L g688 ( 
.A(n_509),
.Y(n_688)
);

INVx1_ASAP7_75t_L g689 ( 
.A(n_459),
.Y(n_689)
);

INVx1_ASAP7_75t_L g690 ( 
.A(n_459),
.Y(n_690)
);

INVxp67_ASAP7_75t_L g691 ( 
.A(n_468),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_583),
.B(n_287),
.Y(n_692)
);

INVx1_ASAP7_75t_L g693 ( 
.A(n_460),
.Y(n_693)
);

AND2x4_ASAP7_75t_L g694 ( 
.A(n_460),
.B(n_414),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_520),
.Y(n_695)
);

A2O1A1Ixp33_ASAP7_75t_L g696 ( 
.A1(n_520),
.A2(n_414),
.B(n_424),
.C(n_417),
.Y(n_696)
);

INVx1_ASAP7_75t_L g697 ( 
.A(n_522),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_SL g698 ( 
.A(n_513),
.B(n_289),
.Y(n_698)
);

INVx1_ASAP7_75t_L g699 ( 
.A(n_522),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_SL g700 ( 
.A(n_578),
.B(n_289),
.Y(n_700)
);

NOR3xp33_ASAP7_75t_L g701 ( 
.A(n_463),
.B(n_264),
.C(n_259),
.Y(n_701)
);

INVx2_ASAP7_75t_L g702 ( 
.A(n_464),
.Y(n_702)
);

NAND2xp5_ASAP7_75t_SL g703 ( 
.A(n_497),
.B(n_298),
.Y(n_703)
);

NAND2xp5_ASAP7_75t_L g704 ( 
.A(n_475),
.B(n_416),
.Y(n_704)
);

INVx2_ASAP7_75t_L g705 ( 
.A(n_464),
.Y(n_705)
);

NAND2xp5_ASAP7_75t_SL g706 ( 
.A(n_555),
.B(n_185),
.Y(n_706)
);

NOR2xp33_ASAP7_75t_L g707 ( 
.A(n_516),
.B(n_298),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_533),
.B(n_256),
.Y(n_708)
);

INVx2_ASAP7_75t_SL g709 ( 
.A(n_521),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_555),
.B(n_525),
.Y(n_710)
);

NAND2xp5_ASAP7_75t_L g711 ( 
.A(n_555),
.B(n_416),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_525),
.B(n_416),
.Y(n_712)
);

NAND2xp33_ASAP7_75t_L g713 ( 
.A(n_466),
.B(n_521),
.Y(n_713)
);

NAND2xp5_ASAP7_75t_SL g714 ( 
.A(n_477),
.B(n_261),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_495),
.B(n_200),
.Y(n_715)
);

NAND2xp5_ASAP7_75t_L g716 ( 
.A(n_537),
.B(n_416),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_SL g717 ( 
.A(n_547),
.B(n_263),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_537),
.Y(n_718)
);

INVx2_ASAP7_75t_L g719 ( 
.A(n_464),
.Y(n_719)
);

AND2x2_ASAP7_75t_SL g720 ( 
.A(n_534),
.B(n_416),
.Y(n_720)
);

NAND2xp5_ASAP7_75t_SL g721 ( 
.A(n_547),
.B(n_266),
.Y(n_721)
);

AND2x2_ASAP7_75t_L g722 ( 
.A(n_466),
.B(n_204),
.Y(n_722)
);

AOI22xp33_ASAP7_75t_L g723 ( 
.A1(n_471),
.A2(n_185),
.B1(n_277),
.B2(n_283),
.Y(n_723)
);

NOR3xp33_ASAP7_75t_L g724 ( 
.A(n_553),
.B(n_243),
.C(n_240),
.Y(n_724)
);

AOI22xp33_ASAP7_75t_L g725 ( 
.A1(n_471),
.A2(n_283),
.B1(n_231),
.B2(n_277),
.Y(n_725)
);

INVxp67_ASAP7_75t_L g726 ( 
.A(n_580),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_563),
.B(n_416),
.Y(n_727)
);

NOR2xp33_ASAP7_75t_L g728 ( 
.A(n_560),
.B(n_211),
.Y(n_728)
);

OAI22xp5_ASAP7_75t_L g729 ( 
.A1(n_570),
.A2(n_275),
.B1(n_272),
.B2(n_244),
.Y(n_729)
);

INVxp67_ASAP7_75t_L g730 ( 
.A(n_580),
.Y(n_730)
);

NAND2xp33_ASAP7_75t_L g731 ( 
.A(n_563),
.B(n_228),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_481),
.Y(n_732)
);

NAND2xp5_ASAP7_75t_SL g733 ( 
.A(n_547),
.B(n_233),
.Y(n_733)
);

NAND2xp5_ASAP7_75t_SL g734 ( 
.A(n_547),
.B(n_250),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_564),
.Y(n_735)
);

O2A1O1Ixp33_ASAP7_75t_L g736 ( 
.A1(n_571),
.A2(n_424),
.B(n_417),
.C(n_414),
.Y(n_736)
);

INVxp67_ASAP7_75t_SL g737 ( 
.A(n_502),
.Y(n_737)
);

NAND2xp5_ASAP7_75t_SL g738 ( 
.A(n_564),
.B(n_427),
.Y(n_738)
);

BUFx6f_ASAP7_75t_L g739 ( 
.A(n_502),
.Y(n_739)
);

INVxp33_ASAP7_75t_L g740 ( 
.A(n_580),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_565),
.Y(n_741)
);

NOR2xp33_ASAP7_75t_L g742 ( 
.A(n_579),
.B(n_308),
.Y(n_742)
);

INVx1_ASAP7_75t_L g743 ( 
.A(n_565),
.Y(n_743)
);

AOI22xp33_ASAP7_75t_L g744 ( 
.A1(n_471),
.A2(n_294),
.B1(n_280),
.B2(n_286),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_527),
.B(n_423),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_481),
.Y(n_746)
);

OR2x2_ASAP7_75t_L g747 ( 
.A(n_527),
.B(n_231),
.Y(n_747)
);

CKINVDCx5p33_ASAP7_75t_R g748 ( 
.A(n_545),
.Y(n_748)
);

BUFx5_ASAP7_75t_L g749 ( 
.A(n_527),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_562),
.Y(n_750)
);

AOI22xp5_ASAP7_75t_L g751 ( 
.A1(n_527),
.A2(n_424),
.B1(n_417),
.B2(n_414),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_585),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_548),
.B(n_427),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_SL g754 ( 
.A(n_548),
.B(n_255),
.Y(n_754)
);

BUFx6f_ASAP7_75t_SL g755 ( 
.A(n_502),
.Y(n_755)
);

NOR2xp33_ASAP7_75t_L g756 ( 
.A(n_549),
.B(n_265),
.Y(n_756)
);

AOI21xp5_ASAP7_75t_L g757 ( 
.A1(n_617),
.A2(n_515),
.B(n_494),
.Y(n_757)
);

INVx2_ASAP7_75t_L g758 ( 
.A(n_624),
.Y(n_758)
);

NAND2xp5_ASAP7_75t_L g759 ( 
.A(n_750),
.B(n_549),
.Y(n_759)
);

NAND2xp33_ASAP7_75t_L g760 ( 
.A(n_749),
.B(n_556),
.Y(n_760)
);

NAND2xp5_ASAP7_75t_L g761 ( 
.A(n_615),
.B(n_556),
.Y(n_761)
);

AOI21xp5_ASAP7_75t_L g762 ( 
.A1(n_665),
.A2(n_515),
.B(n_494),
.Y(n_762)
);

OAI22xp5_ASAP7_75t_L g763 ( 
.A1(n_598),
.A2(n_561),
.B1(n_574),
.B2(n_585),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_597),
.B(n_517),
.Y(n_764)
);

NAND2xp5_ASAP7_75t_L g765 ( 
.A(n_597),
.B(n_585),
.Y(n_765)
);

AOI21xp5_ASAP7_75t_L g766 ( 
.A1(n_737),
.A2(n_515),
.B(n_494),
.Y(n_766)
);

AOI21xp5_ASAP7_75t_L g767 ( 
.A1(n_652),
.A2(n_515),
.B(n_494),
.Y(n_767)
);

AOI21xp5_ASAP7_75t_L g768 ( 
.A1(n_656),
.A2(n_469),
.B(n_536),
.Y(n_768)
);

O2A1O1Ixp33_ASAP7_75t_L g769 ( 
.A1(n_634),
.A2(n_590),
.B(n_577),
.C(n_528),
.Y(n_769)
);

INVx1_ASAP7_75t_L g770 ( 
.A(n_625),
.Y(n_770)
);

AOI21xp5_ASAP7_75t_L g771 ( 
.A1(n_664),
.A2(n_469),
.B(n_536),
.Y(n_771)
);

HB1xp67_ASAP7_75t_L g772 ( 
.A(n_592),
.Y(n_772)
);

AOI21xp5_ASAP7_75t_L g773 ( 
.A1(n_666),
.A2(n_678),
.B(n_667),
.Y(n_773)
);

AOI21xp5_ASAP7_75t_L g774 ( 
.A1(n_679),
.A2(n_469),
.B(n_536),
.Y(n_774)
);

AOI21xp5_ASAP7_75t_L g775 ( 
.A1(n_704),
.A2(n_469),
.B(n_536),
.Y(n_775)
);

INVx2_ASAP7_75t_L g776 ( 
.A(n_625),
.Y(n_776)
);

NAND2xp5_ASAP7_75t_L g777 ( 
.A(n_728),
.B(n_484),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_728),
.B(n_484),
.Y(n_778)
);

OAI21xp5_ASAP7_75t_L g779 ( 
.A1(n_604),
.A2(n_511),
.B(n_505),
.Y(n_779)
);

NAND2xp5_ASAP7_75t_L g780 ( 
.A(n_742),
.B(n_484),
.Y(n_780)
);

INVx2_ASAP7_75t_L g781 ( 
.A(n_628),
.Y(n_781)
);

A2O1A1Ixp33_ASAP7_75t_L g782 ( 
.A1(n_622),
.A2(n_286),
.B(n_280),
.C(n_288),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_742),
.B(n_484),
.Y(n_783)
);

A2O1A1Ixp33_ASAP7_75t_L g784 ( 
.A1(n_622),
.A2(n_288),
.B(n_293),
.C(n_294),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_756),
.B(n_485),
.Y(n_785)
);

INVx3_ASAP7_75t_L g786 ( 
.A(n_636),
.Y(n_786)
);

NAND2xp5_ASAP7_75t_SL g787 ( 
.A(n_636),
.B(n_502),
.Y(n_787)
);

NAND2xp33_ASAP7_75t_L g788 ( 
.A(n_749),
.B(n_502),
.Y(n_788)
);

O2A1O1Ixp33_ASAP7_75t_L g789 ( 
.A1(n_614),
.A2(n_490),
.B(n_447),
.C(n_569),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_609),
.B(n_268),
.Y(n_790)
);

HB1xp67_ASAP7_75t_L g791 ( 
.A(n_596),
.Y(n_791)
);

INVxp67_ASAP7_75t_L g792 ( 
.A(n_630),
.Y(n_792)
);

O2A1O1Ixp33_ASAP7_75t_L g793 ( 
.A1(n_621),
.A2(n_490),
.B(n_447),
.C(n_569),
.Y(n_793)
);

INVx3_ASAP7_75t_L g794 ( 
.A(n_636),
.Y(n_794)
);

NAND2xp5_ASAP7_75t_L g795 ( 
.A(n_756),
.B(n_485),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_654),
.B(n_485),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_747),
.B(n_293),
.Y(n_797)
);

AOI21xp5_ASAP7_75t_L g798 ( 
.A1(n_680),
.A2(n_506),
.B(n_482),
.Y(n_798)
);

O2A1O1Ixp33_ASAP7_75t_L g799 ( 
.A1(n_689),
.A2(n_512),
.B(n_476),
.C(n_479),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_663),
.B(n_485),
.Y(n_800)
);

AND2x2_ASAP7_75t_L g801 ( 
.A(n_648),
.B(n_299),
.Y(n_801)
);

INVxp67_ASAP7_75t_SL g802 ( 
.A(n_739),
.Y(n_802)
);

BUFx3_ASAP7_75t_L g803 ( 
.A(n_626),
.Y(n_803)
);

NOR2xp33_ASAP7_75t_L g804 ( 
.A(n_601),
.B(n_270),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_628),
.Y(n_805)
);

BUFx4f_ASAP7_75t_L g806 ( 
.A(n_683),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_636),
.Y(n_807)
);

INVx2_ASAP7_75t_L g808 ( 
.A(n_651),
.Y(n_808)
);

NAND2xp5_ASAP7_75t_L g809 ( 
.A(n_672),
.B(n_501),
.Y(n_809)
);

NOR2xp33_ASAP7_75t_L g810 ( 
.A(n_601),
.B(n_299),
.Y(n_810)
);

NOR2xp33_ASAP7_75t_L g811 ( 
.A(n_740),
.B(n_726),
.Y(n_811)
);

CKINVDCx5p33_ASAP7_75t_R g812 ( 
.A(n_748),
.Y(n_812)
);

INVx1_ASAP7_75t_L g813 ( 
.A(n_662),
.Y(n_813)
);

A2O1A1Ixp33_ASAP7_75t_L g814 ( 
.A1(n_661),
.A2(n_306),
.B(n_511),
.C(n_505),
.Y(n_814)
);

AOI22xp5_ASAP7_75t_L g815 ( 
.A1(n_616),
.A2(n_587),
.B1(n_573),
.B2(n_567),
.Y(n_815)
);

A2O1A1Ixp33_ASAP7_75t_L g816 ( 
.A1(n_661),
.A2(n_306),
.B(n_511),
.C(n_505),
.Y(n_816)
);

AND2x4_ASAP7_75t_L g817 ( 
.A(n_690),
.B(n_501),
.Y(n_817)
);

OAI22xp5_ASAP7_75t_L g818 ( 
.A1(n_606),
.A2(n_632),
.B1(n_657),
.B2(n_659),
.Y(n_818)
);

HB1xp67_ASAP7_75t_L g819 ( 
.A(n_694),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_662),
.Y(n_820)
);

INVx4_ASAP7_75t_L g821 ( 
.A(n_755),
.Y(n_821)
);

HB1xp67_ASAP7_75t_L g822 ( 
.A(n_694),
.Y(n_822)
);

INVx1_ASAP7_75t_L g823 ( 
.A(n_669),
.Y(n_823)
);

AND2x4_ASAP7_75t_L g824 ( 
.A(n_693),
.B(n_626),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_L g825 ( 
.A(n_673),
.B(n_501),
.Y(n_825)
);

AO21x1_ASAP7_75t_L g826 ( 
.A1(n_708),
.A2(n_506),
.B(n_535),
.Y(n_826)
);

A2O1A1Ixp33_ASAP7_75t_L g827 ( 
.A1(n_668),
.A2(n_530),
.B(n_504),
.C(n_481),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_676),
.B(n_519),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_681),
.B(n_519),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_688),
.B(n_519),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_593),
.B(n_519),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_653),
.B(n_417),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_682),
.A2(n_535),
.B(n_482),
.Y(n_833)
);

OR2x2_ASAP7_75t_L g834 ( 
.A(n_698),
.B(n_15),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_753),
.A2(n_629),
.B(n_745),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_646),
.A2(n_711),
.B(n_710),
.Y(n_836)
);

AND2x4_ASAP7_75t_L g837 ( 
.A(n_709),
.B(n_542),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_595),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_687),
.B(n_542),
.Y(n_839)
);

AOI21xp5_ASAP7_75t_L g840 ( 
.A1(n_613),
.A2(n_535),
.B(n_502),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_695),
.Y(n_841)
);

NAND2xp5_ASAP7_75t_L g842 ( 
.A(n_623),
.B(n_542),
.Y(n_842)
);

AOI22xp5_ASAP7_75t_L g843 ( 
.A1(n_713),
.A2(n_587),
.B1(n_573),
.B2(n_567),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_633),
.A2(n_535),
.B(n_540),
.Y(n_844)
);

AOI21xp5_ASAP7_75t_L g845 ( 
.A1(n_639),
.A2(n_558),
.B(n_540),
.Y(n_845)
);

BUFx3_ASAP7_75t_L g846 ( 
.A(n_683),
.Y(n_846)
);

AOI22xp5_ASAP7_75t_L g847 ( 
.A1(n_677),
.A2(n_587),
.B1(n_573),
.B2(n_567),
.Y(n_847)
);

OAI21xp5_ASAP7_75t_L g848 ( 
.A1(n_675),
.A2(n_559),
.B(n_504),
.Y(n_848)
);

INVx4_ASAP7_75t_L g849 ( 
.A(n_755),
.Y(n_849)
);

NAND2xp33_ASAP7_75t_L g850 ( 
.A(n_749),
.B(n_540),
.Y(n_850)
);

AOI22xp5_ASAP7_75t_L g851 ( 
.A1(n_677),
.A2(n_715),
.B1(n_649),
.B2(n_660),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_697),
.Y(n_852)
);

OAI22xp5_ASAP7_75t_L g853 ( 
.A1(n_606),
.A2(n_557),
.B1(n_552),
.B2(n_546),
.Y(n_853)
);

INVx1_ASAP7_75t_L g854 ( 
.A(n_699),
.Y(n_854)
);

AOI21xp5_ASAP7_75t_L g855 ( 
.A1(n_642),
.A2(n_540),
.B(n_558),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_645),
.B(n_512),
.Y(n_856)
);

AND2x2_ASAP7_75t_L g857 ( 
.A(n_685),
.B(n_543),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_739),
.A2(n_558),
.B(n_540),
.Y(n_858)
);

OAI21xp5_ASAP7_75t_L g859 ( 
.A1(n_657),
.A2(n_559),
.B(n_530),
.Y(n_859)
);

AND2x4_ASAP7_75t_L g860 ( 
.A(n_627),
.B(n_557),
.Y(n_860)
);

NOR3xp33_ASAP7_75t_L g861 ( 
.A(n_635),
.B(n_546),
.C(n_557),
.Y(n_861)
);

INVx2_ASAP7_75t_SL g862 ( 
.A(n_647),
.Y(n_862)
);

INVx3_ASAP7_75t_L g863 ( 
.A(n_627),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_SL g864 ( 
.A(n_749),
.B(n_558),
.Y(n_864)
);

NAND2xp5_ASAP7_75t_L g865 ( 
.A(n_602),
.B(n_546),
.Y(n_865)
);

NAND2xp5_ASAP7_75t_SL g866 ( 
.A(n_749),
.B(n_739),
.Y(n_866)
);

AOI21xp5_ASAP7_75t_L g867 ( 
.A1(n_739),
.A2(n_558),
.B(n_540),
.Y(n_867)
);

AOI21xp5_ASAP7_75t_L g868 ( 
.A1(n_608),
.A2(n_558),
.B(n_557),
.Y(n_868)
);

OAI21xp5_ASAP7_75t_L g869 ( 
.A1(n_611),
.A2(n_559),
.B(n_504),
.Y(n_869)
);

INVx1_ASAP7_75t_L g870 ( 
.A(n_718),
.Y(n_870)
);

NAND2xp5_ASAP7_75t_L g871 ( 
.A(n_603),
.B(n_552),
.Y(n_871)
);

AND2x2_ASAP7_75t_L g872 ( 
.A(n_722),
.B(n_499),
.Y(n_872)
);

NOR2xp67_ASAP7_75t_L g873 ( 
.A(n_715),
.B(n_552),
.Y(n_873)
);

AOI21xp5_ASAP7_75t_L g874 ( 
.A1(n_612),
.A2(n_552),
.B(n_546),
.Y(n_874)
);

OAI21xp5_ASAP7_75t_L g875 ( 
.A1(n_659),
.A2(n_530),
.B(n_543),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_599),
.Y(n_876)
);

NAND2xp5_ASAP7_75t_L g877 ( 
.A(n_618),
.B(n_529),
.Y(n_877)
);

AOI21xp5_ASAP7_75t_L g878 ( 
.A1(n_620),
.A2(n_524),
.B(n_529),
.Y(n_878)
);

NAND2xp5_ASAP7_75t_SL g879 ( 
.A(n_749),
.B(n_499),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_735),
.Y(n_880)
);

O2A1O1Ixp33_ASAP7_75t_SL g881 ( 
.A1(n_696),
.A2(n_476),
.B(n_479),
.C(n_19),
.Y(n_881)
);

AOI22xp5_ASAP7_75t_L g882 ( 
.A1(n_677),
.A2(n_427),
.B1(n_423),
.B2(n_416),
.Y(n_882)
);

INVx2_ASAP7_75t_L g883 ( 
.A(n_605),
.Y(n_883)
);

NAND2xp5_ASAP7_75t_SL g884 ( 
.A(n_605),
.B(n_427),
.Y(n_884)
);

OAI22xp5_ASAP7_75t_L g885 ( 
.A1(n_649),
.A2(n_427),
.B1(n_423),
.B2(n_416),
.Y(n_885)
);

AOI21xp5_ASAP7_75t_L g886 ( 
.A1(n_619),
.A2(n_524),
.B(n_395),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_741),
.Y(n_887)
);

AOI22xp33_ASAP7_75t_L g888 ( 
.A1(n_723),
.A2(n_427),
.B1(n_423),
.B2(n_395),
.Y(n_888)
);

HB1xp67_ASAP7_75t_L g889 ( 
.A(n_730),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_743),
.Y(n_890)
);

AND2x2_ASAP7_75t_L g891 ( 
.A(n_655),
.B(n_423),
.Y(n_891)
);

INVx1_ASAP7_75t_L g892 ( 
.A(n_637),
.Y(n_892)
);

NAND2xp5_ASAP7_75t_L g893 ( 
.A(n_638),
.B(n_427),
.Y(n_893)
);

NAND2xp5_ASAP7_75t_SL g894 ( 
.A(n_752),
.B(n_423),
.Y(n_894)
);

A2O1A1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_668),
.A2(n_423),
.B(n_395),
.C(n_19),
.Y(n_895)
);

HB1xp67_ASAP7_75t_L g896 ( 
.A(n_640),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_644),
.B(n_423),
.Y(n_897)
);

INVx1_ASAP7_75t_L g898 ( 
.A(n_702),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_720),
.B(n_524),
.Y(n_899)
);

NAND2xp5_ASAP7_75t_L g900 ( 
.A(n_607),
.B(n_524),
.Y(n_900)
);

AOI21x1_ASAP7_75t_L g901 ( 
.A1(n_738),
.A2(n_58),
.B(n_136),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_655),
.B(n_15),
.Y(n_902)
);

OAI22xp5_ASAP7_75t_L g903 ( 
.A1(n_660),
.A2(n_60),
.B1(n_128),
.B2(n_127),
.Y(n_903)
);

NOR2xp33_ASAP7_75t_L g904 ( 
.A(n_691),
.B(n_16),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_SL g905 ( 
.A(n_720),
.B(n_724),
.Y(n_905)
);

AOI21xp5_ASAP7_75t_L g906 ( 
.A1(n_712),
.A2(n_716),
.B(n_727),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_705),
.Y(n_907)
);

BUFx6f_ASAP7_75t_L g908 ( 
.A(n_705),
.Y(n_908)
);

AOI21xp5_ASAP7_75t_L g909 ( 
.A1(n_717),
.A2(n_148),
.B(n_125),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_719),
.Y(n_910)
);

AOI22xp5_ASAP7_75t_L g911 ( 
.A1(n_670),
.A2(n_121),
.B1(n_120),
.B2(n_100),
.Y(n_911)
);

NOR2xp33_ASAP7_75t_L g912 ( 
.A(n_594),
.B(n_16),
.Y(n_912)
);

O2A1O1Ixp33_ASAP7_75t_L g913 ( 
.A1(n_723),
.A2(n_20),
.B(n_28),
.C(n_31),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_670),
.B(n_34),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_L g915 ( 
.A(n_671),
.B(n_35),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_721),
.A2(n_53),
.B(n_91),
.Y(n_916)
);

INVx3_ASAP7_75t_L g917 ( 
.A(n_719),
.Y(n_917)
);

OAI21xp5_ASAP7_75t_L g918 ( 
.A1(n_732),
.A2(n_94),
.B(n_89),
.Y(n_918)
);

AOI21xp5_ASAP7_75t_L g919 ( 
.A1(n_706),
.A2(n_734),
.B(n_733),
.Y(n_919)
);

INVx1_ASAP7_75t_L g920 ( 
.A(n_732),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_671),
.B(n_38),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_706),
.A2(n_87),
.B(n_84),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_738),
.A2(n_78),
.B(n_76),
.Y(n_923)
);

NAND2xp5_ASAP7_75t_L g924 ( 
.A(n_707),
.B(n_40),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_703),
.A2(n_70),
.B(n_67),
.Y(n_925)
);

AOI21xp5_ASAP7_75t_L g926 ( 
.A1(n_731),
.A2(n_746),
.B(n_736),
.Y(n_926)
);

OAI21xp5_ASAP7_75t_L g927 ( 
.A1(n_746),
.A2(n_61),
.B(n_45),
.Y(n_927)
);

AOI221xp5_ASAP7_75t_SL g928 ( 
.A1(n_725),
.A2(n_41),
.B1(n_46),
.B2(n_47),
.C(n_48),
.Y(n_928)
);

INVx4_ASAP7_75t_L g929 ( 
.A(n_674),
.Y(n_929)
);

OAI21xp33_ASAP7_75t_L g930 ( 
.A1(n_725),
.A2(n_41),
.B(n_49),
.Y(n_930)
);

INVx1_ASAP7_75t_SL g931 ( 
.A(n_631),
.Y(n_931)
);

AND2x2_ASAP7_75t_L g932 ( 
.A(n_801),
.B(n_707),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_761),
.B(n_744),
.Y(n_933)
);

NAND2xp5_ASAP7_75t_SL g934 ( 
.A(n_851),
.B(n_641),
.Y(n_934)
);

NOR2x1_ASAP7_75t_L g935 ( 
.A(n_821),
.B(n_610),
.Y(n_935)
);

CKINVDCx14_ASAP7_75t_R g936 ( 
.A(n_812),
.Y(n_936)
);

INVx3_ASAP7_75t_L g937 ( 
.A(n_860),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_902),
.A2(n_915),
.B(n_921),
.C(n_914),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_804),
.B(n_744),
.Y(n_939)
);

NAND2xp5_ASAP7_75t_L g940 ( 
.A(n_804),
.B(n_810),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_760),
.A2(n_650),
.B(n_684),
.Y(n_941)
);

INVxp67_ASAP7_75t_SL g942 ( 
.A(n_819),
.Y(n_942)
);

INVx2_ASAP7_75t_SL g943 ( 
.A(n_772),
.Y(n_943)
);

A2O1A1Ixp33_ASAP7_75t_L g944 ( 
.A1(n_810),
.A2(n_912),
.B(n_924),
.C(n_769),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_764),
.A2(n_773),
.B(n_788),
.Y(n_945)
);

NAND2xp5_ASAP7_75t_SL g946 ( 
.A(n_759),
.B(n_658),
.Y(n_946)
);

INVx2_ASAP7_75t_L g947 ( 
.A(n_917),
.Y(n_947)
);

AOI21xp5_ASAP7_75t_L g948 ( 
.A1(n_850),
.A2(n_754),
.B(n_714),
.Y(n_948)
);

NAND2xp5_ASAP7_75t_L g949 ( 
.A(n_832),
.B(n_600),
.Y(n_949)
);

BUFx8_ASAP7_75t_SL g950 ( 
.A(n_806),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_SL g951 ( 
.A(n_824),
.B(n_803),
.Y(n_951)
);

OAI22xp5_ASAP7_75t_L g952 ( 
.A1(n_818),
.A2(n_692),
.B1(n_686),
.B2(n_700),
.Y(n_952)
);

NAND2xp5_ASAP7_75t_L g953 ( 
.A(n_872),
.B(n_729),
.Y(n_953)
);

INVx2_ASAP7_75t_L g954 ( 
.A(n_917),
.Y(n_954)
);

INVxp67_ASAP7_75t_SL g955 ( 
.A(n_819),
.Y(n_955)
);

NAND2xp5_ASAP7_75t_L g956 ( 
.A(n_896),
.B(n_643),
.Y(n_956)
);

O2A1O1Ixp33_ASAP7_75t_L g957 ( 
.A1(n_895),
.A2(n_905),
.B(n_930),
.C(n_913),
.Y(n_957)
);

O2A1O1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_895),
.A2(n_701),
.B(n_751),
.C(n_674),
.Y(n_958)
);

INVxp67_ASAP7_75t_L g959 ( 
.A(n_772),
.Y(n_959)
);

A2O1A1Ixp33_ASAP7_75t_L g960 ( 
.A1(n_912),
.A2(n_683),
.B(n_50),
.C(n_51),
.Y(n_960)
);

A2O1A1Ixp33_ASAP7_75t_L g961 ( 
.A1(n_919),
.A2(n_905),
.B(n_790),
.C(n_927),
.Y(n_961)
);

AOI21xp5_ASAP7_75t_L g962 ( 
.A1(n_835),
.A2(n_778),
.B(n_777),
.Y(n_962)
);

NOR2xp33_ASAP7_75t_L g963 ( 
.A(n_792),
.B(n_49),
.Y(n_963)
);

BUFx6f_ASAP7_75t_L g964 ( 
.A(n_821),
.Y(n_964)
);

OAI22x1_ASAP7_75t_L g965 ( 
.A1(n_904),
.A2(n_50),
.B1(n_52),
.B2(n_889),
.Y(n_965)
);

NAND2xp5_ASAP7_75t_L g966 ( 
.A(n_896),
.B(n_822),
.Y(n_966)
);

OAI22xp5_ASAP7_75t_L g967 ( 
.A1(n_822),
.A2(n_765),
.B1(n_785),
.B2(n_795),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_770),
.Y(n_968)
);

INVx2_ASAP7_75t_L g969 ( 
.A(n_910),
.Y(n_969)
);

INVx3_ASAP7_75t_L g970 ( 
.A(n_860),
.Y(n_970)
);

NOR2xp33_ASAP7_75t_L g971 ( 
.A(n_790),
.B(n_931),
.Y(n_971)
);

O2A1O1Ixp33_ASAP7_75t_L g972 ( 
.A1(n_814),
.A2(n_816),
.B(n_827),
.C(n_782),
.Y(n_972)
);

BUFx2_ASAP7_75t_L g973 ( 
.A(n_889),
.Y(n_973)
);

INVx4_ASAP7_75t_L g974 ( 
.A(n_849),
.Y(n_974)
);

INVx2_ASAP7_75t_L g975 ( 
.A(n_758),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_824),
.B(n_803),
.Y(n_976)
);

NAND2xp5_ASAP7_75t_L g977 ( 
.A(n_892),
.B(n_791),
.Y(n_977)
);

A2O1A1Ixp33_ASAP7_75t_SL g978 ( 
.A1(n_811),
.A2(n_904),
.B(n_918),
.C(n_861),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_791),
.B(n_841),
.Y(n_979)
);

BUFx6f_ASAP7_75t_L g980 ( 
.A(n_786),
.Y(n_980)
);

O2A1O1Ixp5_ASAP7_75t_L g981 ( 
.A1(n_826),
.A2(n_757),
.B(n_767),
.C(n_766),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_814),
.A2(n_816),
.B(n_827),
.C(n_782),
.Y(n_982)
);

AOI22xp33_ASAP7_75t_SL g983 ( 
.A1(n_834),
.A2(n_862),
.B1(n_806),
.B2(n_929),
.Y(n_983)
);

AOI22xp5_ASAP7_75t_L g984 ( 
.A1(n_811),
.A2(n_837),
.B1(n_817),
.B2(n_861),
.Y(n_984)
);

INVx2_ASAP7_75t_L g985 ( 
.A(n_776),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_863),
.B(n_817),
.Y(n_986)
);

NOR2xp33_ASAP7_75t_L g987 ( 
.A(n_797),
.B(n_784),
.Y(n_987)
);

O2A1O1Ixp33_ASAP7_75t_L g988 ( 
.A1(n_784),
.A2(n_881),
.B(n_813),
.C(n_820),
.Y(n_988)
);

INVx2_ASAP7_75t_L g989 ( 
.A(n_781),
.Y(n_989)
);

BUFx6f_ASAP7_75t_L g990 ( 
.A(n_786),
.Y(n_990)
);

OAI22xp33_ASAP7_75t_L g991 ( 
.A1(n_852),
.A2(n_887),
.B1(n_890),
.B2(n_870),
.Y(n_991)
);

BUFx12f_ASAP7_75t_L g992 ( 
.A(n_929),
.Y(n_992)
);

NAND2xp5_ASAP7_75t_SL g993 ( 
.A(n_863),
.B(n_854),
.Y(n_993)
);

OR2x2_ASAP7_75t_L g994 ( 
.A(n_880),
.B(n_837),
.Y(n_994)
);

OAI22xp5_ASAP7_75t_L g995 ( 
.A1(n_780),
.A2(n_783),
.B1(n_847),
.B2(n_802),
.Y(n_995)
);

AOI21xp5_ASAP7_75t_L g996 ( 
.A1(n_891),
.A2(n_762),
.B(n_873),
.Y(n_996)
);

BUFx12f_ASAP7_75t_L g997 ( 
.A(n_846),
.Y(n_997)
);

INVx3_ASAP7_75t_L g998 ( 
.A(n_794),
.Y(n_998)
);

BUFx6f_ASAP7_75t_L g999 ( 
.A(n_794),
.Y(n_999)
);

AOI21xp5_ASAP7_75t_L g1000 ( 
.A1(n_840),
.A2(n_836),
.B(n_831),
.Y(n_1000)
);

A2O1A1Ixp33_ASAP7_75t_L g1001 ( 
.A1(n_926),
.A2(n_823),
.B(n_793),
.C(n_805),
.Y(n_1001)
);

INVx3_ASAP7_75t_L g1002 ( 
.A(n_807),
.Y(n_1002)
);

A2O1A1Ixp33_ASAP7_75t_L g1003 ( 
.A1(n_808),
.A2(n_789),
.B(n_874),
.C(n_906),
.Y(n_1003)
);

OAI22xp5_ASAP7_75t_L g1004 ( 
.A1(n_802),
.A2(n_899),
.B1(n_866),
.B2(n_864),
.Y(n_1004)
);

O2A1O1Ixp33_ASAP7_75t_L g1005 ( 
.A1(n_881),
.A2(n_903),
.B(n_842),
.C(n_763),
.Y(n_1005)
);

BUFx12f_ASAP7_75t_L g1006 ( 
.A(n_846),
.Y(n_1006)
);

INVx2_ASAP7_75t_L g1007 ( 
.A(n_876),
.Y(n_1007)
);

A2O1A1Ixp33_ASAP7_75t_L g1008 ( 
.A1(n_911),
.A2(n_799),
.B(n_868),
.C(n_916),
.Y(n_1008)
);

NOR3xp33_ASAP7_75t_SL g1009 ( 
.A(n_838),
.B(n_925),
.C(n_922),
.Y(n_1009)
);

AOI21xp5_ASAP7_75t_L g1010 ( 
.A1(n_768),
.A2(n_771),
.B(n_774),
.Y(n_1010)
);

OAI21xp5_ASAP7_75t_L g1011 ( 
.A1(n_899),
.A2(n_779),
.B(n_853),
.Y(n_1011)
);

NOR3xp33_ASAP7_75t_L g1012 ( 
.A(n_909),
.B(n_807),
.C(n_928),
.Y(n_1012)
);

OAI22xp5_ASAP7_75t_SL g1013 ( 
.A1(n_843),
.A2(n_815),
.B1(n_920),
.B2(n_898),
.Y(n_1013)
);

O2A1O1Ixp33_ASAP7_75t_L g1014 ( 
.A1(n_877),
.A2(n_865),
.B(n_871),
.C(n_829),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_SL g1015 ( 
.A(n_856),
.B(n_857),
.Y(n_1015)
);

INVx3_ASAP7_75t_SL g1016 ( 
.A(n_866),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_864),
.A2(n_787),
.B1(n_809),
.B2(n_800),
.Y(n_1017)
);

OAI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_859),
.A2(n_875),
.B(n_869),
.Y(n_1018)
);

AND2x2_ASAP7_75t_L g1019 ( 
.A(n_883),
.B(n_907),
.Y(n_1019)
);

BUFx6f_ASAP7_75t_L g1020 ( 
.A(n_908),
.Y(n_1020)
);

AOI22xp33_ASAP7_75t_L g1021 ( 
.A1(n_908),
.A2(n_830),
.B1(n_828),
.B2(n_825),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_775),
.A2(n_833),
.B(n_798),
.Y(n_1022)
);

INVx2_ASAP7_75t_L g1023 ( 
.A(n_908),
.Y(n_1023)
);

O2A1O1Ixp33_ASAP7_75t_SL g1024 ( 
.A1(n_787),
.A2(n_879),
.B(n_900),
.C(n_796),
.Y(n_1024)
);

AOI21xp5_ASAP7_75t_L g1025 ( 
.A1(n_844),
.A2(n_855),
.B(n_845),
.Y(n_1025)
);

INVx4_ASAP7_75t_L g1026 ( 
.A(n_908),
.Y(n_1026)
);

O2A1O1Ixp33_ASAP7_75t_L g1027 ( 
.A1(n_848),
.A2(n_894),
.B(n_839),
.C(n_897),
.Y(n_1027)
);

AND2x2_ASAP7_75t_L g1028 ( 
.A(n_894),
.B(n_884),
.Y(n_1028)
);

OA21x2_ASAP7_75t_L g1029 ( 
.A1(n_888),
.A2(n_893),
.B(n_884),
.Y(n_1029)
);

AND2x2_ASAP7_75t_L g1030 ( 
.A(n_882),
.B(n_879),
.Y(n_1030)
);

O2A1O1Ixp33_ASAP7_75t_L g1031 ( 
.A1(n_885),
.A2(n_923),
.B(n_878),
.C(n_886),
.Y(n_1031)
);

AOI21xp5_ASAP7_75t_L g1032 ( 
.A1(n_858),
.A2(n_867),
.B(n_888),
.Y(n_1032)
);

INVx3_ASAP7_75t_L g1033 ( 
.A(n_901),
.Y(n_1033)
);

AOI21xp5_ASAP7_75t_L g1034 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1034)
);

A2O1A1Ixp33_ASAP7_75t_L g1035 ( 
.A1(n_804),
.A2(n_810),
.B(n_851),
.C(n_902),
.Y(n_1035)
);

NAND3xp33_ASAP7_75t_SL g1036 ( 
.A(n_851),
.B(n_810),
.C(n_804),
.Y(n_1036)
);

AOI21xp5_ASAP7_75t_L g1037 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1037)
);

AOI21x1_ASAP7_75t_L g1038 ( 
.A1(n_873),
.A2(n_795),
.B(n_785),
.Y(n_1038)
);

AOI21xp5_ASAP7_75t_L g1039 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1039)
);

AOI21xp5_ASAP7_75t_L g1040 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_761),
.B(n_615),
.Y(n_1041)
);

INVx4_ASAP7_75t_L g1042 ( 
.A(n_821),
.Y(n_1042)
);

OAI22x1_ASAP7_75t_L g1043 ( 
.A1(n_851),
.A2(n_462),
.B1(n_810),
.B2(n_730),
.Y(n_1043)
);

BUFx10_ASAP7_75t_L g1044 ( 
.A(n_790),
.Y(n_1044)
);

AOI21xp5_ASAP7_75t_L g1045 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1045)
);

NAND2xp5_ASAP7_75t_L g1046 ( 
.A(n_761),
.B(n_615),
.Y(n_1046)
);

AND2x4_ASAP7_75t_L g1047 ( 
.A(n_803),
.B(n_824),
.Y(n_1047)
);

NAND3xp33_ASAP7_75t_L g1048 ( 
.A(n_810),
.B(n_804),
.C(n_851),
.Y(n_1048)
);

AOI21xp5_ASAP7_75t_L g1049 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1049)
);

BUFx3_ASAP7_75t_L g1050 ( 
.A(n_846),
.Y(n_1050)
);

O2A1O1Ixp33_ASAP7_75t_SL g1051 ( 
.A1(n_905),
.A2(n_902),
.B(n_895),
.C(n_621),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_761),
.B(n_615),
.Y(n_1052)
);

A2O1A1Ixp33_ASAP7_75t_L g1053 ( 
.A1(n_804),
.A2(n_810),
.B(n_851),
.C(n_902),
.Y(n_1053)
);

AOI21xp5_ASAP7_75t_L g1054 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1054)
);

O2A1O1Ixp5_ASAP7_75t_L g1055 ( 
.A1(n_804),
.A2(n_764),
.B(n_810),
.C(n_902),
.Y(n_1055)
);

NAND2xp5_ASAP7_75t_L g1056 ( 
.A(n_761),
.B(n_615),
.Y(n_1056)
);

O2A1O1Ixp33_ASAP7_75t_L g1057 ( 
.A1(n_902),
.A2(n_915),
.B(n_921),
.C(n_914),
.Y(n_1057)
);

INVx3_ASAP7_75t_L g1058 ( 
.A(n_860),
.Y(n_1058)
);

AOI21xp5_ASAP7_75t_L g1059 ( 
.A1(n_760),
.A2(n_764),
.B(n_773),
.Y(n_1059)
);

AND2x2_ASAP7_75t_L g1060 ( 
.A(n_801),
.B(n_810),
.Y(n_1060)
);

INVx3_ASAP7_75t_L g1061 ( 
.A(n_860),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_761),
.B(n_615),
.Y(n_1062)
);

INVx3_ASAP7_75t_L g1063 ( 
.A(n_1026),
.Y(n_1063)
);

NAND2xp5_ASAP7_75t_L g1064 ( 
.A(n_940),
.B(n_1041),
.Y(n_1064)
);

BUFx2_ASAP7_75t_L g1065 ( 
.A(n_973),
.Y(n_1065)
);

AOI221xp5_ASAP7_75t_L g1066 ( 
.A1(n_1036),
.A2(n_939),
.B1(n_1048),
.B2(n_987),
.C(n_1043),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1035),
.A2(n_1053),
.B(n_1055),
.Y(n_1067)
);

A2O1A1Ixp33_ASAP7_75t_L g1068 ( 
.A1(n_944),
.A2(n_938),
.B(n_1057),
.C(n_957),
.Y(n_1068)
);

AOI22xp5_ASAP7_75t_L g1069 ( 
.A1(n_1060),
.A2(n_971),
.B1(n_932),
.B2(n_934),
.Y(n_1069)
);

BUFx8_ASAP7_75t_L g1070 ( 
.A(n_992),
.Y(n_1070)
);

OAI22xp5_ASAP7_75t_SL g1071 ( 
.A1(n_965),
.A2(n_983),
.B1(n_963),
.B2(n_936),
.Y(n_1071)
);

NOR2xp33_ASAP7_75t_L g1072 ( 
.A(n_1044),
.B(n_959),
.Y(n_1072)
);

INVx1_ASAP7_75t_SL g1073 ( 
.A(n_943),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_964),
.Y(n_1074)
);

NOR2xp33_ASAP7_75t_L g1075 ( 
.A(n_1044),
.B(n_966),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1034),
.A2(n_1045),
.B(n_1059),
.Y(n_1076)
);

OR2x2_ASAP7_75t_L g1077 ( 
.A(n_1062),
.B(n_1046),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1034),
.A2(n_1049),
.B(n_1045),
.Y(n_1078)
);

HB1xp67_ASAP7_75t_L g1079 ( 
.A(n_1047),
.Y(n_1079)
);

AO31x2_ASAP7_75t_L g1080 ( 
.A1(n_961),
.A2(n_996),
.A3(n_995),
.B(n_1003),
.Y(n_1080)
);

AO32x2_ASAP7_75t_L g1081 ( 
.A1(n_967),
.A2(n_952),
.A3(n_1013),
.B1(n_1004),
.B2(n_1017),
.Y(n_1081)
);

BUFx3_ASAP7_75t_L g1082 ( 
.A(n_997),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1037),
.A2(n_1039),
.B(n_1059),
.Y(n_1083)
);

BUFx3_ASAP7_75t_L g1084 ( 
.A(n_1006),
.Y(n_1084)
);

OAI22x1_ASAP7_75t_L g1085 ( 
.A1(n_1016),
.A2(n_984),
.B1(n_956),
.B2(n_935),
.Y(n_1085)
);

BUFx2_ASAP7_75t_L g1086 ( 
.A(n_1050),
.Y(n_1086)
);

OAI21xp5_ASAP7_75t_L g1087 ( 
.A1(n_938),
.A2(n_1057),
.B(n_953),
.Y(n_1087)
);

O2A1O1Ixp33_ASAP7_75t_SL g1088 ( 
.A1(n_978),
.A2(n_933),
.B(n_1008),
.C(n_949),
.Y(n_1088)
);

A2O1A1Ixp33_ASAP7_75t_L g1089 ( 
.A1(n_957),
.A2(n_941),
.B(n_958),
.C(n_1056),
.Y(n_1089)
);

CKINVDCx20_ASAP7_75t_R g1090 ( 
.A(n_950),
.Y(n_1090)
);

NAND2xp5_ASAP7_75t_L g1091 ( 
.A(n_1052),
.B(n_977),
.Y(n_1091)
);

OAI21xp5_ASAP7_75t_L g1092 ( 
.A1(n_946),
.A2(n_941),
.B(n_1011),
.Y(n_1092)
);

CKINVDCx11_ASAP7_75t_R g1093 ( 
.A(n_964),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_979),
.B(n_1015),
.Y(n_1094)
);

AOI21x1_ASAP7_75t_L g1095 ( 
.A1(n_1038),
.A2(n_945),
.B(n_996),
.Y(n_1095)
);

AO31x2_ASAP7_75t_L g1096 ( 
.A1(n_962),
.A2(n_1049),
.A3(n_1040),
.B(n_1039),
.Y(n_1096)
);

AND2x2_ASAP7_75t_L g1097 ( 
.A(n_942),
.B(n_955),
.Y(n_1097)
);

AO31x2_ASAP7_75t_L g1098 ( 
.A1(n_962),
.A2(n_1054),
.A3(n_1040),
.B(n_1037),
.Y(n_1098)
);

AO31x2_ASAP7_75t_L g1099 ( 
.A1(n_1054),
.A2(n_1022),
.A3(n_1025),
.B(n_945),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_991),
.B(n_994),
.Y(n_1100)
);

AOI21x1_ASAP7_75t_L g1101 ( 
.A1(n_1032),
.A2(n_1022),
.B(n_1010),
.Y(n_1101)
);

AOI221xp5_ASAP7_75t_L g1102 ( 
.A1(n_1051),
.A2(n_960),
.B1(n_958),
.B2(n_982),
.C(n_972),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_951),
.B(n_976),
.Y(n_1103)
);

AOI21xp5_ASAP7_75t_L g1104 ( 
.A1(n_1000),
.A2(n_1018),
.B(n_1010),
.Y(n_1104)
);

OAI21x1_ASAP7_75t_L g1105 ( 
.A1(n_1025),
.A2(n_1032),
.B(n_1000),
.Y(n_1105)
);

O2A1O1Ixp33_ASAP7_75t_SL g1106 ( 
.A1(n_1001),
.A2(n_972),
.B(n_982),
.C(n_993),
.Y(n_1106)
);

AOI221x1_ASAP7_75t_L g1107 ( 
.A1(n_1012),
.A2(n_948),
.B1(n_1033),
.B2(n_1030),
.C(n_968),
.Y(n_1107)
);

NAND2xp5_ASAP7_75t_L g1108 ( 
.A(n_937),
.B(n_1061),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_L g1109 ( 
.A1(n_1014),
.A2(n_1024),
.B(n_1005),
.Y(n_1109)
);

INVx1_ASAP7_75t_L g1110 ( 
.A(n_1019),
.Y(n_1110)
);

AOI21xp5_ASAP7_75t_L g1111 ( 
.A1(n_1014),
.A2(n_1005),
.B(n_1031),
.Y(n_1111)
);

AOI21xp5_ASAP7_75t_L g1112 ( 
.A1(n_1031),
.A2(n_948),
.B(n_1027),
.Y(n_1112)
);

AOI21xp5_ASAP7_75t_L g1113 ( 
.A1(n_1027),
.A2(n_981),
.B(n_1021),
.Y(n_1113)
);

A2O1A1Ixp33_ASAP7_75t_L g1114 ( 
.A1(n_988),
.A2(n_1009),
.B(n_989),
.C(n_985),
.Y(n_1114)
);

NOR2x1_ASAP7_75t_L g1115 ( 
.A(n_1026),
.B(n_1002),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_937),
.B(n_1058),
.Y(n_1116)
);

NAND2xp5_ASAP7_75t_L g1117 ( 
.A(n_970),
.B(n_1061),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_1029),
.A2(n_1033),
.B(n_988),
.Y(n_1118)
);

AOI21xp5_ASAP7_75t_L g1119 ( 
.A1(n_1029),
.A2(n_986),
.B(n_1028),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_969),
.Y(n_1120)
);

AND2x6_ASAP7_75t_L g1121 ( 
.A(n_1020),
.B(n_1058),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_1007),
.Y(n_1122)
);

AO31x2_ASAP7_75t_L g1123 ( 
.A1(n_1023),
.A2(n_947),
.A3(n_954),
.B(n_975),
.Y(n_1123)
);

OAI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_970),
.A2(n_998),
.B(n_974),
.Y(n_1124)
);

A2O1A1Ixp33_ASAP7_75t_L g1125 ( 
.A1(n_1020),
.A2(n_980),
.B(n_990),
.C(n_999),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_1042),
.B(n_980),
.Y(n_1126)
);

OAI22xp5_ASAP7_75t_L g1127 ( 
.A1(n_1020),
.A2(n_999),
.B1(n_980),
.B2(n_990),
.Y(n_1127)
);

AO31x2_ASAP7_75t_L g1128 ( 
.A1(n_990),
.A2(n_961),
.A3(n_944),
.B(n_1035),
.Y(n_1128)
);

OR2x6_ASAP7_75t_L g1129 ( 
.A(n_999),
.B(n_997),
.Y(n_1129)
);

NOR2xp33_ASAP7_75t_SL g1130 ( 
.A(n_1048),
.B(n_940),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_977),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_940),
.B(n_1041),
.Y(n_1132)
);

O2A1O1Ixp33_ASAP7_75t_L g1133 ( 
.A1(n_940),
.A2(n_1053),
.B(n_1035),
.C(n_1036),
.Y(n_1133)
);

CKINVDCx20_ASAP7_75t_R g1134 ( 
.A(n_936),
.Y(n_1134)
);

INVx1_ASAP7_75t_SL g1135 ( 
.A(n_973),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1136)
);

AOI21xp5_ASAP7_75t_L g1137 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1137)
);

OAI21xp5_ASAP7_75t_L g1138 ( 
.A1(n_940),
.A2(n_1053),
.B(n_1035),
.Y(n_1138)
);

AOI21xp5_ASAP7_75t_L g1139 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1139)
);

AND2x4_ASAP7_75t_L g1140 ( 
.A(n_1047),
.B(n_951),
.Y(n_1140)
);

BUFx10_ASAP7_75t_L g1141 ( 
.A(n_971),
.Y(n_1141)
);

NAND2xp5_ASAP7_75t_L g1142 ( 
.A(n_940),
.B(n_1041),
.Y(n_1142)
);

AOI21xp5_ASAP7_75t_L g1143 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_SL g1144 ( 
.A1(n_961),
.A2(n_944),
.B(n_1035),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_940),
.B(n_1041),
.Y(n_1145)
);

NAND2xp5_ASAP7_75t_L g1146 ( 
.A(n_940),
.B(n_1041),
.Y(n_1146)
);

AOI221x1_ASAP7_75t_L g1147 ( 
.A1(n_940),
.A2(n_1036),
.B1(n_1048),
.B2(n_1053),
.C(n_1035),
.Y(n_1147)
);

AO31x2_ASAP7_75t_L g1148 ( 
.A1(n_961),
.A2(n_944),
.A3(n_1053),
.B(n_1035),
.Y(n_1148)
);

AOI21xp5_ASAP7_75t_L g1149 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1149)
);

OA21x2_ASAP7_75t_L g1150 ( 
.A1(n_962),
.A2(n_1011),
.B(n_1018),
.Y(n_1150)
);

OAI21xp33_ASAP7_75t_L g1151 ( 
.A1(n_940),
.A2(n_810),
.B(n_939),
.Y(n_1151)
);

AOI21x1_ASAP7_75t_L g1152 ( 
.A1(n_1038),
.A2(n_945),
.B(n_996),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1153)
);

OAI21x1_ASAP7_75t_L g1154 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_L g1155 ( 
.A(n_940),
.B(n_971),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_977),
.Y(n_1156)
);

OAI21xp5_ASAP7_75t_L g1157 ( 
.A1(n_940),
.A2(n_1053),
.B(n_1035),
.Y(n_1157)
);

OR2x2_ASAP7_75t_L g1158 ( 
.A(n_1060),
.B(n_614),
.Y(n_1158)
);

NAND2xp5_ASAP7_75t_L g1159 ( 
.A(n_940),
.B(n_1041),
.Y(n_1159)
);

OAI21x1_ASAP7_75t_L g1160 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1160)
);

INVx1_ASAP7_75t_L g1161 ( 
.A(n_977),
.Y(n_1161)
);

OAI21x1_ASAP7_75t_L g1162 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1162)
);

INVx1_ASAP7_75t_L g1163 ( 
.A(n_977),
.Y(n_1163)
);

AOI22xp5_ASAP7_75t_L g1164 ( 
.A1(n_940),
.A2(n_1036),
.B1(n_1048),
.B2(n_939),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_940),
.B(n_1041),
.Y(n_1165)
);

OAI21xp5_ASAP7_75t_L g1166 ( 
.A1(n_940),
.A2(n_1053),
.B(n_1035),
.Y(n_1166)
);

AOI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1168)
);

AOI221xp5_ASAP7_75t_L g1169 ( 
.A1(n_940),
.A2(n_810),
.B1(n_1036),
.B2(n_939),
.C(n_1048),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_977),
.Y(n_1171)
);

BUFx4_ASAP7_75t_SL g1172 ( 
.A(n_1050),
.Y(n_1172)
);

OAI21x1_ASAP7_75t_L g1173 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1173)
);

INVx4_ASAP7_75t_L g1174 ( 
.A(n_964),
.Y(n_1174)
);

OAI22x1_ASAP7_75t_L g1175 ( 
.A1(n_1048),
.A2(n_851),
.B1(n_940),
.B2(n_987),
.Y(n_1175)
);

INVx1_ASAP7_75t_L g1176 ( 
.A(n_977),
.Y(n_1176)
);

AND2x2_ASAP7_75t_L g1177 ( 
.A(n_1060),
.B(n_932),
.Y(n_1177)
);

A2O1A1Ixp33_ASAP7_75t_L g1178 ( 
.A1(n_940),
.A2(n_1048),
.B(n_1053),
.C(n_1035),
.Y(n_1178)
);

A2O1A1Ixp33_ASAP7_75t_L g1179 ( 
.A1(n_940),
.A2(n_1048),
.B(n_1053),
.C(n_1035),
.Y(n_1179)
);

AO21x2_ASAP7_75t_L g1180 ( 
.A1(n_996),
.A2(n_962),
.B(n_961),
.Y(n_1180)
);

INVx1_ASAP7_75t_SL g1181 ( 
.A(n_973),
.Y(n_1181)
);

AOI21xp5_ASAP7_75t_L g1182 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1182)
);

OAI21x1_ASAP7_75t_L g1183 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1183)
);

AOI21xp5_ASAP7_75t_L g1184 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1184)
);

NOR2xp33_ASAP7_75t_SL g1185 ( 
.A(n_950),
.B(n_812),
.Y(n_1185)
);

INVx4_ASAP7_75t_L g1186 ( 
.A(n_964),
.Y(n_1186)
);

BUFx2_ASAP7_75t_L g1187 ( 
.A(n_973),
.Y(n_1187)
);

OAI21x1_ASAP7_75t_L g1188 ( 
.A1(n_1022),
.A2(n_1010),
.B(n_1025),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1189)
);

AOI21xp33_ASAP7_75t_L g1190 ( 
.A1(n_940),
.A2(n_1048),
.B(n_939),
.Y(n_1190)
);

NAND2xp5_ASAP7_75t_SL g1191 ( 
.A(n_940),
.B(n_971),
.Y(n_1191)
);

AOI21xp5_ASAP7_75t_L g1192 ( 
.A1(n_1034),
.A2(n_760),
.B(n_1037),
.Y(n_1192)
);

INVx1_ASAP7_75t_L g1193 ( 
.A(n_977),
.Y(n_1193)
);

NAND2xp5_ASAP7_75t_L g1194 ( 
.A(n_940),
.B(n_1041),
.Y(n_1194)
);

BUFx12f_ASAP7_75t_L g1195 ( 
.A(n_1093),
.Y(n_1195)
);

BUFx2_ASAP7_75t_L g1196 ( 
.A(n_1065),
.Y(n_1196)
);

AOI22xp33_ASAP7_75t_SL g1197 ( 
.A1(n_1155),
.A2(n_1071),
.B1(n_1130),
.B2(n_1157),
.Y(n_1197)
);

INVx1_ASAP7_75t_L g1198 ( 
.A(n_1110),
.Y(n_1198)
);

OAI22xp33_ASAP7_75t_L g1199 ( 
.A1(n_1130),
.A2(n_1194),
.B1(n_1165),
.B2(n_1064),
.Y(n_1199)
);

OAI22xp5_ASAP7_75t_L g1200 ( 
.A1(n_1077),
.A2(n_1146),
.B1(n_1145),
.B2(n_1132),
.Y(n_1200)
);

AOI22xp33_ASAP7_75t_SL g1201 ( 
.A1(n_1071),
.A2(n_1166),
.B1(n_1138),
.B2(n_1067),
.Y(n_1201)
);

AOI22xp33_ASAP7_75t_SL g1202 ( 
.A1(n_1087),
.A2(n_1142),
.B1(n_1159),
.B2(n_1141),
.Y(n_1202)
);

BUFx4f_ASAP7_75t_SL g1203 ( 
.A(n_1090),
.Y(n_1203)
);

CKINVDCx11_ASAP7_75t_R g1204 ( 
.A(n_1134),
.Y(n_1204)
);

AOI22xp33_ASAP7_75t_L g1205 ( 
.A1(n_1151),
.A2(n_1169),
.B1(n_1066),
.B2(n_1175),
.Y(n_1205)
);

INVx1_ASAP7_75t_SL g1206 ( 
.A(n_1135),
.Y(n_1206)
);

OAI22xp33_ASAP7_75t_L g1207 ( 
.A1(n_1164),
.A2(n_1069),
.B1(n_1147),
.B2(n_1091),
.Y(n_1207)
);

BUFx10_ASAP7_75t_L g1208 ( 
.A(n_1072),
.Y(n_1208)
);

INVx1_ASAP7_75t_SL g1209 ( 
.A(n_1181),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_1120),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_L g1211 ( 
.A1(n_1151),
.A2(n_1190),
.B1(n_1191),
.B2(n_1102),
.Y(n_1211)
);

CKINVDCx11_ASAP7_75t_R g1212 ( 
.A(n_1141),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_1122),
.Y(n_1213)
);

NAND2xp5_ASAP7_75t_L g1214 ( 
.A(n_1131),
.B(n_1156),
.Y(n_1214)
);

INVx4_ASAP7_75t_L g1215 ( 
.A(n_1074),
.Y(n_1215)
);

AOI22xp33_ASAP7_75t_SL g1216 ( 
.A1(n_1177),
.A2(n_1092),
.B1(n_1163),
.B2(n_1193),
.Y(n_1216)
);

AOI22xp33_ASAP7_75t_L g1217 ( 
.A1(n_1164),
.A2(n_1069),
.B1(n_1158),
.B2(n_1100),
.Y(n_1217)
);

HB1xp67_ASAP7_75t_L g1218 ( 
.A(n_1128),
.Y(n_1218)
);

INVx5_ASAP7_75t_L g1219 ( 
.A(n_1121),
.Y(n_1219)
);

INVx3_ASAP7_75t_L g1220 ( 
.A(n_1121),
.Y(n_1220)
);

OAI22xp33_ASAP7_75t_L g1221 ( 
.A1(n_1161),
.A2(n_1171),
.B1(n_1176),
.B2(n_1094),
.Y(n_1221)
);

BUFx2_ASAP7_75t_L g1222 ( 
.A(n_1187),
.Y(n_1222)
);

AOI22xp33_ASAP7_75t_L g1223 ( 
.A1(n_1111),
.A2(n_1085),
.B1(n_1150),
.B2(n_1109),
.Y(n_1223)
);

CKINVDCx20_ASAP7_75t_R g1224 ( 
.A(n_1070),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_1123),
.Y(n_1225)
);

INVx1_ASAP7_75t_L g1226 ( 
.A(n_1097),
.Y(n_1226)
);

OAI22xp5_ASAP7_75t_L g1227 ( 
.A1(n_1178),
.A2(n_1179),
.B1(n_1075),
.B2(n_1068),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_1172),
.Y(n_1228)
);

CKINVDCx11_ASAP7_75t_R g1229 ( 
.A(n_1082),
.Y(n_1229)
);

OAI22x1_ASAP7_75t_L g1230 ( 
.A1(n_1140),
.A2(n_1079),
.B1(n_1073),
.B2(n_1103),
.Y(n_1230)
);

BUFx3_ASAP7_75t_L g1231 ( 
.A(n_1086),
.Y(n_1231)
);

BUFx3_ASAP7_75t_L g1232 ( 
.A(n_1084),
.Y(n_1232)
);

INVx4_ASAP7_75t_L g1233 ( 
.A(n_1174),
.Y(n_1233)
);

INVx2_ASAP7_75t_L g1234 ( 
.A(n_1116),
.Y(n_1234)
);

INVx2_ASAP7_75t_L g1235 ( 
.A(n_1128),
.Y(n_1235)
);

AOI22xp33_ASAP7_75t_SL g1236 ( 
.A1(n_1185),
.A2(n_1144),
.B1(n_1150),
.B2(n_1133),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1089),
.B(n_1148),
.Y(n_1237)
);

INVx5_ASAP7_75t_L g1238 ( 
.A(n_1121),
.Y(n_1238)
);

INVx6_ASAP7_75t_L g1239 ( 
.A(n_1174),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1070),
.Y(n_1240)
);

OAI21xp33_ASAP7_75t_L g1241 ( 
.A1(n_1114),
.A2(n_1112),
.B(n_1113),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1186),
.Y(n_1242)
);

INVx1_ASAP7_75t_SL g1243 ( 
.A(n_1129),
.Y(n_1243)
);

AOI22xp33_ASAP7_75t_L g1244 ( 
.A1(n_1180),
.A2(n_1104),
.B1(n_1119),
.B2(n_1117),
.Y(n_1244)
);

INVx1_ASAP7_75t_SL g1245 ( 
.A(n_1108),
.Y(n_1245)
);

INVxp67_ASAP7_75t_SL g1246 ( 
.A(n_1118),
.Y(n_1246)
);

NAND2xp5_ASAP7_75t_L g1247 ( 
.A(n_1148),
.B(n_1088),
.Y(n_1247)
);

INVx2_ASAP7_75t_L g1248 ( 
.A(n_1063),
.Y(n_1248)
);

AOI22xp5_ASAP7_75t_L g1249 ( 
.A1(n_1186),
.A2(n_1126),
.B1(n_1124),
.B2(n_1121),
.Y(n_1249)
);

AOI22xp33_ASAP7_75t_L g1250 ( 
.A1(n_1180),
.A2(n_1137),
.B1(n_1192),
.B2(n_1143),
.Y(n_1250)
);

AOI22xp33_ASAP7_75t_L g1251 ( 
.A1(n_1139),
.A2(n_1149),
.B1(n_1168),
.B2(n_1170),
.Y(n_1251)
);

BUFx12f_ASAP7_75t_L g1252 ( 
.A(n_1127),
.Y(n_1252)
);

AOI22xp33_ASAP7_75t_SL g1253 ( 
.A1(n_1081),
.A2(n_1148),
.B1(n_1153),
.B2(n_1167),
.Y(n_1253)
);

AOI22xp33_ASAP7_75t_SL g1254 ( 
.A1(n_1081),
.A2(n_1182),
.B1(n_1184),
.B2(n_1189),
.Y(n_1254)
);

AOI22xp33_ASAP7_75t_SL g1255 ( 
.A1(n_1081),
.A2(n_1106),
.B1(n_1105),
.B2(n_1188),
.Y(n_1255)
);

INVx4_ASAP7_75t_L g1256 ( 
.A(n_1125),
.Y(n_1256)
);

AOI22xp33_ASAP7_75t_L g1257 ( 
.A1(n_1076),
.A2(n_1078),
.B1(n_1083),
.B2(n_1183),
.Y(n_1257)
);

OAI22xp5_ASAP7_75t_L g1258 ( 
.A1(n_1115),
.A2(n_1095),
.B1(n_1152),
.B2(n_1101),
.Y(n_1258)
);

INVx4_ASAP7_75t_L g1259 ( 
.A(n_1107),
.Y(n_1259)
);

AOI22xp33_ASAP7_75t_L g1260 ( 
.A1(n_1136),
.A2(n_1173),
.B1(n_1162),
.B2(n_1160),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1154),
.A2(n_1080),
.B1(n_1096),
.B2(n_1098),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1080),
.A2(n_1096),
.B1(n_1098),
.B2(n_1099),
.Y(n_1262)
);

INVx4_ASAP7_75t_L g1263 ( 
.A(n_1099),
.Y(n_1263)
);

NAND2xp5_ASAP7_75t_L g1264 ( 
.A(n_1080),
.B(n_1096),
.Y(n_1264)
);

CKINVDCx20_ASAP7_75t_R g1265 ( 
.A(n_1098),
.Y(n_1265)
);

AOI22xp33_ASAP7_75t_SL g1266 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_939),
.B2(n_1048),
.Y(n_1266)
);

NAND2xp5_ASAP7_75t_L g1267 ( 
.A(n_1155),
.B(n_1064),
.Y(n_1267)
);

CKINVDCx20_ASAP7_75t_R g1268 ( 
.A(n_1090),
.Y(n_1268)
);

AOI22xp33_ASAP7_75t_SL g1269 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_939),
.B2(n_1048),
.Y(n_1269)
);

BUFx12f_ASAP7_75t_L g1270 ( 
.A(n_1093),
.Y(n_1270)
);

INVx1_ASAP7_75t_SL g1271 ( 
.A(n_1135),
.Y(n_1271)
);

OAI21xp5_ASAP7_75t_SL g1272 ( 
.A1(n_1155),
.A2(n_940),
.B(n_1036),
.Y(n_1272)
);

INVx4_ASAP7_75t_L g1273 ( 
.A(n_1093),
.Y(n_1273)
);

CKINVDCx6p67_ASAP7_75t_R g1274 ( 
.A(n_1093),
.Y(n_1274)
);

CKINVDCx11_ASAP7_75t_R g1275 ( 
.A(n_1090),
.Y(n_1275)
);

BUFx12f_ASAP7_75t_L g1276 ( 
.A(n_1093),
.Y(n_1276)
);

BUFx6f_ASAP7_75t_L g1277 ( 
.A(n_1093),
.Y(n_1277)
);

AOI22xp5_ASAP7_75t_L g1278 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_1036),
.B2(n_591),
.Y(n_1278)
);

AOI22xp33_ASAP7_75t_L g1279 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_1036),
.B2(n_1048),
.Y(n_1279)
);

BUFx12f_ASAP7_75t_L g1280 ( 
.A(n_1093),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_1110),
.Y(n_1281)
);

AND2x2_ASAP7_75t_L g1282 ( 
.A(n_1177),
.B(n_1155),
.Y(n_1282)
);

INVx1_ASAP7_75t_L g1283 ( 
.A(n_1110),
.Y(n_1283)
);

AOI22xp33_ASAP7_75t_L g1284 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_1036),
.B2(n_1048),
.Y(n_1284)
);

AOI22xp33_ASAP7_75t_L g1285 ( 
.A1(n_1169),
.A2(n_1036),
.B1(n_940),
.B2(n_1048),
.Y(n_1285)
);

CKINVDCx20_ASAP7_75t_R g1286 ( 
.A(n_1090),
.Y(n_1286)
);

AOI22xp33_ASAP7_75t_L g1287 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_1036),
.B2(n_1048),
.Y(n_1287)
);

BUFx12f_ASAP7_75t_L g1288 ( 
.A(n_1093),
.Y(n_1288)
);

BUFx4f_ASAP7_75t_SL g1289 ( 
.A(n_1090),
.Y(n_1289)
);

OAI22x1_ASAP7_75t_L g1290 ( 
.A1(n_1155),
.A2(n_1164),
.B1(n_1069),
.B2(n_1048),
.Y(n_1290)
);

BUFx3_ASAP7_75t_L g1291 ( 
.A(n_1093),
.Y(n_1291)
);

INVx2_ASAP7_75t_SL g1292 ( 
.A(n_1172),
.Y(n_1292)
);

INVx2_ASAP7_75t_SL g1293 ( 
.A(n_1172),
.Y(n_1293)
);

BUFx2_ASAP7_75t_L g1294 ( 
.A(n_1065),
.Y(n_1294)
);

INVx2_ASAP7_75t_SL g1295 ( 
.A(n_1172),
.Y(n_1295)
);

INVx1_ASAP7_75t_SL g1296 ( 
.A(n_1135),
.Y(n_1296)
);

AOI22xp5_ASAP7_75t_L g1297 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_1036),
.B2(n_591),
.Y(n_1297)
);

AOI22xp5_ASAP7_75t_L g1298 ( 
.A1(n_1155),
.A2(n_940),
.B1(n_1036),
.B2(n_591),
.Y(n_1298)
);

HB1xp67_ASAP7_75t_L g1299 ( 
.A(n_1128),
.Y(n_1299)
);

BUFx10_ASAP7_75t_L g1300 ( 
.A(n_1072),
.Y(n_1300)
);

OAI21xp5_ASAP7_75t_SL g1301 ( 
.A1(n_1155),
.A2(n_940),
.B(n_1036),
.Y(n_1301)
);

BUFx4f_ASAP7_75t_SL g1302 ( 
.A(n_1090),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_1225),
.Y(n_1303)
);

OAI21x1_ASAP7_75t_L g1304 ( 
.A1(n_1250),
.A2(n_1258),
.B(n_1257),
.Y(n_1304)
);

BUFx6f_ASAP7_75t_SL g1305 ( 
.A(n_1208),
.Y(n_1305)
);

OAI21x1_ASAP7_75t_L g1306 ( 
.A1(n_1250),
.A2(n_1257),
.B(n_1251),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_1218),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1218),
.Y(n_1308)
);

INVx1_ASAP7_75t_L g1309 ( 
.A(n_1299),
.Y(n_1309)
);

OR2x2_ASAP7_75t_L g1310 ( 
.A(n_1264),
.B(n_1237),
.Y(n_1310)
);

AND2x2_ASAP7_75t_L g1311 ( 
.A(n_1201),
.B(n_1299),
.Y(n_1311)
);

AND2x2_ASAP7_75t_L g1312 ( 
.A(n_1201),
.B(n_1259),
.Y(n_1312)
);

NAND2xp5_ASAP7_75t_L g1313 ( 
.A(n_1200),
.B(n_1199),
.Y(n_1313)
);

OA21x2_ASAP7_75t_L g1314 ( 
.A1(n_1251),
.A2(n_1246),
.B(n_1223),
.Y(n_1314)
);

AND2x2_ASAP7_75t_L g1315 ( 
.A(n_1259),
.B(n_1235),
.Y(n_1315)
);

AO21x2_ASAP7_75t_L g1316 ( 
.A1(n_1241),
.A2(n_1247),
.B(n_1207),
.Y(n_1316)
);

INVx1_ASAP7_75t_L g1317 ( 
.A(n_1265),
.Y(n_1317)
);

INVx1_ASAP7_75t_SL g1318 ( 
.A(n_1245),
.Y(n_1318)
);

OA21x2_ASAP7_75t_L g1319 ( 
.A1(n_1223),
.A2(n_1261),
.B(n_1262),
.Y(n_1319)
);

HB1xp67_ASAP7_75t_L g1320 ( 
.A(n_1226),
.Y(n_1320)
);

AND2x4_ASAP7_75t_L g1321 ( 
.A(n_1234),
.B(n_1263),
.Y(n_1321)
);

OA21x2_ASAP7_75t_L g1322 ( 
.A1(n_1261),
.A2(n_1262),
.B(n_1244),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_1210),
.Y(n_1323)
);

AND2x2_ASAP7_75t_L g1324 ( 
.A(n_1205),
.B(n_1290),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1213),
.Y(n_1325)
);

OAI21x1_ASAP7_75t_L g1326 ( 
.A1(n_1260),
.A2(n_1244),
.B(n_1227),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1221),
.Y(n_1327)
);

HB1xp67_ASAP7_75t_L g1328 ( 
.A(n_1230),
.Y(n_1328)
);

BUFx4f_ASAP7_75t_SL g1329 ( 
.A(n_1195),
.Y(n_1329)
);

INVx4_ASAP7_75t_L g1330 ( 
.A(n_1219),
.Y(n_1330)
);

INVx1_ASAP7_75t_L g1331 ( 
.A(n_1221),
.Y(n_1331)
);

HB1xp67_ASAP7_75t_L g1332 ( 
.A(n_1196),
.Y(n_1332)
);

INVx1_ASAP7_75t_L g1333 ( 
.A(n_1255),
.Y(n_1333)
);

CKINVDCx5p33_ASAP7_75t_R g1334 ( 
.A(n_1275),
.Y(n_1334)
);

HB1xp67_ASAP7_75t_L g1335 ( 
.A(n_1222),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1255),
.Y(n_1336)
);

AND2x4_ASAP7_75t_L g1337 ( 
.A(n_1219),
.B(n_1238),
.Y(n_1337)
);

INVxp67_ASAP7_75t_L g1338 ( 
.A(n_1282),
.Y(n_1338)
);

AND2x2_ASAP7_75t_L g1339 ( 
.A(n_1205),
.B(n_1217),
.Y(n_1339)
);

INVx1_ASAP7_75t_L g1340 ( 
.A(n_1253),
.Y(n_1340)
);

AND2x2_ASAP7_75t_L g1341 ( 
.A(n_1217),
.B(n_1216),
.Y(n_1341)
);

INVx1_ASAP7_75t_L g1342 ( 
.A(n_1254),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1199),
.B(n_1266),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1254),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1198),
.Y(n_1345)
);

INVx1_ASAP7_75t_L g1346 ( 
.A(n_1281),
.Y(n_1346)
);

INVx1_ASAP7_75t_L g1347 ( 
.A(n_1283),
.Y(n_1347)
);

INVx6_ASAP7_75t_L g1348 ( 
.A(n_1219),
.Y(n_1348)
);

AND2x2_ASAP7_75t_L g1349 ( 
.A(n_1216),
.B(n_1197),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1207),
.Y(n_1350)
);

AND2x2_ASAP7_75t_L g1351 ( 
.A(n_1197),
.B(n_1202),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1260),
.Y(n_1352)
);

AOI21x1_ASAP7_75t_L g1353 ( 
.A1(n_1214),
.A2(n_1248),
.B(n_1267),
.Y(n_1353)
);

BUFx3_ASAP7_75t_L g1354 ( 
.A(n_1252),
.Y(n_1354)
);

INVx1_ASAP7_75t_L g1355 ( 
.A(n_1236),
.Y(n_1355)
);

HB1xp67_ASAP7_75t_L g1356 ( 
.A(n_1294),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1202),
.B(n_1236),
.Y(n_1357)
);

INVx2_ASAP7_75t_L g1358 ( 
.A(n_1256),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1211),
.Y(n_1359)
);

OAI21x1_ASAP7_75t_L g1360 ( 
.A1(n_1211),
.A2(n_1285),
.B(n_1220),
.Y(n_1360)
);

NOR2x1_ASAP7_75t_SL g1361 ( 
.A(n_1238),
.B(n_1256),
.Y(n_1361)
);

NAND2xp5_ASAP7_75t_L g1362 ( 
.A(n_1266),
.B(n_1269),
.Y(n_1362)
);

AND2x2_ASAP7_75t_L g1363 ( 
.A(n_1269),
.B(n_1284),
.Y(n_1363)
);

INVx1_ASAP7_75t_L g1364 ( 
.A(n_1272),
.Y(n_1364)
);

AO21x2_ASAP7_75t_L g1365 ( 
.A1(n_1301),
.A2(n_1298),
.B(n_1278),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1249),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1297),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1279),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1279),
.Y(n_1369)
);

AND2x2_ASAP7_75t_L g1370 ( 
.A(n_1284),
.B(n_1287),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1287),
.Y(n_1371)
);

BUFx3_ASAP7_75t_L g1372 ( 
.A(n_1208),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1204),
.Y(n_1373)
);

OR2x2_ASAP7_75t_L g1374 ( 
.A(n_1206),
.B(n_1296),
.Y(n_1374)
);

OAI21xp5_ASAP7_75t_L g1375 ( 
.A1(n_1243),
.A2(n_1271),
.B(n_1209),
.Y(n_1375)
);

BUFx2_ASAP7_75t_SL g1376 ( 
.A(n_1242),
.Y(n_1376)
);

INVxp67_ASAP7_75t_L g1377 ( 
.A(n_1332),
.Y(n_1377)
);

AND2x2_ASAP7_75t_L g1378 ( 
.A(n_1317),
.B(n_1231),
.Y(n_1378)
);

INVxp67_ASAP7_75t_L g1379 ( 
.A(n_1335),
.Y(n_1379)
);

INVx2_ASAP7_75t_L g1380 ( 
.A(n_1323),
.Y(n_1380)
);

NAND2xp5_ASAP7_75t_L g1381 ( 
.A(n_1318),
.B(n_1300),
.Y(n_1381)
);

OR2x2_ASAP7_75t_L g1382 ( 
.A(n_1317),
.B(n_1273),
.Y(n_1382)
);

AND2x2_ASAP7_75t_L g1383 ( 
.A(n_1340),
.B(n_1300),
.Y(n_1383)
);

OAI21x1_ASAP7_75t_SL g1384 ( 
.A1(n_1361),
.A2(n_1273),
.B(n_1233),
.Y(n_1384)
);

OR2x2_ASAP7_75t_L g1385 ( 
.A(n_1310),
.B(n_1291),
.Y(n_1385)
);

BUFx5_ASAP7_75t_L g1386 ( 
.A(n_1352),
.Y(n_1386)
);

A2O1A1Ixp33_ASAP7_75t_L g1387 ( 
.A1(n_1351),
.A2(n_1277),
.B(n_1232),
.C(n_1292),
.Y(n_1387)
);

OAI21xp5_ASAP7_75t_L g1388 ( 
.A1(n_1370),
.A2(n_1215),
.B(n_1286),
.Y(n_1388)
);

AOI22xp5_ASAP7_75t_L g1389 ( 
.A1(n_1339),
.A2(n_1212),
.B1(n_1274),
.B2(n_1224),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1333),
.B(n_1277),
.Y(n_1390)
);

OA21x2_ASAP7_75t_L g1391 ( 
.A1(n_1304),
.A2(n_1295),
.B(n_1293),
.Y(n_1391)
);

AO32x2_ASAP7_75t_L g1392 ( 
.A1(n_1330),
.A2(n_1229),
.A3(n_1239),
.B1(n_1270),
.B2(n_1288),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1334),
.Y(n_1393)
);

AND2x4_ASAP7_75t_L g1394 ( 
.A(n_1321),
.B(n_1240),
.Y(n_1394)
);

AOI22xp33_ASAP7_75t_L g1395 ( 
.A1(n_1339),
.A2(n_1363),
.B1(n_1351),
.B2(n_1324),
.Y(n_1395)
);

OAI22xp5_ASAP7_75t_L g1396 ( 
.A1(n_1364),
.A2(n_1239),
.B1(n_1228),
.B2(n_1276),
.Y(n_1396)
);

AND2x2_ASAP7_75t_L g1397 ( 
.A(n_1328),
.B(n_1280),
.Y(n_1397)
);

BUFx2_ASAP7_75t_L g1398 ( 
.A(n_1372),
.Y(n_1398)
);

OAI221xp5_ASAP7_75t_L g1399 ( 
.A1(n_1364),
.A2(n_1203),
.B1(n_1289),
.B2(n_1302),
.C(n_1268),
.Y(n_1399)
);

AND2x2_ASAP7_75t_L g1400 ( 
.A(n_1338),
.B(n_1203),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1318),
.B(n_1289),
.Y(n_1401)
);

OAI22xp5_ASAP7_75t_L g1402 ( 
.A1(n_1362),
.A2(n_1302),
.B1(n_1349),
.B2(n_1359),
.Y(n_1402)
);

OAI21xp5_ASAP7_75t_L g1403 ( 
.A1(n_1343),
.A2(n_1362),
.B(n_1363),
.Y(n_1403)
);

OAI21xp5_ASAP7_75t_L g1404 ( 
.A1(n_1343),
.A2(n_1313),
.B(n_1324),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_SL g1405 ( 
.A1(n_1361),
.A2(n_1313),
.B(n_1353),
.Y(n_1405)
);

INVx1_ASAP7_75t_L g1406 ( 
.A(n_1325),
.Y(n_1406)
);

INVx2_ASAP7_75t_L g1407 ( 
.A(n_1303),
.Y(n_1407)
);

OAI21x1_ASAP7_75t_L g1408 ( 
.A1(n_1304),
.A2(n_1306),
.B(n_1326),
.Y(n_1408)
);

AND2x2_ASAP7_75t_L g1409 ( 
.A(n_1312),
.B(n_1320),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_L g1410 ( 
.A(n_1367),
.B(n_1368),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1336),
.B(n_1342),
.Y(n_1411)
);

BUFx3_ASAP7_75t_L g1412 ( 
.A(n_1372),
.Y(n_1412)
);

AND2x2_ASAP7_75t_L g1413 ( 
.A(n_1336),
.B(n_1342),
.Y(n_1413)
);

A2O1A1Ixp33_ASAP7_75t_L g1414 ( 
.A1(n_1357),
.A2(n_1349),
.B(n_1341),
.C(n_1312),
.Y(n_1414)
);

INVx5_ASAP7_75t_L g1415 ( 
.A(n_1348),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1304),
.A2(n_1306),
.B(n_1352),
.Y(n_1416)
);

AOI22xp5_ASAP7_75t_L g1417 ( 
.A1(n_1367),
.A2(n_1365),
.B1(n_1341),
.B2(n_1369),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1368),
.B(n_1369),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1344),
.B(n_1311),
.Y(n_1419)
);

OR2x2_ASAP7_75t_L g1420 ( 
.A(n_1310),
.B(n_1344),
.Y(n_1420)
);

BUFx3_ASAP7_75t_L g1421 ( 
.A(n_1372),
.Y(n_1421)
);

A2O1A1Ixp33_ASAP7_75t_L g1422 ( 
.A1(n_1357),
.A2(n_1360),
.B(n_1355),
.C(n_1359),
.Y(n_1422)
);

BUFx12f_ASAP7_75t_L g1423 ( 
.A(n_1373),
.Y(n_1423)
);

NAND2x1p5_ASAP7_75t_L g1424 ( 
.A(n_1330),
.B(n_1337),
.Y(n_1424)
);

NOR2x1_ASAP7_75t_SL g1425 ( 
.A(n_1353),
.B(n_1316),
.Y(n_1425)
);

OAI21xp33_ASAP7_75t_L g1426 ( 
.A1(n_1371),
.A2(n_1350),
.B(n_1366),
.Y(n_1426)
);

OAI22xp5_ASAP7_75t_L g1427 ( 
.A1(n_1354),
.A2(n_1371),
.B1(n_1366),
.B2(n_1350),
.Y(n_1427)
);

AND2x2_ASAP7_75t_L g1428 ( 
.A(n_1311),
.B(n_1315),
.Y(n_1428)
);

AO32x2_ASAP7_75t_L g1429 ( 
.A1(n_1330),
.A2(n_1316),
.A3(n_1308),
.B1(n_1309),
.B2(n_1307),
.Y(n_1429)
);

OR2x2_ASAP7_75t_L g1430 ( 
.A(n_1345),
.B(n_1346),
.Y(n_1430)
);

OAI21xp5_ASAP7_75t_L g1431 ( 
.A1(n_1360),
.A2(n_1326),
.B(n_1375),
.Y(n_1431)
);

AND2x2_ASAP7_75t_L g1432 ( 
.A(n_1365),
.B(n_1356),
.Y(n_1432)
);

AND2x2_ASAP7_75t_L g1433 ( 
.A(n_1365),
.B(n_1345),
.Y(n_1433)
);

NAND4xp25_ASAP7_75t_L g1434 ( 
.A(n_1375),
.B(n_1327),
.C(n_1331),
.D(n_1374),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1407),
.Y(n_1435)
);

AND2x2_ASAP7_75t_L g1436 ( 
.A(n_1416),
.B(n_1322),
.Y(n_1436)
);

NOR2xp33_ASAP7_75t_L g1437 ( 
.A(n_1434),
.B(n_1365),
.Y(n_1437)
);

BUFx2_ASAP7_75t_L g1438 ( 
.A(n_1391),
.Y(n_1438)
);

OR2x2_ASAP7_75t_L g1439 ( 
.A(n_1416),
.B(n_1433),
.Y(n_1439)
);

INVxp67_ASAP7_75t_SL g1440 ( 
.A(n_1425),
.Y(n_1440)
);

HB1xp67_ASAP7_75t_L g1441 ( 
.A(n_1391),
.Y(n_1441)
);

INVx2_ASAP7_75t_L g1442 ( 
.A(n_1380),
.Y(n_1442)
);

OAI22xp5_ASAP7_75t_L g1443 ( 
.A1(n_1414),
.A2(n_1355),
.B1(n_1331),
.B2(n_1327),
.Y(n_1443)
);

OR2x2_ASAP7_75t_L g1444 ( 
.A(n_1420),
.B(n_1432),
.Y(n_1444)
);

AOI22xp33_ASAP7_75t_L g1445 ( 
.A1(n_1403),
.A2(n_1404),
.B1(n_1402),
.B2(n_1395),
.Y(n_1445)
);

NAND2xp5_ASAP7_75t_L g1446 ( 
.A(n_1411),
.B(n_1316),
.Y(n_1446)
);

AND2x2_ASAP7_75t_L g1447 ( 
.A(n_1408),
.B(n_1429),
.Y(n_1447)
);

OAI22xp5_ASAP7_75t_SL g1448 ( 
.A1(n_1395),
.A2(n_1314),
.B1(n_1358),
.B2(n_1376),
.Y(n_1448)
);

INVx2_ASAP7_75t_L g1449 ( 
.A(n_1406),
.Y(n_1449)
);

OAI22xp5_ASAP7_75t_L g1450 ( 
.A1(n_1414),
.A2(n_1358),
.B1(n_1374),
.B2(n_1354),
.Y(n_1450)
);

INVx2_ASAP7_75t_L g1451 ( 
.A(n_1429),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_SL g1452 ( 
.A1(n_1431),
.A2(n_1316),
.B1(n_1360),
.B2(n_1376),
.Y(n_1452)
);

INVx1_ASAP7_75t_L g1453 ( 
.A(n_1430),
.Y(n_1453)
);

NOR2xp67_ASAP7_75t_L g1454 ( 
.A(n_1415),
.B(n_1347),
.Y(n_1454)
);

AOI22xp33_ASAP7_75t_L g1455 ( 
.A1(n_1417),
.A2(n_1354),
.B1(n_1314),
.B2(n_1305),
.Y(n_1455)
);

AND2x2_ASAP7_75t_L g1456 ( 
.A(n_1428),
.B(n_1306),
.Y(n_1456)
);

AND2x2_ASAP7_75t_L g1457 ( 
.A(n_1428),
.B(n_1319),
.Y(n_1457)
);

AND2x2_ASAP7_75t_L g1458 ( 
.A(n_1386),
.B(n_1319),
.Y(n_1458)
);

INVx2_ASAP7_75t_L g1459 ( 
.A(n_1405),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1457),
.B(n_1419),
.Y(n_1460)
);

OR2x6_ASAP7_75t_L g1461 ( 
.A(n_1454),
.B(n_1424),
.Y(n_1461)
);

INVxp67_ASAP7_75t_SL g1462 ( 
.A(n_1441),
.Y(n_1462)
);

BUFx3_ASAP7_75t_L g1463 ( 
.A(n_1438),
.Y(n_1463)
);

INVx1_ASAP7_75t_L g1464 ( 
.A(n_1442),
.Y(n_1464)
);

BUFx2_ASAP7_75t_L g1465 ( 
.A(n_1438),
.Y(n_1465)
);

INVxp67_ASAP7_75t_SL g1466 ( 
.A(n_1441),
.Y(n_1466)
);

AND2x2_ASAP7_75t_L g1467 ( 
.A(n_1457),
.B(n_1419),
.Y(n_1467)
);

AOI221xp5_ASAP7_75t_L g1468 ( 
.A1(n_1443),
.A2(n_1422),
.B1(n_1426),
.B2(n_1427),
.C(n_1379),
.Y(n_1468)
);

OR2x2_ASAP7_75t_L g1469 ( 
.A(n_1439),
.B(n_1409),
.Y(n_1469)
);

INVxp67_ASAP7_75t_L g1470 ( 
.A(n_1437),
.Y(n_1470)
);

OAI31xp33_ASAP7_75t_L g1471 ( 
.A1(n_1450),
.A2(n_1422),
.A3(n_1387),
.B(n_1396),
.Y(n_1471)
);

NAND2xp5_ASAP7_75t_L g1472 ( 
.A(n_1446),
.B(n_1453),
.Y(n_1472)
);

OAI221xp5_ASAP7_75t_SL g1473 ( 
.A1(n_1445),
.A2(n_1387),
.B1(n_1389),
.B2(n_1399),
.C(n_1410),
.Y(n_1473)
);

INVx2_ASAP7_75t_L g1474 ( 
.A(n_1447),
.Y(n_1474)
);

AOI221xp5_ASAP7_75t_L g1475 ( 
.A1(n_1443),
.A2(n_1377),
.B1(n_1418),
.B2(n_1413),
.C(n_1381),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1456),
.B(n_1319),
.Y(n_1476)
);

OAI21xp5_ASAP7_75t_L g1477 ( 
.A1(n_1437),
.A2(n_1388),
.B(n_1326),
.Y(n_1477)
);

AND2x2_ASAP7_75t_L g1478 ( 
.A(n_1456),
.B(n_1319),
.Y(n_1478)
);

INVx2_ASAP7_75t_SL g1479 ( 
.A(n_1449),
.Y(n_1479)
);

OAI22xp5_ASAP7_75t_L g1480 ( 
.A1(n_1445),
.A2(n_1385),
.B1(n_1382),
.B2(n_1390),
.Y(n_1480)
);

AND2x2_ASAP7_75t_L g1481 ( 
.A(n_1456),
.B(n_1383),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_1449),
.Y(n_1482)
);

INVx2_ASAP7_75t_L g1483 ( 
.A(n_1447),
.Y(n_1483)
);

BUFx2_ASAP7_75t_L g1484 ( 
.A(n_1438),
.Y(n_1484)
);

HB1xp67_ASAP7_75t_L g1485 ( 
.A(n_1435),
.Y(n_1485)
);

AND2x2_ASAP7_75t_L g1486 ( 
.A(n_1458),
.B(n_1383),
.Y(n_1486)
);

INVx1_ASAP7_75t_SL g1487 ( 
.A(n_1439),
.Y(n_1487)
);

NOR2xp33_ASAP7_75t_L g1488 ( 
.A(n_1459),
.B(n_1390),
.Y(n_1488)
);

HB1xp67_ASAP7_75t_L g1489 ( 
.A(n_1485),
.Y(n_1489)
);

NAND2xp5_ASAP7_75t_L g1490 ( 
.A(n_1470),
.B(n_1453),
.Y(n_1490)
);

OR2x2_ASAP7_75t_L g1491 ( 
.A(n_1487),
.B(n_1451),
.Y(n_1491)
);

NOR2xp33_ASAP7_75t_L g1492 ( 
.A(n_1473),
.B(n_1397),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1463),
.Y(n_1493)
);

AND2x4_ASAP7_75t_L g1494 ( 
.A(n_1461),
.B(n_1454),
.Y(n_1494)
);

AND2x2_ASAP7_75t_L g1495 ( 
.A(n_1474),
.B(n_1483),
.Y(n_1495)
);

INVx2_ASAP7_75t_L g1496 ( 
.A(n_1479),
.Y(n_1496)
);

INVx2_ASAP7_75t_L g1497 ( 
.A(n_1479),
.Y(n_1497)
);

INVx2_ASAP7_75t_L g1498 ( 
.A(n_1479),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1482),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1482),
.Y(n_1500)
);

OR2x2_ASAP7_75t_L g1501 ( 
.A(n_1487),
.B(n_1451),
.Y(n_1501)
);

INVx1_ASAP7_75t_SL g1502 ( 
.A(n_1465),
.Y(n_1502)
);

NOR2x1_ASAP7_75t_L g1503 ( 
.A(n_1463),
.B(n_1459),
.Y(n_1503)
);

AOI22xp33_ASAP7_75t_L g1504 ( 
.A1(n_1468),
.A2(n_1448),
.B1(n_1450),
.B2(n_1452),
.Y(n_1504)
);

AOI22xp33_ASAP7_75t_L g1505 ( 
.A1(n_1468),
.A2(n_1448),
.B1(n_1452),
.B2(n_1455),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1464),
.Y(n_1506)
);

INVx4_ASAP7_75t_L g1507 ( 
.A(n_1461),
.Y(n_1507)
);

AND2x2_ASAP7_75t_L g1508 ( 
.A(n_1476),
.B(n_1447),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1485),
.Y(n_1509)
);

AND2x2_ASAP7_75t_L g1510 ( 
.A(n_1476),
.B(n_1447),
.Y(n_1510)
);

NAND2xp5_ASAP7_75t_L g1511 ( 
.A(n_1470),
.B(n_1453),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1463),
.Y(n_1512)
);

AND2x2_ASAP7_75t_L g1513 ( 
.A(n_1476),
.B(n_1478),
.Y(n_1513)
);

NOR2xp33_ASAP7_75t_L g1514 ( 
.A(n_1473),
.B(n_1401),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1472),
.B(n_1444),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1507),
.B(n_1460),
.Y(n_1516)
);

INVx2_ASAP7_75t_L g1517 ( 
.A(n_1495),
.Y(n_1517)
);

AND2x2_ASAP7_75t_L g1518 ( 
.A(n_1507),
.B(n_1460),
.Y(n_1518)
);

INVx1_ASAP7_75t_L g1519 ( 
.A(n_1489),
.Y(n_1519)
);

OAI21xp5_ASAP7_75t_L g1520 ( 
.A1(n_1492),
.A2(n_1471),
.B(n_1477),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1507),
.B(n_1460),
.Y(n_1521)
);

INVx1_ASAP7_75t_L g1522 ( 
.A(n_1489),
.Y(n_1522)
);

AND2x2_ASAP7_75t_L g1523 ( 
.A(n_1507),
.B(n_1467),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1495),
.Y(n_1524)
);

A2O1A1Ixp33_ASAP7_75t_L g1525 ( 
.A1(n_1492),
.A2(n_1471),
.B(n_1477),
.C(n_1475),
.Y(n_1525)
);

INVx1_ASAP7_75t_L g1526 ( 
.A(n_1509),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1509),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1499),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1495),
.Y(n_1529)
);

NAND2x1p5_ASAP7_75t_L g1530 ( 
.A(n_1503),
.B(n_1415),
.Y(n_1530)
);

INVx2_ASAP7_75t_SL g1531 ( 
.A(n_1503),
.Y(n_1531)
);

INVx2_ASAP7_75t_L g1532 ( 
.A(n_1496),
.Y(n_1532)
);

AND2x4_ASAP7_75t_L g1533 ( 
.A(n_1507),
.B(n_1463),
.Y(n_1533)
);

INVx2_ASAP7_75t_L g1534 ( 
.A(n_1496),
.Y(n_1534)
);

OR2x2_ASAP7_75t_L g1535 ( 
.A(n_1490),
.B(n_1469),
.Y(n_1535)
);

INVxp67_ASAP7_75t_L g1536 ( 
.A(n_1514),
.Y(n_1536)
);

AOI22xp5_ASAP7_75t_L g1537 ( 
.A1(n_1505),
.A2(n_1448),
.B1(n_1455),
.B2(n_1475),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_L g1538 ( 
.A(n_1490),
.B(n_1467),
.Y(n_1538)
);

INVx1_ASAP7_75t_L g1539 ( 
.A(n_1499),
.Y(n_1539)
);

INVxp67_ASAP7_75t_L g1540 ( 
.A(n_1514),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1496),
.Y(n_1541)
);

INVx2_ASAP7_75t_L g1542 ( 
.A(n_1496),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1513),
.B(n_1508),
.Y(n_1543)
);

OR2x2_ASAP7_75t_L g1544 ( 
.A(n_1511),
.B(n_1469),
.Y(n_1544)
);

NOR2xp33_ASAP7_75t_L g1545 ( 
.A(n_1511),
.B(n_1329),
.Y(n_1545)
);

NAND2xp5_ASAP7_75t_L g1546 ( 
.A(n_1515),
.B(n_1467),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1513),
.B(n_1481),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1499),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1513),
.B(n_1481),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1500),
.Y(n_1550)
);

NAND2xp5_ASAP7_75t_L g1551 ( 
.A(n_1515),
.B(n_1472),
.Y(n_1551)
);

AND2x2_ASAP7_75t_L g1552 ( 
.A(n_1508),
.B(n_1481),
.Y(n_1552)
);

INVx1_ASAP7_75t_L g1553 ( 
.A(n_1500),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1508),
.B(n_1486),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1500),
.Y(n_1555)
);

NAND2x1_ASAP7_75t_L g1556 ( 
.A(n_1493),
.B(n_1465),
.Y(n_1556)
);

INVx2_ASAP7_75t_L g1557 ( 
.A(n_1497),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1543),
.Y(n_1558)
);

AND2x2_ASAP7_75t_L g1559 ( 
.A(n_1543),
.B(n_1512),
.Y(n_1559)
);

NAND2xp5_ASAP7_75t_L g1560 ( 
.A(n_1536),
.B(n_1488),
.Y(n_1560)
);

NAND2xp5_ASAP7_75t_L g1561 ( 
.A(n_1536),
.B(n_1488),
.Y(n_1561)
);

AND2x2_ASAP7_75t_L g1562 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1562)
);

NOR2xp33_ASAP7_75t_L g1563 ( 
.A(n_1540),
.B(n_1423),
.Y(n_1563)
);

NAND2xp5_ASAP7_75t_L g1564 ( 
.A(n_1540),
.B(n_1486),
.Y(n_1564)
);

AND2x2_ASAP7_75t_L g1565 ( 
.A(n_1547),
.B(n_1512),
.Y(n_1565)
);

AOI22xp33_ASAP7_75t_SL g1566 ( 
.A1(n_1520),
.A2(n_1480),
.B1(n_1436),
.B2(n_1458),
.Y(n_1566)
);

AOI21xp5_ASAP7_75t_SL g1567 ( 
.A1(n_1525),
.A2(n_1305),
.B(n_1480),
.Y(n_1567)
);

OR2x2_ASAP7_75t_L g1568 ( 
.A(n_1538),
.B(n_1502),
.Y(n_1568)
);

AND2x2_ASAP7_75t_L g1569 ( 
.A(n_1549),
.B(n_1512),
.Y(n_1569)
);

AND2x2_ASAP7_75t_L g1570 ( 
.A(n_1549),
.B(n_1516),
.Y(n_1570)
);

NOR2xp33_ASAP7_75t_L g1571 ( 
.A(n_1545),
.B(n_1423),
.Y(n_1571)
);

NOR2xp67_ASAP7_75t_L g1572 ( 
.A(n_1531),
.B(n_1493),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1528),
.Y(n_1573)
);

OR2x6_ASAP7_75t_L g1574 ( 
.A(n_1520),
.B(n_1384),
.Y(n_1574)
);

INVx2_ASAP7_75t_SL g1575 ( 
.A(n_1556),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1528),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1516),
.B(n_1494),
.Y(n_1577)
);

AOI221xp5_ASAP7_75t_L g1578 ( 
.A1(n_1537),
.A2(n_1504),
.B1(n_1505),
.B2(n_1484),
.C(n_1465),
.Y(n_1578)
);

NOR2x1p5_ASAP7_75t_L g1579 ( 
.A(n_1556),
.B(n_1393),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1518),
.B(n_1521),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1537),
.B(n_1486),
.Y(n_1581)
);

AND3x2_ASAP7_75t_L g1582 ( 
.A(n_1519),
.B(n_1484),
.C(n_1398),
.Y(n_1582)
);

NAND2x1_ASAP7_75t_L g1583 ( 
.A(n_1531),
.B(n_1493),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1551),
.B(n_1504),
.Y(n_1584)
);

AND2x2_ASAP7_75t_L g1585 ( 
.A(n_1518),
.B(n_1494),
.Y(n_1585)
);

NOR2x1_ASAP7_75t_L g1586 ( 
.A(n_1519),
.B(n_1493),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1551),
.B(n_1469),
.Y(n_1587)
);

AND2x2_ASAP7_75t_L g1588 ( 
.A(n_1521),
.B(n_1494),
.Y(n_1588)
);

INVxp67_ASAP7_75t_L g1589 ( 
.A(n_1522),
.Y(n_1589)
);

OAI31xp33_ASAP7_75t_SL g1590 ( 
.A1(n_1533),
.A2(n_1494),
.A3(n_1502),
.B(n_1462),
.Y(n_1590)
);

INVx1_ASAP7_75t_L g1591 ( 
.A(n_1539),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1538),
.B(n_1478),
.Y(n_1592)
);

OR2x2_ASAP7_75t_L g1593 ( 
.A(n_1560),
.B(n_1561),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1573),
.Y(n_1594)
);

INVxp67_ASAP7_75t_L g1595 ( 
.A(n_1563),
.Y(n_1595)
);

OAI22xp33_ASAP7_75t_L g1596 ( 
.A1(n_1578),
.A2(n_1530),
.B1(n_1531),
.B2(n_1535),
.Y(n_1596)
);

INVxp67_ASAP7_75t_L g1597 ( 
.A(n_1586),
.Y(n_1597)
);

AOI32xp33_ASAP7_75t_L g1598 ( 
.A1(n_1566),
.A2(n_1523),
.A3(n_1533),
.B1(n_1522),
.B2(n_1493),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1573),
.Y(n_1599)
);

AOI221xp5_ASAP7_75t_L g1600 ( 
.A1(n_1584),
.A2(n_1527),
.B1(n_1526),
.B2(n_1533),
.C(n_1523),
.Y(n_1600)
);

INVx1_ASAP7_75t_L g1601 ( 
.A(n_1576),
.Y(n_1601)
);

OAI322xp33_ASAP7_75t_SL g1602 ( 
.A1(n_1581),
.A2(n_1546),
.A3(n_1526),
.B1(n_1527),
.B2(n_1529),
.C1(n_1517),
.C2(n_1524),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1589),
.B(n_1552),
.Y(n_1603)
);

OAI22xp5_ASAP7_75t_L g1604 ( 
.A1(n_1567),
.A2(n_1530),
.B1(n_1439),
.B2(n_1484),
.Y(n_1604)
);

AOI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1567),
.A2(n_1533),
.B1(n_1517),
.B2(n_1529),
.C(n_1524),
.Y(n_1605)
);

INVxp67_ASAP7_75t_SL g1606 ( 
.A(n_1572),
.Y(n_1606)
);

AOI31xp33_ASAP7_75t_L g1607 ( 
.A1(n_1571),
.A2(n_1530),
.A3(n_1393),
.B(n_1394),
.Y(n_1607)
);

AOI221x1_ASAP7_75t_L g1608 ( 
.A1(n_1576),
.A2(n_1548),
.B1(n_1539),
.B2(n_1555),
.C(n_1550),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1591),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1591),
.Y(n_1610)
);

AOI22xp5_ASAP7_75t_L g1611 ( 
.A1(n_1579),
.A2(n_1494),
.B1(n_1436),
.B2(n_1459),
.Y(n_1611)
);

INVx3_ASAP7_75t_L g1612 ( 
.A(n_1583),
.Y(n_1612)
);

INVx1_ASAP7_75t_SL g1613 ( 
.A(n_1582),
.Y(n_1613)
);

AND2x2_ASAP7_75t_L g1614 ( 
.A(n_1580),
.B(n_1554),
.Y(n_1614)
);

INVx1_ASAP7_75t_L g1615 ( 
.A(n_1558),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1564),
.B(n_1552),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1580),
.B(n_1554),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1594),
.Y(n_1618)
);

NOR2xp33_ASAP7_75t_L g1619 ( 
.A(n_1595),
.B(n_1593),
.Y(n_1619)
);

OR2x2_ASAP7_75t_L g1620 ( 
.A(n_1603),
.B(n_1558),
.Y(n_1620)
);

INVxp67_ASAP7_75t_L g1621 ( 
.A(n_1606),
.Y(n_1621)
);

OAI21xp5_ASAP7_75t_L g1622 ( 
.A1(n_1596),
.A2(n_1574),
.B(n_1575),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1613),
.A2(n_1574),
.B1(n_1579),
.B2(n_1575),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1599),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1612),
.Y(n_1625)
);

AOI21xp33_ASAP7_75t_SL g1626 ( 
.A1(n_1607),
.A2(n_1590),
.B(n_1574),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_SL g1627 ( 
.A(n_1604),
.B(n_1568),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1600),
.B(n_1570),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1615),
.B(n_1570),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1601),
.Y(n_1630)
);

INVx1_ASAP7_75t_L g1631 ( 
.A(n_1609),
.Y(n_1631)
);

OAI221xp5_ASAP7_75t_L g1632 ( 
.A1(n_1598),
.A2(n_1574),
.B1(n_1530),
.B2(n_1568),
.C(n_1583),
.Y(n_1632)
);

AOI322xp5_ASAP7_75t_L g1633 ( 
.A1(n_1597),
.A2(n_1510),
.A3(n_1587),
.B1(n_1592),
.B2(n_1559),
.C1(n_1569),
.C2(n_1565),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1614),
.B(n_1559),
.Y(n_1634)
);

NOR3xp33_ASAP7_75t_L g1635 ( 
.A(n_1605),
.B(n_1565),
.C(n_1562),
.Y(n_1635)
);

A2O1A1Ixp33_ASAP7_75t_L g1636 ( 
.A1(n_1604),
.A2(n_1494),
.B(n_1585),
.C(n_1577),
.Y(n_1636)
);

AOI221xp5_ASAP7_75t_L g1637 ( 
.A1(n_1626),
.A2(n_1602),
.B1(n_1603),
.B2(n_1610),
.C(n_1616),
.Y(n_1637)
);

INVx1_ASAP7_75t_SL g1638 ( 
.A(n_1620),
.Y(n_1638)
);

INVx2_ASAP7_75t_L g1639 ( 
.A(n_1625),
.Y(n_1639)
);

AOI222xp33_ASAP7_75t_L g1640 ( 
.A1(n_1627),
.A2(n_1616),
.B1(n_1617),
.B2(n_1612),
.C1(n_1562),
.C2(n_1569),
.Y(n_1640)
);

AOI21xp5_ASAP7_75t_SL g1641 ( 
.A1(n_1619),
.A2(n_1608),
.B(n_1305),
.Y(n_1641)
);

NAND2xp5_ASAP7_75t_L g1642 ( 
.A(n_1621),
.B(n_1577),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1629),
.Y(n_1643)
);

INVxp67_ASAP7_75t_SL g1644 ( 
.A(n_1621),
.Y(n_1644)
);

NAND2xp5_ASAP7_75t_L g1645 ( 
.A(n_1619),
.B(n_1585),
.Y(n_1645)
);

OAI21xp5_ASAP7_75t_SL g1646 ( 
.A1(n_1622),
.A2(n_1611),
.B(n_1588),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1618),
.Y(n_1647)
);

NOR2xp33_ASAP7_75t_L g1648 ( 
.A(n_1645),
.B(n_1623),
.Y(n_1648)
);

NAND4xp25_ASAP7_75t_SL g1649 ( 
.A(n_1637),
.B(n_1628),
.C(n_1632),
.D(n_1635),
.Y(n_1649)
);

NAND2xp5_ASAP7_75t_L g1650 ( 
.A(n_1644),
.B(n_1634),
.Y(n_1650)
);

NAND4xp75_ASAP7_75t_L g1651 ( 
.A(n_1639),
.B(n_1631),
.C(n_1630),
.D(n_1624),
.Y(n_1651)
);

INVx1_ASAP7_75t_L g1652 ( 
.A(n_1644),
.Y(n_1652)
);

OAI21xp33_ASAP7_75t_L g1653 ( 
.A1(n_1646),
.A2(n_1633),
.B(n_1635),
.Y(n_1653)
);

NAND2xp5_ASAP7_75t_SL g1654 ( 
.A(n_1640),
.B(n_1636),
.Y(n_1654)
);

NAND2xp5_ASAP7_75t_L g1655 ( 
.A(n_1638),
.B(n_1588),
.Y(n_1655)
);

INVx1_ASAP7_75t_L g1656 ( 
.A(n_1642),
.Y(n_1656)
);

NAND2xp5_ASAP7_75t_L g1657 ( 
.A(n_1643),
.B(n_1535),
.Y(n_1657)
);

OR3x1_ASAP7_75t_L g1658 ( 
.A(n_1647),
.B(n_1550),
.C(n_1548),
.Y(n_1658)
);

NOR3xp33_ASAP7_75t_L g1659 ( 
.A(n_1649),
.B(n_1641),
.C(n_1400),
.Y(n_1659)
);

NOR2x1_ASAP7_75t_L g1660 ( 
.A(n_1652),
.B(n_1532),
.Y(n_1660)
);

OAI211xp5_ASAP7_75t_SL g1661 ( 
.A1(n_1653),
.A2(n_1544),
.B(n_1546),
.C(n_1534),
.Y(n_1661)
);

OAI221xp5_ASAP7_75t_L g1662 ( 
.A1(n_1654),
.A2(n_1544),
.B1(n_1524),
.B2(n_1529),
.C(n_1517),
.Y(n_1662)
);

AOI221x1_ASAP7_75t_L g1663 ( 
.A1(n_1650),
.A2(n_1553),
.B1(n_1555),
.B2(n_1542),
.C(n_1541),
.Y(n_1663)
);

AOI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1661),
.A2(n_1655),
.B(n_1648),
.Y(n_1664)
);

NAND3xp33_ASAP7_75t_L g1665 ( 
.A(n_1659),
.B(n_1656),
.C(n_1657),
.Y(n_1665)
);

NAND4xp25_ASAP7_75t_L g1666 ( 
.A(n_1660),
.B(n_1651),
.C(n_1658),
.D(n_1394),
.Y(n_1666)
);

O2A1O1Ixp33_ASAP7_75t_L g1667 ( 
.A1(n_1662),
.A2(n_1557),
.B(n_1532),
.C(n_1542),
.Y(n_1667)
);

O2A1O1Ixp5_ASAP7_75t_L g1668 ( 
.A1(n_1663),
.A2(n_1557),
.B(n_1532),
.C(n_1542),
.Y(n_1668)
);

AOI221xp5_ASAP7_75t_L g1669 ( 
.A1(n_1661),
.A2(n_1557),
.B1(n_1541),
.B2(n_1534),
.C(n_1553),
.Y(n_1669)
);

INVx2_ASAP7_75t_L g1670 ( 
.A(n_1668),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_SL g1671 ( 
.A(n_1664),
.B(n_1534),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1666),
.B(n_1541),
.Y(n_1672)
);

XOR2xp5_ASAP7_75t_L g1673 ( 
.A(n_1665),
.B(n_1394),
.Y(n_1673)
);

NOR2xp67_ASAP7_75t_L g1674 ( 
.A(n_1667),
.B(n_1497),
.Y(n_1674)
);

BUFx6f_ASAP7_75t_L g1675 ( 
.A(n_1671),
.Y(n_1675)
);

NOR2xp33_ASAP7_75t_L g1676 ( 
.A(n_1673),
.B(n_1669),
.Y(n_1676)
);

NAND3xp33_ASAP7_75t_L g1677 ( 
.A(n_1670),
.B(n_1672),
.C(n_1674),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1675),
.Y(n_1678)
);

AOI22xp5_ASAP7_75t_L g1679 ( 
.A1(n_1678),
.A2(n_1676),
.B1(n_1677),
.B2(n_1305),
.Y(n_1679)
);

AOI21xp5_ASAP7_75t_L g1680 ( 
.A1(n_1679),
.A2(n_1378),
.B(n_1497),
.Y(n_1680)
);

AO22x2_ASAP7_75t_L g1681 ( 
.A1(n_1680),
.A2(n_1497),
.B1(n_1498),
.B2(n_1501),
.Y(n_1681)
);

OA22x2_ASAP7_75t_L g1682 ( 
.A1(n_1681),
.A2(n_1498),
.B1(n_1466),
.B2(n_1462),
.Y(n_1682)
);

AOI22xp33_ASAP7_75t_L g1683 ( 
.A1(n_1682),
.A2(n_1501),
.B1(n_1491),
.B2(n_1459),
.Y(n_1683)
);

AOI21xp33_ASAP7_75t_SL g1684 ( 
.A1(n_1682),
.A2(n_1392),
.B(n_1491),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1684),
.A2(n_1498),
.B(n_1491),
.Y(n_1685)
);

NAND2xp5_ASAP7_75t_L g1686 ( 
.A(n_1683),
.B(n_1498),
.Y(n_1686)
);

OA21x2_ASAP7_75t_L g1687 ( 
.A1(n_1686),
.A2(n_1685),
.B(n_1506),
.Y(n_1687)
);

OAI221xp5_ASAP7_75t_R g1688 ( 
.A1(n_1687),
.A2(n_1392),
.B1(n_1501),
.B2(n_1466),
.C(n_1440),
.Y(n_1688)
);

AOI211xp5_ASAP7_75t_L g1689 ( 
.A1(n_1688),
.A2(n_1421),
.B(n_1412),
.C(n_1392),
.Y(n_1689)
);


endmodule