module fake_jpeg_15304_n_351 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_351);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_351;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_15;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_13;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_14;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_347;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g13 ( 
.A(n_11),
.Y(n_13)
);

BUFx12f_ASAP7_75t_L g14 ( 
.A(n_3),
.Y(n_14)
);

INVx11_ASAP7_75t_L g15 ( 
.A(n_6),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx16_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx2_ASAP7_75t_SL g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_10),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

BUFx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_11),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_6),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

BUFx24_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_23),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_37),
.Y(n_87)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_38),
.Y(n_109)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_39),
.B(n_41),
.Y(n_76)
);

INVx8_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

INVx5_ASAP7_75t_L g74 ( 
.A(n_40),
.Y(n_74)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_24),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_23),
.Y(n_42)
);

BUFx2_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_21),
.Y(n_43)
);

INVx4_ASAP7_75t_L g81 ( 
.A(n_43),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_23),
.Y(n_44)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_12),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_52),
.Y(n_77)
);

BUFx12_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_46),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g47 ( 
.A(n_28),
.B(n_12),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_47),
.B(n_57),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_34),
.Y(n_48)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_48),
.Y(n_93)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_36),
.Y(n_49)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_26),
.Y(n_50)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_50),
.Y(n_102)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_36),
.Y(n_51)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_24),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_34),
.Y(n_54)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_54),
.Y(n_84)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_13),
.B(n_0),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_58),
.B(n_60),
.Y(n_86)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

INVx4_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_13),
.B(n_22),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_36),
.Y(n_61)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_61),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_22),
.B(n_0),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_63),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g63 ( 
.A(n_14),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g64 ( 
.A(n_16),
.B(n_0),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_64),
.A2(n_66),
.B1(n_33),
.B2(n_2),
.Y(n_96)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_65),
.B(n_67),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_16),
.B(n_1),
.Y(n_66)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_47),
.B(n_35),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_68),
.B(n_89),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_15),
.B1(n_29),
.B2(n_19),
.Y(n_72)
);

AOI21xp5_ASAP7_75t_L g133 ( 
.A1(n_72),
.A2(n_75),
.B(n_80),
.Y(n_133)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_56),
.Y(n_73)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_15),
.B1(n_19),
.B2(n_18),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_58),
.A2(n_25),
.B1(n_32),
.B2(n_35),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_78),
.A2(n_79),
.B1(n_85),
.B2(n_100),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_43),
.A2(n_18),
.B1(n_30),
.B2(n_32),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_59),
.A2(n_25),
.B1(n_30),
.B2(n_33),
.Y(n_80)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_46),
.Y(n_82)
);

INVx1_ASAP7_75t_SL g122 ( 
.A(n_82),
.Y(n_122)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_55),
.A2(n_33),
.B1(n_27),
.B2(n_22),
.Y(n_83)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_83),
.A2(n_107),
.B(n_10),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_27),
.B1(n_17),
.B2(n_33),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_14),
.Y(n_89)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_42),
.Y(n_91)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_63),
.B(n_17),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_94),
.B(n_106),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_96),
.B(n_114),
.Y(n_163)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_61),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_99),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_49),
.A2(n_27),
.B1(n_17),
.B2(n_36),
.Y(n_100)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx5_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx4_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g150 ( 
.A(n_105),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_51),
.B(n_1),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_107)
);

BUFx10_ASAP7_75t_L g108 ( 
.A(n_56),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g157 ( 
.A(n_108),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_46),
.B(n_2),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_110),
.B(n_113),
.Y(n_120)
);

INVx6_ASAP7_75t_L g112 ( 
.A(n_53),
.Y(n_112)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_112),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_37),
.B(n_3),
.Y(n_113)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_44),
.B(n_14),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_48),
.B(n_4),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_115),
.B(n_116),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_54),
.B(n_4),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_87),
.Y(n_118)
);

INVx11_ASAP7_75t_L g187 ( 
.A(n_118),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g123 ( 
.A1(n_74),
.A2(n_14),
.B1(n_6),
.B2(n_7),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_123),
.A2(n_134),
.B1(n_137),
.B2(n_141),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_107),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_126),
.A2(n_144),
.B1(n_152),
.B2(n_153),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_77),
.B(n_5),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_127),
.B(n_145),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_74),
.A2(n_5),
.B1(n_7),
.B2(n_9),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_128),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g129 ( 
.A(n_87),
.Y(n_129)
);

INVx3_ASAP7_75t_L g194 ( 
.A(n_129),
.Y(n_194)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_102),
.Y(n_131)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_131),
.Y(n_176)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_78),
.Y(n_132)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_132),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_81),
.A2(n_10),
.B1(n_101),
.B2(n_109),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_SL g186 ( 
.A(n_135),
.B(n_147),
.C(n_136),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_114),
.B(n_96),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_142),
.Y(n_168)
);

OAI22xp33_ASAP7_75t_L g137 ( 
.A1(n_109),
.A2(n_81),
.B1(n_84),
.B2(n_93),
.Y(n_137)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_92),
.Y(n_140)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g141 ( 
.A1(n_84),
.A2(n_69),
.B1(n_90),
.B2(n_86),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_101),
.B(n_88),
.Y(n_142)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_108),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_143),
.B(n_138),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_90),
.A2(n_72),
.B1(n_95),
.B2(n_99),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_76),
.B(n_97),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_80),
.B(n_71),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_147),
.B(n_151),
.Y(n_191)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_97),
.Y(n_148)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_148),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_71),
.B(n_73),
.Y(n_151)
);

OA22x2_ASAP7_75t_L g152 ( 
.A1(n_98),
.A2(n_117),
.B1(n_83),
.B2(n_104),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_L g153 ( 
.A1(n_95),
.A2(n_112),
.B1(n_91),
.B2(n_75),
.Y(n_153)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_103),
.B(n_70),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_154),
.B(n_134),
.Y(n_172)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_71),
.Y(n_155)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_155),
.Y(n_192)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_73),
.Y(n_158)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_158),
.Y(n_202)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_70),
.Y(n_159)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_105),
.A2(n_111),
.B1(n_103),
.B2(n_82),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g175 ( 
.A(n_160),
.B(n_152),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_SL g161 ( 
.A1(n_111),
.A2(n_47),
.B1(n_64),
.B2(n_66),
.Y(n_161)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_161),
.Y(n_174)
);

INVxp67_ASAP7_75t_L g162 ( 
.A(n_82),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_164),
.Y(n_167)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_77),
.B(n_86),
.Y(n_164)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_169),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g171 ( 
.A(n_151),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_171),
.B(n_172),
.Y(n_214)
);

INVx5_ASAP7_75t_L g173 ( 
.A(n_139),
.Y(n_173)
);

INVx3_ASAP7_75t_L g226 ( 
.A(n_173),
.Y(n_226)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_200),
.B1(n_165),
.B2(n_174),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_131),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g231 ( 
.A(n_177),
.B(n_180),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g180 ( 
.A(n_160),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_155),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_182),
.B(n_190),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_140),
.B(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_183),
.Y(n_224)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_185),
.Y(n_234)
);

A2O1A1Ixp33_ASAP7_75t_SL g210 ( 
.A1(n_186),
.A2(n_133),
.B(n_158),
.C(n_137),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g188 ( 
.A(n_121),
.B(n_120),
.Y(n_188)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_188),
.Y(n_205)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_142),
.B(n_163),
.Y(n_189)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_189),
.Y(n_209)
);

INVx5_ASAP7_75t_L g190 ( 
.A(n_139),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_132),
.B(n_163),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_193),
.B(n_196),
.Y(n_213)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_124),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_195),
.B(n_199),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_146),
.B(n_161),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_146),
.B(n_154),
.Y(n_198)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_198),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_157),
.Y(n_199)
);

AND2x2_ASAP7_75t_L g200 ( 
.A(n_152),
.B(n_125),
.Y(n_200)
);

XOR2x2_ASAP7_75t_SL g221 ( 
.A(n_200),
.B(n_150),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_156),
.B(n_148),
.Y(n_203)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_203),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_135),
.B(n_152),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_SL g228 ( 
.A(n_204),
.B(n_170),
.Y(n_228)
);

INVx13_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g243 ( 
.A(n_207),
.B(n_208),
.Y(n_243)
);

BUFx2_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_210),
.B(n_219),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_192),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_212),
.B(n_230),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g251 ( 
.A1(n_215),
.A2(n_216),
.B1(n_233),
.B2(n_197),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_200),
.A2(n_133),
.B1(n_149),
.B2(n_124),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g217 ( 
.A1(n_170),
.A2(n_149),
.B1(n_130),
.B2(n_143),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_217),
.A2(n_220),
.B1(n_194),
.B2(n_202),
.Y(n_260)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_171),
.B(n_130),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_219),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_191),
.B(n_138),
.Y(n_219)
);

OA22x2_ASAP7_75t_L g220 ( 
.A1(n_175),
.A2(n_118),
.B1(n_129),
.B2(n_150),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_221),
.A2(n_228),
.B(n_192),
.Y(n_268)
);

INVx8_ASAP7_75t_L g222 ( 
.A(n_187),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_222),
.Y(n_262)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_193),
.B(n_122),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_223),
.B(n_235),
.Y(n_242)
);

OAI32xp33_ASAP7_75t_L g227 ( 
.A1(n_204),
.A2(n_122),
.A3(n_162),
.B1(n_172),
.B2(n_191),
.Y(n_227)
);

CKINVDCx14_ASAP7_75t_R g247 ( 
.A(n_227),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_199),
.B(n_181),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_168),
.B(n_196),
.C(n_189),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_236),
.C(n_238),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_175),
.A2(n_178),
.B1(n_186),
.B2(n_168),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g235 ( 
.A(n_188),
.B(n_166),
.Y(n_235)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_198),
.B(n_167),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_167),
.B(n_181),
.C(n_202),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_176),
.Y(n_239)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_239),
.Y(n_257)
);

INVxp33_ASAP7_75t_SL g240 ( 
.A(n_221),
.Y(n_240)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_240),
.Y(n_270)
);

OR2x2_ASAP7_75t_L g241 ( 
.A(n_229),
.B(n_178),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_SL g283 ( 
.A(n_241),
.B(n_246),
.Y(n_283)
);

INVx1_ASAP7_75t_SL g244 ( 
.A(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_244),
.B(n_249),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g246 ( 
.A(n_208),
.Y(n_246)
);

XOR2x2_ASAP7_75t_L g248 ( 
.A(n_227),
.B(n_233),
.Y(n_248)
);

OAI21xp33_ASAP7_75t_L g281 ( 
.A1(n_248),
.A2(n_209),
.B(n_237),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_234),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_216),
.A2(n_197),
.B1(n_173),
.B2(n_190),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_250),
.A2(n_254),
.B1(n_259),
.B2(n_260),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g275 ( 
.A1(n_251),
.A2(n_269),
.B1(n_220),
.B2(n_229),
.Y(n_275)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_211),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_253),
.B(n_255),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_215),
.A2(n_201),
.B1(n_177),
.B2(n_176),
.Y(n_254)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_239),
.Y(n_255)
);

HB1xp67_ASAP7_75t_L g256 ( 
.A(n_206),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g290 ( 
.A(n_256),
.Y(n_290)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_210),
.A2(n_201),
.B1(n_184),
.B2(n_203),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_260),
.A2(n_264),
.B1(n_268),
.B2(n_231),
.Y(n_273)
);

INVxp33_ASAP7_75t_L g261 ( 
.A(n_225),
.Y(n_261)
);

INVxp67_ASAP7_75t_L g279 ( 
.A(n_261),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_224),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_263),
.B(n_258),
.Y(n_291)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_210),
.A2(n_184),
.B1(n_166),
.B2(n_194),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g272 ( 
.A1(n_265),
.A2(n_213),
.B(n_214),
.Y(n_272)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_218),
.Y(n_266)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_266),
.Y(n_274)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_226),
.Y(n_267)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_267),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_L g269 ( 
.A1(n_210),
.A2(n_185),
.B1(n_187),
.B2(n_220),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_252),
.B(n_232),
.C(n_236),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_271),
.B(n_276),
.C(n_282),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g294 ( 
.A1(n_272),
.A2(n_275),
.B(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_SL g300 ( 
.A(n_273),
.B(n_281),
.C(n_291),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_252),
.B(n_213),
.C(n_238),
.Y(n_276)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_280),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_265),
.B(n_209),
.C(n_205),
.Y(n_282)
);

HB1xp67_ASAP7_75t_L g284 ( 
.A(n_257),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_292),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_245),
.B(n_205),
.C(n_237),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_285),
.B(n_287),
.C(n_267),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_245),
.B(n_220),
.C(n_226),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_269),
.A2(n_207),
.B1(n_222),
.B2(n_247),
.Y(n_288)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_288),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_248),
.A2(n_266),
.B1(n_250),
.B2(n_244),
.Y(n_289)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_289),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_243),
.Y(n_292)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_293),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_SL g321 ( 
.A(n_294),
.B(n_298),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_270),
.A2(n_268),
.B(n_259),
.Y(n_296)
);

AOI21xp5_ASAP7_75t_L g313 ( 
.A1(n_296),
.A2(n_299),
.B(n_277),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g297 ( 
.A1(n_289),
.A2(n_288),
.B(n_286),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_297),
.A2(n_274),
.B1(n_279),
.B2(n_290),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_SL g298 ( 
.A(n_272),
.B(n_254),
.Y(n_298)
);

XOR2x2_ASAP7_75t_L g299 ( 
.A(n_270),
.B(n_242),
.Y(n_299)
);

OA21x2_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_242),
.B(n_241),
.Y(n_301)
);

AOI31xp67_ASAP7_75t_L g318 ( 
.A1(n_301),
.A2(n_285),
.A3(n_274),
.B(n_293),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_271),
.B(n_262),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_304),
.B(n_308),
.C(n_287),
.Y(n_323)
);

OAI322xp33_ASAP7_75t_L g305 ( 
.A1(n_291),
.A2(n_263),
.A3(n_255),
.B1(n_253),
.B2(n_249),
.C1(n_262),
.C2(n_246),
.Y(n_305)
);

XOR2x2_ASAP7_75t_SL g320 ( 
.A(n_305),
.B(n_283),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_286),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_306),
.B(n_309),
.Y(n_319)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_280),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_276),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_312),
.B(n_323),
.C(n_325),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g327 ( 
.A(n_313),
.B(n_324),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_310),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_314),
.B(n_315),
.Y(n_334)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_297),
.Y(n_315)
);

AOI21xp5_ASAP7_75t_L g316 ( 
.A1(n_294),
.A2(n_275),
.B(n_279),
.Y(n_316)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_316),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_311),
.A2(n_307),
.B1(n_303),
.B2(n_306),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_317),
.A2(n_315),
.B1(n_303),
.B2(n_311),
.Y(n_330)
);

OAI31xp33_ASAP7_75t_L g329 ( 
.A1(n_318),
.A2(n_320),
.A3(n_299),
.B(n_307),
.Y(n_329)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_302),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_322),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_295),
.B(n_290),
.C(n_278),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_318),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_326),
.B(n_296),
.Y(n_340)
);

AOI21xp33_ASAP7_75t_L g341 ( 
.A1(n_329),
.A2(n_300),
.B(n_317),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g338 ( 
.A(n_330),
.B(n_324),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_321),
.B(n_300),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g336 ( 
.A(n_331),
.B(n_332),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_321),
.B(n_298),
.Y(n_332)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_334),
.B(n_319),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_SL g344 ( 
.A(n_337),
.B(n_340),
.Y(n_344)
);

INVxp67_ASAP7_75t_L g342 ( 
.A(n_338),
.Y(n_342)
);

AOI22xp5_ASAP7_75t_L g339 ( 
.A1(n_328),
.A2(n_320),
.B1(n_302),
.B2(n_308),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_339),
.B(n_326),
.Y(n_343)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_341),
.A2(n_327),
.B(n_331),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g347 ( 
.A1(n_343),
.A2(n_345),
.B(n_336),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g346 ( 
.A(n_344),
.B(n_337),
.Y(n_346)
);

OR2x2_ASAP7_75t_L g348 ( 
.A(n_346),
.B(n_347),
.Y(n_348)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_348),
.A2(n_342),
.B1(n_335),
.B2(n_323),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_349),
.B(n_325),
.C(n_333),
.Y(n_350)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_350),
.B(n_327),
.Y(n_351)
);


endmodule