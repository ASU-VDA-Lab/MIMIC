module fake_ariane_2373_n_1788 (n_83, n_8, n_56, n_60, n_160, n_64, n_119, n_124, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_149, n_34, n_158, n_69, n_95, n_92, n_143, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_152, n_120, n_106, n_12, n_53, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_52, n_157, n_135, n_73, n_77, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_125, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1788);

input n_83;
input n_8;
input n_56;
input n_60;
input n_160;
input n_64;
input n_119;
input n_124;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_149;
input n_34;
input n_158;
input n_69;
input n_95;
input n_92;
input n_143;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_152;
input n_120;
input n_106;
input n_12;
input n_53;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_52;
input n_157;
input n_135;
input n_73;
input n_77;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_125;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1788;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_1214;
wire n_634;
wire n_1246;
wire n_1138;
wire n_214;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1457;
wire n_377;
wire n_1682;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_945;
wire n_958;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_167;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_267;
wire n_495;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1006;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_182;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_460;
wire n_1555;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_179;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_337;
wire n_437;
wire n_274;
wire n_1083;
wire n_967;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_824;
wire n_428;
wire n_892;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_172;
wire n_1058;
wire n_347;
wire n_1042;
wire n_183;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_348;
wire n_552;
wire n_670;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1163;
wire n_186;
wire n_1384;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_727;
wire n_699;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_163;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_888;
wire n_845;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_178;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_982;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_642;
wire n_211;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_180;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_169;
wire n_1201;
wire n_1288;
wire n_173;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_166;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1023;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_168;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_181;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_601;
wire n_683;
wire n_236;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_532;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1183;
wire n_1326;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_185;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_164;
wire n_184;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_170;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_176;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_908;
wire n_788;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_898;
wire n_857;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_761;
wire n_733;
wire n_731;
wire n_336;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1409;
wire n_1148;
wire n_1588;
wire n_1684;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1497;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_175;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_948;
wire n_922;
wire n_1004;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_252;
wire n_664;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1126;
wire n_195;
wire n_938;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_174;
wire n_275;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_165;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_177;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1228;
wire n_1244;
wire n_484;
wire n_411;
wire n_849;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g163 ( 
.A(n_116),
.Y(n_163)
);

CKINVDCx5p33_ASAP7_75t_R g164 ( 
.A(n_42),
.Y(n_164)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_141),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_6),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_73),
.Y(n_167)
);

CKINVDCx5p33_ASAP7_75t_R g168 ( 
.A(n_72),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_121),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_71),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_38),
.Y(n_171)
);

CKINVDCx5p33_ASAP7_75t_R g172 ( 
.A(n_82),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_44),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g174 ( 
.A(n_63),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_38),
.Y(n_175)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_23),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_96),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_15),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_124),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_114),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_48),
.Y(n_181)
);

BUFx10_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_36),
.Y(n_183)
);

CKINVDCx5p33_ASAP7_75t_R g184 ( 
.A(n_36),
.Y(n_184)
);

BUFx10_ASAP7_75t_L g185 ( 
.A(n_78),
.Y(n_185)
);

BUFx10_ASAP7_75t_L g186 ( 
.A(n_68),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_17),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_127),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_30),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_107),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_136),
.Y(n_191)
);

CKINVDCx5p33_ASAP7_75t_R g192 ( 
.A(n_77),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g193 ( 
.A(n_64),
.Y(n_193)
);

CKINVDCx20_ASAP7_75t_R g194 ( 
.A(n_44),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_152),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_143),
.Y(n_196)
);

INVx2_ASAP7_75t_L g197 ( 
.A(n_51),
.Y(n_197)
);

CKINVDCx5p33_ASAP7_75t_R g198 ( 
.A(n_46),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g199 ( 
.A(n_21),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_148),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_144),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_39),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_32),
.Y(n_203)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_86),
.Y(n_204)
);

CKINVDCx5p33_ASAP7_75t_R g205 ( 
.A(n_80),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_147),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_43),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_6),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_134),
.Y(n_209)
);

CKINVDCx5p33_ASAP7_75t_R g210 ( 
.A(n_84),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_156),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_109),
.B(n_8),
.Y(n_212)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_120),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_2),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_92),
.Y(n_215)
);

BUFx3_ASAP7_75t_L g216 ( 
.A(n_19),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_131),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_106),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_46),
.Y(n_219)
);

CKINVDCx20_ASAP7_75t_R g220 ( 
.A(n_85),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_130),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_90),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_129),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_108),
.Y(n_224)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_27),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_87),
.Y(n_226)
);

CKINVDCx16_ASAP7_75t_R g227 ( 
.A(n_18),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_17),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_91),
.Y(n_229)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_111),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

BUFx6f_ASAP7_75t_L g232 ( 
.A(n_149),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_32),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_157),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g235 ( 
.A(n_158),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_135),
.Y(n_236)
);

CKINVDCx5p33_ASAP7_75t_R g237 ( 
.A(n_88),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_140),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_94),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_54),
.Y(n_240)
);

CKINVDCx5p33_ASAP7_75t_R g241 ( 
.A(n_7),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_13),
.Y(n_242)
);

CKINVDCx5p33_ASAP7_75t_R g243 ( 
.A(n_3),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_138),
.Y(n_244)
);

HB1xp67_ASAP7_75t_L g245 ( 
.A(n_66),
.Y(n_245)
);

CKINVDCx5p33_ASAP7_75t_R g246 ( 
.A(n_50),
.Y(n_246)
);

HB1xp67_ASAP7_75t_L g247 ( 
.A(n_0),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_39),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_21),
.Y(n_249)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_2),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_139),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_25),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_126),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_65),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_101),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_146),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_115),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g258 ( 
.A(n_70),
.Y(n_258)
);

BUFx10_ASAP7_75t_L g259 ( 
.A(n_62),
.Y(n_259)
);

CKINVDCx12_ASAP7_75t_R g260 ( 
.A(n_13),
.Y(n_260)
);

INVx1_ASAP7_75t_SL g261 ( 
.A(n_47),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_4),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_11),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_151),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_29),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_14),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_83),
.Y(n_267)
);

BUFx10_ASAP7_75t_L g268 ( 
.A(n_95),
.Y(n_268)
);

INVxp67_ASAP7_75t_SL g269 ( 
.A(n_48),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_19),
.Y(n_270)
);

CKINVDCx5p33_ASAP7_75t_R g271 ( 
.A(n_93),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_58),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_4),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_28),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_119),
.Y(n_275)
);

INVx1_ASAP7_75t_SL g276 ( 
.A(n_1),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_110),
.Y(n_277)
);

CKINVDCx20_ASAP7_75t_R g278 ( 
.A(n_55),
.Y(n_278)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_7),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_45),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_27),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_58),
.Y(n_282)
);

INVx2_ASAP7_75t_L g283 ( 
.A(n_67),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_161),
.Y(n_284)
);

CKINVDCx5p33_ASAP7_75t_R g285 ( 
.A(n_8),
.Y(n_285)
);

CKINVDCx5p33_ASAP7_75t_R g286 ( 
.A(n_59),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_14),
.Y(n_287)
);

CKINVDCx5p33_ASAP7_75t_R g288 ( 
.A(n_154),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_133),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_100),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_98),
.Y(n_291)
);

CKINVDCx5p33_ASAP7_75t_R g292 ( 
.A(n_29),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_81),
.Y(n_293)
);

CKINVDCx5p33_ASAP7_75t_R g294 ( 
.A(n_162),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_76),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_122),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_150),
.Y(n_297)
);

CKINVDCx5p33_ASAP7_75t_R g298 ( 
.A(n_113),
.Y(n_298)
);

CKINVDCx5p33_ASAP7_75t_R g299 ( 
.A(n_43),
.Y(n_299)
);

CKINVDCx5p33_ASAP7_75t_R g300 ( 
.A(n_54),
.Y(n_300)
);

BUFx10_ASAP7_75t_L g301 ( 
.A(n_102),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_160),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_45),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_30),
.Y(n_304)
);

CKINVDCx5p33_ASAP7_75t_R g305 ( 
.A(n_28),
.Y(n_305)
);

CKINVDCx5p33_ASAP7_75t_R g306 ( 
.A(n_55),
.Y(n_306)
);

CKINVDCx5p33_ASAP7_75t_R g307 ( 
.A(n_35),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_97),
.Y(n_308)
);

INVx2_ASAP7_75t_L g309 ( 
.A(n_33),
.Y(n_309)
);

INVx2_ASAP7_75t_SL g310 ( 
.A(n_53),
.Y(n_310)
);

CKINVDCx5p33_ASAP7_75t_R g311 ( 
.A(n_155),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_153),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_128),
.Y(n_313)
);

BUFx6f_ASAP7_75t_L g314 ( 
.A(n_89),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_9),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_142),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_1),
.Y(n_317)
);

CKINVDCx5p33_ASAP7_75t_R g318 ( 
.A(n_105),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_3),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_59),
.Y(n_320)
);

HB1xp67_ASAP7_75t_L g321 ( 
.A(n_57),
.Y(n_321)
);

CKINVDCx5p33_ASAP7_75t_R g322 ( 
.A(n_10),
.Y(n_322)
);

CKINVDCx5p33_ASAP7_75t_R g323 ( 
.A(n_50),
.Y(n_323)
);

CKINVDCx5p33_ASAP7_75t_R g324 ( 
.A(n_10),
.Y(n_324)
);

CKINVDCx20_ASAP7_75t_R g325 ( 
.A(n_99),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_11),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_40),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_165),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_165),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_167),
.Y(n_330)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_167),
.Y(n_331)
);

OR2x2_ASAP7_75t_L g332 ( 
.A(n_247),
.B(n_0),
.Y(n_332)
);

HB1xp67_ASAP7_75t_L g333 ( 
.A(n_321),
.Y(n_333)
);

CKINVDCx5p33_ASAP7_75t_R g334 ( 
.A(n_227),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_169),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_169),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_174),
.Y(n_337)
);

CKINVDCx14_ASAP7_75t_R g338 ( 
.A(n_182),
.Y(n_338)
);

INVxp67_ASAP7_75t_L g339 ( 
.A(n_310),
.Y(n_339)
);

INVxp67_ASAP7_75t_SL g340 ( 
.A(n_199),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_170),
.Y(n_341)
);

CKINVDCx5p33_ASAP7_75t_R g342 ( 
.A(n_209),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_213),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_220),
.Y(n_344)
);

HB1xp67_ASAP7_75t_L g345 ( 
.A(n_260),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_230),
.B(n_5),
.Y(n_346)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_170),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g348 ( 
.A(n_251),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g349 ( 
.A(n_310),
.Y(n_349)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_166),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g351 ( 
.A(n_230),
.B(n_5),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_319),
.Y(n_352)
);

CKINVDCx5p33_ASAP7_75t_R g353 ( 
.A(n_258),
.Y(n_353)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_177),
.Y(n_354)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_177),
.Y(n_355)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_179),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_179),
.Y(n_357)
);

INVxp67_ASAP7_75t_L g358 ( 
.A(n_319),
.Y(n_358)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_188),
.Y(n_359)
);

CKINVDCx5p33_ASAP7_75t_R g360 ( 
.A(n_325),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_188),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_204),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g363 ( 
.A(n_256),
.B(n_9),
.Y(n_363)
);

INVxp33_ASAP7_75t_SL g364 ( 
.A(n_164),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_171),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_204),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_206),
.Y(n_367)
);

INVxp33_ASAP7_75t_SL g368 ( 
.A(n_175),
.Y(n_368)
);

CKINVDCx5p33_ASAP7_75t_R g369 ( 
.A(n_181),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_206),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g371 ( 
.A(n_194),
.Y(n_371)
);

CKINVDCx5p33_ASAP7_75t_R g372 ( 
.A(n_184),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_198),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_203),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_217),
.Y(n_375)
);

CKINVDCx5p33_ASAP7_75t_R g376 ( 
.A(n_208),
.Y(n_376)
);

CKINVDCx5p33_ASAP7_75t_R g377 ( 
.A(n_214),
.Y(n_377)
);

CKINVDCx5p33_ASAP7_75t_R g378 ( 
.A(n_228),
.Y(n_378)
);

HB1xp67_ASAP7_75t_L g379 ( 
.A(n_260),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_199),
.Y(n_380)
);

INVx2_ASAP7_75t_L g381 ( 
.A(n_217),
.Y(n_381)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_218),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_202),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_218),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_222),
.Y(n_385)
);

INVxp67_ASAP7_75t_SL g386 ( 
.A(n_216),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_222),
.Y(n_387)
);

CKINVDCx5p33_ASAP7_75t_R g388 ( 
.A(n_233),
.Y(n_388)
);

CKINVDCx20_ASAP7_75t_R g389 ( 
.A(n_278),
.Y(n_389)
);

INVx1_ASAP7_75t_L g390 ( 
.A(n_223),
.Y(n_390)
);

INVxp67_ASAP7_75t_SL g391 ( 
.A(n_216),
.Y(n_391)
);

CKINVDCx20_ASAP7_75t_R g392 ( 
.A(n_326),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_182),
.Y(n_393)
);

INVx2_ASAP7_75t_L g394 ( 
.A(n_223),
.Y(n_394)
);

CKINVDCx5p33_ASAP7_75t_R g395 ( 
.A(n_241),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_224),
.Y(n_396)
);

CKINVDCx5p33_ASAP7_75t_R g397 ( 
.A(n_243),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_224),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_185),
.Y(n_399)
);

INVxp67_ASAP7_75t_SL g400 ( 
.A(n_166),
.Y(n_400)
);

NOR2xp67_ASAP7_75t_L g401 ( 
.A(n_256),
.B(n_12),
.Y(n_401)
);

CKINVDCx5p33_ASAP7_75t_R g402 ( 
.A(n_246),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_226),
.Y(n_403)
);

INVx4_ASAP7_75t_R g404 ( 
.A(n_193),
.Y(n_404)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_226),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_185),
.Y(n_406)
);

CKINVDCx5p33_ASAP7_75t_R g407 ( 
.A(n_248),
.Y(n_407)
);

INVx1_ASAP7_75t_L g408 ( 
.A(n_229),
.Y(n_408)
);

CKINVDCx20_ASAP7_75t_R g409 ( 
.A(n_185),
.Y(n_409)
);

CKINVDCx5p33_ASAP7_75t_R g410 ( 
.A(n_337),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_L g411 ( 
.A(n_328),
.B(n_245),
.Y(n_411)
);

AND2x4_ASAP7_75t_L g412 ( 
.A(n_328),
.B(n_330),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g413 ( 
.A(n_330),
.B(n_229),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_329),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_329),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g416 ( 
.A(n_342),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_331),
.B(n_231),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_329),
.Y(n_418)
);

INVxp67_ASAP7_75t_L g419 ( 
.A(n_380),
.Y(n_419)
);

OR2x2_ASAP7_75t_L g420 ( 
.A(n_333),
.B(n_173),
.Y(n_420)
);

INVx5_ASAP7_75t_L g421 ( 
.A(n_347),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_347),
.Y(n_422)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_331),
.B(n_335),
.Y(n_423)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_347),
.Y(n_424)
);

INVx1_ASAP7_75t_L g425 ( 
.A(n_381),
.Y(n_425)
);

BUFx3_ASAP7_75t_L g426 ( 
.A(n_335),
.Y(n_426)
);

AND2x6_ASAP7_75t_L g427 ( 
.A(n_381),
.B(n_256),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_381),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g429 ( 
.A(n_336),
.B(n_197),
.Y(n_429)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_385),
.Y(n_430)
);

INVx2_ASAP7_75t_L g431 ( 
.A(n_385),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g432 ( 
.A(n_340),
.B(n_231),
.Y(n_432)
);

AND2x4_ASAP7_75t_L g433 ( 
.A(n_336),
.B(n_197),
.Y(n_433)
);

BUFx6f_ASAP7_75t_L g434 ( 
.A(n_385),
.Y(n_434)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_387),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_341),
.B(n_257),
.Y(n_436)
);

INVx2_ASAP7_75t_L g437 ( 
.A(n_387),
.Y(n_437)
);

AND2x2_ASAP7_75t_L g438 ( 
.A(n_341),
.B(n_309),
.Y(n_438)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_354),
.B(n_309),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g440 ( 
.A1(n_387),
.A2(n_267),
.B(n_257),
.Y(n_440)
);

BUFx6f_ASAP7_75t_L g441 ( 
.A(n_394),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_394),
.Y(n_442)
);

INVx2_ASAP7_75t_L g443 ( 
.A(n_394),
.Y(n_443)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_354),
.Y(n_444)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_355),
.Y(n_445)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_355),
.Y(n_446)
);

INVx1_ASAP7_75t_L g447 ( 
.A(n_356),
.Y(n_447)
);

AND2x2_ASAP7_75t_L g448 ( 
.A(n_356),
.B(n_186),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_357),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_357),
.Y(n_450)
);

INVx2_ASAP7_75t_L g451 ( 
.A(n_359),
.Y(n_451)
);

INVx3_ASAP7_75t_L g452 ( 
.A(n_359),
.Y(n_452)
);

AND2x4_ASAP7_75t_L g453 ( 
.A(n_361),
.B(n_173),
.Y(n_453)
);

AND2x4_ASAP7_75t_L g454 ( 
.A(n_361),
.B(n_176),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_362),
.Y(n_455)
);

INVx2_ASAP7_75t_L g456 ( 
.A(n_362),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_366),
.Y(n_457)
);

BUFx6f_ASAP7_75t_L g458 ( 
.A(n_366),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_367),
.Y(n_459)
);

BUFx6f_ASAP7_75t_L g460 ( 
.A(n_367),
.Y(n_460)
);

INVx1_ASAP7_75t_L g461 ( 
.A(n_370),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g462 ( 
.A(n_363),
.B(n_255),
.Y(n_462)
);

INVx2_ASAP7_75t_L g463 ( 
.A(n_370),
.Y(n_463)
);

BUFx3_ASAP7_75t_L g464 ( 
.A(n_375),
.Y(n_464)
);

INVx2_ASAP7_75t_L g465 ( 
.A(n_375),
.Y(n_465)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_382),
.B(n_267),
.Y(n_466)
);

AND2x4_ASAP7_75t_L g467 ( 
.A(n_382),
.B(n_176),
.Y(n_467)
);

AO22x1_ASAP7_75t_L g468 ( 
.A1(n_346),
.A2(n_269),
.B1(n_289),
.B2(n_290),
.Y(n_468)
);

BUFx6f_ASAP7_75t_L g469 ( 
.A(n_384),
.Y(n_469)
);

INVx2_ASAP7_75t_L g470 ( 
.A(n_384),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_390),
.Y(n_471)
);

NAND2xp5_ASAP7_75t_SL g472 ( 
.A(n_363),
.B(n_401),
.Y(n_472)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_390),
.Y(n_473)
);

AND2x4_ASAP7_75t_L g474 ( 
.A(n_396),
.B(n_178),
.Y(n_474)
);

INVx2_ASAP7_75t_L g475 ( 
.A(n_396),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_398),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_398),
.Y(n_477)
);

INVx2_ASAP7_75t_L g478 ( 
.A(n_403),
.Y(n_478)
);

INVx2_ASAP7_75t_L g479 ( 
.A(n_403),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_405),
.Y(n_480)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_405),
.Y(n_481)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_408),
.Y(n_482)
);

INVx2_ASAP7_75t_L g483 ( 
.A(n_408),
.Y(n_483)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_401),
.Y(n_484)
);

INVx1_ASAP7_75t_L g485 ( 
.A(n_400),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_458),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_458),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_458),
.Y(n_488)
);

BUFx2_ASAP7_75t_L g489 ( 
.A(n_419),
.Y(n_489)
);

BUFx10_ASAP7_75t_L g490 ( 
.A(n_410),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_448),
.B(n_365),
.Y(n_491)
);

AND2x2_ASAP7_75t_L g492 ( 
.A(n_448),
.B(n_386),
.Y(n_492)
);

BUFx10_ASAP7_75t_L g493 ( 
.A(n_432),
.Y(n_493)
);

AND3x2_ASAP7_75t_L g494 ( 
.A(n_448),
.B(n_351),
.C(n_345),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_447),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g496 ( 
.A1(n_420),
.A2(n_332),
.B1(n_352),
.B2(n_339),
.Y(n_496)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_447),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_412),
.B(n_369),
.Y(n_498)
);

OR2x6_ASAP7_75t_L g499 ( 
.A(n_468),
.B(n_332),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_434),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_484),
.B(n_338),
.Y(n_501)
);

INVx4_ASAP7_75t_L g502 ( 
.A(n_412),
.Y(n_502)
);

INVx2_ASAP7_75t_L g503 ( 
.A(n_434),
.Y(n_503)
);

INVx6_ASAP7_75t_L g504 ( 
.A(n_412),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_412),
.B(n_372),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_L g506 ( 
.A(n_458),
.B(n_373),
.Y(n_506)
);

INVx1_ASAP7_75t_SL g507 ( 
.A(n_416),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_L g508 ( 
.A(n_485),
.B(n_364),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g509 ( 
.A(n_484),
.B(n_374),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_412),
.B(n_376),
.Y(n_510)
);

AOI22xp33_ASAP7_75t_L g511 ( 
.A1(n_432),
.A2(n_368),
.B1(n_187),
.B2(n_279),
.Y(n_511)
);

INVx2_ASAP7_75t_L g512 ( 
.A(n_434),
.Y(n_512)
);

INVx2_ASAP7_75t_L g513 ( 
.A(n_434),
.Y(n_513)
);

BUFx3_ASAP7_75t_L g514 ( 
.A(n_426),
.Y(n_514)
);

INVx4_ASAP7_75t_L g515 ( 
.A(n_412),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_L g516 ( 
.A(n_484),
.B(n_377),
.Y(n_516)
);

NOR2xp33_ASAP7_75t_L g517 ( 
.A(n_485),
.B(n_378),
.Y(n_517)
);

INVx3_ASAP7_75t_L g518 ( 
.A(n_460),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_SL g519 ( 
.A(n_485),
.B(n_388),
.Y(n_519)
);

AND2x6_ASAP7_75t_L g520 ( 
.A(n_423),
.B(n_453),
.Y(n_520)
);

INVx4_ASAP7_75t_L g521 ( 
.A(n_452),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g522 ( 
.A(n_423),
.B(n_395),
.Y(n_522)
);

INVx1_ASAP7_75t_L g523 ( 
.A(n_447),
.Y(n_523)
);

AND2x6_ASAP7_75t_L g524 ( 
.A(n_423),
.B(n_453),
.Y(n_524)
);

BUFx6f_ASAP7_75t_L g525 ( 
.A(n_434),
.Y(n_525)
);

INVx3_ASAP7_75t_L g526 ( 
.A(n_460),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_449),
.Y(n_527)
);

INVx2_ASAP7_75t_L g528 ( 
.A(n_434),
.Y(n_528)
);

INVx2_ASAP7_75t_L g529 ( 
.A(n_434),
.Y(n_529)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_449),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_449),
.Y(n_531)
);

HB1xp67_ASAP7_75t_L g532 ( 
.A(n_419),
.Y(n_532)
);

NOR2xp33_ASAP7_75t_L g533 ( 
.A(n_472),
.B(n_397),
.Y(n_533)
);

BUFx10_ASAP7_75t_L g534 ( 
.A(n_453),
.Y(n_534)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_472),
.B(n_402),
.Y(n_535)
);

NOR2x1p5_ASAP7_75t_L g536 ( 
.A(n_420),
.B(n_334),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_L g537 ( 
.A(n_446),
.B(n_407),
.Y(n_537)
);

INVx3_ASAP7_75t_L g538 ( 
.A(n_460),
.Y(n_538)
);

INVx2_ASAP7_75t_SL g539 ( 
.A(n_411),
.Y(n_539)
);

INVx1_ASAP7_75t_L g540 ( 
.A(n_450),
.Y(n_540)
);

INVx2_ASAP7_75t_L g541 ( 
.A(n_434),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_L g542 ( 
.A(n_426),
.B(n_391),
.Y(n_542)
);

INVx5_ASAP7_75t_L g543 ( 
.A(n_427),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_434),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g545 ( 
.A(n_446),
.B(n_379),
.Y(n_545)
);

AOI22xp5_ASAP7_75t_L g546 ( 
.A1(n_468),
.A2(n_250),
.B1(n_261),
.B2(n_276),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_411),
.B(n_393),
.Y(n_547)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_450),
.Y(n_548)
);

INVx2_ASAP7_75t_L g549 ( 
.A(n_441),
.Y(n_549)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_460),
.Y(n_550)
);

INVx3_ASAP7_75t_L g551 ( 
.A(n_460),
.Y(n_551)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_460),
.Y(n_552)
);

NOR3xp33_ASAP7_75t_L g553 ( 
.A(n_468),
.B(n_350),
.C(n_273),
.Y(n_553)
);

NAND2xp5_ASAP7_75t_SL g554 ( 
.A(n_426),
.B(n_343),
.Y(n_554)
);

HB1xp67_ASAP7_75t_L g555 ( 
.A(n_416),
.Y(n_555)
);

INVx2_ASAP7_75t_SL g556 ( 
.A(n_464),
.Y(n_556)
);

AOI22xp5_ASAP7_75t_L g557 ( 
.A1(n_462),
.A2(n_320),
.B1(n_287),
.B2(n_286),
.Y(n_557)
);

AND2x2_ASAP7_75t_L g558 ( 
.A(n_429),
.B(n_339),
.Y(n_558)
);

INVx2_ASAP7_75t_L g559 ( 
.A(n_441),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_464),
.B(n_349),
.Y(n_560)
);

BUFx3_ASAP7_75t_L g561 ( 
.A(n_464),
.Y(n_561)
);

BUFx2_ASAP7_75t_L g562 ( 
.A(n_420),
.Y(n_562)
);

INVx2_ASAP7_75t_L g563 ( 
.A(n_441),
.Y(n_563)
);

BUFx6f_ASAP7_75t_L g564 ( 
.A(n_441),
.Y(n_564)
);

INVx2_ASAP7_75t_L g565 ( 
.A(n_441),
.Y(n_565)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_450),
.Y(n_566)
);

INVxp67_ASAP7_75t_SL g567 ( 
.A(n_452),
.Y(n_567)
);

INVx4_ASAP7_75t_L g568 ( 
.A(n_452),
.Y(n_568)
);

INVx2_ASAP7_75t_L g569 ( 
.A(n_441),
.Y(n_569)
);

INVx2_ASAP7_75t_SL g570 ( 
.A(n_464),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_429),
.B(n_349),
.Y(n_571)
);

INVx8_ASAP7_75t_L g572 ( 
.A(n_427),
.Y(n_572)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_457),
.Y(n_573)
);

NOR2xp33_ASAP7_75t_L g574 ( 
.A(n_462),
.B(n_457),
.Y(n_574)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_452),
.B(n_352),
.Y(n_575)
);

INVx1_ASAP7_75t_L g576 ( 
.A(n_457),
.Y(n_576)
);

INVx1_ASAP7_75t_SL g577 ( 
.A(n_429),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_459),
.Y(n_578)
);

AOI22xp33_ASAP7_75t_L g579 ( 
.A1(n_440),
.A2(n_207),
.B1(n_219),
.B2(n_225),
.Y(n_579)
);

NOR2xp33_ASAP7_75t_L g580 ( 
.A(n_459),
.B(n_399),
.Y(n_580)
);

INVx4_ASAP7_75t_L g581 ( 
.A(n_452),
.Y(n_581)
);

INVx2_ASAP7_75t_SL g582 ( 
.A(n_453),
.Y(n_582)
);

INVx1_ASAP7_75t_L g583 ( 
.A(n_459),
.Y(n_583)
);

BUFx6f_ASAP7_75t_L g584 ( 
.A(n_441),
.Y(n_584)
);

INVx4_ASAP7_75t_L g585 ( 
.A(n_460),
.Y(n_585)
);

AOI22xp33_ASAP7_75t_L g586 ( 
.A1(n_440),
.A2(n_207),
.B1(n_219),
.B2(n_225),
.Y(n_586)
);

NOR2xp33_ASAP7_75t_L g587 ( 
.A(n_461),
.B(n_406),
.Y(n_587)
);

OR2x6_ASAP7_75t_L g588 ( 
.A(n_438),
.B(n_358),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_461),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_SL g590 ( 
.A(n_453),
.B(n_344),
.Y(n_590)
);

NAND2xp5_ASAP7_75t_SL g591 ( 
.A(n_453),
.B(n_353),
.Y(n_591)
);

OAI22xp33_ASAP7_75t_L g592 ( 
.A1(n_413),
.A2(n_358),
.B1(n_272),
.B2(n_281),
.Y(n_592)
);

INVx4_ASAP7_75t_L g593 ( 
.A(n_469),
.Y(n_593)
);

BUFx6f_ASAP7_75t_L g594 ( 
.A(n_469),
.Y(n_594)
);

OR2x6_ASAP7_75t_L g595 ( 
.A(n_438),
.B(n_178),
.Y(n_595)
);

BUFx2_ASAP7_75t_L g596 ( 
.A(n_454),
.Y(n_596)
);

INVxp67_ASAP7_75t_L g597 ( 
.A(n_438),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_454),
.Y(n_598)
);

INVx1_ASAP7_75t_L g599 ( 
.A(n_473),
.Y(n_599)
);

INVx2_ASAP7_75t_SL g600 ( 
.A(n_454),
.Y(n_600)
);

INVx1_ASAP7_75t_L g601 ( 
.A(n_473),
.Y(n_601)
);

OR2x6_ASAP7_75t_L g602 ( 
.A(n_439),
.B(n_183),
.Y(n_602)
);

INVx1_ASAP7_75t_L g603 ( 
.A(n_473),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_477),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_414),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_414),
.Y(n_606)
);

BUFx3_ASAP7_75t_L g607 ( 
.A(n_477),
.Y(n_607)
);

INVx2_ASAP7_75t_SL g608 ( 
.A(n_454),
.Y(n_608)
);

NOR2x1p5_ASAP7_75t_L g609 ( 
.A(n_413),
.B(n_360),
.Y(n_609)
);

INVx2_ASAP7_75t_L g610 ( 
.A(n_414),
.Y(n_610)
);

AOI22xp33_ASAP7_75t_L g611 ( 
.A1(n_440),
.A2(n_454),
.B1(n_467),
.B2(n_474),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_469),
.Y(n_612)
);

OAI22xp33_ASAP7_75t_SL g613 ( 
.A1(n_417),
.A2(n_306),
.B1(n_327),
.B2(n_324),
.Y(n_613)
);

INVx4_ASAP7_75t_L g614 ( 
.A(n_469),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_414),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_SL g616 ( 
.A(n_454),
.B(n_467),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_431),
.Y(n_617)
);

AOI22xp33_ASAP7_75t_L g618 ( 
.A1(n_440),
.A2(n_280),
.B1(n_187),
.B2(n_189),
.Y(n_618)
);

NAND2xp5_ASAP7_75t_SL g619 ( 
.A(n_467),
.B(n_409),
.Y(n_619)
);

NAND2xp33_ASAP7_75t_L g620 ( 
.A(n_469),
.B(n_289),
.Y(n_620)
);

AND2x2_ASAP7_75t_L g621 ( 
.A(n_439),
.B(n_183),
.Y(n_621)
);

INVx1_ASAP7_75t_L g622 ( 
.A(n_469),
.Y(n_622)
);

INVx1_ASAP7_75t_L g623 ( 
.A(n_469),
.Y(n_623)
);

NOR2xp33_ASAP7_75t_L g624 ( 
.A(n_477),
.B(n_348),
.Y(n_624)
);

BUFx3_ASAP7_75t_L g625 ( 
.A(n_480),
.Y(n_625)
);

CKINVDCx20_ASAP7_75t_R g626 ( 
.A(n_439),
.Y(n_626)
);

AOI22xp33_ASAP7_75t_L g627 ( 
.A1(n_499),
.A2(n_440),
.B1(n_467),
.B2(n_474),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_539),
.B(n_480),
.Y(n_628)
);

INVx8_ASAP7_75t_L g629 ( 
.A(n_520),
.Y(n_629)
);

INVxp67_ASAP7_75t_L g630 ( 
.A(n_555),
.Y(n_630)
);

BUFx10_ASAP7_75t_L g631 ( 
.A(n_547),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_605),
.Y(n_632)
);

INVxp67_ASAP7_75t_L g633 ( 
.A(n_507),
.Y(n_633)
);

BUFx8_ASAP7_75t_L g634 ( 
.A(n_489),
.Y(n_634)
);

AOI21xp5_ASAP7_75t_L g635 ( 
.A1(n_567),
.A2(n_570),
.B(n_556),
.Y(n_635)
);

NAND2xp33_ASAP7_75t_L g636 ( 
.A(n_520),
.B(n_469),
.Y(n_636)
);

NAND2xp5_ASAP7_75t_L g637 ( 
.A(n_539),
.B(n_480),
.Y(n_637)
);

NAND2xp5_ASAP7_75t_SL g638 ( 
.A(n_534),
.B(n_502),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_534),
.B(n_469),
.Y(n_639)
);

INVx2_ASAP7_75t_L g640 ( 
.A(n_605),
.Y(n_640)
);

INVx2_ASAP7_75t_L g641 ( 
.A(n_606),
.Y(n_641)
);

NAND2xp5_ASAP7_75t_L g642 ( 
.A(n_517),
.B(n_467),
.Y(n_642)
);

NAND2xp5_ASAP7_75t_L g643 ( 
.A(n_508),
.B(n_467),
.Y(n_643)
);

AND2x4_ASAP7_75t_L g644 ( 
.A(n_502),
.B(n_474),
.Y(n_644)
);

HB1xp67_ASAP7_75t_L g645 ( 
.A(n_489),
.Y(n_645)
);

NAND2xp5_ASAP7_75t_SL g646 ( 
.A(n_534),
.B(n_444),
.Y(n_646)
);

INVx3_ASAP7_75t_L g647 ( 
.A(n_502),
.Y(n_647)
);

NAND2xp33_ASAP7_75t_L g648 ( 
.A(n_520),
.B(n_524),
.Y(n_648)
);

INVx2_ASAP7_75t_L g649 ( 
.A(n_606),
.Y(n_649)
);

NAND2xp5_ASAP7_75t_L g650 ( 
.A(n_537),
.B(n_474),
.Y(n_650)
);

NOR2xp33_ASAP7_75t_L g651 ( 
.A(n_493),
.B(n_417),
.Y(n_651)
);

NAND2xp5_ASAP7_75t_SL g652 ( 
.A(n_515),
.B(n_444),
.Y(n_652)
);

NAND2xp5_ASAP7_75t_L g653 ( 
.A(n_492),
.B(n_474),
.Y(n_653)
);

NOR2xp33_ASAP7_75t_L g654 ( 
.A(n_493),
.B(n_436),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_SL g655 ( 
.A(n_515),
.B(n_444),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_L g656 ( 
.A(n_492),
.B(n_474),
.Y(n_656)
);

HB1xp67_ASAP7_75t_L g657 ( 
.A(n_588),
.Y(n_657)
);

NOR2xp33_ASAP7_75t_R g658 ( 
.A(n_490),
.B(n_371),
.Y(n_658)
);

INVx2_ASAP7_75t_L g659 ( 
.A(n_610),
.Y(n_659)
);

NAND2xp5_ASAP7_75t_L g660 ( 
.A(n_596),
.B(n_444),
.Y(n_660)
);

INVx2_ASAP7_75t_L g661 ( 
.A(n_610),
.Y(n_661)
);

O2A1O1Ixp33_ASAP7_75t_L g662 ( 
.A1(n_597),
.A2(n_470),
.B(n_482),
.C(n_481),
.Y(n_662)
);

NOR2xp33_ASAP7_75t_L g663 ( 
.A(n_493),
.B(n_522),
.Y(n_663)
);

AND2x2_ASAP7_75t_L g664 ( 
.A(n_562),
.B(n_383),
.Y(n_664)
);

BUFx6f_ASAP7_75t_L g665 ( 
.A(n_504),
.Y(n_665)
);

NAND2xp5_ASAP7_75t_SL g666 ( 
.A(n_515),
.B(n_582),
.Y(n_666)
);

NOR2xp33_ASAP7_75t_L g667 ( 
.A(n_509),
.B(n_436),
.Y(n_667)
);

INVxp67_ASAP7_75t_L g668 ( 
.A(n_580),
.Y(n_668)
);

AND2x6_ASAP7_75t_L g669 ( 
.A(n_607),
.B(n_625),
.Y(n_669)
);

BUFx3_ASAP7_75t_L g670 ( 
.A(n_520),
.Y(n_670)
);

INVxp67_ASAP7_75t_L g671 ( 
.A(n_587),
.Y(n_671)
);

NAND2xp5_ASAP7_75t_L g672 ( 
.A(n_596),
.B(n_445),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_L g673 ( 
.A(n_582),
.B(n_445),
.Y(n_673)
);

NAND2xp5_ASAP7_75t_L g674 ( 
.A(n_598),
.B(n_445),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_625),
.Y(n_675)
);

NAND2xp5_ASAP7_75t_L g676 ( 
.A(n_598),
.B(n_445),
.Y(n_676)
);

NAND3xp33_ASAP7_75t_L g677 ( 
.A(n_624),
.B(n_466),
.C(n_455),
.Y(n_677)
);

NAND2xp5_ASAP7_75t_L g678 ( 
.A(n_600),
.B(n_451),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_600),
.B(n_451),
.Y(n_679)
);

NAND2xp5_ASAP7_75t_SL g680 ( 
.A(n_533),
.B(n_466),
.Y(n_680)
);

NAND3xp33_ASAP7_75t_L g681 ( 
.A(n_532),
.B(n_455),
.C(n_451),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_608),
.B(n_455),
.Y(n_682)
);

NAND2xp5_ASAP7_75t_SL g683 ( 
.A(n_608),
.B(n_455),
.Y(n_683)
);

INVx1_ASAP7_75t_L g684 ( 
.A(n_504),
.Y(n_684)
);

INVx2_ASAP7_75t_SL g685 ( 
.A(n_558),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_504),
.Y(n_686)
);

NAND2xp5_ASAP7_75t_L g687 ( 
.A(n_542),
.B(n_456),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_L g688 ( 
.A(n_520),
.B(n_524),
.Y(n_688)
);

INVx2_ASAP7_75t_L g689 ( 
.A(n_615),
.Y(n_689)
);

NAND2xp5_ASAP7_75t_L g690 ( 
.A(n_575),
.B(n_456),
.Y(n_690)
);

A2O1A1Ixp33_ASAP7_75t_L g691 ( 
.A1(n_574),
.A2(n_483),
.B(n_482),
.C(n_481),
.Y(n_691)
);

NAND2xp5_ASAP7_75t_SL g692 ( 
.A(n_521),
.B(n_456),
.Y(n_692)
);

AOI221xp5_ASAP7_75t_L g693 ( 
.A1(n_496),
.A2(n_280),
.B1(n_240),
.B2(n_279),
.C(n_249),
.Y(n_693)
);

NAND2xp5_ASAP7_75t_L g694 ( 
.A(n_577),
.B(n_456),
.Y(n_694)
);

NOR2xp33_ASAP7_75t_L g695 ( 
.A(n_516),
.B(n_463),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_520),
.B(n_524),
.Y(n_696)
);

INVx4_ASAP7_75t_L g697 ( 
.A(n_524),
.Y(n_697)
);

AOI22xp33_ASAP7_75t_L g698 ( 
.A1(n_499),
.A2(n_553),
.B1(n_546),
.B2(n_611),
.Y(n_698)
);

AND2x2_ASAP7_75t_L g699 ( 
.A(n_562),
.B(n_389),
.Y(n_699)
);

NAND2xp33_ASAP7_75t_L g700 ( 
.A(n_524),
.B(n_427),
.Y(n_700)
);

INVx2_ASAP7_75t_L g701 ( 
.A(n_615),
.Y(n_701)
);

OR2x2_ASAP7_75t_L g702 ( 
.A(n_588),
.B(n_433),
.Y(n_702)
);

OR2x6_ASAP7_75t_L g703 ( 
.A(n_499),
.B(n_433),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_L g704 ( 
.A(n_524),
.B(n_427),
.Y(n_704)
);

NAND3xp33_ASAP7_75t_L g705 ( 
.A(n_511),
.B(n_465),
.C(n_463),
.Y(n_705)
);

INVx2_ASAP7_75t_L g706 ( 
.A(n_617),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_588),
.B(n_392),
.Y(n_707)
);

CKINVDCx5p33_ASAP7_75t_R g708 ( 
.A(n_490),
.Y(n_708)
);

INVx3_ASAP7_75t_L g709 ( 
.A(n_504),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_SL g710 ( 
.A(n_535),
.B(n_463),
.Y(n_710)
);

INVxp67_ASAP7_75t_L g711 ( 
.A(n_545),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_560),
.B(n_463),
.Y(n_712)
);

NAND2xp5_ASAP7_75t_L g713 ( 
.A(n_556),
.B(n_465),
.Y(n_713)
);

NOR2xp33_ASAP7_75t_L g714 ( 
.A(n_519),
.B(n_491),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_570),
.B(n_465),
.Y(n_715)
);

NOR2xp33_ASAP7_75t_L g716 ( 
.A(n_498),
.B(n_465),
.Y(n_716)
);

INVx2_ASAP7_75t_L g717 ( 
.A(n_617),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_495),
.Y(n_718)
);

INVx2_ASAP7_75t_SL g719 ( 
.A(n_558),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_497),
.Y(n_720)
);

OR2x6_ASAP7_75t_L g721 ( 
.A(n_499),
.B(n_433),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_571),
.Y(n_722)
);

INVx2_ASAP7_75t_L g723 ( 
.A(n_523),
.Y(n_723)
);

NOR2xp67_ASAP7_75t_L g724 ( 
.A(n_501),
.B(n_471),
.Y(n_724)
);

INVx2_ASAP7_75t_L g725 ( 
.A(n_527),
.Y(n_725)
);

NAND2xp5_ASAP7_75t_SL g726 ( 
.A(n_568),
.B(n_471),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_568),
.B(n_581),
.Y(n_727)
);

INVx1_ASAP7_75t_L g728 ( 
.A(n_530),
.Y(n_728)
);

NAND2xp33_ASAP7_75t_L g729 ( 
.A(n_594),
.B(n_427),
.Y(n_729)
);

NAND2xp5_ASAP7_75t_L g730 ( 
.A(n_581),
.B(n_471),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_531),
.Y(n_731)
);

INVx2_ASAP7_75t_L g732 ( 
.A(n_540),
.Y(n_732)
);

NOR2xp33_ASAP7_75t_L g733 ( 
.A(n_505),
.B(n_475),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_571),
.Y(n_734)
);

INVx2_ASAP7_75t_L g735 ( 
.A(n_548),
.Y(n_735)
);

BUFx2_ASAP7_75t_R g736 ( 
.A(n_619),
.Y(n_736)
);

INVxp67_ASAP7_75t_L g737 ( 
.A(n_588),
.Y(n_737)
);

OR2x2_ASAP7_75t_L g738 ( 
.A(n_595),
.B(n_433),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_581),
.B(n_475),
.Y(n_739)
);

INVx1_ASAP7_75t_L g740 ( 
.A(n_566),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_616),
.B(n_475),
.Y(n_741)
);

NAND2xp5_ASAP7_75t_L g742 ( 
.A(n_621),
.B(n_475),
.Y(n_742)
);

AND2x2_ASAP7_75t_L g743 ( 
.A(n_490),
.B(n_433),
.Y(n_743)
);

O2A1O1Ixp33_ASAP7_75t_L g744 ( 
.A1(n_573),
.A2(n_482),
.B(n_481),
.C(n_479),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_SL g745 ( 
.A(n_594),
.B(n_476),
.Y(n_745)
);

NAND2xp5_ASAP7_75t_L g746 ( 
.A(n_621),
.B(n_476),
.Y(n_746)
);

NOR3xp33_ASAP7_75t_L g747 ( 
.A(n_510),
.B(n_274),
.C(n_242),
.Y(n_747)
);

INVx2_ASAP7_75t_L g748 ( 
.A(n_576),
.Y(n_748)
);

NAND2xp5_ASAP7_75t_L g749 ( 
.A(n_578),
.B(n_476),
.Y(n_749)
);

NAND3xp33_ASAP7_75t_L g750 ( 
.A(n_557),
.B(n_478),
.C(n_476),
.Y(n_750)
);

HB1xp67_ASAP7_75t_L g751 ( 
.A(n_626),
.Y(n_751)
);

INVx1_ASAP7_75t_L g752 ( 
.A(n_583),
.Y(n_752)
);

BUFx6f_ASAP7_75t_L g753 ( 
.A(n_572),
.Y(n_753)
);

NAND2xp5_ASAP7_75t_L g754 ( 
.A(n_589),
.B(n_478),
.Y(n_754)
);

NAND2xp5_ASAP7_75t_SL g755 ( 
.A(n_594),
.B(n_478),
.Y(n_755)
);

AOI221xp5_ASAP7_75t_L g756 ( 
.A1(n_592),
.A2(n_189),
.B1(n_240),
.B2(n_249),
.C(n_263),
.Y(n_756)
);

AOI22xp5_ASAP7_75t_L g757 ( 
.A1(n_626),
.A2(n_433),
.B1(n_482),
.B2(n_481),
.Y(n_757)
);

BUFx6f_ASAP7_75t_L g758 ( 
.A(n_572),
.Y(n_758)
);

INVxp67_ASAP7_75t_L g759 ( 
.A(n_536),
.Y(n_759)
);

OAI22xp5_ASAP7_75t_L g760 ( 
.A1(n_514),
.A2(n_483),
.B1(n_479),
.B2(n_307),
.Y(n_760)
);

AND2x4_ASAP7_75t_L g761 ( 
.A(n_595),
.B(n_479),
.Y(n_761)
);

INVx1_ASAP7_75t_L g762 ( 
.A(n_599),
.Y(n_762)
);

AOI22xp33_ASAP7_75t_L g763 ( 
.A1(n_579),
.A2(n_440),
.B1(n_479),
.B2(n_483),
.Y(n_763)
);

BUFx3_ASAP7_75t_L g764 ( 
.A(n_514),
.Y(n_764)
);

XNOR2xp5_ASAP7_75t_L g765 ( 
.A(n_494),
.B(n_404),
.Y(n_765)
);

AOI22xp33_ASAP7_75t_L g766 ( 
.A1(n_586),
.A2(n_483),
.B1(n_442),
.B2(n_443),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_601),
.Y(n_767)
);

BUFx3_ASAP7_75t_L g768 ( 
.A(n_561),
.Y(n_768)
);

NAND2xp5_ASAP7_75t_L g769 ( 
.A(n_603),
.B(n_442),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_SL g770 ( 
.A(n_594),
.B(n_415),
.Y(n_770)
);

NOR3xp33_ASAP7_75t_L g771 ( 
.A(n_590),
.B(n_265),
.C(n_263),
.Y(n_771)
);

INVx2_ASAP7_75t_SL g772 ( 
.A(n_609),
.Y(n_772)
);

AND2x4_ASAP7_75t_L g773 ( 
.A(n_595),
.B(n_265),
.Y(n_773)
);

NAND2xp33_ASAP7_75t_SL g774 ( 
.A(n_591),
.B(n_252),
.Y(n_774)
);

NAND2xp5_ASAP7_75t_L g775 ( 
.A(n_604),
.B(n_415),
.Y(n_775)
);

NAND2xp5_ASAP7_75t_L g776 ( 
.A(n_561),
.B(n_595),
.Y(n_776)
);

INVx1_ASAP7_75t_L g777 ( 
.A(n_602),
.Y(n_777)
);

NAND2xp5_ASAP7_75t_L g778 ( 
.A(n_602),
.B(n_415),
.Y(n_778)
);

NAND2xp5_ASAP7_75t_SL g779 ( 
.A(n_554),
.B(n_262),
.Y(n_779)
);

INVx2_ASAP7_75t_SL g780 ( 
.A(n_602),
.Y(n_780)
);

AOI22xp33_ASAP7_75t_L g781 ( 
.A1(n_618),
.A2(n_443),
.B1(n_437),
.B2(n_431),
.Y(n_781)
);

NOR2xp33_ASAP7_75t_L g782 ( 
.A(n_602),
.B(n_418),
.Y(n_782)
);

INVx1_ASAP7_75t_L g783 ( 
.A(n_486),
.Y(n_783)
);

INVx2_ASAP7_75t_L g784 ( 
.A(n_518),
.Y(n_784)
);

AND2x2_ASAP7_75t_L g785 ( 
.A(n_620),
.B(n_418),
.Y(n_785)
);

NAND2xp5_ASAP7_75t_SL g786 ( 
.A(n_525),
.B(n_418),
.Y(n_786)
);

AOI22xp5_ASAP7_75t_L g787 ( 
.A1(n_506),
.A2(n_212),
.B1(n_424),
.B2(n_435),
.Y(n_787)
);

NAND2xp5_ASAP7_75t_SL g788 ( 
.A(n_697),
.B(n_525),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_642),
.A2(n_650),
.B1(n_697),
.B2(n_643),
.Y(n_789)
);

AO21x1_ASAP7_75t_L g790 ( 
.A1(n_695),
.A2(n_710),
.B(n_654),
.Y(n_790)
);

INVx2_ASAP7_75t_L g791 ( 
.A(n_632),
.Y(n_791)
);

AO21x1_ASAP7_75t_L g792 ( 
.A1(n_695),
.A2(n_506),
.B(n_293),
.Y(n_792)
);

NAND2xp33_ASAP7_75t_L g793 ( 
.A(n_669),
.B(n_572),
.Y(n_793)
);

BUFx6f_ASAP7_75t_L g794 ( 
.A(n_753),
.Y(n_794)
);

INVx2_ASAP7_75t_L g795 ( 
.A(n_632),
.Y(n_795)
);

NAND2xp5_ASAP7_75t_L g796 ( 
.A(n_651),
.B(n_585),
.Y(n_796)
);

CKINVDCx8_ASAP7_75t_R g797 ( 
.A(n_708),
.Y(n_797)
);

NOR2xp33_ASAP7_75t_SL g798 ( 
.A(n_633),
.B(n_613),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_654),
.B(n_585),
.Y(n_799)
);

AOI21xp5_ASAP7_75t_L g800 ( 
.A1(n_727),
.A2(n_488),
.B(n_487),
.Y(n_800)
);

AO21x1_ASAP7_75t_L g801 ( 
.A1(n_667),
.A2(n_293),
.B(n_290),
.Y(n_801)
);

HB1xp67_ASAP7_75t_L g802 ( 
.A(n_645),
.Y(n_802)
);

AND2x2_ASAP7_75t_L g803 ( 
.A(n_668),
.B(n_422),
.Y(n_803)
);

INVx1_ASAP7_75t_L g804 ( 
.A(n_720),
.Y(n_804)
);

INVx2_ASAP7_75t_L g805 ( 
.A(n_640),
.Y(n_805)
);

NOR2xp67_ASAP7_75t_L g806 ( 
.A(n_671),
.B(n_422),
.Y(n_806)
);

INVx3_ASAP7_75t_L g807 ( 
.A(n_753),
.Y(n_807)
);

OAI22xp5_ASAP7_75t_L g808 ( 
.A1(n_670),
.A2(n_696),
.B1(n_667),
.B2(n_628),
.Y(n_808)
);

O2A1O1Ixp33_ASAP7_75t_L g809 ( 
.A1(n_711),
.A2(n_620),
.B(n_270),
.C(n_266),
.Y(n_809)
);

OAI22xp5_ASAP7_75t_L g810 ( 
.A1(n_628),
.A2(n_614),
.B1(n_593),
.B2(n_551),
.Y(n_810)
);

BUFx2_ASAP7_75t_L g811 ( 
.A(n_634),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_L g812 ( 
.A(n_663),
.B(n_614),
.Y(n_812)
);

NAND2xp5_ASAP7_75t_L g813 ( 
.A(n_663),
.B(n_526),
.Y(n_813)
);

AND2x2_ASAP7_75t_L g814 ( 
.A(n_630),
.B(n_422),
.Y(n_814)
);

NOR2xp33_ASAP7_75t_L g815 ( 
.A(n_722),
.B(n_526),
.Y(n_815)
);

AND2x2_ASAP7_75t_L g816 ( 
.A(n_734),
.B(n_424),
.Y(n_816)
);

INVx4_ASAP7_75t_L g817 ( 
.A(n_629),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_653),
.B(n_526),
.Y(n_818)
);

AOI21xp33_ASAP7_75t_L g819 ( 
.A1(n_698),
.A2(n_503),
.B(n_500),
.Y(n_819)
);

HB1xp67_ASAP7_75t_L g820 ( 
.A(n_644),
.Y(n_820)
);

A2O1A1Ixp33_ASAP7_75t_L g821 ( 
.A1(n_756),
.A2(n_424),
.B(n_425),
.C(n_428),
.Y(n_821)
);

BUFx3_ASAP7_75t_L g822 ( 
.A(n_665),
.Y(n_822)
);

BUFx4f_ASAP7_75t_L g823 ( 
.A(n_665),
.Y(n_823)
);

NOR3xp33_ASAP7_75t_L g824 ( 
.A(n_693),
.B(n_270),
.C(n_266),
.Y(n_824)
);

AOI21xp5_ASAP7_75t_L g825 ( 
.A1(n_730),
.A2(n_739),
.B(n_726),
.Y(n_825)
);

A2O1A1Ixp33_ASAP7_75t_L g826 ( 
.A1(n_656),
.A2(n_428),
.B(n_435),
.C(n_430),
.Y(n_826)
);

INVx4_ASAP7_75t_L g827 ( 
.A(n_629),
.Y(n_827)
);

NAND2xp5_ASAP7_75t_L g828 ( 
.A(n_637),
.B(n_680),
.Y(n_828)
);

OR2x2_ASAP7_75t_L g829 ( 
.A(n_664),
.B(n_425),
.Y(n_829)
);

NAND2xp5_ASAP7_75t_L g830 ( 
.A(n_685),
.B(n_538),
.Y(n_830)
);

NAND2xp5_ASAP7_75t_L g831 ( 
.A(n_719),
.B(n_538),
.Y(n_831)
);

AND2x4_ASAP7_75t_L g832 ( 
.A(n_780),
.B(n_543),
.Y(n_832)
);

AOI21xp5_ASAP7_75t_L g833 ( 
.A1(n_692),
.A2(n_552),
.B(n_550),
.Y(n_833)
);

INVx2_ASAP7_75t_L g834 ( 
.A(n_641),
.Y(n_834)
);

AOI21xp5_ASAP7_75t_L g835 ( 
.A1(n_635),
.A2(n_622),
.B(n_612),
.Y(n_835)
);

AOI21xp5_ASAP7_75t_L g836 ( 
.A1(n_712),
.A2(n_690),
.B(n_713),
.Y(n_836)
);

AND2x2_ASAP7_75t_L g837 ( 
.A(n_699),
.B(n_425),
.Y(n_837)
);

OAI21x1_ASAP7_75t_L g838 ( 
.A1(n_763),
.A2(n_512),
.B(n_503),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_694),
.B(n_782),
.Y(n_839)
);

INVx3_ASAP7_75t_L g840 ( 
.A(n_753),
.Y(n_840)
);

NAND2xp5_ASAP7_75t_L g841 ( 
.A(n_782),
.B(n_538),
.Y(n_841)
);

AOI21xp5_ASAP7_75t_L g842 ( 
.A1(n_715),
.A2(n_623),
.B(n_622),
.Y(n_842)
);

INVxp67_ASAP7_75t_SL g843 ( 
.A(n_648),
.Y(n_843)
);

AOI21xp5_ASAP7_75t_L g844 ( 
.A1(n_784),
.A2(n_513),
.B(n_512),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_761),
.B(n_428),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_641),
.Y(n_846)
);

OAI321xp33_ASAP7_75t_L g847 ( 
.A1(n_677),
.A2(n_317),
.A3(n_304),
.B1(n_308),
.B2(n_296),
.C(n_313),
.Y(n_847)
);

NAND2xp5_ASAP7_75t_SL g848 ( 
.A(n_647),
.B(n_525),
.Y(n_848)
);

A2O1A1Ixp33_ASAP7_75t_L g849 ( 
.A1(n_716),
.A2(n_430),
.B(n_435),
.C(n_317),
.Y(n_849)
);

OAI21xp5_ASAP7_75t_L g850 ( 
.A1(n_691),
.A2(n_529),
.B(n_528),
.Y(n_850)
);

AO21x1_ASAP7_75t_L g851 ( 
.A1(n_716),
.A2(n_308),
.B(n_296),
.Y(n_851)
);

AOI21xp5_ASAP7_75t_L g852 ( 
.A1(n_784),
.A2(n_529),
.B(n_528),
.Y(n_852)
);

A2O1A1Ixp33_ASAP7_75t_L g853 ( 
.A1(n_733),
.A2(n_430),
.B(n_304),
.C(n_443),
.Y(n_853)
);

NAND2xp5_ASAP7_75t_L g854 ( 
.A(n_761),
.B(n_541),
.Y(n_854)
);

AOI22xp33_ASAP7_75t_L g855 ( 
.A1(n_627),
.A2(n_437),
.B1(n_431),
.B2(n_443),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_631),
.B(n_431),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_SL g857 ( 
.A(n_647),
.B(n_525),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_636),
.A2(n_755),
.B(n_745),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_745),
.A2(n_755),
.B(n_646),
.Y(n_859)
);

O2A1O1Ixp33_ASAP7_75t_L g860 ( 
.A1(n_660),
.A2(n_672),
.B(n_746),
.C(n_742),
.Y(n_860)
);

INVx1_ASAP7_75t_L g861 ( 
.A(n_720),
.Y(n_861)
);

INVx1_ASAP7_75t_SL g862 ( 
.A(n_707),
.Y(n_862)
);

AOI22xp5_ASAP7_75t_L g863 ( 
.A1(n_688),
.A2(n_714),
.B1(n_669),
.B2(n_737),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_761),
.B(n_541),
.Y(n_864)
);

INVx2_ASAP7_75t_L g865 ( 
.A(n_649),
.Y(n_865)
);

AOI22xp5_ASAP7_75t_L g866 ( 
.A1(n_714),
.A2(n_572),
.B1(n_563),
.B2(n_569),
.Y(n_866)
);

NAND2x1p5_ASAP7_75t_L g867 ( 
.A(n_753),
.B(n_543),
.Y(n_867)
);

NAND2xp5_ASAP7_75t_L g868 ( 
.A(n_644),
.B(n_544),
.Y(n_868)
);

AOI22xp5_ASAP7_75t_L g869 ( 
.A1(n_669),
.A2(n_565),
.B1(n_563),
.B2(n_559),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_649),
.Y(n_870)
);

NOR2xp33_ASAP7_75t_L g871 ( 
.A(n_709),
.B(n_657),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_644),
.B(n_549),
.Y(n_872)
);

NAND2xp5_ASAP7_75t_SL g873 ( 
.A(n_665),
.B(n_629),
.Y(n_873)
);

NOR3xp33_ASAP7_75t_L g874 ( 
.A(n_779),
.B(n_292),
.C(n_299),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_723),
.Y(n_875)
);

INVx2_ASAP7_75t_L g876 ( 
.A(n_659),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_639),
.A2(n_683),
.B(n_749),
.Y(n_877)
);

NOR2xp33_ASAP7_75t_L g878 ( 
.A(n_709),
.B(n_549),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_652),
.A2(n_655),
.B(n_750),
.Y(n_879)
);

NOR2xp33_ASAP7_75t_L g880 ( 
.A(n_631),
.B(n_564),
.Y(n_880)
);

INVx1_ASAP7_75t_L g881 ( 
.A(n_723),
.Y(n_881)
);

INVx3_ASAP7_75t_L g882 ( 
.A(n_758),
.Y(n_882)
);

NAND2xp5_ASAP7_75t_L g883 ( 
.A(n_773),
.B(n_437),
.Y(n_883)
);

AOI21xp5_ASAP7_75t_L g884 ( 
.A1(n_754),
.A2(n_584),
.B(n_564),
.Y(n_884)
);

NAND2xp5_ASAP7_75t_L g885 ( 
.A(n_773),
.B(n_437),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_659),
.Y(n_886)
);

NOR2xp33_ASAP7_75t_L g887 ( 
.A(n_684),
.B(n_686),
.Y(n_887)
);

A2O1A1Ixp33_ASAP7_75t_L g888 ( 
.A1(n_733),
.A2(n_313),
.B(n_275),
.C(n_255),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_661),
.Y(n_889)
);

AOI21xp5_ASAP7_75t_L g890 ( 
.A1(n_786),
.A2(n_584),
.B(n_564),
.Y(n_890)
);

INVx2_ASAP7_75t_L g891 ( 
.A(n_661),
.Y(n_891)
);

AND2x4_ASAP7_75t_L g892 ( 
.A(n_777),
.B(n_543),
.Y(n_892)
);

OAI22xp5_ASAP7_75t_L g893 ( 
.A1(n_725),
.A2(n_584),
.B1(n_305),
.B2(n_303),
.Y(n_893)
);

A2O1A1Ixp33_ASAP7_75t_L g894 ( 
.A1(n_705),
.A2(n_283),
.B(n_315),
.C(n_282),
.Y(n_894)
);

OAI21xp5_ASAP7_75t_L g895 ( 
.A1(n_652),
.A2(n_543),
.B(n_427),
.Y(n_895)
);

NOR2xp33_ASAP7_75t_L g896 ( 
.A(n_702),
.B(n_584),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_718),
.B(n_728),
.Y(n_897)
);

NAND2xp5_ASAP7_75t_L g898 ( 
.A(n_740),
.B(n_285),
.Y(n_898)
);

NAND2xp5_ASAP7_75t_SL g899 ( 
.A(n_758),
.B(n_421),
.Y(n_899)
);

AOI21xp5_ASAP7_75t_L g900 ( 
.A1(n_673),
.A2(n_192),
.B(n_195),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_674),
.A2(n_191),
.B(n_196),
.Y(n_901)
);

NAND2xp5_ASAP7_75t_L g902 ( 
.A(n_752),
.B(n_300),
.Y(n_902)
);

INVx3_ASAP7_75t_L g903 ( 
.A(n_758),
.Y(n_903)
);

NOR3xp33_ASAP7_75t_L g904 ( 
.A(n_759),
.B(n_323),
.C(n_322),
.Y(n_904)
);

O2A1O1Ixp33_ASAP7_75t_L g905 ( 
.A1(n_741),
.A2(n_283),
.B(n_193),
.C(n_16),
.Y(n_905)
);

OAI21xp5_ASAP7_75t_L g906 ( 
.A1(n_655),
.A2(n_427),
.B(n_421),
.Y(n_906)
);

INVx2_ASAP7_75t_L g907 ( 
.A(n_689),
.Y(n_907)
);

NAND2xp5_ASAP7_75t_L g908 ( 
.A(n_762),
.B(n_421),
.Y(n_908)
);

NOR2xp67_ASAP7_75t_L g909 ( 
.A(n_765),
.B(n_421),
.Y(n_909)
);

NOR3xp33_ASAP7_75t_L g910 ( 
.A(n_774),
.B(n_180),
.C(n_318),
.Y(n_910)
);

AOI21xp5_ASAP7_75t_L g911 ( 
.A1(n_676),
.A2(n_172),
.B(n_163),
.Y(n_911)
);

AOI22xp5_ASAP7_75t_L g912 ( 
.A1(n_669),
.A2(n_427),
.B1(n_316),
.B2(n_312),
.Y(n_912)
);

AND2x2_ASAP7_75t_L g913 ( 
.A(n_751),
.B(n_186),
.Y(n_913)
);

NOR3xp33_ASAP7_75t_L g914 ( 
.A(n_743),
.B(n_168),
.C(n_311),
.Y(n_914)
);

NAND2xp5_ASAP7_75t_SL g915 ( 
.A(n_758),
.B(n_421),
.Y(n_915)
);

BUFx2_ASAP7_75t_L g916 ( 
.A(n_634),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_L g917 ( 
.A(n_757),
.B(n_421),
.Y(n_917)
);

NAND2xp5_ASAP7_75t_SL g918 ( 
.A(n_638),
.B(n_421),
.Y(n_918)
);

AO21x1_ASAP7_75t_L g919 ( 
.A1(n_687),
.A2(n_427),
.B(n_421),
.Y(n_919)
);

INVx2_ASAP7_75t_SL g920 ( 
.A(n_658),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_778),
.B(n_421),
.Y(n_921)
);

AND2x4_ASAP7_75t_L g922 ( 
.A(n_703),
.B(n_421),
.Y(n_922)
);

NAND2xp5_ASAP7_75t_L g923 ( 
.A(n_725),
.B(n_427),
.Y(n_923)
);

INVx5_ASAP7_75t_L g924 ( 
.A(n_669),
.Y(n_924)
);

AOI21xp5_ASAP7_75t_L g925 ( 
.A1(n_678),
.A2(n_253),
.B(n_210),
.Y(n_925)
);

NAND2xp5_ASAP7_75t_L g926 ( 
.A(n_731),
.B(n_427),
.Y(n_926)
);

INVx2_ASAP7_75t_L g927 ( 
.A(n_689),
.Y(n_927)
);

NAND2xp33_ASAP7_75t_L g928 ( 
.A(n_731),
.B(n_190),
.Y(n_928)
);

OAI22xp5_ASAP7_75t_L g929 ( 
.A1(n_732),
.A2(n_298),
.B1(n_236),
.B2(n_235),
.Y(n_929)
);

AND2x2_ASAP7_75t_L g930 ( 
.A(n_658),
.B(n_186),
.Y(n_930)
);

AOI21x1_ASAP7_75t_L g931 ( 
.A1(n_770),
.A2(n_404),
.B(n_314),
.Y(n_931)
);

NAND2xp5_ASAP7_75t_L g932 ( 
.A(n_732),
.B(n_259),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_735),
.B(n_259),
.Y(n_933)
);

OAI22xp5_ASAP7_75t_L g934 ( 
.A1(n_735),
.A2(n_244),
.B1(n_302),
.B2(n_297),
.Y(n_934)
);

OAI22xp5_ASAP7_75t_L g935 ( 
.A1(n_748),
.A2(n_767),
.B1(n_679),
.B2(n_682),
.Y(n_935)
);

NAND2x1p5_ASAP7_75t_L g936 ( 
.A(n_764),
.B(n_314),
.Y(n_936)
);

NAND2xp5_ASAP7_75t_L g937 ( 
.A(n_748),
.B(n_259),
.Y(n_937)
);

AOI21xp5_ASAP7_75t_L g938 ( 
.A1(n_770),
.A2(n_254),
.B(n_201),
.Y(n_938)
);

AOI21xp5_ASAP7_75t_L g939 ( 
.A1(n_783),
.A2(n_264),
.B(n_205),
.Y(n_939)
);

NAND3xp33_ASAP7_75t_L g940 ( 
.A(n_666),
.B(n_239),
.C(n_295),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_666),
.A2(n_200),
.B(n_211),
.Y(n_941)
);

INVx1_ASAP7_75t_L g942 ( 
.A(n_767),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_769),
.Y(n_943)
);

AOI21xp5_ASAP7_75t_L g944 ( 
.A1(n_775),
.A2(n_271),
.B(n_215),
.Y(n_944)
);

NOR2xp33_ASAP7_75t_L g945 ( 
.A(n_776),
.B(n_738),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_638),
.A2(n_277),
.B(n_221),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_SL g947 ( 
.A(n_764),
.B(n_314),
.Y(n_947)
);

INVx2_ASAP7_75t_L g948 ( 
.A(n_701),
.Y(n_948)
);

INVx3_ASAP7_75t_L g949 ( 
.A(n_768),
.Y(n_949)
);

NAND2xp5_ASAP7_75t_L g950 ( 
.A(n_675),
.B(n_301),
.Y(n_950)
);

NAND2xp5_ASAP7_75t_L g951 ( 
.A(n_724),
.B(n_301),
.Y(n_951)
);

INVx1_ASAP7_75t_L g952 ( 
.A(n_701),
.Y(n_952)
);

NOR2xp33_ASAP7_75t_L g953 ( 
.A(n_736),
.B(n_268),
.Y(n_953)
);

NAND2xp5_ASAP7_75t_L g954 ( 
.A(n_785),
.B(n_301),
.Y(n_954)
);

NOR2x1_ASAP7_75t_L g955 ( 
.A(n_703),
.B(n_232),
.Y(n_955)
);

AOI21xp5_ASAP7_75t_L g956 ( 
.A1(n_789),
.A2(n_704),
.B(n_700),
.Y(n_956)
);

AOI21xp5_ASAP7_75t_L g957 ( 
.A1(n_836),
.A2(n_662),
.B(n_744),
.Y(n_957)
);

A2O1A1Ixp33_ASAP7_75t_L g958 ( 
.A1(n_808),
.A2(n_681),
.B(n_747),
.C(n_771),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_804),
.Y(n_959)
);

NOR2xp33_ASAP7_75t_L g960 ( 
.A(n_802),
.B(n_703),
.Y(n_960)
);

HB1xp67_ASAP7_75t_L g961 ( 
.A(n_802),
.Y(n_961)
);

INVx1_ASAP7_75t_SL g962 ( 
.A(n_862),
.Y(n_962)
);

AOI21xp5_ASAP7_75t_L g963 ( 
.A1(n_812),
.A2(n_768),
.B(n_729),
.Y(n_963)
);

HB1xp67_ASAP7_75t_L g964 ( 
.A(n_820),
.Y(n_964)
);

AND2x2_ASAP7_75t_L g965 ( 
.A(n_837),
.B(n_721),
.Y(n_965)
);

INVx2_ASAP7_75t_SL g966 ( 
.A(n_811),
.Y(n_966)
);

NAND2xp33_ASAP7_75t_L g967 ( 
.A(n_924),
.B(n_772),
.Y(n_967)
);

OAI22xp5_ASAP7_75t_L g968 ( 
.A1(n_943),
.A2(n_897),
.B1(n_839),
.B2(n_828),
.Y(n_968)
);

NOR2xp33_ASAP7_75t_L g969 ( 
.A(n_945),
.B(n_721),
.Y(n_969)
);

NOR2xp33_ASAP7_75t_R g970 ( 
.A(n_797),
.B(n_706),
.Y(n_970)
);

AND2x2_ASAP7_75t_L g971 ( 
.A(n_930),
.B(n_721),
.Y(n_971)
);

BUFx6f_ASAP7_75t_L g972 ( 
.A(n_823),
.Y(n_972)
);

OAI22xp5_ASAP7_75t_L g973 ( 
.A1(n_863),
.A2(n_787),
.B1(n_766),
.B2(n_760),
.Y(n_973)
);

NOR2xp67_ASAP7_75t_L g974 ( 
.A(n_920),
.B(n_717),
.Y(n_974)
);

INVx2_ASAP7_75t_SL g975 ( 
.A(n_916),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_L g976 ( 
.A(n_945),
.B(n_781),
.Y(n_976)
);

AND2x2_ASAP7_75t_L g977 ( 
.A(n_814),
.B(n_268),
.Y(n_977)
);

BUFx5_ASAP7_75t_L g978 ( 
.A(n_822),
.Y(n_978)
);

NAND2xp5_ASAP7_75t_L g979 ( 
.A(n_803),
.B(n_12),
.Y(n_979)
);

AOI21xp5_ASAP7_75t_L g980 ( 
.A1(n_796),
.A2(n_284),
.B(n_294),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_861),
.Y(n_981)
);

INVx3_ASAP7_75t_L g982 ( 
.A(n_817),
.Y(n_982)
);

BUFx6f_ASAP7_75t_L g983 ( 
.A(n_823),
.Y(n_983)
);

INVx1_ASAP7_75t_L g984 ( 
.A(n_875),
.Y(n_984)
);

NAND2xp5_ASAP7_75t_L g985 ( 
.A(n_820),
.B(n_15),
.Y(n_985)
);

NAND2xp5_ASAP7_75t_SL g986 ( 
.A(n_924),
.B(n_268),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_799),
.A2(n_825),
.B(n_813),
.Y(n_987)
);

AND2x2_ASAP7_75t_L g988 ( 
.A(n_824),
.B(n_16),
.Y(n_988)
);

NOR2xp33_ASAP7_75t_R g989 ( 
.A(n_924),
.B(n_234),
.Y(n_989)
);

O2A1O1Ixp33_ASAP7_75t_SL g990 ( 
.A1(n_848),
.A2(n_18),
.B(n_20),
.C(n_22),
.Y(n_990)
);

OAI21xp33_ASAP7_75t_L g991 ( 
.A1(n_824),
.A2(n_291),
.B(n_288),
.Y(n_991)
);

INVx2_ASAP7_75t_L g992 ( 
.A(n_791),
.Y(n_992)
);

NOR2xp33_ASAP7_75t_L g993 ( 
.A(n_871),
.B(n_238),
.Y(n_993)
);

BUFx6f_ASAP7_75t_L g994 ( 
.A(n_822),
.Y(n_994)
);

O2A1O1Ixp33_ASAP7_75t_L g995 ( 
.A1(n_860),
.A2(n_20),
.B(n_22),
.C(n_23),
.Y(n_995)
);

NOR2xp33_ASAP7_75t_L g996 ( 
.A(n_871),
.B(n_237),
.Y(n_996)
);

AOI22xp33_ASAP7_75t_L g997 ( 
.A1(n_953),
.A2(n_314),
.B1(n_232),
.B2(n_26),
.Y(n_997)
);

NAND2xp5_ASAP7_75t_SL g998 ( 
.A(n_924),
.B(n_314),
.Y(n_998)
);

AOI22xp5_ASAP7_75t_L g999 ( 
.A1(n_914),
.A2(n_232),
.B1(n_25),
.B2(n_26),
.Y(n_999)
);

AND2x2_ASAP7_75t_L g1000 ( 
.A(n_829),
.B(n_24),
.Y(n_1000)
);

BUFx2_ASAP7_75t_L g1001 ( 
.A(n_856),
.Y(n_1001)
);

INVx1_ASAP7_75t_SL g1002 ( 
.A(n_913),
.Y(n_1002)
);

OAI22xp5_ASAP7_75t_L g1003 ( 
.A1(n_843),
.A2(n_232),
.B1(n_31),
.B2(n_33),
.Y(n_1003)
);

NAND2xp5_ASAP7_75t_L g1004 ( 
.A(n_816),
.B(n_24),
.Y(n_1004)
);

OAI21xp5_ASAP7_75t_L g1005 ( 
.A1(n_877),
.A2(n_31),
.B(n_34),
.Y(n_1005)
);

AND2x4_ASAP7_75t_L g1006 ( 
.A(n_817),
.B(n_34),
.Y(n_1006)
);

BUFx6f_ASAP7_75t_L g1007 ( 
.A(n_794),
.Y(n_1007)
);

NOR2xp33_ASAP7_75t_L g1008 ( 
.A(n_954),
.B(n_35),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_SL g1009 ( 
.A(n_806),
.B(n_37),
.Y(n_1009)
);

INVx2_ASAP7_75t_SL g1010 ( 
.A(n_922),
.Y(n_1010)
);

OAI22x1_ASAP7_75t_L g1011 ( 
.A1(n_953),
.A2(n_37),
.B1(n_40),
.B2(n_41),
.Y(n_1011)
);

O2A1O1Ixp33_ASAP7_75t_L g1012 ( 
.A1(n_898),
.A2(n_41),
.B(n_42),
.C(n_47),
.Y(n_1012)
);

A2O1A1Ixp33_ASAP7_75t_L g1013 ( 
.A1(n_888),
.A2(n_49),
.B(n_51),
.C(n_52),
.Y(n_1013)
);

NAND2xp5_ASAP7_75t_L g1014 ( 
.A(n_843),
.B(n_49),
.Y(n_1014)
);

NAND3xp33_ASAP7_75t_L g1015 ( 
.A(n_914),
.B(n_52),
.C(n_53),
.Y(n_1015)
);

BUFx3_ASAP7_75t_L g1016 ( 
.A(n_922),
.Y(n_1016)
);

NAND2xp5_ASAP7_75t_L g1017 ( 
.A(n_881),
.B(n_56),
.Y(n_1017)
);

NAND2xp5_ASAP7_75t_L g1018 ( 
.A(n_942),
.B(n_56),
.Y(n_1018)
);

AND2x6_ASAP7_75t_L g1019 ( 
.A(n_955),
.B(n_794),
.Y(n_1019)
);

NAND2xp5_ASAP7_75t_L g1020 ( 
.A(n_818),
.B(n_57),
.Y(n_1020)
);

OAI21xp33_ASAP7_75t_L g1021 ( 
.A1(n_902),
.A2(n_60),
.B(n_61),
.Y(n_1021)
);

AOI21xp5_ASAP7_75t_L g1022 ( 
.A1(n_884),
.A2(n_793),
.B(n_935),
.Y(n_1022)
);

NAND2xp5_ASAP7_75t_L g1023 ( 
.A(n_896),
.B(n_60),
.Y(n_1023)
);

NOR2xp33_ASAP7_75t_L g1024 ( 
.A(n_798),
.B(n_69),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_952),
.Y(n_1025)
);

AOI21xp5_ASAP7_75t_L g1026 ( 
.A1(n_800),
.A2(n_74),
.B(n_75),
.Y(n_1026)
);

BUFx2_ASAP7_75t_L g1027 ( 
.A(n_949),
.Y(n_1027)
);

NAND2xp5_ASAP7_75t_SL g1028 ( 
.A(n_827),
.B(n_79),
.Y(n_1028)
);

INVx1_ASAP7_75t_L g1029 ( 
.A(n_795),
.Y(n_1029)
);

NAND3xp33_ASAP7_75t_SL g1030 ( 
.A(n_904),
.B(n_104),
.C(n_112),
.Y(n_1030)
);

NAND2xp5_ASAP7_75t_SL g1031 ( 
.A(n_827),
.B(n_117),
.Y(n_1031)
);

NAND2xp5_ASAP7_75t_SL g1032 ( 
.A(n_949),
.B(n_896),
.Y(n_1032)
);

NAND2xp5_ASAP7_75t_L g1033 ( 
.A(n_815),
.B(n_118),
.Y(n_1033)
);

NAND2xp5_ASAP7_75t_L g1034 ( 
.A(n_815),
.B(n_123),
.Y(n_1034)
);

O2A1O1Ixp5_ASAP7_75t_L g1035 ( 
.A1(n_792),
.A2(n_790),
.B(n_801),
.C(n_851),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_835),
.A2(n_125),
.B(n_132),
.Y(n_1036)
);

AOI22xp33_ASAP7_75t_L g1037 ( 
.A1(n_904),
.A2(n_889),
.B1(n_834),
.B2(n_907),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_805),
.Y(n_1038)
);

NAND2xp5_ASAP7_75t_L g1039 ( 
.A(n_841),
.B(n_137),
.Y(n_1039)
);

CKINVDCx5p33_ASAP7_75t_R g1040 ( 
.A(n_880),
.Y(n_1040)
);

NAND2xp5_ASAP7_75t_L g1041 ( 
.A(n_865),
.B(n_145),
.Y(n_1041)
);

NAND2xp5_ASAP7_75t_L g1042 ( 
.A(n_865),
.B(n_870),
.Y(n_1042)
);

O2A1O1Ixp33_ASAP7_75t_L g1043 ( 
.A1(n_888),
.A2(n_874),
.B(n_894),
.C(n_826),
.Y(n_1043)
);

NAND2xp5_ASAP7_75t_L g1044 ( 
.A(n_870),
.B(n_886),
.Y(n_1044)
);

NAND2xp5_ASAP7_75t_L g1045 ( 
.A(n_886),
.B(n_846),
.Y(n_1045)
);

O2A1O1Ixp33_ASAP7_75t_L g1046 ( 
.A1(n_874),
.A2(n_894),
.B(n_826),
.C(n_910),
.Y(n_1046)
);

OAI22xp5_ASAP7_75t_L g1047 ( 
.A1(n_849),
.A2(n_853),
.B1(n_868),
.B2(n_872),
.Y(n_1047)
);

O2A1O1Ixp33_ASAP7_75t_L g1048 ( 
.A1(n_910),
.A2(n_905),
.B(n_809),
.C(n_887),
.Y(n_1048)
);

CKINVDCx5p33_ASAP7_75t_R g1049 ( 
.A(n_880),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_950),
.Y(n_1050)
);

AOI22xp33_ASAP7_75t_L g1051 ( 
.A1(n_876),
.A2(n_948),
.B1(n_927),
.B2(n_891),
.Y(n_1051)
);

AND2x2_ASAP7_75t_L g1052 ( 
.A(n_932),
.B(n_933),
.Y(n_1052)
);

INVx4_ASAP7_75t_L g1053 ( 
.A(n_794),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_937),
.B(n_909),
.Y(n_1054)
);

INVx1_ASAP7_75t_L g1055 ( 
.A(n_883),
.Y(n_1055)
);

INVx2_ASAP7_75t_L g1056 ( 
.A(n_885),
.Y(n_1056)
);

AOI22xp5_ASAP7_75t_L g1057 ( 
.A1(n_928),
.A2(n_934),
.B1(n_929),
.B2(n_887),
.Y(n_1057)
);

BUFx2_ASAP7_75t_L g1058 ( 
.A(n_892),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_845),
.Y(n_1059)
);

OR2x2_ASAP7_75t_L g1060 ( 
.A(n_893),
.B(n_854),
.Y(n_1060)
);

A2O1A1Ixp33_ASAP7_75t_SL g1061 ( 
.A1(n_879),
.A2(n_878),
.B(n_944),
.C(n_911),
.Y(n_1061)
);

BUFx2_ASAP7_75t_L g1062 ( 
.A(n_892),
.Y(n_1062)
);

NOR2xp67_ASAP7_75t_SL g1063 ( 
.A(n_794),
.B(n_847),
.Y(n_1063)
);

OAI22xp5_ASAP7_75t_L g1064 ( 
.A1(n_849),
.A2(n_853),
.B1(n_821),
.B2(n_831),
.Y(n_1064)
);

NOR2xp33_ASAP7_75t_L g1065 ( 
.A(n_830),
.B(n_951),
.Y(n_1065)
);

OR2x6_ASAP7_75t_SL g1066 ( 
.A(n_940),
.B(n_864),
.Y(n_1066)
);

NAND2xp5_ASAP7_75t_L g1067 ( 
.A(n_832),
.B(n_821),
.Y(n_1067)
);

OAI21xp33_ASAP7_75t_L g1068 ( 
.A1(n_939),
.A2(n_941),
.B(n_878),
.Y(n_1068)
);

INVx1_ASAP7_75t_L g1069 ( 
.A(n_908),
.Y(n_1069)
);

INVx2_ASAP7_75t_L g1070 ( 
.A(n_838),
.Y(n_1070)
);

BUFx6f_ASAP7_75t_L g1071 ( 
.A(n_832),
.Y(n_1071)
);

NAND2xp5_ASAP7_75t_SL g1072 ( 
.A(n_807),
.B(n_840),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_L g1073 ( 
.A1(n_842),
.A2(n_858),
.B(n_859),
.Y(n_1073)
);

AOI21xp5_ASAP7_75t_L g1074 ( 
.A1(n_844),
.A2(n_852),
.B(n_890),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_923),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_926),
.Y(n_1076)
);

O2A1O1Ixp33_ASAP7_75t_L g1077 ( 
.A1(n_918),
.A2(n_857),
.B(n_848),
.C(n_810),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_850),
.A2(n_833),
.B(n_788),
.Y(n_1078)
);

O2A1O1Ixp33_ASAP7_75t_L g1079 ( 
.A1(n_857),
.A2(n_925),
.B(n_901),
.C(n_900),
.Y(n_1079)
);

BUFx2_ASAP7_75t_L g1080 ( 
.A(n_936),
.Y(n_1080)
);

A2O1A1Ixp33_ASAP7_75t_L g1081 ( 
.A1(n_866),
.A2(n_819),
.B(n_917),
.C(n_869),
.Y(n_1081)
);

NOR2xp33_ASAP7_75t_L g1082 ( 
.A(n_873),
.B(n_921),
.Y(n_1082)
);

NAND2xp5_ASAP7_75t_L g1083 ( 
.A(n_855),
.B(n_903),
.Y(n_1083)
);

BUFx2_ASAP7_75t_L g1084 ( 
.A(n_936),
.Y(n_1084)
);

OAI22xp5_ASAP7_75t_SL g1085 ( 
.A1(n_912),
.A2(n_807),
.B1(n_903),
.B2(n_840),
.Y(n_1085)
);

NAND2xp5_ASAP7_75t_L g1086 ( 
.A(n_855),
.B(n_882),
.Y(n_1086)
);

OAI22xp5_ASAP7_75t_L g1087 ( 
.A1(n_882),
.A2(n_906),
.B1(n_895),
.B2(n_899),
.Y(n_1087)
);

NAND2xp5_ASAP7_75t_L g1088 ( 
.A(n_867),
.B(n_899),
.Y(n_1088)
);

INVx4_ASAP7_75t_L g1089 ( 
.A(n_867),
.Y(n_1089)
);

NOR3xp33_ASAP7_75t_L g1090 ( 
.A(n_946),
.B(n_915),
.C(n_938),
.Y(n_1090)
);

BUFx2_ASAP7_75t_L g1091 ( 
.A(n_919),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_947),
.Y(n_1092)
);

NOR2xp67_ASAP7_75t_L g1093 ( 
.A(n_947),
.B(n_931),
.Y(n_1093)
);

NAND2xp5_ASAP7_75t_L g1094 ( 
.A(n_839),
.B(n_539),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_804),
.Y(n_1095)
);

INVx8_ASAP7_75t_L g1096 ( 
.A(n_924),
.Y(n_1096)
);

AO32x1_ASAP7_75t_L g1097 ( 
.A1(n_935),
.A2(n_893),
.A3(n_804),
.B1(n_881),
.B2(n_875),
.Y(n_1097)
);

NAND2xp5_ASAP7_75t_L g1098 ( 
.A(n_839),
.B(n_539),
.Y(n_1098)
);

HB1xp67_ASAP7_75t_L g1099 ( 
.A(n_961),
.Y(n_1099)
);

NAND2xp5_ASAP7_75t_L g1100 ( 
.A(n_1094),
.B(n_1098),
.Y(n_1100)
);

INVx6_ASAP7_75t_L g1101 ( 
.A(n_972),
.Y(n_1101)
);

NOR2xp33_ASAP7_75t_L g1102 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1102)
);

OR2x2_ASAP7_75t_L g1103 ( 
.A(n_1002),
.B(n_962),
.Y(n_1103)
);

AOI22xp33_ASAP7_75t_L g1104 ( 
.A1(n_1008),
.A2(n_988),
.B1(n_977),
.B2(n_1024),
.Y(n_1104)
);

AO32x2_ASAP7_75t_L g1105 ( 
.A1(n_968),
.A2(n_1003),
.A3(n_1064),
.B1(n_1047),
.B2(n_973),
.Y(n_1105)
);

BUFx3_ASAP7_75t_L g1106 ( 
.A(n_966),
.Y(n_1106)
);

AOI21xp5_ASAP7_75t_L g1107 ( 
.A1(n_987),
.A2(n_956),
.B(n_968),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_1033),
.A2(n_1034),
.B(n_1039),
.Y(n_1108)
);

AOI21xp5_ASAP7_75t_SL g1109 ( 
.A1(n_1081),
.A2(n_976),
.B(n_1067),
.Y(n_1109)
);

INVx2_ASAP7_75t_SL g1110 ( 
.A(n_970),
.Y(n_1110)
);

AO31x2_ASAP7_75t_L g1111 ( 
.A1(n_1070),
.A2(n_1091),
.A3(n_1064),
.B(n_1078),
.Y(n_1111)
);

BUFx10_ASAP7_75t_L g1112 ( 
.A(n_1006),
.Y(n_1112)
);

NAND2xp5_ASAP7_75t_L g1113 ( 
.A(n_964),
.B(n_1052),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_959),
.Y(n_1114)
);

OAI21xp5_ASAP7_75t_L g1115 ( 
.A1(n_1035),
.A2(n_973),
.B(n_957),
.Y(n_1115)
);

AND2x2_ASAP7_75t_L g1116 ( 
.A(n_1000),
.B(n_960),
.Y(n_1116)
);

AO22x2_ASAP7_75t_L g1117 ( 
.A1(n_1003),
.A2(n_1005),
.B1(n_1015),
.B2(n_1069),
.Y(n_1117)
);

BUFx12f_ASAP7_75t_L g1118 ( 
.A(n_975),
.Y(n_1118)
);

OAI22x1_ASAP7_75t_L g1119 ( 
.A1(n_999),
.A2(n_1001),
.B1(n_969),
.B2(n_1057),
.Y(n_1119)
);

AOI21xp5_ASAP7_75t_L g1120 ( 
.A1(n_1039),
.A2(n_963),
.B(n_1061),
.Y(n_1120)
);

AOI21xp5_ASAP7_75t_L g1121 ( 
.A1(n_1079),
.A2(n_1077),
.B(n_1068),
.Y(n_1121)
);

INVx1_ASAP7_75t_L g1122 ( 
.A(n_981),
.Y(n_1122)
);

NAND2xp5_ASAP7_75t_L g1123 ( 
.A(n_1059),
.B(n_965),
.Y(n_1123)
);

AOI21xp5_ASAP7_75t_L g1124 ( 
.A1(n_1014),
.A2(n_1036),
.B(n_1026),
.Y(n_1124)
);

INVx3_ASAP7_75t_L g1125 ( 
.A(n_1089),
.Y(n_1125)
);

NOR2xp67_ASAP7_75t_L g1126 ( 
.A(n_1053),
.B(n_982),
.Y(n_1126)
);

NOR2xp33_ASAP7_75t_L g1127 ( 
.A(n_1050),
.B(n_1010),
.Y(n_1127)
);

AND2x2_ASAP7_75t_L g1128 ( 
.A(n_1016),
.B(n_971),
.Y(n_1128)
);

BUFx6f_ASAP7_75t_L g1129 ( 
.A(n_972),
.Y(n_1129)
);

INVx1_ASAP7_75t_SL g1130 ( 
.A(n_1058),
.Y(n_1130)
);

INVx3_ASAP7_75t_L g1131 ( 
.A(n_1096),
.Y(n_1131)
);

INVx1_ASAP7_75t_L g1132 ( 
.A(n_984),
.Y(n_1132)
);

NAND2xp5_ASAP7_75t_L g1133 ( 
.A(n_1062),
.B(n_993),
.Y(n_1133)
);

A2O1A1Ixp33_ASAP7_75t_L g1134 ( 
.A1(n_1046),
.A2(n_1043),
.B(n_1048),
.C(n_1021),
.Y(n_1134)
);

AOI21xp5_ASAP7_75t_SL g1135 ( 
.A1(n_1060),
.A2(n_1082),
.B(n_1014),
.Y(n_1135)
);

NAND2xp5_ASAP7_75t_L g1136 ( 
.A(n_996),
.B(n_1065),
.Y(n_1136)
);

O2A1O1Ixp5_ASAP7_75t_SL g1137 ( 
.A1(n_1005),
.A2(n_1092),
.B(n_1009),
.C(n_1032),
.Y(n_1137)
);

INVx2_ASAP7_75t_L g1138 ( 
.A(n_992),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_1047),
.A2(n_1041),
.A3(n_1042),
.B(n_1044),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1023),
.A2(n_1020),
.B(n_1087),
.Y(n_1140)
);

INVx1_ASAP7_75t_SL g1141 ( 
.A(n_1027),
.Y(n_1141)
);

AOI21xp5_ASAP7_75t_L g1142 ( 
.A1(n_1023),
.A2(n_1020),
.B(n_1087),
.Y(n_1142)
);

OAI21x1_ASAP7_75t_L g1143 ( 
.A1(n_1041),
.A2(n_1093),
.B(n_1042),
.Y(n_1143)
);

BUFx12f_ASAP7_75t_L g1144 ( 
.A(n_972),
.Y(n_1144)
);

OAI21x1_ASAP7_75t_L g1145 ( 
.A1(n_1088),
.A2(n_1086),
.B(n_1083),
.Y(n_1145)
);

AOI21xp5_ASAP7_75t_L g1146 ( 
.A1(n_958),
.A2(n_1096),
.B(n_1090),
.Y(n_1146)
);

AOI22xp33_ASAP7_75t_L g1147 ( 
.A1(n_991),
.A2(n_997),
.B1(n_1054),
.B2(n_1056),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_L g1148 ( 
.A1(n_1096),
.A2(n_1083),
.B(n_1075),
.Y(n_1148)
);

AO21x1_ASAP7_75t_L g1149 ( 
.A1(n_995),
.A2(n_1012),
.B(n_1018),
.Y(n_1149)
);

INVx1_ASAP7_75t_L g1150 ( 
.A(n_1095),
.Y(n_1150)
);

NAND2xp5_ASAP7_75t_L g1151 ( 
.A(n_1071),
.B(n_979),
.Y(n_1151)
);

OAI21xp5_ASAP7_75t_L g1152 ( 
.A1(n_1004),
.A2(n_980),
.B(n_985),
.Y(n_1152)
);

AOI21xp5_ASAP7_75t_L g1153 ( 
.A1(n_1076),
.A2(n_1028),
.B(n_1031),
.Y(n_1153)
);

A2O1A1Ixp33_ASAP7_75t_L g1154 ( 
.A1(n_1013),
.A2(n_1063),
.B(n_1017),
.C(n_1018),
.Y(n_1154)
);

NOR2xp33_ASAP7_75t_SL g1155 ( 
.A(n_1006),
.B(n_1030),
.Y(n_1155)
);

OAI21xp5_ASAP7_75t_L g1156 ( 
.A1(n_1017),
.A2(n_1055),
.B(n_1037),
.Y(n_1156)
);

AOI22xp33_ASAP7_75t_L g1157 ( 
.A1(n_1029),
.A2(n_1038),
.B1(n_1011),
.B2(n_1025),
.Y(n_1157)
);

AOI21xp5_ASAP7_75t_L g1158 ( 
.A1(n_1085),
.A2(n_1097),
.B(n_1072),
.Y(n_1158)
);

INVx1_ASAP7_75t_L g1159 ( 
.A(n_1045),
.Y(n_1159)
);

OAI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_998),
.A2(n_1045),
.B(n_1051),
.Y(n_1160)
);

AOI221xp5_ASAP7_75t_SL g1161 ( 
.A1(n_986),
.A2(n_967),
.B1(n_990),
.B2(n_994),
.C(n_1007),
.Y(n_1161)
);

NAND2xp5_ASAP7_75t_L g1162 ( 
.A(n_1071),
.B(n_983),
.Y(n_1162)
);

INVx1_ASAP7_75t_SL g1163 ( 
.A(n_994),
.Y(n_1163)
);

AOI21xp5_ASAP7_75t_L g1164 ( 
.A1(n_1097),
.A2(n_982),
.B(n_1007),
.Y(n_1164)
);

AOI221x1_ASAP7_75t_L g1165 ( 
.A1(n_1053),
.A2(n_994),
.B1(n_1097),
.B2(n_1007),
.C(n_1066),
.Y(n_1165)
);

BUFx6f_ASAP7_75t_L g1166 ( 
.A(n_983),
.Y(n_1166)
);

OAI22xp5_ASAP7_75t_L g1167 ( 
.A1(n_974),
.A2(n_983),
.B1(n_1080),
.B2(n_1084),
.Y(n_1167)
);

AOI21xp5_ASAP7_75t_L g1168 ( 
.A1(n_978),
.A2(n_1019),
.B(n_989),
.Y(n_1168)
);

OR2x2_ASAP7_75t_L g1169 ( 
.A(n_978),
.B(n_1019),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_978),
.A2(n_987),
.B(n_1022),
.Y(n_1170)
);

BUFx6f_ASAP7_75t_L g1171 ( 
.A(n_1019),
.Y(n_1171)
);

NAND2xp5_ASAP7_75t_L g1172 ( 
.A(n_978),
.B(n_1019),
.Y(n_1172)
);

INVx3_ASAP7_75t_L g1173 ( 
.A(n_1019),
.Y(n_1173)
);

AND2x2_ASAP7_75t_L g1174 ( 
.A(n_978),
.B(n_664),
.Y(n_1174)
);

AND2x2_ASAP7_75t_L g1175 ( 
.A(n_988),
.B(n_664),
.Y(n_1175)
);

INVx4_ASAP7_75t_L g1176 ( 
.A(n_972),
.Y(n_1176)
);

BUFx4_ASAP7_75t_SL g1177 ( 
.A(n_1040),
.Y(n_1177)
);

NOR2xp67_ASAP7_75t_L g1178 ( 
.A(n_968),
.B(n_924),
.Y(n_1178)
);

BUFx2_ASAP7_75t_L g1179 ( 
.A(n_970),
.Y(n_1179)
);

A2O1A1Ixp33_ASAP7_75t_L g1180 ( 
.A1(n_1008),
.A2(n_663),
.B(n_1046),
.C(n_667),
.Y(n_1180)
);

AOI21xp5_ASAP7_75t_L g1181 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1181)
);

BUFx6f_ASAP7_75t_L g1182 ( 
.A(n_972),
.Y(n_1182)
);

OAI22xp5_ASAP7_75t_L g1183 ( 
.A1(n_1057),
.A2(n_668),
.B1(n_671),
.B2(n_711),
.Y(n_1183)
);

NAND2xp5_ASAP7_75t_L g1184 ( 
.A(n_1094),
.B(n_668),
.Y(n_1184)
);

OAI21xp5_ASAP7_75t_L g1185 ( 
.A1(n_968),
.A2(n_654),
.B(n_651),
.Y(n_1185)
);

AOI221xp5_ASAP7_75t_SL g1186 ( 
.A1(n_995),
.A2(n_1005),
.B1(n_1003),
.B2(n_1046),
.C(n_1013),
.Y(n_1186)
);

CKINVDCx11_ASAP7_75t_R g1187 ( 
.A(n_1066),
.Y(n_1187)
);

AOI21xp5_ASAP7_75t_SL g1188 ( 
.A1(n_968),
.A2(n_789),
.B(n_808),
.Y(n_1188)
);

BUFx10_ASAP7_75t_L g1189 ( 
.A(n_1006),
.Y(n_1189)
);

AOI21xp5_ASAP7_75t_L g1190 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1190)
);

AOI21xp5_ASAP7_75t_L g1191 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1191)
);

NAND2xp5_ASAP7_75t_SL g1192 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1192)
);

OAI22xp5_ASAP7_75t_L g1193 ( 
.A1(n_1057),
.A2(n_668),
.B1(n_671),
.B2(n_711),
.Y(n_1193)
);

AOI21xp5_ASAP7_75t_L g1194 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1194)
);

INVx1_ASAP7_75t_L g1195 ( 
.A(n_959),
.Y(n_1195)
);

O2A1O1Ixp33_ASAP7_75t_SL g1196 ( 
.A1(n_1061),
.A2(n_808),
.B(n_1020),
.C(n_812),
.Y(n_1196)
);

AND2x2_ASAP7_75t_SL g1197 ( 
.A(n_1024),
.B(n_988),
.Y(n_1197)
);

NAND2xp5_ASAP7_75t_SL g1198 ( 
.A(n_1040),
.B(n_1049),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_959),
.Y(n_1199)
);

INVx2_ASAP7_75t_SL g1200 ( 
.A(n_970),
.Y(n_1200)
);

INVx5_ASAP7_75t_L g1201 ( 
.A(n_972),
.Y(n_1201)
);

BUFx6f_ASAP7_75t_L g1202 ( 
.A(n_972),
.Y(n_1202)
);

NOR2xp33_ASAP7_75t_L g1203 ( 
.A(n_1040),
.B(n_668),
.Y(n_1203)
);

INVx1_ASAP7_75t_L g1204 ( 
.A(n_959),
.Y(n_1204)
);

OAI22x1_ASAP7_75t_L g1205 ( 
.A1(n_999),
.A2(n_1024),
.B1(n_546),
.B2(n_671),
.Y(n_1205)
);

NAND2xp5_ASAP7_75t_L g1206 ( 
.A(n_1094),
.B(n_668),
.Y(n_1206)
);

OAI21xp33_ASAP7_75t_L g1207 ( 
.A1(n_1005),
.A2(n_671),
.B(n_668),
.Y(n_1207)
);

AOI21xp5_ASAP7_75t_L g1208 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_959),
.Y(n_1209)
);

AOI21xp5_ASAP7_75t_SL g1210 ( 
.A1(n_968),
.A2(n_789),
.B(n_808),
.Y(n_1210)
);

NAND2xp5_ASAP7_75t_L g1211 ( 
.A(n_1094),
.B(n_668),
.Y(n_1211)
);

INVxp67_ASAP7_75t_SL g1212 ( 
.A(n_961),
.Y(n_1212)
);

INVx3_ASAP7_75t_L g1213 ( 
.A(n_1089),
.Y(n_1213)
);

A2O1A1Ixp33_ASAP7_75t_L g1214 ( 
.A1(n_1008),
.A2(n_663),
.B(n_1046),
.C(n_667),
.Y(n_1214)
);

NOR2xp67_ASAP7_75t_SL g1215 ( 
.A(n_972),
.B(n_797),
.Y(n_1215)
);

AOI21xp5_ASAP7_75t_L g1216 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1216)
);

AND2x4_ASAP7_75t_L g1217 ( 
.A(n_1016),
.B(n_1010),
.Y(n_1217)
);

BUFx10_ASAP7_75t_L g1218 ( 
.A(n_1006),
.Y(n_1218)
);

NAND2xp5_ASAP7_75t_L g1219 ( 
.A(n_1094),
.B(n_668),
.Y(n_1219)
);

INVxp67_ASAP7_75t_SL g1220 ( 
.A(n_961),
.Y(n_1220)
);

AOI21xp5_ASAP7_75t_L g1221 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_962),
.Y(n_1222)
);

A2O1A1Ixp33_ASAP7_75t_L g1223 ( 
.A1(n_1008),
.A2(n_663),
.B(n_1046),
.C(n_667),
.Y(n_1223)
);

BUFx2_ASAP7_75t_L g1224 ( 
.A(n_970),
.Y(n_1224)
);

OR2x2_ASAP7_75t_L g1225 ( 
.A(n_961),
.B(n_802),
.Y(n_1225)
);

NOR2xp67_ASAP7_75t_L g1226 ( 
.A(n_968),
.B(n_924),
.Y(n_1226)
);

OAI21x1_ASAP7_75t_L g1227 ( 
.A1(n_1022),
.A2(n_1073),
.B(n_1074),
.Y(n_1227)
);

NOR2xp33_ASAP7_75t_L g1228 ( 
.A(n_1040),
.B(n_668),
.Y(n_1228)
);

O2A1O1Ixp33_ASAP7_75t_L g1229 ( 
.A1(n_1008),
.A2(n_668),
.B(n_671),
.C(n_711),
.Y(n_1229)
);

AOI21xp5_ASAP7_75t_L g1230 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1230)
);

O2A1O1Ixp33_ASAP7_75t_SL g1231 ( 
.A1(n_1061),
.A2(n_808),
.B(n_1020),
.C(n_812),
.Y(n_1231)
);

INVx1_ASAP7_75t_L g1232 ( 
.A(n_959),
.Y(n_1232)
);

AOI21xp5_ASAP7_75t_L g1233 ( 
.A1(n_987),
.A2(n_1022),
.B(n_956),
.Y(n_1233)
);

A2O1A1Ixp33_ASAP7_75t_L g1234 ( 
.A1(n_1008),
.A2(n_663),
.B(n_1046),
.C(n_667),
.Y(n_1234)
);

OAI21x1_ASAP7_75t_L g1235 ( 
.A1(n_1022),
.A2(n_1073),
.B(n_1074),
.Y(n_1235)
);

NAND3xp33_ASAP7_75t_L g1236 ( 
.A(n_995),
.B(n_671),
.C(n_668),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_972),
.Y(n_1237)
);

INVx8_ASAP7_75t_L g1238 ( 
.A(n_1096),
.Y(n_1238)
);

OAI21xp5_ASAP7_75t_L g1239 ( 
.A1(n_968),
.A2(n_654),
.B(n_651),
.Y(n_1239)
);

CKINVDCx20_ASAP7_75t_R g1240 ( 
.A(n_1179),
.Y(n_1240)
);

BUFx4f_ASAP7_75t_SL g1241 ( 
.A(n_1144),
.Y(n_1241)
);

AOI22xp33_ASAP7_75t_L g1242 ( 
.A1(n_1197),
.A2(n_1104),
.B1(n_1205),
.B2(n_1187),
.Y(n_1242)
);

BUFx2_ASAP7_75t_L g1243 ( 
.A(n_1225),
.Y(n_1243)
);

INVx2_ASAP7_75t_L g1244 ( 
.A(n_1138),
.Y(n_1244)
);

INVx1_ASAP7_75t_L g1245 ( 
.A(n_1114),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_1122),
.Y(n_1246)
);

CKINVDCx11_ASAP7_75t_R g1247 ( 
.A(n_1112),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1132),
.Y(n_1248)
);

BUFx2_ASAP7_75t_SL g1249 ( 
.A(n_1110),
.Y(n_1249)
);

INVx1_ASAP7_75t_SL g1250 ( 
.A(n_1177),
.Y(n_1250)
);

BUFx3_ASAP7_75t_L g1251 ( 
.A(n_1224),
.Y(n_1251)
);

BUFx2_ASAP7_75t_L g1252 ( 
.A(n_1118),
.Y(n_1252)
);

AOI21xp5_ASAP7_75t_L g1253 ( 
.A1(n_1108),
.A2(n_1210),
.B(n_1188),
.Y(n_1253)
);

INVx1_ASAP7_75t_L g1254 ( 
.A(n_1150),
.Y(n_1254)
);

BUFx12f_ASAP7_75t_L g1255 ( 
.A(n_1200),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1195),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1199),
.Y(n_1257)
);

AOI22xp33_ASAP7_75t_L g1258 ( 
.A1(n_1136),
.A2(n_1175),
.B1(n_1207),
.B2(n_1117),
.Y(n_1258)
);

INVx1_ASAP7_75t_L g1259 ( 
.A(n_1204),
.Y(n_1259)
);

BUFx8_ASAP7_75t_L g1260 ( 
.A(n_1116),
.Y(n_1260)
);

INVx1_ASAP7_75t_L g1261 ( 
.A(n_1209),
.Y(n_1261)
);

AOI22xp33_ASAP7_75t_L g1262 ( 
.A1(n_1207),
.A2(n_1117),
.B1(n_1239),
.B2(n_1185),
.Y(n_1262)
);

BUFx2_ASAP7_75t_SL g1263 ( 
.A(n_1201),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1180),
.A2(n_1234),
.B1(n_1223),
.B2(n_1214),
.Y(n_1264)
);

AOI22xp33_ASAP7_75t_SL g1265 ( 
.A1(n_1155),
.A2(n_1115),
.B1(n_1193),
.B2(n_1183),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1232),
.Y(n_1266)
);

CKINVDCx11_ASAP7_75t_R g1267 ( 
.A(n_1112),
.Y(n_1267)
);

CKINVDCx11_ASAP7_75t_R g1268 ( 
.A(n_1189),
.Y(n_1268)
);

OAI22xp33_ASAP7_75t_R g1269 ( 
.A1(n_1203),
.A2(n_1228),
.B1(n_1102),
.B2(n_1099),
.Y(n_1269)
);

INVx6_ASAP7_75t_L g1270 ( 
.A(n_1201),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1159),
.Y(n_1271)
);

INVx2_ASAP7_75t_SL g1272 ( 
.A(n_1101),
.Y(n_1272)
);

CKINVDCx6p67_ASAP7_75t_R g1273 ( 
.A(n_1106),
.Y(n_1273)
);

CKINVDCx20_ASAP7_75t_R g1274 ( 
.A(n_1192),
.Y(n_1274)
);

AOI22xp33_ASAP7_75t_L g1275 ( 
.A1(n_1119),
.A2(n_1236),
.B1(n_1149),
.B2(n_1157),
.Y(n_1275)
);

AOI22xp33_ASAP7_75t_L g1276 ( 
.A1(n_1236),
.A2(n_1115),
.B1(n_1156),
.B2(n_1147),
.Y(n_1276)
);

AOI22xp33_ASAP7_75t_SL g1277 ( 
.A1(n_1155),
.A2(n_1174),
.B1(n_1156),
.B2(n_1105),
.Y(n_1277)
);

OAI22xp33_ASAP7_75t_L g1278 ( 
.A1(n_1113),
.A2(n_1100),
.B1(n_1133),
.B2(n_1219),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_L g1279 ( 
.A(n_1184),
.B(n_1206),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_1198),
.Y(n_1280)
);

OAI22xp33_ASAP7_75t_SL g1281 ( 
.A1(n_1103),
.A2(n_1222),
.B1(n_1123),
.B2(n_1151),
.Y(n_1281)
);

INVx1_ASAP7_75t_L g1282 ( 
.A(n_1212),
.Y(n_1282)
);

AOI22xp33_ASAP7_75t_L g1283 ( 
.A1(n_1152),
.A2(n_1140),
.B1(n_1142),
.B2(n_1211),
.Y(n_1283)
);

BUFx3_ASAP7_75t_L g1284 ( 
.A(n_1101),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1220),
.Y(n_1285)
);

AOI22xp33_ASAP7_75t_L g1286 ( 
.A1(n_1222),
.A2(n_1128),
.B1(n_1127),
.B2(n_1130),
.Y(n_1286)
);

NAND2xp5_ASAP7_75t_L g1287 ( 
.A(n_1130),
.B(n_1141),
.Y(n_1287)
);

INVx1_ASAP7_75t_SL g1288 ( 
.A(n_1141),
.Y(n_1288)
);

AOI22xp5_ASAP7_75t_L g1289 ( 
.A1(n_1186),
.A2(n_1134),
.B1(n_1215),
.B2(n_1218),
.Y(n_1289)
);

AOI22xp33_ASAP7_75t_SL g1290 ( 
.A1(n_1105),
.A2(n_1186),
.B1(n_1189),
.B2(n_1218),
.Y(n_1290)
);

OAI22x1_ASAP7_75t_L g1291 ( 
.A1(n_1217),
.A2(n_1163),
.B1(n_1105),
.B2(n_1173),
.Y(n_1291)
);

OAI22xp5_ASAP7_75t_SL g1292 ( 
.A1(n_1229),
.A2(n_1176),
.B1(n_1162),
.B2(n_1202),
.Y(n_1292)
);

AOI22xp33_ASAP7_75t_L g1293 ( 
.A1(n_1178),
.A2(n_1226),
.B1(n_1217),
.B2(n_1158),
.Y(n_1293)
);

CKINVDCx20_ASAP7_75t_R g1294 ( 
.A(n_1163),
.Y(n_1294)
);

INVx6_ASAP7_75t_L g1295 ( 
.A(n_1238),
.Y(n_1295)
);

BUFx2_ASAP7_75t_L g1296 ( 
.A(n_1129),
.Y(n_1296)
);

CKINVDCx5p33_ASAP7_75t_R g1297 ( 
.A(n_1129),
.Y(n_1297)
);

AOI22xp33_ASAP7_75t_L g1298 ( 
.A1(n_1178),
.A2(n_1226),
.B1(n_1121),
.B2(n_1146),
.Y(n_1298)
);

OAI22xp5_ASAP7_75t_L g1299 ( 
.A1(n_1154),
.A2(n_1135),
.B1(n_1109),
.B2(n_1107),
.Y(n_1299)
);

INVx4_ASAP7_75t_SL g1300 ( 
.A(n_1171),
.Y(n_1300)
);

BUFx8_ASAP7_75t_L g1301 ( 
.A(n_1129),
.Y(n_1301)
);

CKINVDCx20_ASAP7_75t_R g1302 ( 
.A(n_1166),
.Y(n_1302)
);

AOI22xp33_ASAP7_75t_L g1303 ( 
.A1(n_1160),
.A2(n_1145),
.B1(n_1167),
.B2(n_1148),
.Y(n_1303)
);

INVx6_ASAP7_75t_L g1304 ( 
.A(n_1238),
.Y(n_1304)
);

CKINVDCx20_ASAP7_75t_R g1305 ( 
.A(n_1166),
.Y(n_1305)
);

AOI22xp33_ASAP7_75t_L g1306 ( 
.A1(n_1160),
.A2(n_1124),
.B1(n_1202),
.B2(n_1166),
.Y(n_1306)
);

AOI22xp33_ASAP7_75t_L g1307 ( 
.A1(n_1182),
.A2(n_1237),
.B1(n_1202),
.B2(n_1153),
.Y(n_1307)
);

CKINVDCx20_ASAP7_75t_R g1308 ( 
.A(n_1182),
.Y(n_1308)
);

AOI22xp5_ASAP7_75t_L g1309 ( 
.A1(n_1161),
.A2(n_1176),
.B1(n_1182),
.B2(n_1237),
.Y(n_1309)
);

OAI22xp5_ASAP7_75t_L g1310 ( 
.A1(n_1126),
.A2(n_1131),
.B1(n_1216),
.B2(n_1208),
.Y(n_1310)
);

INVx6_ASAP7_75t_L g1311 ( 
.A(n_1238),
.Y(n_1311)
);

AOI22xp33_ASAP7_75t_L g1312 ( 
.A1(n_1237),
.A2(n_1168),
.B1(n_1164),
.B2(n_1213),
.Y(n_1312)
);

INVx6_ASAP7_75t_L g1313 ( 
.A(n_1169),
.Y(n_1313)
);

BUFx2_ASAP7_75t_SL g1314 ( 
.A(n_1126),
.Y(n_1314)
);

AOI22xp33_ASAP7_75t_L g1315 ( 
.A1(n_1125),
.A2(n_1172),
.B1(n_1120),
.B2(n_1143),
.Y(n_1315)
);

NAND2xp5_ASAP7_75t_L g1316 ( 
.A(n_1139),
.B(n_1131),
.Y(n_1316)
);

INVx4_ASAP7_75t_L g1317 ( 
.A(n_1161),
.Y(n_1317)
);

CKINVDCx11_ASAP7_75t_R g1318 ( 
.A(n_1137),
.Y(n_1318)
);

OAI22xp5_ASAP7_75t_SL g1319 ( 
.A1(n_1165),
.A2(n_1231),
.B1(n_1196),
.B2(n_1139),
.Y(n_1319)
);

CKINVDCx6p67_ASAP7_75t_R g1320 ( 
.A(n_1139),
.Y(n_1320)
);

NOR2x1_ASAP7_75t_R g1321 ( 
.A(n_1111),
.B(n_1170),
.Y(n_1321)
);

INVx1_ASAP7_75t_SL g1322 ( 
.A(n_1181),
.Y(n_1322)
);

OAI22xp33_ASAP7_75t_L g1323 ( 
.A1(n_1190),
.A2(n_1233),
.B1(n_1221),
.B2(n_1230),
.Y(n_1323)
);

BUFx2_ASAP7_75t_SL g1324 ( 
.A(n_1191),
.Y(n_1324)
);

BUFx12f_ASAP7_75t_L g1325 ( 
.A(n_1194),
.Y(n_1325)
);

INVx6_ASAP7_75t_L g1326 ( 
.A(n_1227),
.Y(n_1326)
);

INVx3_ASAP7_75t_SL g1327 ( 
.A(n_1235),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1114),
.Y(n_1328)
);

OAI22xp33_ASAP7_75t_L g1329 ( 
.A1(n_1136),
.A2(n_499),
.B1(n_999),
.B2(n_1003),
.Y(n_1329)
);

AOI22xp33_ASAP7_75t_SL g1330 ( 
.A1(n_1197),
.A2(n_348),
.B1(n_1136),
.B2(n_1117),
.Y(n_1330)
);

BUFx3_ASAP7_75t_L g1331 ( 
.A(n_1144),
.Y(n_1331)
);

OAI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_1136),
.A2(n_1180),
.B1(n_1223),
.B2(n_1214),
.Y(n_1332)
);

AND2x2_ASAP7_75t_L g1333 ( 
.A(n_1175),
.B(n_1116),
.Y(n_1333)
);

HB1xp67_ASAP7_75t_L g1334 ( 
.A(n_1111),
.Y(n_1334)
);

AOI22xp33_ASAP7_75t_L g1335 ( 
.A1(n_1197),
.A2(n_1104),
.B1(n_1205),
.B2(n_1187),
.Y(n_1335)
);

AOI22xp5_ASAP7_75t_L g1336 ( 
.A1(n_1197),
.A2(n_1136),
.B1(n_547),
.B2(n_671),
.Y(n_1336)
);

BUFx4f_ASAP7_75t_SL g1337 ( 
.A(n_1144),
.Y(n_1337)
);

OAI22x1_ASAP7_75t_L g1338 ( 
.A1(n_1136),
.A2(n_1024),
.B1(n_999),
.B2(n_1175),
.Y(n_1338)
);

OAI22xp5_ASAP7_75t_L g1339 ( 
.A1(n_1136),
.A2(n_1180),
.B1(n_1223),
.B2(n_1214),
.Y(n_1339)
);

AOI22xp33_ASAP7_75t_SL g1340 ( 
.A1(n_1197),
.A2(n_348),
.B1(n_1136),
.B2(n_1117),
.Y(n_1340)
);

OAI22xp5_ASAP7_75t_L g1341 ( 
.A1(n_1136),
.A2(n_1180),
.B1(n_1223),
.B2(n_1214),
.Y(n_1341)
);

AOI22xp33_ASAP7_75t_L g1342 ( 
.A1(n_1197),
.A2(n_1104),
.B1(n_1205),
.B2(n_1187),
.Y(n_1342)
);

AOI22xp33_ASAP7_75t_L g1343 ( 
.A1(n_1197),
.A2(n_1104),
.B1(n_1205),
.B2(n_1187),
.Y(n_1343)
);

INVx4_ASAP7_75t_L g1344 ( 
.A(n_1201),
.Y(n_1344)
);

CKINVDCx14_ASAP7_75t_R g1345 ( 
.A(n_1102),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1177),
.Y(n_1346)
);

NAND2xp5_ASAP7_75t_L g1347 ( 
.A(n_1136),
.B(n_1184),
.Y(n_1347)
);

HB1xp67_ASAP7_75t_L g1348 ( 
.A(n_1111),
.Y(n_1348)
);

BUFx2_ASAP7_75t_L g1349 ( 
.A(n_1225),
.Y(n_1349)
);

AOI22xp33_ASAP7_75t_L g1350 ( 
.A1(n_1197),
.A2(n_1104),
.B1(n_1205),
.B2(n_1187),
.Y(n_1350)
);

AOI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1253),
.A2(n_1299),
.B(n_1310),
.Y(n_1351)
);

HB1xp67_ASAP7_75t_L g1352 ( 
.A(n_1316),
.Y(n_1352)
);

AND2x2_ASAP7_75t_L g1353 ( 
.A(n_1320),
.B(n_1291),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_1326),
.Y(n_1354)
);

INVx1_ASAP7_75t_SL g1355 ( 
.A(n_1288),
.Y(n_1355)
);

AND2x2_ASAP7_75t_L g1356 ( 
.A(n_1334),
.B(n_1348),
.Y(n_1356)
);

BUFx6f_ASAP7_75t_L g1357 ( 
.A(n_1325),
.Y(n_1357)
);

AND2x4_ASAP7_75t_L g1358 ( 
.A(n_1322),
.B(n_1317),
.Y(n_1358)
);

AOI22xp33_ASAP7_75t_L g1359 ( 
.A1(n_1330),
.A2(n_1340),
.B1(n_1277),
.B2(n_1329),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_1271),
.Y(n_1360)
);

AOI21xp33_ASAP7_75t_L g1361 ( 
.A1(n_1276),
.A2(n_1329),
.B(n_1262),
.Y(n_1361)
);

AND2x2_ASAP7_75t_L g1362 ( 
.A(n_1334),
.B(n_1348),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1282),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1285),
.Y(n_1364)
);

BUFx2_ASAP7_75t_SL g1365 ( 
.A(n_1317),
.Y(n_1365)
);

NOR2xp33_ASAP7_75t_L g1366 ( 
.A(n_1347),
.B(n_1279),
.Y(n_1366)
);

BUFx2_ASAP7_75t_L g1367 ( 
.A(n_1321),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_1245),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1246),
.Y(n_1369)
);

BUFx2_ASAP7_75t_L g1370 ( 
.A(n_1327),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1248),
.Y(n_1371)
);

INVx1_ASAP7_75t_L g1372 ( 
.A(n_1254),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_1256),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1257),
.Y(n_1374)
);

OA21x2_ASAP7_75t_L g1375 ( 
.A1(n_1283),
.A2(n_1262),
.B(n_1303),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1259),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1261),
.Y(n_1377)
);

OAI21x1_ASAP7_75t_L g1378 ( 
.A1(n_1315),
.A2(n_1298),
.B(n_1264),
.Y(n_1378)
);

OAI21x1_ASAP7_75t_L g1379 ( 
.A1(n_1298),
.A2(n_1283),
.B(n_1312),
.Y(n_1379)
);

HB1xp67_ASAP7_75t_L g1380 ( 
.A(n_1243),
.Y(n_1380)
);

OR2x6_ASAP7_75t_L g1381 ( 
.A(n_1313),
.B(n_1324),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1303),
.A2(n_1312),
.B(n_1306),
.Y(n_1382)
);

INVx1_ASAP7_75t_L g1383 ( 
.A(n_1266),
.Y(n_1383)
);

INVx1_ASAP7_75t_L g1384 ( 
.A(n_1328),
.Y(n_1384)
);

HB1xp67_ASAP7_75t_L g1385 ( 
.A(n_1349),
.Y(n_1385)
);

OAI21x1_ASAP7_75t_L g1386 ( 
.A1(n_1306),
.A2(n_1293),
.B(n_1332),
.Y(n_1386)
);

HB1xp67_ASAP7_75t_L g1387 ( 
.A(n_1319),
.Y(n_1387)
);

INVx3_ASAP7_75t_L g1388 ( 
.A(n_1313),
.Y(n_1388)
);

INVx2_ASAP7_75t_L g1389 ( 
.A(n_1244),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1277),
.B(n_1333),
.Y(n_1390)
);

CKINVDCx20_ASAP7_75t_R g1391 ( 
.A(n_1240),
.Y(n_1391)
);

AOI21x1_ASAP7_75t_L g1392 ( 
.A1(n_1339),
.A2(n_1341),
.B(n_1338),
.Y(n_1392)
);

AND2x4_ASAP7_75t_L g1393 ( 
.A(n_1300),
.B(n_1293),
.Y(n_1393)
);

NAND2xp5_ASAP7_75t_L g1394 ( 
.A(n_1278),
.B(n_1258),
.Y(n_1394)
);

HB1xp67_ASAP7_75t_SL g1395 ( 
.A(n_1260),
.Y(n_1395)
);

HB1xp67_ASAP7_75t_L g1396 ( 
.A(n_1287),
.Y(n_1396)
);

BUFx2_ASAP7_75t_L g1397 ( 
.A(n_1251),
.Y(n_1397)
);

AND2x2_ASAP7_75t_L g1398 ( 
.A(n_1258),
.B(n_1290),
.Y(n_1398)
);

INVx1_ASAP7_75t_L g1399 ( 
.A(n_1323),
.Y(n_1399)
);

INVx1_ASAP7_75t_L g1400 ( 
.A(n_1323),
.Y(n_1400)
);

OAI21x1_ASAP7_75t_SL g1401 ( 
.A1(n_1276),
.A2(n_1289),
.B(n_1275),
.Y(n_1401)
);

HB1xp67_ASAP7_75t_L g1402 ( 
.A(n_1296),
.Y(n_1402)
);

HB1xp67_ASAP7_75t_L g1403 ( 
.A(n_1251),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1278),
.Y(n_1404)
);

INVx2_ASAP7_75t_SL g1405 ( 
.A(n_1270),
.Y(n_1405)
);

HB1xp67_ASAP7_75t_L g1406 ( 
.A(n_1275),
.Y(n_1406)
);

AOI22xp33_ASAP7_75t_L g1407 ( 
.A1(n_1330),
.A2(n_1340),
.B1(n_1265),
.B2(n_1335),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1307),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1265),
.A2(n_1336),
.B(n_1290),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1307),
.Y(n_1410)
);

INVx1_ASAP7_75t_L g1411 ( 
.A(n_1281),
.Y(n_1411)
);

AO21x2_ASAP7_75t_L g1412 ( 
.A1(n_1309),
.A2(n_1318),
.B(n_1242),
.Y(n_1412)
);

OAI22xp5_ASAP7_75t_L g1413 ( 
.A1(n_1242),
.A2(n_1350),
.B1(n_1343),
.B2(n_1342),
.Y(n_1413)
);

OAI21xp5_ASAP7_75t_L g1414 ( 
.A1(n_1335),
.A2(n_1350),
.B(n_1342),
.Y(n_1414)
);

AO21x2_ASAP7_75t_L g1415 ( 
.A1(n_1343),
.A2(n_1286),
.B(n_1292),
.Y(n_1415)
);

HB1xp67_ASAP7_75t_L g1416 ( 
.A(n_1314),
.Y(n_1416)
);

INVxp33_ASAP7_75t_L g1417 ( 
.A(n_1247),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1286),
.B(n_1345),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1260),
.Y(n_1419)
);

OA21x2_ASAP7_75t_L g1420 ( 
.A1(n_1378),
.A2(n_1297),
.B(n_1272),
.Y(n_1420)
);

AND2x2_ASAP7_75t_L g1421 ( 
.A(n_1368),
.B(n_1345),
.Y(n_1421)
);

AND2x2_ASAP7_75t_L g1422 ( 
.A(n_1368),
.B(n_1273),
.Y(n_1422)
);

BUFx3_ASAP7_75t_L g1423 ( 
.A(n_1397),
.Y(n_1423)
);

OAI21xp5_ASAP7_75t_L g1424 ( 
.A1(n_1409),
.A2(n_1280),
.B(n_1274),
.Y(n_1424)
);

OAI21xp5_ASAP7_75t_L g1425 ( 
.A1(n_1409),
.A2(n_1294),
.B(n_1252),
.Y(n_1425)
);

OAI21xp5_ASAP7_75t_L g1426 ( 
.A1(n_1392),
.A2(n_1344),
.B(n_1308),
.Y(n_1426)
);

BUFx2_ASAP7_75t_L g1427 ( 
.A(n_1397),
.Y(n_1427)
);

OR2x2_ASAP7_75t_L g1428 ( 
.A(n_1396),
.B(n_1249),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_1363),
.Y(n_1429)
);

AND2x2_ASAP7_75t_L g1430 ( 
.A(n_1369),
.B(n_1284),
.Y(n_1430)
);

AND2x4_ASAP7_75t_L g1431 ( 
.A(n_1381),
.B(n_1302),
.Y(n_1431)
);

NAND2xp5_ASAP7_75t_L g1432 ( 
.A(n_1396),
.B(n_1284),
.Y(n_1432)
);

O2A1O1Ixp5_ASAP7_75t_L g1433 ( 
.A1(n_1392),
.A2(n_1269),
.B(n_1247),
.C(n_1267),
.Y(n_1433)
);

NOR2xp33_ASAP7_75t_L g1434 ( 
.A(n_1391),
.B(n_1346),
.Y(n_1434)
);

HB1xp67_ASAP7_75t_L g1435 ( 
.A(n_1380),
.Y(n_1435)
);

NOR2xp33_ASAP7_75t_L g1436 ( 
.A(n_1366),
.B(n_1250),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1357),
.Y(n_1437)
);

A2O1A1Ixp33_ASAP7_75t_L g1438 ( 
.A1(n_1361),
.A2(n_1305),
.B(n_1263),
.C(n_1331),
.Y(n_1438)
);

INVx1_ASAP7_75t_L g1439 ( 
.A(n_1363),
.Y(n_1439)
);

CKINVDCx20_ASAP7_75t_R g1440 ( 
.A(n_1419),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1389),
.Y(n_1441)
);

AND2x2_ASAP7_75t_L g1442 ( 
.A(n_1369),
.B(n_1371),
.Y(n_1442)
);

NOR2x1_ASAP7_75t_SL g1443 ( 
.A(n_1365),
.B(n_1255),
.Y(n_1443)
);

INVx1_ASAP7_75t_L g1444 ( 
.A(n_1364),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1364),
.Y(n_1445)
);

AND2x4_ASAP7_75t_L g1446 ( 
.A(n_1381),
.B(n_1331),
.Y(n_1446)
);

OR2x2_ASAP7_75t_L g1447 ( 
.A(n_1380),
.B(n_1267),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1385),
.B(n_1301),
.Y(n_1448)
);

AND2x4_ASAP7_75t_L g1449 ( 
.A(n_1381),
.B(n_1301),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1371),
.Y(n_1450)
);

NOR2xp33_ASAP7_75t_L g1451 ( 
.A(n_1419),
.B(n_1241),
.Y(n_1451)
);

AND2x2_ASAP7_75t_L g1452 ( 
.A(n_1372),
.B(n_1268),
.Y(n_1452)
);

O2A1O1Ixp33_ASAP7_75t_SL g1453 ( 
.A1(n_1387),
.A2(n_1295),
.B(n_1304),
.C(n_1311),
.Y(n_1453)
);

NOR2x1_ASAP7_75t_SL g1454 ( 
.A(n_1365),
.B(n_1304),
.Y(n_1454)
);

AND2x2_ASAP7_75t_L g1455 ( 
.A(n_1372),
.B(n_1268),
.Y(n_1455)
);

AND2x2_ASAP7_75t_SL g1456 ( 
.A(n_1387),
.B(n_1304),
.Y(n_1456)
);

OAI22xp33_ASAP7_75t_L g1457 ( 
.A1(n_1413),
.A2(n_1241),
.B1(n_1337),
.B2(n_1311),
.Y(n_1457)
);

BUFx6f_ASAP7_75t_L g1458 ( 
.A(n_1357),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1395),
.Y(n_1459)
);

AND2x2_ASAP7_75t_L g1460 ( 
.A(n_1373),
.B(n_1337),
.Y(n_1460)
);

INVx1_ASAP7_75t_SL g1461 ( 
.A(n_1355),
.Y(n_1461)
);

AND2x2_ASAP7_75t_L g1462 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1462)
);

AND2x2_ASAP7_75t_L g1463 ( 
.A(n_1374),
.B(n_1376),
.Y(n_1463)
);

OAI21xp5_ASAP7_75t_L g1464 ( 
.A1(n_1361),
.A2(n_1386),
.B(n_1407),
.Y(n_1464)
);

AND2x4_ASAP7_75t_L g1465 ( 
.A(n_1381),
.B(n_1393),
.Y(n_1465)
);

AO32x2_ASAP7_75t_L g1466 ( 
.A1(n_1413),
.A2(n_1354),
.A3(n_1405),
.B1(n_1385),
.B2(n_1411),
.Y(n_1466)
);

OR2x2_ASAP7_75t_L g1467 ( 
.A(n_1403),
.B(n_1377),
.Y(n_1467)
);

BUFx2_ASAP7_75t_L g1468 ( 
.A(n_1403),
.Y(n_1468)
);

AND2x2_ASAP7_75t_L g1469 ( 
.A(n_1377),
.B(n_1383),
.Y(n_1469)
);

INVx1_ASAP7_75t_L g1470 ( 
.A(n_1383),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1384),
.Y(n_1471)
);

OA21x2_ASAP7_75t_L g1472 ( 
.A1(n_1378),
.A2(n_1379),
.B(n_1386),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1417),
.B(n_1395),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1355),
.B(n_1404),
.Y(n_1474)
);

AND2x4_ASAP7_75t_L g1475 ( 
.A(n_1393),
.B(n_1388),
.Y(n_1475)
);

AOI22xp33_ASAP7_75t_L g1476 ( 
.A1(n_1359),
.A2(n_1406),
.B1(n_1398),
.B2(n_1414),
.Y(n_1476)
);

NAND2xp5_ASAP7_75t_L g1477 ( 
.A(n_1404),
.B(n_1360),
.Y(n_1477)
);

AO32x2_ASAP7_75t_L g1478 ( 
.A1(n_1354),
.A2(n_1405),
.A3(n_1411),
.B1(n_1352),
.B2(n_1394),
.Y(n_1478)
);

OAI22xp5_ASAP7_75t_L g1479 ( 
.A1(n_1406),
.A2(n_1394),
.B1(n_1414),
.B2(n_1375),
.Y(n_1479)
);

AO21x2_ASAP7_75t_L g1480 ( 
.A1(n_1401),
.A2(n_1408),
.B(n_1410),
.Y(n_1480)
);

A2O1A1Ixp33_ASAP7_75t_L g1481 ( 
.A1(n_1398),
.A2(n_1386),
.B(n_1378),
.C(n_1379),
.Y(n_1481)
);

OR2x2_ASAP7_75t_L g1482 ( 
.A(n_1352),
.B(n_1356),
.Y(n_1482)
);

INVxp67_ASAP7_75t_SL g1483 ( 
.A(n_1358),
.Y(n_1483)
);

NAND3xp33_ASAP7_75t_L g1484 ( 
.A(n_1375),
.B(n_1399),
.C(n_1400),
.Y(n_1484)
);

OAI21xp5_ASAP7_75t_L g1485 ( 
.A1(n_1379),
.A2(n_1375),
.B(n_1398),
.Y(n_1485)
);

HB1xp67_ASAP7_75t_L g1486 ( 
.A(n_1402),
.Y(n_1486)
);

INVxp67_ASAP7_75t_L g1487 ( 
.A(n_1435),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_1450),
.Y(n_1488)
);

AND2x2_ASAP7_75t_L g1489 ( 
.A(n_1483),
.B(n_1421),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1470),
.Y(n_1490)
);

AND2x2_ASAP7_75t_L g1491 ( 
.A(n_1421),
.B(n_1353),
.Y(n_1491)
);

INVx2_ASAP7_75t_L g1492 ( 
.A(n_1441),
.Y(n_1492)
);

NAND2xp5_ASAP7_75t_L g1493 ( 
.A(n_1461),
.B(n_1358),
.Y(n_1493)
);

OR2x2_ASAP7_75t_L g1494 ( 
.A(n_1482),
.B(n_1399),
.Y(n_1494)
);

AND2x4_ASAP7_75t_L g1495 ( 
.A(n_1465),
.B(n_1353),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1429),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_1471),
.Y(n_1497)
);

INVxp67_ASAP7_75t_SL g1498 ( 
.A(n_1482),
.Y(n_1498)
);

AOI22xp5_ASAP7_75t_L g1499 ( 
.A1(n_1479),
.A2(n_1415),
.B1(n_1412),
.B2(n_1375),
.Y(n_1499)
);

CKINVDCx14_ASAP7_75t_R g1500 ( 
.A(n_1440),
.Y(n_1500)
);

AND2x2_ASAP7_75t_L g1501 ( 
.A(n_1427),
.B(n_1358),
.Y(n_1501)
);

OR2x2_ASAP7_75t_L g1502 ( 
.A(n_1486),
.B(n_1467),
.Y(n_1502)
);

NOR2xp67_ASAP7_75t_L g1503 ( 
.A(n_1473),
.B(n_1416),
.Y(n_1503)
);

NAND2xp5_ASAP7_75t_L g1504 ( 
.A(n_1474),
.B(n_1358),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1423),
.B(n_1370),
.Y(n_1505)
);

INVx1_ASAP7_75t_L g1506 ( 
.A(n_1439),
.Y(n_1506)
);

AND2x2_ASAP7_75t_L g1507 ( 
.A(n_1423),
.B(n_1370),
.Y(n_1507)
);

AND2x4_ASAP7_75t_L g1508 ( 
.A(n_1465),
.B(n_1475),
.Y(n_1508)
);

INVx11_ASAP7_75t_L g1509 ( 
.A(n_1459),
.Y(n_1509)
);

AOI22xp33_ASAP7_75t_SL g1510 ( 
.A1(n_1464),
.A2(n_1401),
.B1(n_1415),
.B2(n_1412),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_1444),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1445),
.Y(n_1512)
);

AO22x1_ASAP7_75t_L g1513 ( 
.A1(n_1485),
.A2(n_1393),
.B1(n_1418),
.B2(n_1390),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1442),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1462),
.B(n_1463),
.Y(n_1515)
);

AND2x2_ASAP7_75t_L g1516 ( 
.A(n_1468),
.B(n_1400),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1462),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1463),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1469),
.B(n_1354),
.Y(n_1519)
);

NOR2x1_ASAP7_75t_L g1520 ( 
.A(n_1440),
.B(n_1428),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1475),
.B(n_1418),
.Y(n_1521)
);

AOI22xp33_ASAP7_75t_L g1522 ( 
.A1(n_1476),
.A2(n_1412),
.B1(n_1415),
.B2(n_1390),
.Y(n_1522)
);

OR2x2_ASAP7_75t_L g1523 ( 
.A(n_1477),
.B(n_1356),
.Y(n_1523)
);

HB1xp67_ASAP7_75t_L g1524 ( 
.A(n_1430),
.Y(n_1524)
);

AND2x4_ASAP7_75t_L g1525 ( 
.A(n_1475),
.B(n_1356),
.Y(n_1525)
);

OR2x2_ASAP7_75t_L g1526 ( 
.A(n_1484),
.B(n_1362),
.Y(n_1526)
);

INVx1_ASAP7_75t_L g1527 ( 
.A(n_1506),
.Y(n_1527)
);

HB1xp67_ASAP7_75t_L g1528 ( 
.A(n_1487),
.Y(n_1528)
);

INVx2_ASAP7_75t_L g1529 ( 
.A(n_1492),
.Y(n_1529)
);

HB1xp67_ASAP7_75t_L g1530 ( 
.A(n_1502),
.Y(n_1530)
);

INVx1_ASAP7_75t_L g1531 ( 
.A(n_1506),
.Y(n_1531)
);

INVx2_ASAP7_75t_SL g1532 ( 
.A(n_1525),
.Y(n_1532)
);

OR2x2_ASAP7_75t_L g1533 ( 
.A(n_1494),
.B(n_1472),
.Y(n_1533)
);

OAI33xp33_ASAP7_75t_L g1534 ( 
.A1(n_1526),
.A2(n_1432),
.A3(n_1428),
.B1(n_1457),
.B2(n_1447),
.B3(n_1360),
.Y(n_1534)
);

INVx2_ASAP7_75t_L g1535 ( 
.A(n_1492),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1525),
.B(n_1478),
.Y(n_1536)
);

INVx1_ASAP7_75t_L g1537 ( 
.A(n_1511),
.Y(n_1537)
);

NAND2xp5_ASAP7_75t_SL g1538 ( 
.A(n_1503),
.B(n_1456),
.Y(n_1538)
);

OR2x2_ASAP7_75t_L g1539 ( 
.A(n_1494),
.B(n_1472),
.Y(n_1539)
);

HB1xp67_ASAP7_75t_L g1540 ( 
.A(n_1502),
.Y(n_1540)
);

INVx1_ASAP7_75t_L g1541 ( 
.A(n_1511),
.Y(n_1541)
);

OR2x2_ASAP7_75t_L g1542 ( 
.A(n_1526),
.B(n_1472),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1525),
.B(n_1478),
.Y(n_1543)
);

BUFx2_ASAP7_75t_L g1544 ( 
.A(n_1500),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1512),
.Y(n_1545)
);

AOI211xp5_ASAP7_75t_L g1546 ( 
.A1(n_1513),
.A2(n_1424),
.B(n_1425),
.C(n_1481),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1491),
.B(n_1478),
.Y(n_1547)
);

BUFx3_ASAP7_75t_L g1548 ( 
.A(n_1505),
.Y(n_1548)
);

NAND2x1_ASAP7_75t_L g1549 ( 
.A(n_1508),
.B(n_1449),
.Y(n_1549)
);

BUFx3_ASAP7_75t_L g1550 ( 
.A(n_1505),
.Y(n_1550)
);

INVx1_ASAP7_75t_L g1551 ( 
.A(n_1512),
.Y(n_1551)
);

OR2x2_ASAP7_75t_L g1552 ( 
.A(n_1498),
.B(n_1481),
.Y(n_1552)
);

BUFx3_ASAP7_75t_L g1553 ( 
.A(n_1507),
.Y(n_1553)
);

HB1xp67_ASAP7_75t_L g1554 ( 
.A(n_1516),
.Y(n_1554)
);

HB1xp67_ASAP7_75t_L g1555 ( 
.A(n_1516),
.Y(n_1555)
);

AND2x4_ASAP7_75t_SL g1556 ( 
.A(n_1508),
.B(n_1449),
.Y(n_1556)
);

INVx1_ASAP7_75t_L g1557 ( 
.A(n_1488),
.Y(n_1557)
);

AOI21xp33_ASAP7_75t_L g1558 ( 
.A1(n_1510),
.A2(n_1415),
.B(n_1480),
.Y(n_1558)
);

HB1xp67_ASAP7_75t_L g1559 ( 
.A(n_1496),
.Y(n_1559)
);

OAI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1522),
.A2(n_1375),
.B1(n_1456),
.B2(n_1438),
.Y(n_1560)
);

INVx1_ASAP7_75t_L g1561 ( 
.A(n_1488),
.Y(n_1561)
);

AOI33xp33_ASAP7_75t_L g1562 ( 
.A1(n_1499),
.A2(n_1452),
.A3(n_1455),
.B1(n_1422),
.B2(n_1460),
.B3(n_1430),
.Y(n_1562)
);

OAI221xp5_ASAP7_75t_L g1563 ( 
.A1(n_1520),
.A2(n_1433),
.B1(n_1438),
.B2(n_1390),
.C(n_1426),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1491),
.B(n_1478),
.Y(n_1564)
);

INVx3_ASAP7_75t_L g1565 ( 
.A(n_1508),
.Y(n_1565)
);

NAND2xp5_ASAP7_75t_L g1566 ( 
.A(n_1523),
.B(n_1480),
.Y(n_1566)
);

AOI22xp33_ASAP7_75t_L g1567 ( 
.A1(n_1504),
.A2(n_1412),
.B1(n_1480),
.B2(n_1382),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1519),
.B(n_1466),
.Y(n_1568)
);

INVx2_ASAP7_75t_L g1569 ( 
.A(n_1529),
.Y(n_1569)
);

INVx2_ASAP7_75t_L g1570 ( 
.A(n_1529),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1530),
.B(n_1523),
.Y(n_1571)
);

INVx2_ASAP7_75t_L g1572 ( 
.A(n_1529),
.Y(n_1572)
);

INVx1_ASAP7_75t_L g1573 ( 
.A(n_1557),
.Y(n_1573)
);

NOR2x1_ASAP7_75t_L g1574 ( 
.A(n_1544),
.B(n_1447),
.Y(n_1574)
);

OR2x2_ASAP7_75t_L g1575 ( 
.A(n_1530),
.B(n_1515),
.Y(n_1575)
);

INVx2_ASAP7_75t_SL g1576 ( 
.A(n_1549),
.Y(n_1576)
);

OR2x2_ASAP7_75t_L g1577 ( 
.A(n_1540),
.B(n_1514),
.Y(n_1577)
);

NOR2x1p5_ASAP7_75t_L g1578 ( 
.A(n_1549),
.B(n_1459),
.Y(n_1578)
);

INVx2_ASAP7_75t_L g1579 ( 
.A(n_1535),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1557),
.Y(n_1581)
);

INVx1_ASAP7_75t_L g1582 ( 
.A(n_1561),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1561),
.Y(n_1583)
);

BUFx6f_ASAP7_75t_L g1584 ( 
.A(n_1544),
.Y(n_1584)
);

HB1xp67_ASAP7_75t_L g1585 ( 
.A(n_1540),
.Y(n_1585)
);

AND2x4_ASAP7_75t_L g1586 ( 
.A(n_1565),
.B(n_1495),
.Y(n_1586)
);

AND2x2_ASAP7_75t_L g1587 ( 
.A(n_1536),
.B(n_1489),
.Y(n_1587)
);

OR2x2_ASAP7_75t_L g1588 ( 
.A(n_1552),
.B(n_1514),
.Y(n_1588)
);

HB1xp67_ASAP7_75t_L g1589 ( 
.A(n_1559),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1559),
.B(n_1490),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1527),
.B(n_1490),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_SL g1592 ( 
.A(n_1546),
.B(n_1495),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1527),
.B(n_1497),
.Y(n_1593)
);

AND2x2_ASAP7_75t_L g1594 ( 
.A(n_1536),
.B(n_1524),
.Y(n_1594)
);

AND2x2_ASAP7_75t_SL g1595 ( 
.A(n_1552),
.B(n_1420),
.Y(n_1595)
);

AND2x2_ASAP7_75t_L g1596 ( 
.A(n_1543),
.B(n_1507),
.Y(n_1596)
);

OAI31xp33_ASAP7_75t_L g1597 ( 
.A1(n_1563),
.A2(n_1367),
.A3(n_1422),
.B(n_1455),
.Y(n_1597)
);

INVx2_ASAP7_75t_SL g1598 ( 
.A(n_1556),
.Y(n_1598)
);

OR2x2_ASAP7_75t_L g1599 ( 
.A(n_1552),
.B(n_1517),
.Y(n_1599)
);

OR2x2_ASAP7_75t_L g1600 ( 
.A(n_1566),
.B(n_1517),
.Y(n_1600)
);

AND2x2_ASAP7_75t_L g1601 ( 
.A(n_1543),
.B(n_1518),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1543),
.B(n_1518),
.Y(n_1602)
);

INVx2_ASAP7_75t_L g1603 ( 
.A(n_1535),
.Y(n_1603)
);

OR2x2_ASAP7_75t_L g1604 ( 
.A(n_1566),
.B(n_1554),
.Y(n_1604)
);

OAI221xp5_ASAP7_75t_L g1605 ( 
.A1(n_1546),
.A2(n_1420),
.B1(n_1382),
.B2(n_1351),
.C(n_1436),
.Y(n_1605)
);

AND2x2_ASAP7_75t_L g1606 ( 
.A(n_1547),
.B(n_1501),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1531),
.B(n_1497),
.Y(n_1607)
);

INVx1_ASAP7_75t_L g1608 ( 
.A(n_1573),
.Y(n_1608)
);

INVx1_ASAP7_75t_L g1609 ( 
.A(n_1573),
.Y(n_1609)
);

INVx2_ASAP7_75t_SL g1610 ( 
.A(n_1584),
.Y(n_1610)
);

INVx2_ASAP7_75t_L g1611 ( 
.A(n_1569),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1581),
.Y(n_1612)
);

NAND2xp5_ASAP7_75t_L g1613 ( 
.A(n_1585),
.B(n_1528),
.Y(n_1613)
);

NAND2xp5_ASAP7_75t_L g1614 ( 
.A(n_1585),
.B(n_1528),
.Y(n_1614)
);

NAND2x1_ASAP7_75t_L g1615 ( 
.A(n_1576),
.B(n_1565),
.Y(n_1615)
);

INVx2_ASAP7_75t_L g1616 ( 
.A(n_1569),
.Y(n_1616)
);

AND2x2_ASAP7_75t_L g1617 ( 
.A(n_1598),
.B(n_1565),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1581),
.Y(n_1618)
);

INVx2_ASAP7_75t_L g1619 ( 
.A(n_1569),
.Y(n_1619)
);

INVx1_ASAP7_75t_L g1620 ( 
.A(n_1582),
.Y(n_1620)
);

NAND2xp5_ASAP7_75t_L g1621 ( 
.A(n_1589),
.B(n_1562),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1589),
.B(n_1554),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1570),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1574),
.B(n_1555),
.Y(n_1624)
);

INVx2_ASAP7_75t_L g1625 ( 
.A(n_1570),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1574),
.B(n_1555),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1570),
.Y(n_1627)
);

AND2x2_ASAP7_75t_L g1628 ( 
.A(n_1598),
.B(n_1565),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1572),
.Y(n_1629)
);

OR2x2_ASAP7_75t_L g1630 ( 
.A(n_1571),
.B(n_1542),
.Y(n_1630)
);

OR2x2_ASAP7_75t_L g1631 ( 
.A(n_1571),
.B(n_1542),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1632)
);

AOI22xp5_ASAP7_75t_L g1633 ( 
.A1(n_1605),
.A2(n_1560),
.B1(n_1563),
.B2(n_1558),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1582),
.Y(n_1634)
);

INVx2_ASAP7_75t_SL g1635 ( 
.A(n_1584),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1583),
.Y(n_1636)
);

INVx3_ASAP7_75t_L g1637 ( 
.A(n_1586),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1597),
.B(n_1568),
.Y(n_1638)
);

INVx1_ASAP7_75t_L g1639 ( 
.A(n_1583),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1591),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1584),
.B(n_1509),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1572),
.Y(n_1642)
);

OR2x2_ASAP7_75t_L g1643 ( 
.A(n_1575),
.B(n_1542),
.Y(n_1643)
);

NAND4xp25_ASAP7_75t_L g1644 ( 
.A(n_1605),
.B(n_1460),
.C(n_1590),
.D(n_1592),
.Y(n_1644)
);

BUFx2_ASAP7_75t_L g1645 ( 
.A(n_1584),
.Y(n_1645)
);

AND2x2_ASAP7_75t_L g1646 ( 
.A(n_1598),
.B(n_1580),
.Y(n_1646)
);

AND2x4_ASAP7_75t_L g1647 ( 
.A(n_1578),
.B(n_1532),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1591),
.Y(n_1648)
);

NOR2xp33_ASAP7_75t_SL g1649 ( 
.A(n_1584),
.B(n_1451),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1572),
.Y(n_1650)
);

INVx1_ASAP7_75t_SL g1651 ( 
.A(n_1649),
.Y(n_1651)
);

AND2x2_ASAP7_75t_L g1652 ( 
.A(n_1646),
.B(n_1584),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1608),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1608),
.Y(n_1654)
);

OAI221xp5_ASAP7_75t_L g1655 ( 
.A1(n_1633),
.A2(n_1558),
.B1(n_1560),
.B2(n_1567),
.C(n_1539),
.Y(n_1655)
);

AND2x2_ASAP7_75t_L g1656 ( 
.A(n_1646),
.B(n_1578),
.Y(n_1656)
);

NAND2x1_ASAP7_75t_L g1657 ( 
.A(n_1637),
.B(n_1576),
.Y(n_1657)
);

AND2x2_ASAP7_75t_L g1658 ( 
.A(n_1641),
.B(n_1580),
.Y(n_1658)
);

AND2x2_ASAP7_75t_L g1659 ( 
.A(n_1617),
.B(n_1580),
.Y(n_1659)
);

OR2x2_ASAP7_75t_L g1660 ( 
.A(n_1621),
.B(n_1588),
.Y(n_1660)
);

NOR2xp33_ASAP7_75t_L g1661 ( 
.A(n_1644),
.B(n_1509),
.Y(n_1661)
);

NAND2x1p5_ASAP7_75t_L g1662 ( 
.A(n_1615),
.B(n_1538),
.Y(n_1662)
);

OR2x2_ASAP7_75t_L g1663 ( 
.A(n_1613),
.B(n_1588),
.Y(n_1663)
);

NOR2xp33_ASAP7_75t_L g1664 ( 
.A(n_1614),
.B(n_1534),
.Y(n_1664)
);

OR2x6_ASAP7_75t_L g1665 ( 
.A(n_1610),
.B(n_1357),
.Y(n_1665)
);

OR2x2_ASAP7_75t_L g1666 ( 
.A(n_1622),
.B(n_1599),
.Y(n_1666)
);

OR2x2_ASAP7_75t_L g1667 ( 
.A(n_1643),
.B(n_1599),
.Y(n_1667)
);

INVx1_ASAP7_75t_L g1668 ( 
.A(n_1609),
.Y(n_1668)
);

NOR2xp33_ASAP7_75t_L g1669 ( 
.A(n_1610),
.B(n_1534),
.Y(n_1669)
);

NOR2xp67_ASAP7_75t_SL g1670 ( 
.A(n_1645),
.B(n_1576),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1633),
.B(n_1568),
.Y(n_1671)
);

NOR2x1_ASAP7_75t_L g1672 ( 
.A(n_1645),
.B(n_1434),
.Y(n_1672)
);

OR2x2_ASAP7_75t_L g1673 ( 
.A(n_1643),
.B(n_1575),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1609),
.Y(n_1674)
);

OR2x2_ASAP7_75t_L g1675 ( 
.A(n_1632),
.B(n_1577),
.Y(n_1675)
);

NAND2x1p5_ASAP7_75t_L g1676 ( 
.A(n_1615),
.B(n_1595),
.Y(n_1676)
);

INVxp67_ASAP7_75t_L g1677 ( 
.A(n_1635),
.Y(n_1677)
);

INVx2_ASAP7_75t_SL g1678 ( 
.A(n_1637),
.Y(n_1678)
);

INVx1_ASAP7_75t_SL g1679 ( 
.A(n_1635),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1640),
.B(n_1547),
.Y(n_1680)
);

BUFx2_ASAP7_75t_L g1681 ( 
.A(n_1647),
.Y(n_1681)
);

AND2x4_ASAP7_75t_L g1682 ( 
.A(n_1647),
.B(n_1586),
.Y(n_1682)
);

AOI322xp5_ASAP7_75t_L g1683 ( 
.A1(n_1638),
.A2(n_1547),
.A3(n_1564),
.B1(n_1595),
.B2(n_1587),
.C1(n_1567),
.C2(n_1601),
.Y(n_1683)
);

NAND2xp5_ASAP7_75t_L g1684 ( 
.A(n_1640),
.B(n_1564),
.Y(n_1684)
);

OAI21xp33_ASAP7_75t_L g1685 ( 
.A1(n_1624),
.A2(n_1604),
.B(n_1595),
.Y(n_1685)
);

INVx1_ASAP7_75t_SL g1686 ( 
.A(n_1617),
.Y(n_1686)
);

OAI22xp5_ASAP7_75t_L g1687 ( 
.A1(n_1671),
.A2(n_1637),
.B1(n_1647),
.B2(n_1626),
.Y(n_1687)
);

INVxp67_ASAP7_75t_L g1688 ( 
.A(n_1681),
.Y(n_1688)
);

NAND3xp33_ASAP7_75t_L g1689 ( 
.A(n_1683),
.B(n_1648),
.C(n_1618),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1653),
.Y(n_1690)
);

OAI32xp33_ASAP7_75t_L g1691 ( 
.A1(n_1664),
.A2(n_1637),
.A3(n_1630),
.B1(n_1631),
.B2(n_1604),
.Y(n_1691)
);

OR2x2_ASAP7_75t_L g1692 ( 
.A(n_1675),
.B(n_1630),
.Y(n_1692)
);

AOI21xp33_ASAP7_75t_L g1693 ( 
.A1(n_1655),
.A2(n_1623),
.B(n_1619),
.Y(n_1693)
);

OAI321xp33_ASAP7_75t_L g1694 ( 
.A1(n_1685),
.A2(n_1631),
.A3(n_1648),
.B1(n_1628),
.B2(n_1623),
.C(n_1625),
.Y(n_1694)
);

OAI22xp33_ASAP7_75t_L g1695 ( 
.A1(n_1651),
.A2(n_1533),
.B1(n_1539),
.B2(n_1564),
.Y(n_1695)
);

NAND2xp5_ASAP7_75t_L g1696 ( 
.A(n_1686),
.B(n_1587),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1654),
.Y(n_1697)
);

NOR2xp33_ASAP7_75t_L g1698 ( 
.A(n_1686),
.B(n_1647),
.Y(n_1698)
);

NOR2x1p5_ASAP7_75t_L g1699 ( 
.A(n_1657),
.B(n_1628),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1669),
.B(n_1587),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1683),
.B(n_1606),
.Y(n_1701)
);

AOI21xp33_ASAP7_75t_L g1702 ( 
.A1(n_1685),
.A2(n_1623),
.B(n_1619),
.Y(n_1702)
);

INVxp67_ASAP7_75t_SL g1703 ( 
.A(n_1672),
.Y(n_1703)
);

OAI31xp33_ASAP7_75t_L g1704 ( 
.A1(n_1676),
.A2(n_1539),
.A3(n_1533),
.B(n_1625),
.Y(n_1704)
);

NOR2xp33_ASAP7_75t_L g1705 ( 
.A(n_1652),
.B(n_1590),
.Y(n_1705)
);

OAI32xp33_ASAP7_75t_L g1706 ( 
.A1(n_1676),
.A2(n_1612),
.A3(n_1618),
.B1(n_1634),
.B2(n_1639),
.Y(n_1706)
);

NAND2xp5_ASAP7_75t_L g1707 ( 
.A(n_1663),
.B(n_1679),
.Y(n_1707)
);

OAI21xp33_ASAP7_75t_SL g1708 ( 
.A1(n_1659),
.A2(n_1596),
.B(n_1606),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1658),
.B(n_1596),
.Y(n_1709)
);

INVx2_ASAP7_75t_L g1710 ( 
.A(n_1678),
.Y(n_1710)
);

INVx1_ASAP7_75t_L g1711 ( 
.A(n_1668),
.Y(n_1711)
);

NOR2xp67_ASAP7_75t_L g1712 ( 
.A(n_1682),
.B(n_1586),
.Y(n_1712)
);

OAI22xp5_ASAP7_75t_L g1713 ( 
.A1(n_1703),
.A2(n_1662),
.B1(n_1660),
.B2(n_1682),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1690),
.Y(n_1714)
);

INVxp67_ASAP7_75t_L g1715 ( 
.A(n_1703),
.Y(n_1715)
);

O2A1O1Ixp5_ASAP7_75t_L g1716 ( 
.A1(n_1691),
.A2(n_1670),
.B(n_1674),
.C(n_1661),
.Y(n_1716)
);

AND2x2_ASAP7_75t_L g1717 ( 
.A(n_1709),
.B(n_1656),
.Y(n_1717)
);

INVx1_ASAP7_75t_L g1718 ( 
.A(n_1697),
.Y(n_1718)
);

AOI322xp5_ASAP7_75t_L g1719 ( 
.A1(n_1701),
.A2(n_1684),
.A3(n_1680),
.B1(n_1619),
.B2(n_1625),
.C1(n_1627),
.C2(n_1650),
.Y(n_1719)
);

AOI21xp5_ASAP7_75t_L g1720 ( 
.A1(n_1694),
.A2(n_1679),
.B(n_1662),
.Y(n_1720)
);

HB1xp67_ASAP7_75t_L g1721 ( 
.A(n_1688),
.Y(n_1721)
);

OAI31xp33_ASAP7_75t_L g1722 ( 
.A1(n_1689),
.A2(n_1667),
.A3(n_1673),
.B(n_1666),
.Y(n_1722)
);

INVxp33_ASAP7_75t_L g1723 ( 
.A(n_1698),
.Y(n_1723)
);

AOI21xp5_ASAP7_75t_L g1724 ( 
.A1(n_1706),
.A2(n_1702),
.B(n_1693),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_SL g1725 ( 
.A(n_1688),
.B(n_1677),
.Y(n_1725)
);

AOI22xp33_ASAP7_75t_L g1726 ( 
.A1(n_1700),
.A2(n_1650),
.B1(n_1627),
.B2(n_1642),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_L g1727 ( 
.A(n_1707),
.B(n_1665),
.Y(n_1727)
);

INVx1_ASAP7_75t_SL g1728 ( 
.A(n_1692),
.Y(n_1728)
);

INVx1_ASAP7_75t_L g1729 ( 
.A(n_1711),
.Y(n_1729)
);

AND2x4_ASAP7_75t_L g1730 ( 
.A(n_1712),
.B(n_1665),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1696),
.Y(n_1731)
);

OAI21xp33_ASAP7_75t_SL g1732 ( 
.A1(n_1704),
.A2(n_1665),
.B(n_1594),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1721),
.Y(n_1733)
);

AOI21xp5_ASAP7_75t_L g1734 ( 
.A1(n_1724),
.A2(n_1687),
.B(n_1695),
.Y(n_1734)
);

INVx1_ASAP7_75t_L g1735 ( 
.A(n_1728),
.Y(n_1735)
);

OAI31xp33_ASAP7_75t_L g1736 ( 
.A1(n_1722),
.A2(n_1720),
.A3(n_1695),
.B(n_1713),
.Y(n_1736)
);

AOI31xp33_ASAP7_75t_L g1737 ( 
.A1(n_1723),
.A2(n_1710),
.A3(n_1705),
.B(n_1708),
.Y(n_1737)
);

AOI221xp5_ASAP7_75t_L g1738 ( 
.A1(n_1715),
.A2(n_1705),
.B1(n_1650),
.B2(n_1627),
.C(n_1642),
.Y(n_1738)
);

OAI21xp33_ASAP7_75t_SL g1739 ( 
.A1(n_1719),
.A2(n_1699),
.B(n_1620),
.Y(n_1739)
);

OA22x2_ASAP7_75t_L g1740 ( 
.A1(n_1725),
.A2(n_1639),
.B1(n_1636),
.B2(n_1634),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1717),
.B(n_1594),
.Y(n_1741)
);

A2O1A1Ixp33_ASAP7_75t_L g1742 ( 
.A1(n_1716),
.A2(n_1533),
.B(n_1616),
.C(n_1629),
.Y(n_1742)
);

XNOR2xp5_ASAP7_75t_L g1743 ( 
.A(n_1725),
.B(n_1452),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1714),
.Y(n_1744)
);

NAND2xp5_ASAP7_75t_L g1745 ( 
.A(n_1741),
.B(n_1731),
.Y(n_1745)
);

NAND2xp5_ASAP7_75t_L g1746 ( 
.A(n_1735),
.B(n_1718),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1733),
.B(n_1729),
.Y(n_1747)
);

NAND2xp5_ASAP7_75t_L g1748 ( 
.A(n_1734),
.B(n_1727),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1743),
.B(n_1727),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1737),
.B(n_1726),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1736),
.B(n_1730),
.Y(n_1751)
);

NAND2xp5_ASAP7_75t_L g1752 ( 
.A(n_1744),
.B(n_1726),
.Y(n_1752)
);

OAI22xp5_ASAP7_75t_SL g1753 ( 
.A1(n_1739),
.A2(n_1730),
.B1(n_1732),
.B2(n_1448),
.Y(n_1753)
);

NOR3xp33_ASAP7_75t_L g1754 ( 
.A(n_1739),
.B(n_1730),
.C(n_1616),
.Y(n_1754)
);

AOI221xp5_ASAP7_75t_L g1755 ( 
.A1(n_1742),
.A2(n_1629),
.B1(n_1611),
.B2(n_1620),
.C(n_1612),
.Y(n_1755)
);

OAI211xp5_ASAP7_75t_L g1756 ( 
.A1(n_1750),
.A2(n_1754),
.B(n_1748),
.C(n_1752),
.Y(n_1756)
);

A2O1A1Ixp33_ASAP7_75t_L g1757 ( 
.A1(n_1751),
.A2(n_1738),
.B(n_1740),
.C(n_1611),
.Y(n_1757)
);

OAI222xp33_ASAP7_75t_L g1758 ( 
.A1(n_1753),
.A2(n_1636),
.B1(n_1600),
.B2(n_1603),
.C1(n_1579),
.C2(n_1416),
.Y(n_1758)
);

OAI221xp5_ASAP7_75t_L g1759 ( 
.A1(n_1755),
.A2(n_1579),
.B1(n_1603),
.B2(n_1600),
.C(n_1577),
.Y(n_1759)
);

OAI211xp5_ASAP7_75t_L g1760 ( 
.A1(n_1746),
.A2(n_1550),
.B(n_1553),
.C(n_1548),
.Y(n_1760)
);

AOI21xp5_ASAP7_75t_L g1761 ( 
.A1(n_1745),
.A2(n_1607),
.B(n_1593),
.Y(n_1761)
);

XNOR2xp5_ASAP7_75t_L g1762 ( 
.A(n_1756),
.B(n_1749),
.Y(n_1762)
);

CKINVDCx20_ASAP7_75t_R g1763 ( 
.A(n_1761),
.Y(n_1763)
);

AOI221xp5_ASAP7_75t_L g1764 ( 
.A1(n_1757),
.A2(n_1747),
.B1(n_1513),
.B2(n_1603),
.C(n_1579),
.Y(n_1764)
);

AOI321xp33_ASAP7_75t_L g1765 ( 
.A1(n_1759),
.A2(n_1602),
.A3(n_1601),
.B1(n_1446),
.B2(n_1431),
.C(n_1521),
.Y(n_1765)
);

AOI211xp5_ASAP7_75t_L g1766 ( 
.A1(n_1758),
.A2(n_1602),
.B(n_1601),
.C(n_1453),
.Y(n_1766)
);

AOI22xp5_ASAP7_75t_L g1767 ( 
.A1(n_1760),
.A2(n_1602),
.B1(n_1586),
.B2(n_1532),
.Y(n_1767)
);

INVx1_ASAP7_75t_L g1768 ( 
.A(n_1762),
.Y(n_1768)
);

INVx1_ASAP7_75t_L g1769 ( 
.A(n_1763),
.Y(n_1769)
);

AND3x4_ASAP7_75t_L g1770 ( 
.A(n_1766),
.B(n_1548),
.C(n_1550),
.Y(n_1770)
);

AOI22xp5_ASAP7_75t_L g1771 ( 
.A1(n_1764),
.A2(n_1767),
.B1(n_1765),
.B2(n_1532),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1762),
.B(n_1593),
.Y(n_1772)
);

NOR3xp33_ASAP7_75t_SL g1773 ( 
.A(n_1768),
.B(n_1607),
.C(n_1443),
.Y(n_1773)
);

NOR3xp33_ASAP7_75t_L g1774 ( 
.A(n_1769),
.B(n_1453),
.C(n_1493),
.Y(n_1774)
);

AND2x4_ASAP7_75t_L g1775 ( 
.A(n_1772),
.B(n_1548),
.Y(n_1775)
);

NAND2x1_ASAP7_75t_SL g1776 ( 
.A(n_1775),
.B(n_1771),
.Y(n_1776)
);

INVx2_ASAP7_75t_L g1777 ( 
.A(n_1776),
.Y(n_1777)
);

INVx2_ASAP7_75t_L g1778 ( 
.A(n_1777),
.Y(n_1778)
);

INVx2_ASAP7_75t_L g1779 ( 
.A(n_1777),
.Y(n_1779)
);

INVx1_ASAP7_75t_L g1780 ( 
.A(n_1778),
.Y(n_1780)
);

OAI22xp5_ASAP7_75t_L g1781 ( 
.A1(n_1779),
.A2(n_1770),
.B1(n_1773),
.B2(n_1774),
.Y(n_1781)
);

OAI22xp5_ASAP7_75t_L g1782 ( 
.A1(n_1780),
.A2(n_1550),
.B1(n_1553),
.B2(n_1537),
.Y(n_1782)
);

OAI22xp5_ASAP7_75t_L g1783 ( 
.A1(n_1781),
.A2(n_1553),
.B1(n_1531),
.B2(n_1537),
.Y(n_1783)
);

XNOR2xp5_ASAP7_75t_L g1784 ( 
.A(n_1783),
.B(n_1446),
.Y(n_1784)
);

AOI21x1_ASAP7_75t_L g1785 ( 
.A1(n_1784),
.A2(n_1782),
.B(n_1551),
.Y(n_1785)
);

AO21x2_ASAP7_75t_L g1786 ( 
.A1(n_1785),
.A2(n_1551),
.B(n_1545),
.Y(n_1786)
);

OAI221xp5_ASAP7_75t_R g1787 ( 
.A1(n_1786),
.A2(n_1454),
.B1(n_1556),
.B2(n_1545),
.C(n_1541),
.Y(n_1787)
);

AOI211xp5_ASAP7_75t_L g1788 ( 
.A1(n_1787),
.A2(n_1458),
.B(n_1437),
.C(n_1357),
.Y(n_1788)
);


endmodule