module real_aes_6281_n_222 (n_17, n_28, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_165, n_51, n_195, n_176, n_27, n_163, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_169, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_86, n_93, n_182, n_154, n_127, n_199, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_145, n_62, n_105, n_84, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_16, n_116, n_94, n_39, n_5, n_45, n_60, n_38, n_155, n_118, n_143, n_139, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_107, n_184, n_53, n_36, n_222);
input n_17;
input n_28;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_165;
input n_51;
input n_195;
input n_176;
input n_27;
input n_163;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_169;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_145;
input n_62;
input n_105;
input n_84;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_16;
input n_116;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_155;
input n_118;
input n_143;
input n_139;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_107;
input n_184;
input n_53;
input n_36;
output n_222;
wire n_480;
wire n_476;
wire n_599;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_362;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_461;
wire n_242;
wire n_571;
wire n_376;
wire n_549;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_372;
wire n_578;
wire n_528;
wire n_495;
wire n_370;
wire n_384;
wire n_352;
wire n_467;
wire n_327;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_517;
wire n_683;
wire n_570;
wire n_675;
wire n_530;
wire n_535;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_234;
wire n_284;
wire n_532;
wire n_316;
wire n_656;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_671;
wire n_231;
wire n_659;
wire n_547;
wire n_682;
wire n_634;
wire n_454;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_236;
wire n_278;
wire n_367;
wire n_267;
wire n_581;
wire n_610;
wire n_620;
wire n_582;
wire n_641;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_600;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_361;
wire n_632;
wire n_246;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_604;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_588;
wire n_536;
wire n_707;
wire n_622;
wire n_470;
wire n_494;
wire n_377;
wire n_273;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_481;
wire n_498;
wire n_691;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_282;
wire n_389;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_482;
wire n_679;
wire n_520;
wire n_633;
wire n_472;
wire n_452;
wire n_262;
wire n_630;
wire n_689;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_438;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_623;
wire n_249;
wire n_446;
wire n_681;
wire n_359;
wire n_456;
wire n_312;
wire n_266;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_705;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_541;
wire n_224;
wire n_546;
wire n_587;
wire n_639;
wire n_253;
wire n_459;
wire n_558;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_228;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_566;
wire n_474;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_241;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_424;
wire n_225;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
AOI22xp33_ASAP7_75t_L g378 ( .A1(n_0), .A2(n_179), .B1(n_379), .B2(n_380), .Y(n_378) );
AOI222xp33_ASAP7_75t_L g482 ( .A1(n_1), .A2(n_64), .B1(n_202), .B2(n_399), .C1(n_402), .C2(n_442), .Y(n_482) );
INVx1_ASAP7_75t_L g485 ( .A(n_2), .Y(n_485) );
AOI22xp33_ASAP7_75t_L g341 ( .A1(n_3), .A2(n_11), .B1(n_342), .B2(n_343), .Y(n_341) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_4), .A2(n_40), .B1(n_273), .B2(n_286), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_5), .B(n_266), .Y(n_479) );
AOI22xp33_ASAP7_75t_L g670 ( .A1(n_6), .A2(n_138), .B1(n_272), .B2(n_279), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g431 ( .A1(n_7), .A2(n_119), .B1(n_306), .B2(n_432), .Y(n_431) );
AOI22xp33_ASAP7_75t_L g581 ( .A1(n_8), .A2(n_93), .B1(n_301), .B2(n_380), .Y(n_581) );
AOI222xp33_ASAP7_75t_L g537 ( .A1(n_9), .A2(n_94), .B1(n_169), .B2(n_295), .C1(n_401), .C2(n_538), .Y(n_537) );
AOI22xp33_ASAP7_75t_L g392 ( .A1(n_10), .A2(n_112), .B1(n_393), .B2(n_394), .Y(n_392) );
AOI222xp33_ASAP7_75t_L g364 ( .A1(n_12), .A2(n_62), .B1(n_111), .B2(n_242), .C1(n_365), .C2(n_366), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g439 ( .A(n_13), .B(n_394), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g555 ( .A1(n_14), .A2(n_133), .B1(n_311), .B2(n_556), .Y(n_555) );
CKINVDCx20_ASAP7_75t_R g514 ( .A(n_15), .Y(n_514) );
AO22x2_ASAP7_75t_L g245 ( .A1(n_16), .A2(n_68), .B1(n_246), .B2(n_247), .Y(n_245) );
INVx1_ASAP7_75t_L g639 ( .A(n_16), .Y(n_639) );
NAND2xp5_ASAP7_75t_SL g550 ( .A(n_17), .B(n_551), .Y(n_550) );
AOI22xp33_ASAP7_75t_L g529 ( .A1(n_18), .A2(n_158), .B1(n_452), .B2(n_530), .Y(n_529) );
AOI22xp33_ASAP7_75t_SL g494 ( .A1(n_19), .A2(n_105), .B1(n_303), .B2(n_495), .Y(n_494) );
CKINVDCx20_ASAP7_75t_R g573 ( .A(n_20), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_21), .A2(n_35), .B1(n_354), .B2(n_686), .Y(n_685) );
AOI22xp5_ASAP7_75t_L g453 ( .A1(n_22), .A2(n_220), .B1(n_432), .B2(n_454), .Y(n_453) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_23), .A2(n_130), .B1(n_345), .B2(n_560), .Y(n_618) );
AOI22xp5_ASAP7_75t_L g422 ( .A1(n_24), .A2(n_201), .B1(n_423), .B2(n_424), .Y(n_422) );
CKINVDCx20_ASAP7_75t_R g698 ( .A(n_25), .Y(n_698) );
AOI222xp33_ASAP7_75t_L g398 ( .A1(n_26), .A2(n_154), .B1(n_195), .B2(n_399), .C1(n_401), .C2(n_402), .Y(n_398) );
CKINVDCx20_ASAP7_75t_R g658 ( .A(n_27), .Y(n_658) );
AOI22xp33_ASAP7_75t_L g467 ( .A1(n_28), .A2(n_193), .B1(n_303), .B2(n_468), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_29), .B(n_393), .Y(n_535) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_30), .Y(n_291) );
INVx1_ASAP7_75t_L g416 ( .A(n_31), .Y(n_416) );
AOI22xp33_ASAP7_75t_SL g552 ( .A1(n_32), .A2(n_139), .B1(n_273), .B2(n_447), .Y(n_552) );
AO22x2_ASAP7_75t_L g249 ( .A1(n_33), .A2(n_71), .B1(n_246), .B2(n_250), .Y(n_249) );
INVx1_ASAP7_75t_L g640 ( .A(n_33), .Y(n_640) );
CKINVDCx20_ASAP7_75t_R g327 ( .A(n_34), .Y(n_327) );
AOI22xp33_ASAP7_75t_L g353 ( .A1(n_36), .A2(n_63), .B1(n_354), .B2(n_355), .Y(n_353) );
CKINVDCx20_ASAP7_75t_R g546 ( .A(n_37), .Y(n_546) );
AOI22xp33_ASAP7_75t_L g693 ( .A1(n_38), .A2(n_72), .B1(n_620), .B2(n_694), .Y(n_693) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_39), .A2(n_97), .B1(n_350), .B2(n_651), .Y(n_650) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_41), .A2(n_51), .B1(n_303), .B2(n_427), .Y(n_459) );
CKINVDCx20_ASAP7_75t_R g589 ( .A(n_42), .Y(n_589) );
CKINVDCx20_ASAP7_75t_R g318 ( .A(n_43), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g604 ( .A(n_44), .Y(n_604) );
AOI22xp33_ASAP7_75t_L g465 ( .A1(n_45), .A2(n_172), .B1(n_386), .B2(n_466), .Y(n_465) );
CKINVDCx20_ASAP7_75t_R g614 ( .A(n_46), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g621 ( .A1(n_47), .A2(n_215), .B1(n_379), .B2(n_490), .Y(n_621) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_48), .A2(n_122), .B1(n_279), .B2(n_443), .Y(n_536) );
AOI22xp33_ASAP7_75t_L g310 ( .A1(n_49), .A2(n_153), .B1(n_311), .B2(n_315), .Y(n_310) );
AOI22xp33_ASAP7_75t_SL g554 ( .A1(n_50), .A2(n_159), .B1(n_379), .B2(n_432), .Y(n_554) );
CKINVDCx20_ASAP7_75t_R g500 ( .A(n_52), .Y(n_500) );
XNOR2x2_ASAP7_75t_L g462 ( .A(n_53), .B(n_463), .Y(n_462) );
CKINVDCx20_ASAP7_75t_R g609 ( .A(n_54), .Y(n_609) );
AO22x2_ASAP7_75t_L g600 ( .A1(n_55), .A2(n_601), .B1(n_623), .B2(n_624), .Y(n_600) );
CKINVDCx20_ASAP7_75t_R g624 ( .A(n_55), .Y(n_624) );
AOI22xp33_ASAP7_75t_L g619 ( .A1(n_56), .A2(n_184), .B1(n_556), .B2(n_620), .Y(n_619) );
AOI22xp33_ASAP7_75t_SL g663 ( .A1(n_57), .A2(n_132), .B1(n_571), .B2(n_664), .Y(n_663) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_58), .Y(n_257) );
AOI211xp5_ASAP7_75t_L g241 ( .A1(n_59), .A2(n_242), .B(n_256), .C(n_283), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_60), .A2(n_190), .B1(n_647), .B2(n_648), .Y(n_646) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_61), .A2(n_174), .B1(n_359), .B2(n_361), .Y(n_358) );
INVx1_ASAP7_75t_L g434 ( .A(n_65), .Y(n_434) );
AOI22xp5_ASAP7_75t_SL g488 ( .A1(n_66), .A2(n_120), .B1(n_345), .B2(n_424), .Y(n_488) );
AOI22xp33_ASAP7_75t_L g692 ( .A1(n_67), .A2(n_118), .B1(n_375), .B2(n_384), .Y(n_692) );
AOI22xp33_ASAP7_75t_L g570 ( .A1(n_69), .A2(n_109), .B1(n_365), .B2(n_571), .Y(n_570) );
AOI22xp33_ASAP7_75t_L g382 ( .A1(n_70), .A2(n_212), .B1(n_383), .B2(n_384), .Y(n_382) );
INVx1_ASAP7_75t_L g230 ( .A(n_73), .Y(n_230) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_74), .A2(n_207), .B1(n_388), .B2(n_390), .Y(n_387) );
INVx1_ASAP7_75t_L g460 ( .A(n_75), .Y(n_460) );
AOI22xp33_ASAP7_75t_L g470 ( .A1(n_76), .A2(n_100), .B1(n_330), .B2(n_471), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_77), .A2(n_107), .B1(n_301), .B2(n_306), .Y(n_356) );
AOI22xp5_ASAP7_75t_SL g492 ( .A1(n_78), .A2(n_189), .B1(n_454), .B2(n_493), .Y(n_492) );
AOI22xp33_ASAP7_75t_L g300 ( .A1(n_79), .A2(n_161), .B1(n_301), .B2(n_306), .Y(n_300) );
AOI22xp5_ASAP7_75t_L g510 ( .A1(n_80), .A2(n_147), .B1(n_279), .B2(n_402), .Y(n_510) );
INVx1_ASAP7_75t_L g228 ( .A(n_81), .Y(n_228) );
AOI22xp33_ASAP7_75t_SL g547 ( .A1(n_82), .A2(n_117), .B1(n_296), .B2(n_442), .Y(n_547) );
CKINVDCx20_ASAP7_75t_R g653 ( .A(n_83), .Y(n_653) );
XOR2x2_ASAP7_75t_L g370 ( .A(n_84), .B(n_371), .Y(n_370) );
AOI22xp33_ASAP7_75t_L g473 ( .A1(n_85), .A2(n_148), .B1(n_311), .B2(n_474), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_86), .B(n_413), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_87), .A2(n_192), .B1(n_426), .B2(n_532), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g441 ( .A1(n_88), .A2(n_170), .B1(n_442), .B2(n_443), .Y(n_441) );
CKINVDCx20_ASAP7_75t_R g567 ( .A(n_89), .Y(n_567) );
AOI22xp5_ASAP7_75t_L g489 ( .A1(n_90), .A2(n_134), .B1(n_325), .B2(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_91), .B(n_393), .Y(n_440) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_92), .A2(n_141), .B1(n_451), .B2(n_452), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_95), .B(n_669), .Y(n_668) );
CKINVDCx20_ASAP7_75t_R g662 ( .A(n_96), .Y(n_662) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_98), .B(n_413), .Y(n_667) );
INVx1_ASAP7_75t_L g445 ( .A(n_99), .Y(n_445) );
CKINVDCx20_ASAP7_75t_R g702 ( .A(n_101), .Y(n_702) );
AOI22xp33_ASAP7_75t_L g527 ( .A1(n_102), .A2(n_185), .B1(n_351), .B2(n_458), .Y(n_527) );
AOI22xp33_ASAP7_75t_L g395 ( .A1(n_103), .A2(n_188), .B1(n_279), .B2(n_396), .Y(n_395) );
CKINVDCx20_ASAP7_75t_R g578 ( .A(n_104), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g271 ( .A1(n_106), .A2(n_166), .B1(n_272), .B2(n_277), .Y(n_271) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_108), .A2(n_213), .B1(n_350), .B2(n_388), .Y(n_582) );
AOI22xp5_ASAP7_75t_SL g562 ( .A1(n_110), .A2(n_563), .B1(n_593), .B2(n_594), .Y(n_562) );
INVx1_ASAP7_75t_L g594 ( .A(n_110), .Y(n_594) );
CKINVDCx20_ASAP7_75t_R g655 ( .A(n_113), .Y(n_655) );
CKINVDCx20_ASAP7_75t_R g539 ( .A(n_114), .Y(n_539) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_115), .B(n_266), .Y(n_265) );
INVx2_ASAP7_75t_L g231 ( .A(n_116), .Y(n_231) );
CKINVDCx20_ASAP7_75t_R g708 ( .A(n_121), .Y(n_708) );
AOI22xp33_ASAP7_75t_L g363 ( .A1(n_123), .A2(n_181), .B1(n_272), .B2(n_280), .Y(n_363) );
CKINVDCx20_ASAP7_75t_R g284 ( .A(n_124), .Y(n_284) );
AOI22xp33_ASAP7_75t_L g480 ( .A1(n_125), .A2(n_163), .B1(n_396), .B2(n_481), .Y(n_480) );
CKINVDCx20_ASAP7_75t_R g566 ( .A(n_126), .Y(n_566) );
CKINVDCx16_ASAP7_75t_R g239 ( .A(n_127), .Y(n_239) );
AND2x6_ASAP7_75t_L g227 ( .A(n_128), .B(n_228), .Y(n_227) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_128), .Y(n_633) );
AO22x2_ASAP7_75t_L g253 ( .A1(n_129), .A2(n_180), .B1(n_246), .B2(n_250), .Y(n_253) );
AOI22xp33_ASAP7_75t_L g526 ( .A1(n_131), .A2(n_199), .B1(n_429), .B2(n_490), .Y(n_526) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_135), .Y(n_509) );
AOI22xp33_ASAP7_75t_SL g428 ( .A1(n_136), .A2(n_204), .B1(n_345), .B2(n_429), .Y(n_428) );
CKINVDCx20_ASAP7_75t_R g534 ( .A(n_137), .Y(n_534) );
CKINVDCx20_ASAP7_75t_R g512 ( .A(n_140), .Y(n_512) );
AOI22xp33_ASAP7_75t_SL g456 ( .A1(n_142), .A2(n_157), .B1(n_457), .B2(n_458), .Y(n_456) );
AOI211xp5_ASAP7_75t_L g222 ( .A1(n_143), .A2(n_223), .B(n_232), .C(n_641), .Y(n_222) );
AOI22xp5_ASAP7_75t_SL g642 ( .A1(n_144), .A2(n_643), .B1(n_671), .B2(n_672), .Y(n_642) );
CKINVDCx20_ASAP7_75t_R g672 ( .A(n_144), .Y(n_672) );
AOI22xp33_ASAP7_75t_L g622 ( .A1(n_145), .A2(n_203), .B1(n_451), .B2(n_532), .Y(n_622) );
AOI22xp33_ASAP7_75t_SL g558 ( .A1(n_146), .A2(n_196), .B1(n_452), .B2(n_454), .Y(n_558) );
CKINVDCx20_ASAP7_75t_R g561 ( .A(n_149), .Y(n_561) );
AO22x2_ASAP7_75t_L g255 ( .A1(n_150), .A2(n_194), .B1(n_246), .B2(n_247), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g446 ( .A1(n_151), .A2(n_211), .B1(n_295), .B2(n_447), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g587 ( .A(n_152), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g611 ( .A1(n_155), .A2(n_198), .B1(n_293), .B2(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g332 ( .A(n_156), .Y(n_332) );
CKINVDCx20_ASAP7_75t_R g659 ( .A(n_160), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g418 ( .A1(n_162), .A2(n_218), .B1(n_419), .B2(n_420), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_164), .B(n_393), .Y(n_411) );
AOI22xp33_ASAP7_75t_SL g559 ( .A1(n_165), .A2(n_197), .B1(n_320), .B2(n_560), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g347 ( .A1(n_167), .A2(n_219), .B1(n_348), .B2(n_350), .Y(n_347) );
CKINVDCx20_ASAP7_75t_R g592 ( .A(n_168), .Y(n_592) );
CKINVDCx20_ASAP7_75t_R g616 ( .A(n_171), .Y(n_616) );
CKINVDCx20_ASAP7_75t_R g476 ( .A(n_173), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_175), .B(n_571), .Y(n_704) );
CKINVDCx20_ASAP7_75t_R g323 ( .A(n_176), .Y(n_323) );
AOI22xp33_ASAP7_75t_SL g425 ( .A1(n_177), .A2(n_187), .B1(n_426), .B2(n_427), .Y(n_425) );
CKINVDCx20_ASAP7_75t_R g569 ( .A(n_178), .Y(n_569) );
NOR2xp33_ASAP7_75t_L g637 ( .A(n_180), .B(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_182), .B(n_413), .Y(n_549) );
CKINVDCx20_ASAP7_75t_R g706 ( .A(n_183), .Y(n_706) );
CKINVDCx20_ASAP7_75t_R g584 ( .A(n_186), .Y(n_584) );
CKINVDCx20_ASAP7_75t_R g607 ( .A(n_191), .Y(n_607) );
INVx1_ASAP7_75t_L g636 ( .A(n_194), .Y(n_636) );
CKINVDCx20_ASAP7_75t_R g697 ( .A(n_200), .Y(n_697) );
INVx1_ASAP7_75t_L g680 ( .A(n_205), .Y(n_680) );
AOI22xp5_ASAP7_75t_L g681 ( .A1(n_205), .A2(n_680), .B1(n_682), .B2(n_709), .Y(n_681) );
CKINVDCx20_ASAP7_75t_R g504 ( .A(n_206), .Y(n_504) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_208), .A2(n_210), .B1(n_374), .B2(n_375), .Y(n_373) );
INVx1_ASAP7_75t_L g246 ( .A(n_209), .Y(n_246) );
INVx1_ASAP7_75t_L g248 ( .A(n_209), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g703 ( .A(n_214), .Y(n_703) );
AOI22xp33_ASAP7_75t_L g687 ( .A1(n_216), .A2(n_221), .B1(n_688), .B2(n_690), .Y(n_687) );
OA22x2_ASAP7_75t_L g337 ( .A1(n_217), .A2(n_338), .B1(n_339), .B2(n_367), .Y(n_337) );
INVx1_ASAP7_75t_L g338 ( .A(n_217), .Y(n_338) );
CKINVDCx20_ASAP7_75t_R g223 ( .A(n_224), .Y(n_223) );
CKINVDCx20_ASAP7_75t_R g224 ( .A(n_225), .Y(n_224) );
HB1xp67_ASAP7_75t_L g225 ( .A(n_226), .Y(n_225) );
AND2x4_ASAP7_75t_L g226 ( .A(n_227), .B(n_229), .Y(n_226) );
HB1xp67_ASAP7_75t_L g632 ( .A(n_228), .Y(n_632) );
OAI21xp5_ASAP7_75t_L g678 ( .A1(n_229), .A2(n_631), .B(n_679), .Y(n_678) );
AND2x2_ASAP7_75t_L g229 ( .A(n_230), .B(n_231), .Y(n_229) );
AOI221xp5_ASAP7_75t_L g232 ( .A1(n_233), .A2(n_520), .B1(n_626), .B2(n_627), .C(n_628), .Y(n_232) );
INVx1_ASAP7_75t_L g626 ( .A(n_233), .Y(n_626) );
AOI22xp5_ASAP7_75t_L g233 ( .A1(n_234), .A2(n_235), .B1(n_369), .B2(n_519), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_235), .Y(n_234) );
AOI22xp5_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_336), .B1(n_337), .B2(n_368), .Y(n_235) );
INVx1_ASAP7_75t_SL g368 ( .A(n_236), .Y(n_368) );
INVx1_ASAP7_75t_L g236 ( .A(n_237), .Y(n_236) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
XNOR2xp5_ASAP7_75t_L g238 ( .A(n_239), .B(n_240), .Y(n_238) );
AND2x2_ASAP7_75t_L g240 ( .A(n_241), .B(n_298), .Y(n_240) );
INVx3_ASAP7_75t_L g610 ( .A(n_242), .Y(n_610) );
BUFx3_ASAP7_75t_L g242 ( .A(n_243), .Y(n_242) );
INVx4_ASAP7_75t_L g400 ( .A(n_243), .Y(n_400) );
INVx2_ASAP7_75t_L g417 ( .A(n_243), .Y(n_417) );
BUFx6f_ASAP7_75t_L g538 ( .A(n_243), .Y(n_538) );
AND2x6_ASAP7_75t_L g243 ( .A(n_244), .B(n_251), .Y(n_243) );
AND2x4_ASAP7_75t_L g280 ( .A(n_244), .B(n_281), .Y(n_280) );
INVx1_ASAP7_75t_L g576 ( .A(n_244), .Y(n_576) );
AND2x2_ASAP7_75t_L g244 ( .A(n_245), .B(n_249), .Y(n_244) );
INVx2_ASAP7_75t_L g263 ( .A(n_245), .Y(n_263) );
AND2x2_ASAP7_75t_L g276 ( .A(n_245), .B(n_253), .Y(n_276) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
INVx1_ASAP7_75t_L g250 ( .A(n_248), .Y(n_250) );
AND2x2_ASAP7_75t_L g262 ( .A(n_249), .B(n_263), .Y(n_262) );
OR2x2_ASAP7_75t_L g270 ( .A(n_249), .B(n_263), .Y(n_270) );
INVx1_ASAP7_75t_L g275 ( .A(n_249), .Y(n_275) );
INVx2_ASAP7_75t_L g290 ( .A(n_249), .Y(n_290) );
AND2x6_ASAP7_75t_L g322 ( .A(n_251), .B(n_269), .Y(n_322) );
AND2x4_ASAP7_75t_L g325 ( .A(n_251), .B(n_262), .Y(n_325) );
AND2x2_ASAP7_75t_L g331 ( .A(n_251), .B(n_305), .Y(n_331) );
AND2x2_ASAP7_75t_L g251 ( .A(n_252), .B(n_254), .Y(n_251) );
AND2x2_ASAP7_75t_L g264 ( .A(n_252), .B(n_255), .Y(n_264) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_253), .B(n_255), .Y(n_309) );
AND2x2_ASAP7_75t_L g314 ( .A(n_253), .B(n_282), .Y(n_314) );
INVx1_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
INVx1_ASAP7_75t_L g282 ( .A(n_255), .Y(n_282) );
INVx1_ASAP7_75t_L g289 ( .A(n_255), .Y(n_289) );
OAI211xp5_ASAP7_75t_L g256 ( .A1(n_257), .A2(n_258), .B(n_265), .C(n_271), .Y(n_256) );
INVx2_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
INVx2_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
OA211x2_ASAP7_75t_L g533 ( .A1(n_260), .A2(n_534), .B(n_535), .C(n_536), .Y(n_533) );
OAI22xp5_ASAP7_75t_SL g565 ( .A1(n_260), .A2(n_507), .B1(n_566), .B2(n_567), .Y(n_565) );
BUFx3_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
INVx1_ASAP7_75t_L g478 ( .A(n_261), .Y(n_478) );
NAND2x1p5_ASAP7_75t_L g261 ( .A(n_262), .B(n_264), .Y(n_261) );
AND2x2_ASAP7_75t_L g313 ( .A(n_262), .B(n_314), .Y(n_313) );
AND2x6_ASAP7_75t_L g362 ( .A(n_262), .B(n_264), .Y(n_362) );
AND2x2_ASAP7_75t_L g305 ( .A(n_263), .B(n_290), .Y(n_305) );
AND2x4_ASAP7_75t_L g268 ( .A(n_264), .B(n_269), .Y(n_268) );
AND2x4_ASAP7_75t_L g304 ( .A(n_264), .B(n_305), .Y(n_304) );
INVx1_ASAP7_75t_L g508 ( .A(n_264), .Y(n_508) );
INVx2_ASAP7_75t_L g266 ( .A(n_267), .Y(n_266) );
INVx5_ASAP7_75t_L g360 ( .A(n_267), .Y(n_360) );
INVx2_ASAP7_75t_L g393 ( .A(n_267), .Y(n_393) );
INVx2_ASAP7_75t_L g551 ( .A(n_267), .Y(n_551) );
INVx4_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
INVx2_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
OR2x2_ASAP7_75t_L g507 ( .A(n_270), .B(n_508), .Y(n_507) );
BUFx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
INVx1_ASAP7_75t_L g397 ( .A(n_273), .Y(n_397) );
BUFx3_ASAP7_75t_L g443 ( .A(n_273), .Y(n_443) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
OR2x6_ASAP7_75t_L g316 ( .A(n_275), .B(n_309), .Y(n_316) );
AND2x4_ASAP7_75t_L g287 ( .A(n_276), .B(n_288), .Y(n_287) );
AND2x4_ASAP7_75t_L g296 ( .A(n_276), .B(n_297), .Y(n_296) );
NAND2x1p5_ASAP7_75t_L g503 ( .A(n_276), .B(n_496), .Y(n_503) );
INVx2_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_SL g278 ( .A(n_279), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_280), .Y(n_279) );
BUFx2_ASAP7_75t_SL g420 ( .A(n_280), .Y(n_420) );
BUFx3_ASAP7_75t_L g447 ( .A(n_280), .Y(n_447) );
BUFx2_ASAP7_75t_SL g481 ( .A(n_280), .Y(n_481) );
INVx1_ASAP7_75t_L g577 ( .A(n_281), .Y(n_577) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI22xp5_ASAP7_75t_L g283 ( .A1(n_284), .A2(n_285), .B1(n_291), .B2(n_292), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
BUFx6f_ASAP7_75t_L g286 ( .A(n_287), .Y(n_286) );
BUFx4f_ASAP7_75t_SL g365 ( .A(n_287), .Y(n_365) );
BUFx6f_ASAP7_75t_L g401 ( .A(n_287), .Y(n_401) );
BUFx6f_ASAP7_75t_L g442 ( .A(n_287), .Y(n_442) );
BUFx2_ASAP7_75t_L g612 ( .A(n_287), .Y(n_612) );
AND2x2_ASAP7_75t_L g288 ( .A(n_289), .B(n_290), .Y(n_288) );
INVx1_ASAP7_75t_L g297 ( .A(n_289), .Y(n_297) );
INVx1_ASAP7_75t_L g496 ( .A(n_290), .Y(n_496) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx3_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
BUFx4f_ASAP7_75t_SL g366 ( .A(n_295), .Y(n_366) );
BUFx12f_ASAP7_75t_L g295 ( .A(n_296), .Y(n_295) );
BUFx6f_ASAP7_75t_L g402 ( .A(n_296), .Y(n_402) );
BUFx6f_ASAP7_75t_L g419 ( .A(n_296), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g298 ( .A(n_299), .B(n_317), .C(n_326), .Y(n_298) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_300), .B(n_310), .Y(n_299) );
INVx3_ASAP7_75t_L g301 ( .A(n_302), .Y(n_301) );
INVx4_ASAP7_75t_L g647 ( .A(n_302), .Y(n_647) );
INVx4_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
BUFx6f_ASAP7_75t_L g303 ( .A(n_304), .Y(n_303) );
BUFx3_ASAP7_75t_L g379 ( .A(n_304), .Y(n_379) );
BUFx3_ASAP7_75t_L g426 ( .A(n_304), .Y(n_426) );
INVx2_ASAP7_75t_L g689 ( .A(n_304), .Y(n_689) );
AND2x4_ASAP7_75t_L g307 ( .A(n_305), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g335 ( .A(n_305), .B(n_314), .Y(n_335) );
AND2x2_ASAP7_75t_L g346 ( .A(n_305), .B(n_314), .Y(n_346) );
BUFx2_ASAP7_75t_L g306 ( .A(n_307), .Y(n_306) );
BUFx3_ASAP7_75t_L g380 ( .A(n_307), .Y(n_380) );
BUFx3_ASAP7_75t_L g454 ( .A(n_307), .Y(n_454) );
BUFx2_ASAP7_75t_SL g468 ( .A(n_307), .Y(n_468) );
BUFx3_ASAP7_75t_L g532 ( .A(n_307), .Y(n_532) );
AND2x2_ASAP7_75t_L g495 ( .A(n_308), .B(n_496), .Y(n_495) );
INVx1_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx1_ASAP7_75t_L g311 ( .A(n_312), .Y(n_311) );
INVx4_ASAP7_75t_L g349 ( .A(n_312), .Y(n_349) );
INVx3_ASAP7_75t_L g424 ( .A(n_312), .Y(n_424) );
INVx5_ASAP7_75t_L g458 ( .A(n_312), .Y(n_458) );
INVx2_ASAP7_75t_L g620 ( .A(n_312), .Y(n_620) );
INVx8_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
INVx1_ASAP7_75t_SL g315 ( .A(n_316), .Y(n_315) );
INVx6_ASAP7_75t_SL g351 ( .A(n_316), .Y(n_351) );
INVx1_ASAP7_75t_SL g427 ( .A(n_316), .Y(n_427) );
INVx1_ASAP7_75t_L g474 ( .A(n_316), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_319), .B1(n_323), .B2(n_324), .Y(n_317) );
INVx1_ASAP7_75t_L g319 ( .A(n_320), .Y(n_319) );
INVx3_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
INVx2_ASAP7_75t_SL g355 ( .A(n_321), .Y(n_355) );
INVx4_ASAP7_75t_L g374 ( .A(n_321), .Y(n_374) );
INVx4_ASAP7_75t_L g493 ( .A(n_321), .Y(n_493) );
INVx11_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx11_ASAP7_75t_L g430 ( .A(n_322), .Y(n_430) );
INVx2_ASAP7_75t_L g342 ( .A(n_324), .Y(n_342) );
INVx2_ASAP7_75t_L g423 ( .A(n_324), .Y(n_423) );
INVx3_ASAP7_75t_L g530 ( .A(n_324), .Y(n_530) );
OAI22xp5_ASAP7_75t_L g583 ( .A1(n_324), .A2(n_584), .B1(n_585), .B2(n_587), .Y(n_583) );
INVx6_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
BUFx3_ASAP7_75t_L g386 ( .A(n_325), .Y(n_386) );
BUFx3_ASAP7_75t_L g457 ( .A(n_325), .Y(n_457) );
BUFx3_ASAP7_75t_L g560 ( .A(n_325), .Y(n_560) );
OAI22xp5_ASAP7_75t_L g326 ( .A1(n_327), .A2(n_328), .B1(n_332), .B2(n_333), .Y(n_326) );
INVx1_ASAP7_75t_SL g328 ( .A(n_329), .Y(n_328) );
BUFx6f_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
BUFx3_ASAP7_75t_L g354 ( .A(n_330), .Y(n_354) );
BUFx6f_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
BUFx2_ASAP7_75t_SL g383 ( .A(n_331), .Y(n_383) );
INVx2_ASAP7_75t_L g433 ( .A(n_331), .Y(n_433) );
BUFx2_ASAP7_75t_SL g591 ( .A(n_331), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g588 ( .A1(n_333), .A2(n_589), .B1(n_590), .B2(n_592), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_333), .A2(n_590), .B1(n_658), .B2(n_659), .Y(n_657) );
INVx1_ASAP7_75t_L g333 ( .A(n_334), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
INVx1_ASAP7_75t_L g336 ( .A(n_337), .Y(n_336) );
INVx1_ASAP7_75t_SL g367 ( .A(n_339), .Y(n_367) );
NAND4xp75_ASAP7_75t_L g339 ( .A(n_340), .B(n_352), .C(n_357), .D(n_364), .Y(n_339) );
AND2x2_ASAP7_75t_L g340 ( .A(n_341), .B(n_347), .Y(n_340) );
INVx2_ASAP7_75t_L g343 ( .A(n_344), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
BUFx3_ASAP7_75t_L g345 ( .A(n_346), .Y(n_345) );
BUFx3_ASAP7_75t_L g377 ( .A(n_346), .Y(n_377) );
BUFx3_ASAP7_75t_L g452 ( .A(n_346), .Y(n_452) );
BUFx3_ASAP7_75t_L g472 ( .A(n_346), .Y(n_472) );
BUFx2_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx2_ASAP7_75t_L g389 ( .A(n_349), .Y(n_389) );
BUFx6f_ASAP7_75t_L g651 ( .A(n_349), .Y(n_651) );
BUFx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
BUFx2_ASAP7_75t_L g390 ( .A(n_351), .Y(n_390) );
BUFx2_ASAP7_75t_L g556 ( .A(n_351), .Y(n_556) );
BUFx2_ASAP7_75t_L g694 ( .A(n_351), .Y(n_694) );
AND2x2_ASAP7_75t_L g352 ( .A(n_353), .B(n_356), .Y(n_352) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_358), .B(n_363), .Y(n_357) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
HB1xp67_ASAP7_75t_L g669 ( .A(n_360), .Y(n_669) );
BUFx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
BUFx2_ASAP7_75t_L g394 ( .A(n_362), .Y(n_394) );
BUFx4f_ASAP7_75t_L g413 ( .A(n_362), .Y(n_413) );
INVx1_ASAP7_75t_L g519 ( .A(n_369), .Y(n_519) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_370), .A2(n_403), .B1(n_404), .B2(n_518), .Y(n_369) );
INVx1_ASAP7_75t_L g518 ( .A(n_370), .Y(n_518) );
NAND4xp75_ASAP7_75t_L g371 ( .A(n_372), .B(n_381), .C(n_391), .D(n_398), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_373), .B(n_378), .Y(n_372) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
INVx2_ASAP7_75t_L g649 ( .A(n_380), .Y(n_649) );
AND2x2_ASAP7_75t_L g381 ( .A(n_382), .B(n_387), .Y(n_381) );
INVx2_ASAP7_75t_L g384 ( .A(n_385), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx3_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
AND2x2_ASAP7_75t_SL g391 ( .A(n_392), .B(n_395), .Y(n_391) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g701 ( .A(n_399), .Y(n_701) );
INVx4_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
OAI22xp5_ASAP7_75t_SL g511 ( .A1(n_400), .A2(n_512), .B1(n_513), .B2(n_514), .Y(n_511) );
OAI21xp5_ASAP7_75t_SL g568 ( .A1(n_400), .A2(n_569), .B(n_570), .Y(n_568) );
OAI21xp5_ASAP7_75t_SL g661 ( .A1(n_400), .A2(n_662), .B(n_663), .Y(n_661) );
BUFx4f_ASAP7_75t_L g571 ( .A(n_402), .Y(n_571) );
INVx1_ASAP7_75t_L g403 ( .A(n_404), .Y(n_403) );
OAI22xp5_ASAP7_75t_L g404 ( .A1(n_405), .A2(n_406), .B1(n_461), .B2(n_517), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
XOR2x2_ASAP7_75t_L g406 ( .A(n_407), .B(n_435), .Y(n_406) );
XOR2x2_ASAP7_75t_L g407 ( .A(n_408), .B(n_434), .Y(n_407) );
NAND4xp75_ASAP7_75t_SL g408 ( .A(n_409), .B(n_421), .C(n_428), .D(n_431), .Y(n_408) );
NOR2xp67_ASAP7_75t_SL g409 ( .A(n_410), .B(n_415), .Y(n_409) );
NAND3xp33_ASAP7_75t_L g410 ( .A(n_411), .B(n_412), .C(n_414), .Y(n_410) );
OAI21xp5_ASAP7_75t_L g415 ( .A1(n_416), .A2(n_417), .B(n_418), .Y(n_415) );
OAI21xp5_ASAP7_75t_SL g444 ( .A1(n_417), .A2(n_445), .B(n_446), .Y(n_444) );
OAI21xp5_ASAP7_75t_SL g545 ( .A1(n_417), .A2(n_546), .B(n_547), .Y(n_545) );
AND2x2_ASAP7_75t_L g421 ( .A(n_422), .B(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g654 ( .A(n_429), .Y(n_654) );
INVx5_ASAP7_75t_SL g429 ( .A(n_430), .Y(n_429) );
INVx2_ASAP7_75t_SL g451 ( .A(n_430), .Y(n_451) );
INVx1_ASAP7_75t_L g466 ( .A(n_430), .Y(n_466) );
INVx4_ASAP7_75t_L g586 ( .A(n_430), .Y(n_586) );
INVx3_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx3_ASAP7_75t_L g490 ( .A(n_433), .Y(n_490) );
XOR2x2_ASAP7_75t_SL g435 ( .A(n_436), .B(n_460), .Y(n_435) );
NAND2x1p5_ASAP7_75t_L g436 ( .A(n_437), .B(n_448), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g437 ( .A(n_438), .B(n_444), .Y(n_437) );
NAND3xp33_ASAP7_75t_L g438 ( .A(n_439), .B(n_440), .C(n_441), .Y(n_438) );
INVx2_ASAP7_75t_L g513 ( .A(n_442), .Y(n_513) );
INVx4_ASAP7_75t_L g665 ( .A(n_442), .Y(n_665) );
NOR2x1_ASAP7_75t_L g448 ( .A(n_449), .B(n_455), .Y(n_448) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .Y(n_449) );
BUFx2_ASAP7_75t_L g690 ( .A(n_454), .Y(n_690) );
NAND2xp5_ASAP7_75t_L g455 ( .A(n_456), .B(n_459), .Y(n_455) );
INVx1_ASAP7_75t_L g656 ( .A(n_457), .Y(n_656) );
INVx1_ASAP7_75t_L g517 ( .A(n_461), .Y(n_517) );
OAI22xp5_ASAP7_75t_SL g461 ( .A1(n_462), .A2(n_483), .B1(n_515), .B2(n_516), .Y(n_461) );
INVx1_ASAP7_75t_L g515 ( .A(n_462), .Y(n_515) );
NAND4xp75_ASAP7_75t_L g463 ( .A(n_464), .B(n_469), .C(n_475), .D(n_482), .Y(n_463) );
AND2x2_ASAP7_75t_L g464 ( .A(n_465), .B(n_467), .Y(n_464) );
AND2x2_ASAP7_75t_L g469 ( .A(n_470), .B(n_473), .Y(n_469) );
BUFx4f_ASAP7_75t_SL g471 ( .A(n_472), .Y(n_471) );
OA211x2_ASAP7_75t_L g475 ( .A1(n_476), .A2(n_477), .B(n_479), .C(n_480), .Y(n_475) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_L g499 ( .A(n_478), .Y(n_499) );
INVx1_ASAP7_75t_SL g699 ( .A(n_478), .Y(n_699) );
INVx1_ASAP7_75t_SL g516 ( .A(n_483), .Y(n_516) );
HB1xp67_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
XNOR2xp5_ASAP7_75t_L g484 ( .A(n_485), .B(n_486), .Y(n_484) );
NAND3x1_ASAP7_75t_SL g486 ( .A(n_487), .B(n_491), .C(n_497), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_488), .B(n_489), .Y(n_487) );
AND2x2_ASAP7_75t_L g491 ( .A(n_492), .B(n_494), .Y(n_491) );
NOR3xp33_ASAP7_75t_L g497 ( .A(n_498), .B(n_505), .C(n_511), .Y(n_497) );
OAI22xp5_ASAP7_75t_SL g498 ( .A1(n_499), .A2(n_500), .B1(n_501), .B2(n_504), .Y(n_498) );
OAI22xp5_ASAP7_75t_L g603 ( .A1(n_499), .A2(n_604), .B1(n_605), .B2(n_607), .Y(n_603) );
OAI22xp5_ASAP7_75t_SL g572 ( .A1(n_501), .A2(n_573), .B1(n_574), .B2(n_578), .Y(n_572) );
INVx3_ASAP7_75t_SL g501 ( .A(n_502), .Y(n_501) );
INVx2_ASAP7_75t_L g615 ( .A(n_502), .Y(n_615) );
INVx4_ASAP7_75t_L g502 ( .A(n_503), .Y(n_502) );
BUFx3_ASAP7_75t_L g707 ( .A(n_503), .Y(n_707) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_506), .A2(n_509), .B(n_510), .Y(n_505) );
OAI22xp5_ASAP7_75t_L g696 ( .A1(n_506), .A2(n_697), .B1(n_698), .B2(n_699), .Y(n_696) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_507), .Y(n_506) );
INVx2_ASAP7_75t_L g606 ( .A(n_507), .Y(n_606) );
OAI221xp5_ASAP7_75t_L g700 ( .A1(n_513), .A2(n_701), .B1(n_702), .B2(n_703), .C(n_704), .Y(n_700) );
INVx1_ASAP7_75t_L g627 ( .A(n_520), .Y(n_627) );
AOI22xp5_ASAP7_75t_SL g520 ( .A1(n_521), .A2(n_598), .B1(n_599), .B2(n_625), .Y(n_520) );
INVx1_ASAP7_75t_L g625 ( .A(n_521), .Y(n_625) );
INVx1_ASAP7_75t_L g521 ( .A(n_522), .Y(n_521) );
AO22x1_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_540), .B1(n_541), .B2(n_597), .Y(n_522) );
INVx2_ASAP7_75t_SL g597 ( .A(n_523), .Y(n_597) );
XOR2x2_ASAP7_75t_L g523 ( .A(n_524), .B(n_539), .Y(n_523) );
NAND4xp75_ASAP7_75t_L g524 ( .A(n_525), .B(n_528), .C(n_533), .D(n_537), .Y(n_524) );
AND2x2_ASAP7_75t_L g525 ( .A(n_526), .B(n_527), .Y(n_525) );
AND2x2_ASAP7_75t_L g528 ( .A(n_529), .B(n_531), .Y(n_528) );
INVx1_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AO22x2_ASAP7_75t_SL g541 ( .A1(n_542), .A2(n_562), .B1(n_595), .B2(n_596), .Y(n_541) );
INVx4_ASAP7_75t_SL g595 ( .A(n_542), .Y(n_595) );
XOR2x2_ASAP7_75t_L g542 ( .A(n_543), .B(n_561), .Y(n_542) );
NAND3x1_ASAP7_75t_L g543 ( .A(n_544), .B(n_553), .C(n_557), .Y(n_543) );
NOR2xp33_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
NAND3xp33_ASAP7_75t_L g548 ( .A(n_549), .B(n_550), .C(n_552), .Y(n_548) );
AND2x2_ASAP7_75t_L g553 ( .A(n_554), .B(n_555), .Y(n_553) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g596 ( .A(n_562), .Y(n_596) );
INVx1_ASAP7_75t_L g593 ( .A(n_563), .Y(n_593) );
AND2x2_ASAP7_75t_L g563 ( .A(n_564), .B(n_579), .Y(n_563) );
NOR3xp33_ASAP7_75t_L g564 ( .A(n_565), .B(n_568), .C(n_572), .Y(n_564) );
OAI22xp5_ASAP7_75t_L g705 ( .A1(n_574), .A2(n_706), .B1(n_707), .B2(n_708), .Y(n_705) );
BUFx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
OAI22xp5_ASAP7_75t_L g613 ( .A1(n_575), .A2(n_614), .B1(n_615), .B2(n_616), .Y(n_613) );
OR2x6_ASAP7_75t_L g575 ( .A(n_576), .B(n_577), .Y(n_575) );
NOR3xp33_ASAP7_75t_L g579 ( .A(n_580), .B(n_583), .C(n_588), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_581), .B(n_582), .Y(n_580) );
INVx1_ASAP7_75t_SL g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
INVx1_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx1_ASAP7_75t_SL g623 ( .A(n_601), .Y(n_623) );
AND2x2_ASAP7_75t_SL g601 ( .A(n_602), .B(n_617), .Y(n_601) );
NOR3xp33_ASAP7_75t_L g602 ( .A(n_603), .B(n_608), .C(n_613), .Y(n_602) );
INVx2_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
OAI21xp33_ASAP7_75t_L g608 ( .A1(n_609), .A2(n_610), .B(n_611), .Y(n_608) );
AND4x1_ASAP7_75t_L g617 ( .A(n_618), .B(n_619), .C(n_621), .D(n_622), .Y(n_617) );
INVx1_ASAP7_75t_SL g628 ( .A(n_629), .Y(n_628) );
NOR2x1_ASAP7_75t_L g629 ( .A(n_630), .B(n_634), .Y(n_629) );
OR2x2_ASAP7_75t_SL g710 ( .A(n_630), .B(n_635), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
HB1xp67_ASAP7_75t_L g673 ( .A(n_632), .Y(n_673) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_632), .B(n_676), .Y(n_679) );
CKINVDCx16_ASAP7_75t_R g676 ( .A(n_633), .Y(n_676) );
CKINVDCx20_ASAP7_75t_R g634 ( .A(n_635), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_636), .B(n_637), .Y(n_635) );
NAND2xp5_ASAP7_75t_L g638 ( .A(n_639), .B(n_640), .Y(n_638) );
OAI322xp33_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_673), .A3(n_674), .B1(n_677), .B2(n_680), .C1(n_681), .C2(n_710), .Y(n_641) );
INVx1_ASAP7_75t_L g671 ( .A(n_643), .Y(n_671) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_644), .B(n_660), .Y(n_643) );
NOR3xp33_ASAP7_75t_L g644 ( .A(n_645), .B(n_652), .C(n_657), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_646), .B(n_650), .Y(n_645) );
INVx2_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OAI22xp5_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_654), .B1(n_655), .B2(n_656), .Y(n_652) );
INVx2_ASAP7_75t_L g686 ( .A(n_654), .Y(n_686) );
NOR2xp33_ASAP7_75t_L g660 ( .A(n_661), .B(n_666), .Y(n_660) );
INVx3_ASAP7_75t_L g664 ( .A(n_665), .Y(n_664) );
NAND3xp33_ASAP7_75t_L g666 ( .A(n_667), .B(n_668), .C(n_670), .Y(n_666) );
HB1xp67_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
CKINVDCx20_ASAP7_75t_R g677 ( .A(n_678), .Y(n_677) );
INVx2_ASAP7_75t_L g709 ( .A(n_682), .Y(n_709) );
AND2x2_ASAP7_75t_SL g682 ( .A(n_683), .B(n_695), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_684), .B(n_691), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_685), .B(n_687), .Y(n_684) );
INVx2_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_692), .B(n_693), .Y(n_691) );
NOR3xp33_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .C(n_705), .Y(n_695) );
endmodule