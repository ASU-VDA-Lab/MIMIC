module fake_jpeg_2684_n_440 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_440);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_440;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx5_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx13_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_15),
.Y(n_24)
);

BUFx10_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_0),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_4),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_10),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_10),
.Y(n_34)
);

INVx13_ASAP7_75t_L g35 ( 
.A(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_11),
.B(n_13),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_5),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_6),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_9),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_1),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_15),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_11),
.Y(n_42)
);

BUFx10_ASAP7_75t_L g43 ( 
.A(n_6),
.Y(n_43)
);

BUFx5_ASAP7_75t_L g44 ( 
.A(n_11),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_10),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_4),
.Y(n_46)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_2),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_9),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_14),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_17),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_13),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_12),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_36),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_54),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g55 ( 
.A(n_39),
.B(n_17),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_55),
.B(n_59),
.Y(n_150)
);

INVx4_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx3_ASAP7_75t_L g135 ( 
.A(n_56),
.Y(n_135)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_22),
.Y(n_57)
);

NAND2xp33_ASAP7_75t_SL g184 ( 
.A(n_57),
.B(n_68),
.Y(n_184)
);

BUFx5_ASAP7_75t_L g58 ( 
.A(n_49),
.Y(n_58)
);

INVx4_ASAP7_75t_L g143 ( 
.A(n_58),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_39),
.B(n_52),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_8),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_60),
.B(n_63),
.Y(n_173)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_26),
.Y(n_61)
);

INVx5_ASAP7_75t_L g132 ( 
.A(n_61),
.Y(n_132)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_48),
.Y(n_62)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_62),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_24),
.B(n_8),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_64),
.Y(n_116)
);

AND2x2_ASAP7_75t_SL g65 ( 
.A(n_26),
.B(n_32),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_65),
.B(n_83),
.C(n_115),
.Y(n_161)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_20),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_46),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_67),
.Y(n_120)
);

CKINVDCx14_ASAP7_75t_R g68 ( 
.A(n_22),
.Y(n_68)
);

INVx1_ASAP7_75t_SL g69 ( 
.A(n_22),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_69),
.B(n_109),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_46),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_70),
.Y(n_174)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g126 ( 
.A(n_71),
.Y(n_126)
);

BUFx4f_ASAP7_75t_SL g72 ( 
.A(n_26),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g124 ( 
.A(n_72),
.Y(n_124)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_73),
.Y(n_129)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_74),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_20),
.Y(n_75)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_75),
.Y(n_147)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_18),
.Y(n_76)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_20),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_77),
.B(n_88),
.Y(n_125)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_27),
.Y(n_78)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_27),
.Y(n_79)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_79),
.Y(n_178)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx8_ASAP7_75t_L g159 ( 
.A(n_80),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_24),
.B(n_16),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g122 ( 
.A(n_81),
.B(n_89),
.Y(n_122)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_28),
.Y(n_82)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_82),
.Y(n_164)
);

CKINVDCx14_ASAP7_75t_R g83 ( 
.A(n_47),
.Y(n_83)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_83),
.Y(n_128)
);

BUFx16f_ASAP7_75t_L g84 ( 
.A(n_35),
.Y(n_84)
);

INVx13_ASAP7_75t_L g190 ( 
.A(n_84),
.Y(n_190)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_85),
.Y(n_133)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_28),
.Y(n_86)
);

BUFx2_ASAP7_75t_L g136 ( 
.A(n_86),
.Y(n_136)
);

BUFx10_ASAP7_75t_L g87 ( 
.A(n_32),
.Y(n_87)
);

BUFx2_ASAP7_75t_L g191 ( 
.A(n_87),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_38),
.B(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_38),
.B(n_16),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_23),
.Y(n_90)
);

INVx5_ASAP7_75t_L g165 ( 
.A(n_90),
.Y(n_165)
);

INVx3_ASAP7_75t_L g91 ( 
.A(n_32),
.Y(n_91)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_91),
.Y(n_162)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_29),
.Y(n_92)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_92),
.Y(n_138)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_32),
.Y(n_93)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_93),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_51),
.B(n_7),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_94),
.B(n_95),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_23),
.Y(n_95)
);

INVx4_ASAP7_75t_L g96 ( 
.A(n_21),
.Y(n_96)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_96),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_33),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_97),
.B(n_105),
.Y(n_172)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_33),
.Y(n_98)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_98),
.Y(n_142)
);

INVx8_ASAP7_75t_L g99 ( 
.A(n_33),
.Y(n_99)
);

INVx3_ASAP7_75t_L g140 ( 
.A(n_99),
.Y(n_140)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_34),
.Y(n_100)
);

INVx4_ASAP7_75t_L g160 ( 
.A(n_100),
.Y(n_160)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_34),
.Y(n_101)
);

BUFx12f_ASAP7_75t_L g186 ( 
.A(n_101),
.Y(n_186)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_34),
.Y(n_102)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_102),
.Y(n_151)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_41),
.Y(n_103)
);

INVx4_ASAP7_75t_L g169 ( 
.A(n_103),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_41),
.Y(n_104)
);

INVx3_ASAP7_75t_L g145 ( 
.A(n_104),
.Y(n_145)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_41),
.Y(n_105)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

INVx4_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

HB1xp67_ASAP7_75t_L g181 ( 
.A(n_107),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g108 ( 
.A(n_42),
.B(n_45),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_108),
.B(n_112),
.Y(n_176)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_45),
.Y(n_109)
);

INVx3_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

INVx3_ASAP7_75t_L g185 ( 
.A(n_110),
.Y(n_185)
);

INVx11_ASAP7_75t_SL g111 ( 
.A(n_47),
.Y(n_111)
);

CKINVDCx14_ASAP7_75t_R g158 ( 
.A(n_111),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_51),
.B(n_7),
.Y(n_112)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_35),
.Y(n_113)
);

INVx4_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_47),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_114),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_25),
.Y(n_115)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_115),
.B(n_57),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_56),
.A2(n_53),
.B1(n_52),
.B2(n_37),
.Y(n_117)
);

OAI21xp5_ASAP7_75t_SL g211 ( 
.A1(n_117),
.A2(n_184),
.B(n_134),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g119 ( 
.A1(n_108),
.A2(n_53),
.B1(n_19),
.B2(n_50),
.Y(n_119)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_119),
.A2(n_123),
.B1(n_130),
.B2(n_149),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_19),
.B1(n_31),
.B2(n_40),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_96),
.A2(n_50),
.B1(n_31),
.B2(n_40),
.Y(n_127)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_127),
.A2(n_134),
.B1(n_137),
.B2(n_148),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_65),
.A2(n_43),
.B1(n_25),
.B2(n_44),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_57),
.A2(n_35),
.B1(n_44),
.B2(n_30),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_69),
.A2(n_30),
.B1(n_25),
.B2(n_43),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_68),
.B(n_12),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_139),
.B(n_182),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_64),
.A2(n_67),
.B1(n_70),
.B2(n_104),
.Y(n_144)
);

OAI22xp33_ASAP7_75t_L g215 ( 
.A1(n_144),
.A2(n_166),
.B1(n_179),
.B2(n_163),
.Y(n_215)
);

AOI22xp33_ASAP7_75t_SL g148 ( 
.A1(n_71),
.A2(n_25),
.B1(n_43),
.B2(n_3),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g149 ( 
.A1(n_75),
.A2(n_43),
.B1(n_25),
.B2(n_9),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_82),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g237 ( 
.A1(n_152),
.A2(n_153),
.B1(n_156),
.B2(n_157),
.Y(n_237)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_82),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_153)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_80),
.A2(n_13),
.B1(n_14),
.B2(n_16),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_L g217 ( 
.A1(n_154),
.A2(n_177),
.B1(n_124),
.B2(n_143),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_84),
.A2(n_0),
.B1(n_4),
.B2(n_5),
.Y(n_156)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_111),
.B1(n_61),
.B2(n_103),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_161),
.B(n_156),
.Y(n_236)
);

AOI22xp33_ASAP7_75t_SL g163 ( 
.A1(n_103),
.A2(n_100),
.B1(n_99),
.B2(n_106),
.Y(n_163)
);

AOI22xp33_ASAP7_75t_SL g250 ( 
.A1(n_163),
.A2(n_175),
.B1(n_179),
.B2(n_157),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_90),
.A2(n_101),
.B1(n_72),
.B2(n_86),
.Y(n_166)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_87),
.A2(n_49),
.B1(n_96),
.B2(n_56),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_87),
.A2(n_108),
.B1(n_60),
.B2(n_48),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_56),
.A2(n_49),
.B1(n_96),
.B2(n_28),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_54),
.B(n_59),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_54),
.B(n_59),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_SL g246 ( 
.A(n_183),
.B(n_187),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_54),
.B(n_59),
.Y(n_187)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_189),
.Y(n_233)
);

INVx13_ASAP7_75t_L g192 ( 
.A(n_190),
.Y(n_192)
);

INVx13_ASAP7_75t_L g287 ( 
.A(n_192),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_150),
.B(n_173),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_SL g298 ( 
.A(n_194),
.B(n_199),
.Y(n_298)
);

INVx3_ASAP7_75t_L g195 ( 
.A(n_132),
.Y(n_195)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_195),
.Y(n_259)
);

INVx8_ASAP7_75t_L g196 ( 
.A(n_186),
.Y(n_196)
);

INVx3_ASAP7_75t_L g268 ( 
.A(n_196),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g197 ( 
.A(n_158),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g255 ( 
.A(n_197),
.B(n_200),
.Y(n_255)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_129),
.Y(n_198)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_198),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_118),
.B(n_138),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_122),
.B(n_125),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_172),
.Y(n_201)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_201),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_128),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_202),
.B(n_204),
.Y(n_257)
);

INVx3_ASAP7_75t_L g203 ( 
.A(n_132),
.Y(n_203)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_203),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_171),
.B(n_176),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g205 ( 
.A(n_116),
.Y(n_205)
);

INVx6_ASAP7_75t_L g258 ( 
.A(n_205),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_141),
.B(n_133),
.Y(n_206)
);

OAI21x1_ASAP7_75t_L g276 ( 
.A1(n_206),
.A2(n_211),
.B(n_225),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g207 ( 
.A(n_181),
.Y(n_207)
);

HB1xp67_ASAP7_75t_L g286 ( 
.A(n_207),
.Y(n_286)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_142),
.Y(n_208)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_208),
.Y(n_280)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_151),
.Y(n_209)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_209),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_155),
.B(n_162),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_210),
.B(n_226),
.Y(n_263)
);

INVx3_ASAP7_75t_L g212 ( 
.A(n_140),
.Y(n_212)
);

INVx3_ASAP7_75t_L g297 ( 
.A(n_212),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_185),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g264 ( 
.A(n_213),
.Y(n_264)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_121),
.Y(n_214)
);

INVx2_ASAP7_75t_L g278 ( 
.A(n_214),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_215),
.B(n_238),
.Y(n_284)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_131),
.B(n_167),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_216),
.B(n_236),
.C(n_241),
.Y(n_292)
);

OA22x2_ASAP7_75t_L g285 ( 
.A1(n_217),
.A2(n_234),
.B1(n_195),
.B2(n_203),
.Y(n_285)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_178),
.Y(n_219)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_219),
.Y(n_256)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_145),
.Y(n_220)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_220),
.Y(n_299)
);

INVx13_ASAP7_75t_L g221 ( 
.A(n_190),
.Y(n_221)
);

INVx13_ASAP7_75t_L g300 ( 
.A(n_221),
.Y(n_300)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_116),
.Y(n_222)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_222),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g223 ( 
.A(n_191),
.Y(n_223)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_223),
.Y(n_273)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_146),
.Y(n_224)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_224),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_180),
.B(n_146),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_135),
.B(n_168),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_127),
.B(n_189),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_227),
.B(n_228),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_145),
.B(n_188),
.Y(n_228)
);

BUFx6f_ASAP7_75t_L g229 ( 
.A(n_120),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_229),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_188),
.B(n_191),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_232),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_169),
.B(n_126),
.Y(n_232)
);

AOI22xp33_ASAP7_75t_L g234 ( 
.A1(n_144),
.A2(n_166),
.B1(n_136),
.B2(n_170),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_137),
.A2(n_175),
.B(n_152),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_235),
.A2(n_248),
.B(n_251),
.Y(n_295)
);

INVx3_ASAP7_75t_L g238 ( 
.A(n_140),
.Y(n_238)
);

INVx2_ASAP7_75t_L g239 ( 
.A(n_147),
.Y(n_239)
);

AND2x2_ASAP7_75t_L g290 ( 
.A(n_239),
.B(n_243),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_169),
.B(n_126),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_240),
.B(n_242),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_136),
.B(n_148),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_170),
.B(n_165),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_160),
.Y(n_243)
);

BUFx12f_ASAP7_75t_L g244 ( 
.A(n_159),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g267 ( 
.A(n_244),
.Y(n_267)
);

INVx2_ASAP7_75t_L g245 ( 
.A(n_147),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g262 ( 
.A1(n_245),
.A2(n_247),
.B1(n_248),
.B2(n_250),
.Y(n_262)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_160),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_186),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_143),
.B(n_165),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_251),
.Y(n_269)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_164),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_252),
.B(n_254),
.Y(n_272)
);

INVx4_ASAP7_75t_L g253 ( 
.A(n_159),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_253),
.B(n_244),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g254 ( 
.A(n_120),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g261 ( 
.A1(n_218),
.A2(n_153),
.B1(n_174),
.B2(n_164),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g326 ( 
.A1(n_261),
.A2(n_281),
.B1(n_294),
.B2(n_289),
.Y(n_326)
);

AND2x4_ASAP7_75t_L g271 ( 
.A(n_235),
.B(n_164),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g322 ( 
.A(n_271),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_218),
.A2(n_174),
.B1(n_215),
.B2(n_241),
.Y(n_274)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_274),
.A2(n_284),
.B1(n_295),
.B2(n_265),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g281 ( 
.A1(n_193),
.A2(n_237),
.B1(n_250),
.B2(n_236),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_SL g282 ( 
.A1(n_193),
.A2(n_233),
.B(n_237),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g334 ( 
.A1(n_282),
.A2(n_283),
.B(n_295),
.Y(n_334)
);

OAI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_233),
.A2(n_216),
.B(n_212),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g310 ( 
.A(n_285),
.B(n_284),
.Y(n_310)
);

AOI32xp33_ASAP7_75t_L g291 ( 
.A1(n_230),
.A2(n_239),
.A3(n_245),
.B1(n_220),
.B2(n_253),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_291),
.B(n_271),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_238),
.A2(n_229),
.B1(n_254),
.B2(n_205),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_222),
.B(n_244),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_296),
.B(n_223),
.Y(n_304)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_301),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_290),
.Y(n_302)
);

NOR3xp33_ASAP7_75t_L g362 ( 
.A(n_302),
.B(n_303),
.C(n_309),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_255),
.B(n_246),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g341 ( 
.A(n_304),
.B(n_305),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_SL g305 ( 
.A(n_283),
.B(n_192),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_292),
.B(n_221),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_306),
.B(n_307),
.Y(n_346)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_257),
.B(n_298),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_196),
.C(n_281),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_308),
.B(n_314),
.Y(n_348)
);

CKINVDCx20_ASAP7_75t_R g309 ( 
.A(n_290),
.Y(n_309)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_310),
.B(n_324),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_311),
.A2(n_336),
.B1(n_285),
.B2(n_297),
.Y(n_337)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_263),
.B(n_270),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g340 ( 
.A(n_312),
.B(n_315),
.Y(n_340)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_266),
.Y(n_313)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_313),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g314 ( 
.A(n_275),
.B(n_276),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_L g315 ( 
.A(n_288),
.B(n_279),
.Y(n_315)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_259),
.Y(n_316)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_316),
.Y(n_342)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_290),
.Y(n_318)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_318),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_274),
.B(n_269),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_319),
.B(n_320),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_SL g320 ( 
.A(n_269),
.B(n_288),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_282),
.B(n_271),
.C(n_293),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_321),
.B(n_323),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_272),
.B(n_301),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g325 ( 
.A1(n_271),
.A2(n_284),
.B(n_262),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_325),
.A2(n_331),
.B(n_332),
.Y(n_353)
);

OAI22xp5_ASAP7_75t_L g344 ( 
.A1(n_326),
.A2(n_328),
.B1(n_299),
.B2(n_278),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_272),
.B(n_296),
.Y(n_327)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_261),
.A2(n_285),
.B1(n_294),
.B2(n_266),
.Y(n_328)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_286),
.B(n_280),
.Y(n_329)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_329),
.Y(n_354)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_256),
.Y(n_330)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_330),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_L g331 ( 
.A1(n_256),
.A2(n_267),
.B(n_260),
.Y(n_331)
);

AOI21xp5_ASAP7_75t_L g332 ( 
.A1(n_287),
.A2(n_300),
.B(n_297),
.Y(n_332)
);

CKINVDCx14_ASAP7_75t_R g333 ( 
.A(n_287),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g352 ( 
.A(n_333),
.Y(n_352)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_299),
.Y(n_335)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_335),
.Y(n_359)
);

OAI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_285),
.A2(n_258),
.B1(n_259),
.B2(n_277),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g380 ( 
.A1(n_337),
.A2(n_344),
.B1(n_357),
.B2(n_360),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g343 ( 
.A1(n_319),
.A2(n_277),
.B1(n_264),
.B2(n_268),
.Y(n_343)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_343),
.A2(n_345),
.B1(n_358),
.B2(n_302),
.Y(n_372)
);

AOI22xp5_ASAP7_75t_L g345 ( 
.A1(n_311),
.A2(n_268),
.B1(n_278),
.B2(n_273),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g355 ( 
.A(n_329),
.Y(n_355)
);

NOR3xp33_ASAP7_75t_L g379 ( 
.A(n_355),
.B(n_314),
.C(n_305),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_328),
.A2(n_258),
.B1(n_273),
.B2(n_300),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_326),
.A2(n_310),
.B1(n_317),
.B2(n_327),
.Y(n_358)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_312),
.A2(n_310),
.B1(n_317),
.B2(n_320),
.Y(n_360)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_330),
.Y(n_361)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_361),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_L g363 ( 
.A1(n_334),
.A2(n_322),
.B(n_325),
.Y(n_363)
);

INVxp67_ASAP7_75t_L g365 ( 
.A(n_363),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g364 ( 
.A(n_352),
.B(n_303),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_364),
.B(n_366),
.Y(n_395)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_356),
.B(n_315),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_338),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_368),
.B(n_372),
.Y(n_389)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_347),
.B(n_323),
.Y(n_369)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_369),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_308),
.C(n_306),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_382),
.C(n_350),
.Y(n_386)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_349),
.Y(n_371)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_371),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_356),
.B(n_304),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_373),
.B(n_375),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_347),
.B(n_309),
.Y(n_374)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_374),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_354),
.B(n_339),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_349),
.Y(n_376)
);

CKINVDCx16_ASAP7_75t_R g392 ( 
.A(n_376),
.Y(n_392)
);

NOR2xp33_ASAP7_75t_L g377 ( 
.A(n_340),
.B(n_307),
.Y(n_377)
);

XOR2xp5_ASAP7_75t_L g390 ( 
.A(n_377),
.B(n_381),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_338),
.Y(n_378)
);

INVx4_ASAP7_75t_L g387 ( 
.A(n_378),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_379),
.A2(n_351),
.B1(n_346),
.B2(n_322),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_362),
.B(n_331),
.Y(n_381)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_348),
.B(n_321),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g394 ( 
.A(n_382),
.B(n_384),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g383 ( 
.A(n_341),
.Y(n_383)
);

OAI22xp5_ASAP7_75t_L g388 ( 
.A1(n_383),
.A2(n_341),
.B1(n_346),
.B2(n_345),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g384 ( 
.A(n_358),
.B(n_318),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g407 ( 
.A1(n_385),
.A2(n_381),
.B(n_375),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g409 ( 
.A(n_386),
.B(n_391),
.C(n_398),
.Y(n_409)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_388),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_370),
.B(n_351),
.C(n_373),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g393 ( 
.A1(n_380),
.A2(n_337),
.B1(n_353),
.B2(n_351),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_374),
.B(n_363),
.C(n_334),
.Y(n_398)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_387),
.Y(n_402)
);

NOR2xp33_ASAP7_75t_L g413 ( 
.A(n_402),
.B(n_403),
.Y(n_413)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_400),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_399),
.B(n_378),
.Y(n_404)
);

XNOR2xp5_ASAP7_75t_L g415 ( 
.A(n_404),
.B(n_405),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_399),
.B(n_368),
.Y(n_405)
);

OAI21xp5_ASAP7_75t_L g406 ( 
.A1(n_389),
.A2(n_365),
.B(n_383),
.Y(n_406)
);

AOI21xp5_ASAP7_75t_L g420 ( 
.A1(n_406),
.A2(n_407),
.B(n_404),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_369),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_386),
.B(n_366),
.C(n_380),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g417 ( 
.A(n_410),
.B(n_391),
.C(n_394),
.Y(n_417)
);

BUFx12_ASAP7_75t_L g411 ( 
.A(n_392),
.Y(n_411)
);

OAI21xp5_ASAP7_75t_SL g416 ( 
.A1(n_411),
.A2(n_412),
.B(n_385),
.Y(n_416)
);

AOI322xp5_ASAP7_75t_L g412 ( 
.A1(n_389),
.A2(n_377),
.A3(n_364),
.B1(n_376),
.B2(n_371),
.C1(n_367),
.C2(n_359),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_L g414 ( 
.A1(n_401),
.A2(n_393),
.B1(n_390),
.B2(n_396),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_418),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g421 ( 
.A(n_416),
.B(n_407),
.Y(n_421)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_417),
.B(n_409),
.C(n_410),
.Y(n_425)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_401),
.A2(n_390),
.B1(n_396),
.B2(n_395),
.Y(n_418)
);

MAJIxp5_ASAP7_75t_L g419 ( 
.A(n_409),
.B(n_394),
.C(n_342),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_L g424 ( 
.A(n_419),
.B(n_420),
.Y(n_424)
);

NAND2xp5_ASAP7_75t_L g427 ( 
.A(n_421),
.B(n_422),
.Y(n_427)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_418),
.B(n_395),
.Y(n_422)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_425),
.B(n_417),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_420),
.B(n_408),
.Y(n_426)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g432 ( 
.A1(n_429),
.A2(n_430),
.B(n_424),
.Y(n_432)
);

OAI21xp5_ASAP7_75t_SL g430 ( 
.A1(n_421),
.A2(n_414),
.B(n_406),
.Y(n_430)
);

CKINVDCx20_ASAP7_75t_R g431 ( 
.A(n_423),
.Y(n_431)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_431),
.Y(n_433)
);

AOI21xp5_ASAP7_75t_L g436 ( 
.A1(n_432),
.A2(n_427),
.B(n_430),
.Y(n_436)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_428),
.Y(n_434)
);

AOI322xp5_ASAP7_75t_L g435 ( 
.A1(n_434),
.A2(n_411),
.A3(n_413),
.B1(n_405),
.B2(n_403),
.C1(n_397),
.C2(n_367),
.Y(n_435)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_435),
.Y(n_437)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_437),
.Y(n_438)
);

OAI221xp5_ASAP7_75t_L g439 ( 
.A1(n_438),
.A2(n_436),
.B1(n_433),
.B2(n_412),
.C(n_397),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_439),
.B(n_415),
.Y(n_440)
);


endmodule