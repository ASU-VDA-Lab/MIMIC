module fake_jpeg_17104_n_240 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_240);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_240;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

INVx11_ASAP7_75t_L g17 ( 
.A(n_14),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_12),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_9),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_10),
.Y(n_24)
);

INVx4_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_2),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_2),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_7),
.B(n_12),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_9),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_8),
.Y(n_36)
);

BUFx10_ASAP7_75t_L g37 ( 
.A(n_5),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_0),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_38),
.B(n_50),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_22),
.Y(n_39)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_39),
.Y(n_106)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_22),
.Y(n_40)
);

INVx5_ASAP7_75t_L g82 ( 
.A(n_40),
.Y(n_82)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_17),
.Y(n_41)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_41),
.Y(n_74)
);

INVx5_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_28),
.B(n_0),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_43),
.B(n_48),
.Y(n_87)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_22),
.Y(n_45)
);

BUFx12f_ASAP7_75t_L g78 ( 
.A(n_45),
.Y(n_78)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_34),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_46),
.B(n_52),
.Y(n_94)
);

INVx11_ASAP7_75t_L g47 ( 
.A(n_15),
.Y(n_47)
);

INVx6_ASAP7_75t_L g67 ( 
.A(n_47),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g48 ( 
.A(n_18),
.B(n_1),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_49),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_21),
.B(n_1),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_31),
.Y(n_51)
);

BUFx4f_ASAP7_75t_SL g92 ( 
.A(n_51),
.Y(n_92)
);

INVx3_ASAP7_75t_SL g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g53 ( 
.A(n_32),
.Y(n_53)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_53),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_18),
.B(n_1),
.Y(n_54)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_54),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_19),
.B(n_3),
.Y(n_55)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_55),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_32),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_56),
.Y(n_86)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_16),
.Y(n_57)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_57),
.Y(n_90)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_37),
.Y(n_58)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_59),
.B(n_60),
.Y(n_97)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g61 ( 
.A(n_21),
.B(n_4),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_61),
.B(n_50),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_19),
.B(n_4),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_62),
.B(n_63),
.Y(n_100)
);

BUFx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_64),
.B(n_5),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_34),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g95 ( 
.A(n_65),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_25),
.B1(n_15),
.B2(n_17),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_L g137 ( 
.A1(n_66),
.A2(n_68),
.B1(n_75),
.B2(n_80),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_44),
.A2(n_25),
.B1(n_23),
.B2(n_26),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_58),
.B(n_20),
.C(n_15),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g138 ( 
.A(n_70),
.B(n_88),
.C(n_103),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_72),
.B(n_79),
.Y(n_118)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_57),
.A2(n_29),
.B1(n_36),
.B2(n_35),
.Y(n_75)
);

CKINVDCx14_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_76),
.B(n_81),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_L g77 ( 
.A1(n_41),
.A2(n_15),
.B(n_23),
.C(n_30),
.Y(n_77)
);

OAI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_77),
.A2(n_85),
.B1(n_53),
.B2(n_74),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_39),
.B(n_24),
.Y(n_79)
);

OAI22xp33_ASAP7_75t_L g80 ( 
.A1(n_52),
.A2(n_37),
.B1(n_30),
.B2(n_26),
.Y(n_80)
);

CKINVDCx5p33_ASAP7_75t_R g81 ( 
.A(n_47),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_42),
.A2(n_36),
.B1(n_35),
.B2(n_29),
.Y(n_85)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_64),
.B(n_20),
.C(n_37),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_46),
.A2(n_27),
.B1(n_24),
.B2(n_7),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g120 ( 
.A1(n_93),
.A2(n_96),
.B1(n_56),
.B2(n_49),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_60),
.A2(n_27),
.B1(n_5),
.B2(n_8),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_65),
.B(n_4),
.Y(n_98)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_98),
.B(n_13),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_45),
.B(n_20),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_99),
.B(n_102),
.Y(n_111)
);

OR2x2_ASAP7_75t_L g102 ( 
.A(n_63),
.B(n_33),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_40),
.B(n_20),
.C(n_33),
.Y(n_103)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_104),
.Y(n_115)
);

XOR2xp5_ASAP7_75t_L g105 ( 
.A(n_40),
.B(n_8),
.Y(n_105)
);

XOR2xp5_ASAP7_75t_L g113 ( 
.A(n_105),
.B(n_9),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_105),
.B(n_90),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_107),
.B(n_126),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_73),
.B(n_13),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g139 ( 
.A(n_108),
.B(n_122),
.Y(n_139)
);

BUFx2_ASAP7_75t_L g110 ( 
.A(n_78),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_110),
.B(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_69),
.Y(n_112)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_112),
.Y(n_140)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_113),
.B(n_123),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_91),
.B(n_10),
.Y(n_114)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_114),
.Y(n_154)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_106),
.Y(n_116)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_116),
.Y(n_156)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_77),
.Y(n_117)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_117),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_89),
.B(n_11),
.Y(n_119)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_119),
.Y(n_160)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_120),
.A2(n_71),
.B1(n_82),
.B2(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_94),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_92),
.Y(n_122)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_97),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_124),
.B(n_129),
.Y(n_146)
);

INVxp67_ASAP7_75t_L g125 ( 
.A(n_93),
.Y(n_125)
);

OAI32xp33_ASAP7_75t_L g126 ( 
.A1(n_100),
.A2(n_51),
.A3(n_53),
.B1(n_102),
.B2(n_96),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g127 ( 
.A(n_80),
.B(n_51),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_127),
.B(n_130),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g151 ( 
.A(n_128),
.Y(n_151)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_84),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_87),
.B(n_81),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_87),
.B(n_74),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_131),
.B(n_132),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_84),
.B(n_86),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_78),
.Y(n_133)
);

INVx2_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_86),
.B(n_66),
.Y(n_134)
);

INVxp33_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_67),
.B(n_101),
.Y(n_135)
);

INVxp33_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_78),
.B(n_98),
.Y(n_136)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_136),
.B(n_107),
.C(n_113),
.Y(n_143)
);

AND2x2_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_136),
.Y(n_171)
);

INVx13_ASAP7_75t_L g145 ( 
.A(n_110),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_145),
.B(n_149),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_117),
.A2(n_71),
.B1(n_82),
.B2(n_67),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_148),
.A2(n_153),
.B1(n_129),
.B2(n_122),
.Y(n_166)
);

INVxp33_ASAP7_75t_L g149 ( 
.A(n_132),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_138),
.B(n_92),
.C(n_83),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_150),
.B(n_161),
.C(n_121),
.Y(n_182)
);

INVxp33_ASAP7_75t_L g152 ( 
.A(n_135),
.Y(n_152)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_152),
.Y(n_170)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_138),
.B(n_83),
.C(n_95),
.Y(n_161)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_164),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_142),
.A2(n_137),
.B1(n_134),
.B2(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g196 ( 
.A1(n_165),
.A2(n_169),
.B1(n_158),
.B2(n_160),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_166),
.A2(n_157),
.B1(n_158),
.B2(n_109),
.Y(n_195)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_162),
.Y(n_167)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_167),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_143),
.B(n_111),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_168),
.B(n_179),
.C(n_182),
.Y(n_186)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_142),
.A2(n_111),
.B1(n_127),
.B2(n_126),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_171),
.B(n_123),
.Y(n_197)
);

OR2x6_ASAP7_75t_L g172 ( 
.A(n_141),
.B(n_127),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g193 ( 
.A1(n_172),
.A2(n_184),
.B(n_147),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_163),
.B(n_118),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_174),
.B(n_181),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g198 ( 
.A(n_176),
.B(n_178),
.Y(n_198)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_156),
.Y(n_177)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_159),
.B(n_130),
.Y(n_179)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_162),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_180),
.B(n_183),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_163),
.B(n_118),
.Y(n_181)
);

BUFx24_ASAP7_75t_SL g183 ( 
.A(n_154),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_151),
.A2(n_115),
.B1(n_124),
.B2(n_123),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_150),
.C(n_161),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_187),
.B(n_188),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_168),
.B(n_179),
.C(n_159),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_169),
.B(n_155),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_194),
.Y(n_201)
);

NOR3xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_147),
.C(n_109),
.Y(n_191)
);

NOR3xp33_ASAP7_75t_L g203 ( 
.A(n_191),
.B(n_172),
.C(n_160),
.Y(n_203)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_193),
.A2(n_172),
.B(n_171),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_155),
.Y(n_194)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_195),
.A2(n_189),
.B1(n_194),
.B2(n_193),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_196),
.B(n_172),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_199),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_170),
.B(n_140),
.Y(n_199)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_198),
.Y(n_202)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_202),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_203),
.B(n_210),
.Y(n_217)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_199),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_204),
.B(n_148),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g220 ( 
.A1(n_205),
.A2(n_211),
.B(n_119),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_206),
.B(n_208),
.Y(n_214)
);

OAI322xp33_ASAP7_75t_L g209 ( 
.A1(n_190),
.A2(n_154),
.A3(n_184),
.B1(n_144),
.B2(n_139),
.C1(n_146),
.C2(n_114),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_209),
.B(n_197),
.C(n_196),
.Y(n_213)
);

NOR3xp33_ASAP7_75t_L g210 ( 
.A(n_200),
.B(n_139),
.C(n_173),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_188),
.A2(n_146),
.B(n_112),
.Y(n_211)
);

FAx1_ASAP7_75t_SL g227 ( 
.A(n_213),
.B(n_110),
.CI(n_145),
.CON(n_227),
.SN(n_227)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_186),
.C(n_187),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g222 ( 
.A(n_215),
.B(n_207),
.C(n_205),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_220),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_204),
.B(n_192),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_218),
.B(n_116),
.Y(n_228)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_212),
.A2(n_186),
.B1(n_167),
.B2(n_175),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_221),
.B(n_185),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g232 ( 
.A(n_222),
.B(n_223),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_215),
.B(n_211),
.C(n_201),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_224),
.B(n_226),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_219),
.B(n_164),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_227),
.B(n_213),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g230 ( 
.A(n_228),
.B(n_217),
.Y(n_230)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_230),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_231),
.A2(n_233),
.B(n_214),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_225),
.B(n_221),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g239 ( 
.A1(n_235),
.A2(n_234),
.B(n_236),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_232),
.A2(n_222),
.B1(n_223),
.B2(n_227),
.Y(n_236)
);

OAI21x1_ASAP7_75t_SL g238 ( 
.A1(n_236),
.A2(n_237),
.B(n_229),
.Y(n_238)
);

OAI22xp5_ASAP7_75t_L g237 ( 
.A1(n_230),
.A2(n_145),
.B1(n_133),
.B2(n_95),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_238),
.B(n_239),
.Y(n_240)
);


endmodule