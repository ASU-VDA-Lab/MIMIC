module fake_netlist_1_12541_n_754 (n_44, n_81, n_69, n_22, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_97, n_80, n_107, n_60, n_41, n_35, n_94, n_65, n_9, n_10, n_103, n_19, n_87, n_104, n_98, n_74, n_7, n_29, n_45, n_85, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_16, n_13, n_95, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_84, n_55, n_12, n_86, n_75, n_105, n_72, n_43, n_76, n_89, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_83, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_3, n_18, n_110, n_66, n_1, n_82, n_106, n_15, n_61, n_21, n_99, n_109, n_93, n_51, n_96, n_39, n_754);
input n_44;
input n_81;
input n_69;
input n_22;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_97;
input n_80;
input n_107;
input n_60;
input n_41;
input n_35;
input n_94;
input n_65;
input n_9;
input n_10;
input n_103;
input n_19;
input n_87;
input n_104;
input n_98;
input n_74;
input n_7;
input n_29;
input n_45;
input n_85;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_16;
input n_13;
input n_95;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_84;
input n_55;
input n_12;
input n_86;
input n_75;
input n_105;
input n_72;
input n_43;
input n_76;
input n_89;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_83;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_110;
input n_66;
input n_1;
input n_82;
input n_106;
input n_15;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_51;
input n_96;
input n_39;
output n_754;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_732;
wire n_752;
wire n_199;
wire n_351;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_724;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_623;
wire n_167;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_711;
wire n_238;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_533;
wire n_506;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_746;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_751;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_450;
wire n_579;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_649;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_621;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_409;
wire n_363;
wire n_733;
wire n_295;
wire n_143;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_749;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_449;
wire n_115;
wire n_300;
wire n_158;
wire n_734;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_180;
wire n_441;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_146;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_736;
wire n_194;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_739;
wire n_145;
wire n_740;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_2), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_19), .Y(n_112) );
CKINVDCx5p33_ASAP7_75t_R g113 ( .A(n_29), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_79), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_52), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_81), .Y(n_116) );
CKINVDCx20_ASAP7_75t_R g117 ( .A(n_25), .Y(n_117) );
BUFx3_ASAP7_75t_L g118 ( .A(n_3), .Y(n_118) );
CKINVDCx5p33_ASAP7_75t_R g119 ( .A(n_73), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_40), .Y(n_120) );
CKINVDCx16_ASAP7_75t_R g121 ( .A(n_103), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_82), .Y(n_122) );
BUFx3_ASAP7_75t_L g123 ( .A(n_45), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_49), .Y(n_124) );
HB1xp67_ASAP7_75t_L g125 ( .A(n_14), .Y(n_125) );
NOR2xp67_ASAP7_75t_L g126 ( .A(n_15), .B(n_110), .Y(n_126) );
BUFx2_ASAP7_75t_L g127 ( .A(n_62), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_70), .Y(n_128) );
CKINVDCx5p33_ASAP7_75t_R g129 ( .A(n_23), .Y(n_129) );
INVx1_ASAP7_75t_L g130 ( .A(n_89), .Y(n_130) );
CKINVDCx5p33_ASAP7_75t_R g131 ( .A(n_18), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_63), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_59), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_27), .Y(n_134) );
INVxp33_ASAP7_75t_SL g135 ( .A(n_24), .Y(n_135) );
INVx1_ASAP7_75t_L g136 ( .A(n_22), .Y(n_136) );
INVx2_ASAP7_75t_L g137 ( .A(n_101), .Y(n_137) );
CKINVDCx5p33_ASAP7_75t_R g138 ( .A(n_75), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_92), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_7), .Y(n_140) );
INVx1_ASAP7_75t_L g141 ( .A(n_71), .Y(n_141) );
BUFx10_ASAP7_75t_L g142 ( .A(n_32), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_56), .Y(n_143) );
BUFx5_ASAP7_75t_L g144 ( .A(n_42), .Y(n_144) );
INVx1_ASAP7_75t_L g145 ( .A(n_11), .Y(n_145) );
INVx1_ASAP7_75t_L g146 ( .A(n_48), .Y(n_146) );
BUFx3_ASAP7_75t_L g147 ( .A(n_87), .Y(n_147) );
HB1xp67_ASAP7_75t_L g148 ( .A(n_44), .Y(n_148) );
CKINVDCx5p33_ASAP7_75t_R g149 ( .A(n_6), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g150 ( .A(n_105), .Y(n_150) );
INVx1_ASAP7_75t_L g151 ( .A(n_38), .Y(n_151) );
NOR2xp67_ASAP7_75t_L g152 ( .A(n_88), .B(n_7), .Y(n_152) );
CKINVDCx5p33_ASAP7_75t_R g153 ( .A(n_69), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_34), .Y(n_154) );
CKINVDCx5p33_ASAP7_75t_R g155 ( .A(n_43), .Y(n_155) );
CKINVDCx5p33_ASAP7_75t_R g156 ( .A(n_57), .Y(n_156) );
INVx1_ASAP7_75t_L g157 ( .A(n_68), .Y(n_157) );
NAND2xp5_ASAP7_75t_L g158 ( .A(n_125), .B(n_0), .Y(n_158) );
CKINVDCx5p33_ASAP7_75t_R g159 ( .A(n_121), .Y(n_159) );
NAND2xp5_ASAP7_75t_SL g160 ( .A(n_127), .B(n_0), .Y(n_160) );
BUFx8_ASAP7_75t_L g161 ( .A(n_144), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g162 ( .A1(n_135), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_162) );
OA21x2_ASAP7_75t_L g163 ( .A1(n_137), .A2(n_58), .B(n_108), .Y(n_163) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_148), .B(n_1), .Y(n_164) );
INVx2_ASAP7_75t_L g165 ( .A(n_144), .Y(n_165) );
INVx2_ASAP7_75t_L g166 ( .A(n_144), .Y(n_166) );
INVx2_ASAP7_75t_SL g167 ( .A(n_142), .Y(n_167) );
BUFx2_ASAP7_75t_L g168 ( .A(n_118), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_118), .Y(n_169) );
INVx2_ASAP7_75t_L g170 ( .A(n_144), .Y(n_170) );
BUFx6f_ASAP7_75t_L g171 ( .A(n_123), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_140), .B(n_4), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_123), .Y(n_174) );
INVx2_ASAP7_75t_L g175 ( .A(n_144), .Y(n_175) );
NAND2xp5_ASAP7_75t_L g176 ( .A(n_145), .B(n_4), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_135), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_177) );
INVx2_ASAP7_75t_SL g178 ( .A(n_161), .Y(n_178) );
INVx2_ASAP7_75t_L g179 ( .A(n_165), .Y(n_179) );
INVx2_ASAP7_75t_L g180 ( .A(n_165), .Y(n_180) );
INVx3_ASAP7_75t_L g181 ( .A(n_166), .Y(n_181) );
NAND2xp5_ASAP7_75t_SL g182 ( .A(n_167), .B(n_142), .Y(n_182) );
OAI22xp33_ASAP7_75t_SL g183 ( .A1(n_162), .A2(n_153), .B1(n_156), .B2(n_155), .Y(n_183) );
INVx3_ASAP7_75t_L g184 ( .A(n_166), .Y(n_184) );
BUFx6f_ASAP7_75t_L g185 ( .A(n_163), .Y(n_185) );
NOR2xp67_ASAP7_75t_L g186 ( .A(n_169), .B(n_119), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_170), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_170), .Y(n_188) );
NAND2xp33_ASAP7_75t_L g189 ( .A(n_167), .B(n_144), .Y(n_189) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_168), .B(n_112), .Y(n_190) );
AOI21x1_ASAP7_75t_L g191 ( .A1(n_172), .A2(n_137), .B(n_139), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_168), .B(n_112), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_172), .Y(n_193) );
NAND3xp33_ASAP7_75t_L g194 ( .A(n_161), .B(n_111), .C(n_149), .Y(n_194) );
INVx3_ASAP7_75t_L g195 ( .A(n_175), .Y(n_195) );
INVx1_ASAP7_75t_L g196 ( .A(n_175), .Y(n_196) );
INVx2_ASAP7_75t_L g197 ( .A(n_171), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_169), .B(n_113), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_171), .Y(n_199) );
NOR2xp33_ASAP7_75t_L g200 ( .A(n_159), .B(n_115), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_171), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_161), .B(n_113), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g203 ( .A(n_159), .B(n_114), .Y(n_203) );
INVx2_ASAP7_75t_L g204 ( .A(n_171), .Y(n_204) );
INVx2_ASAP7_75t_SL g205 ( .A(n_171), .Y(n_205) );
NAND2xp5_ASAP7_75t_L g206 ( .A(n_190), .B(n_164), .Y(n_206) );
INVx2_ASAP7_75t_SL g207 ( .A(n_178), .Y(n_207) );
INVx2_ASAP7_75t_L g208 ( .A(n_191), .Y(n_208) );
NOR2xp33_ASAP7_75t_L g209 ( .A(n_182), .B(n_203), .Y(n_209) );
INVx2_ASAP7_75t_L g210 ( .A(n_191), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_179), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_179), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g213 ( .A(n_192), .B(n_158), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_188), .Y(n_214) );
NAND2xp5_ASAP7_75t_SL g215 ( .A(n_178), .B(n_114), .Y(n_215) );
NAND2xp33_ASAP7_75t_L g216 ( .A(n_185), .B(n_153), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_179), .Y(n_217) );
INVx3_ASAP7_75t_L g218 ( .A(n_181), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_180), .Y(n_219) );
INVx2_ASAP7_75t_L g220 ( .A(n_180), .Y(n_220) );
AO221x1_ASAP7_75t_L g221 ( .A1(n_185), .A2(n_174), .B1(n_141), .B2(n_151), .C(n_136), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_188), .Y(n_222) );
NOR3xp33_ASAP7_75t_L g223 ( .A(n_183), .B(n_160), .C(n_177), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_198), .B(n_155), .Y(n_224) );
INVx2_ASAP7_75t_SL g225 ( .A(n_202), .Y(n_225) );
NAND2xp5_ASAP7_75t_SL g226 ( .A(n_194), .B(n_156), .Y(n_226) );
INVx3_ASAP7_75t_L g227 ( .A(n_181), .Y(n_227) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_200), .B(n_173), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_186), .B(n_176), .Y(n_229) );
INVx2_ASAP7_75t_L g230 ( .A(n_181), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_193), .Y(n_231) );
NOR2xp33_ASAP7_75t_L g232 ( .A(n_183), .B(n_142), .Y(n_232) );
INVx2_ASAP7_75t_SL g233 ( .A(n_185), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_193), .Y(n_234) );
INVx2_ASAP7_75t_SL g235 ( .A(n_185), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_186), .B(n_117), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_185), .B(n_126), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_180), .Y(n_238) );
INVx1_ASAP7_75t_L g239 ( .A(n_196), .Y(n_239) );
NAND2xp5_ASAP7_75t_L g240 ( .A(n_196), .B(n_124), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_189), .B(n_129), .Y(n_241) );
NAND2xp5_ASAP7_75t_SL g242 ( .A(n_181), .B(n_131), .Y(n_242) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_213), .B(n_187), .Y(n_243) );
OAI21xp5_ASAP7_75t_L g244 ( .A1(n_208), .A2(n_187), .B(n_184), .Y(n_244) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_206), .B(n_185), .Y(n_245) );
NAND2xp5_ASAP7_75t_L g246 ( .A(n_228), .B(n_187), .Y(n_246) );
INVx3_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_214), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_233), .A2(n_163), .B(n_184), .Y(n_249) );
INVx1_ASAP7_75t_L g250 ( .A(n_214), .Y(n_250) );
INVx4_ASAP7_75t_L g251 ( .A(n_218), .Y(n_251) );
NOR3xp33_ASAP7_75t_L g252 ( .A(n_223), .B(n_146), .C(n_120), .Y(n_252) );
AOI21xp5_ASAP7_75t_L g253 ( .A1(n_233), .A2(n_163), .B(n_184), .Y(n_253) );
INVx2_ASAP7_75t_L g254 ( .A(n_211), .Y(n_254) );
AOI21xp5_ASAP7_75t_L g255 ( .A1(n_235), .A2(n_195), .B(n_184), .Y(n_255) );
BUFx3_ASAP7_75t_L g256 ( .A(n_211), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_225), .B(n_195), .Y(n_257) );
OAI21xp5_ASAP7_75t_L g258 ( .A1(n_208), .A2(n_195), .B(n_205), .Y(n_258) );
INVx3_ASAP7_75t_L g259 ( .A(n_218), .Y(n_259) );
NAND2xp5_ASAP7_75t_L g260 ( .A(n_225), .B(n_195), .Y(n_260) );
AOI21xp5_ASAP7_75t_L g261 ( .A1(n_235), .A2(n_210), .B(n_208), .Y(n_261) );
BUFx3_ASAP7_75t_L g262 ( .A(n_211), .Y(n_262) );
AOI21xp5_ASAP7_75t_L g263 ( .A1(n_210), .A2(n_205), .B(n_204), .Y(n_263) );
AOI21xp5_ASAP7_75t_L g264 ( .A1(n_210), .A2(n_204), .B(n_201), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_229), .B(n_117), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g266 ( .A1(n_216), .A2(n_204), .B(n_201), .Y(n_266) );
INVx3_ASAP7_75t_L g267 ( .A(n_218), .Y(n_267) );
NOR2xp33_ASAP7_75t_L g268 ( .A(n_209), .B(n_116), .Y(n_268) );
INVxp67_ASAP7_75t_L g269 ( .A(n_236), .Y(n_269) );
AOI21xp5_ASAP7_75t_L g270 ( .A1(n_224), .A2(n_201), .B(n_199), .Y(n_270) );
NAND2xp5_ASAP7_75t_SL g271 ( .A(n_212), .B(n_122), .Y(n_271) );
INVx1_ASAP7_75t_L g272 ( .A(n_222), .Y(n_272) );
INVx11_ASAP7_75t_L g273 ( .A(n_226), .Y(n_273) );
NAND2xp5_ASAP7_75t_SL g274 ( .A(n_212), .B(n_128), .Y(n_274) );
O2A1O1Ixp33_ASAP7_75t_L g275 ( .A1(n_232), .A2(n_130), .B(n_132), .C(n_157), .Y(n_275) );
AOI31xp67_ASAP7_75t_L g276 ( .A1(n_271), .A2(n_199), .A3(n_197), .B(n_154), .Y(n_276) );
OAI21x1_ASAP7_75t_L g277 ( .A1(n_249), .A2(n_231), .B(n_222), .Y(n_277) );
AOI21x1_ASAP7_75t_SL g278 ( .A1(n_257), .A2(n_229), .B(n_236), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_248), .Y(n_279) );
BUFx10_ASAP7_75t_L g280 ( .A(n_245), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_250), .B(n_231), .Y(n_281) );
BUFx6f_ASAP7_75t_L g282 ( .A(n_256), .Y(n_282) );
A2O1A1Ixp33_ASAP7_75t_L g283 ( .A1(n_268), .A2(n_234), .B(n_239), .C(n_227), .Y(n_283) );
AOI21xp5_ASAP7_75t_L g284 ( .A1(n_253), .A2(n_237), .B(n_234), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_272), .B(n_239), .Y(n_285) );
OAI21x1_ASAP7_75t_L g286 ( .A1(n_261), .A2(n_264), .B(n_244), .Y(n_286) );
AOI22xp5_ASAP7_75t_L g287 ( .A1(n_265), .A2(n_207), .B1(n_215), .B2(n_240), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_243), .Y(n_288) );
AND2x2_ASAP7_75t_L g289 ( .A(n_269), .B(n_252), .Y(n_289) );
OAI21x1_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_212), .B(n_217), .Y(n_290) );
BUFx6f_ASAP7_75t_L g291 ( .A(n_256), .Y(n_291) );
BUFx3_ASAP7_75t_L g292 ( .A(n_262), .Y(n_292) );
NAND3xp33_ASAP7_75t_L g293 ( .A(n_268), .B(n_237), .C(n_207), .Y(n_293) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_245), .B(n_217), .Y(n_294) );
INVx1_ASAP7_75t_SL g295 ( .A(n_260), .Y(n_295) );
AOI21xp5_ASAP7_75t_L g296 ( .A1(n_263), .A2(n_237), .B(n_220), .Y(n_296) );
AOI221x1_ASAP7_75t_L g297 ( .A1(n_266), .A2(n_221), .B1(n_174), .B2(n_133), .C(n_197), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_246), .B(n_217), .Y(n_298) );
AO31x2_ASAP7_75t_L g299 ( .A1(n_254), .A2(n_221), .A3(n_199), .B(n_197), .Y(n_299) );
NAND2xp33_ASAP7_75t_L g300 ( .A(n_254), .B(n_219), .Y(n_300) );
A2O1A1Ixp33_ASAP7_75t_L g301 ( .A1(n_275), .A2(n_227), .B(n_219), .C(n_238), .Y(n_301) );
AOI21xp5_ASAP7_75t_SL g302 ( .A1(n_298), .A2(n_262), .B(n_237), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_288), .B(n_247), .Y(n_303) );
OAI21x1_ASAP7_75t_L g304 ( .A1(n_284), .A2(n_270), .B(n_255), .Y(n_304) );
AO21x2_ASAP7_75t_L g305 ( .A1(n_284), .A2(n_274), .B(n_271), .Y(n_305) );
AOI21xp5_ASAP7_75t_L g306 ( .A1(n_300), .A2(n_237), .B(n_274), .Y(n_306) );
INVx2_ASAP7_75t_L g307 ( .A(n_277), .Y(n_307) );
OAI21x1_ASAP7_75t_L g308 ( .A1(n_286), .A2(n_296), .B(n_297), .Y(n_308) );
AND2x2_ASAP7_75t_L g309 ( .A(n_298), .B(n_219), .Y(n_309) );
INVx2_ASAP7_75t_L g310 ( .A(n_290), .Y(n_310) );
OAI21x1_ASAP7_75t_L g311 ( .A1(n_296), .A2(n_247), .B(n_267), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g312 ( .A(n_281), .B(n_247), .Y(n_312) );
INVx4_ASAP7_75t_SL g313 ( .A(n_282), .Y(n_313) );
AOI21x1_ASAP7_75t_L g314 ( .A1(n_293), .A2(n_139), .B(n_154), .Y(n_314) );
INVx1_ASAP7_75t_L g315 ( .A(n_281), .Y(n_315) );
OAI21x1_ASAP7_75t_L g316 ( .A1(n_278), .A2(n_267), .B(n_259), .Y(n_316) );
INVx1_ASAP7_75t_L g317 ( .A(n_285), .Y(n_317) );
NOR2xp67_ASAP7_75t_L g318 ( .A(n_279), .B(n_251), .Y(n_318) );
AOI22xp33_ASAP7_75t_L g319 ( .A1(n_289), .A2(n_251), .B1(n_259), .B2(n_227), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_294), .Y(n_320) );
INVxp67_ASAP7_75t_SL g321 ( .A(n_282), .Y(n_321) );
INVx1_ASAP7_75t_SL g322 ( .A(n_292), .Y(n_322) );
OA21x2_ASAP7_75t_L g323 ( .A1(n_283), .A2(n_152), .B(n_230), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_320), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_320), .Y(n_325) );
INVx1_ASAP7_75t_L g326 ( .A(n_320), .Y(n_326) );
BUFx2_ASAP7_75t_L g327 ( .A(n_321), .Y(n_327) );
OAI21x1_ASAP7_75t_L g328 ( .A1(n_308), .A2(n_294), .B(n_285), .Y(n_328) );
INVx3_ASAP7_75t_L g329 ( .A(n_309), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_309), .B(n_280), .Y(n_330) );
AND2x4_ASAP7_75t_L g331 ( .A(n_313), .B(n_282), .Y(n_331) );
INVx2_ASAP7_75t_L g332 ( .A(n_307), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_315), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_315), .Y(n_334) );
INVx6_ASAP7_75t_L g335 ( .A(n_313), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_307), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_317), .Y(n_337) );
AND2x2_ASAP7_75t_L g338 ( .A(n_317), .B(n_280), .Y(n_338) );
INVx4_ASAP7_75t_L g339 ( .A(n_313), .Y(n_339) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_322), .Y(n_340) );
AND2x2_ASAP7_75t_L g341 ( .A(n_312), .B(n_291), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_307), .Y(n_342) );
OR2x6_ASAP7_75t_L g343 ( .A(n_302), .B(n_318), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_312), .Y(n_344) );
HB1xp67_ASAP7_75t_L g345 ( .A(n_322), .Y(n_345) );
NAND2x1_ASAP7_75t_L g346 ( .A(n_318), .B(n_291), .Y(n_346) );
INVx1_ASAP7_75t_L g347 ( .A(n_311), .Y(n_347) );
INVxp67_ASAP7_75t_SL g348 ( .A(n_321), .Y(n_348) );
BUFx2_ASAP7_75t_L g349 ( .A(n_311), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_303), .Y(n_350) );
INVx1_ASAP7_75t_L g351 ( .A(n_311), .Y(n_351) );
AND2x2_ASAP7_75t_L g352 ( .A(n_329), .B(n_323), .Y(n_352) );
AND2x4_ASAP7_75t_L g353 ( .A(n_343), .B(n_313), .Y(n_353) );
OR2x6_ASAP7_75t_L g354 ( .A(n_343), .B(n_308), .Y(n_354) );
INVx2_ASAP7_75t_SL g355 ( .A(n_327), .Y(n_355) );
OAI21x1_ASAP7_75t_L g356 ( .A1(n_328), .A2(n_308), .B(n_304), .Y(n_356) );
AND2x2_ASAP7_75t_L g357 ( .A(n_329), .B(n_323), .Y(n_357) );
NOR2xp33_ASAP7_75t_L g358 ( .A(n_338), .B(n_295), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_329), .B(n_323), .Y(n_359) );
INVx1_ASAP7_75t_L g360 ( .A(n_333), .Y(n_360) );
INVx1_ASAP7_75t_L g361 ( .A(n_333), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_332), .Y(n_362) );
OR2x2_ASAP7_75t_L g363 ( .A(n_324), .B(n_323), .Y(n_363) );
AND2x2_ASAP7_75t_L g364 ( .A(n_325), .B(n_324), .Y(n_364) );
OAI21x1_ASAP7_75t_L g365 ( .A1(n_328), .A2(n_304), .B(n_314), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_326), .B(n_323), .Y(n_366) );
OR2x2_ASAP7_75t_L g367 ( .A(n_326), .B(n_299), .Y(n_367) );
HB1xp67_ASAP7_75t_L g368 ( .A(n_327), .Y(n_368) );
BUFx3_ASAP7_75t_L g369 ( .A(n_335), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_334), .Y(n_370) );
INVx2_ASAP7_75t_L g371 ( .A(n_332), .Y(n_371) );
BUFx3_ASAP7_75t_L g372 ( .A(n_335), .Y(n_372) );
AND2x2_ASAP7_75t_L g373 ( .A(n_325), .B(n_305), .Y(n_373) );
NAND2xp5_ASAP7_75t_SL g374 ( .A(n_339), .B(n_313), .Y(n_374) );
BUFx12f_ASAP7_75t_L g375 ( .A(n_335), .Y(n_375) );
INVx2_ASAP7_75t_L g376 ( .A(n_336), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_334), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_337), .Y(n_378) );
NOR2x1_ASAP7_75t_L g379 ( .A(n_339), .B(n_305), .Y(n_379) );
INVx2_ASAP7_75t_L g380 ( .A(n_336), .Y(n_380) );
OR2x2_ASAP7_75t_L g381 ( .A(n_350), .B(n_299), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_337), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_341), .B(n_305), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_342), .Y(n_384) );
AND2x2_ASAP7_75t_L g385 ( .A(n_341), .B(n_305), .Y(n_385) );
AND2x2_ASAP7_75t_L g386 ( .A(n_344), .B(n_299), .Y(n_386) );
BUFx2_ASAP7_75t_L g387 ( .A(n_343), .Y(n_387) );
AND2x2_ASAP7_75t_L g388 ( .A(n_342), .B(n_310), .Y(n_388) );
INVx2_ASAP7_75t_L g389 ( .A(n_347), .Y(n_389) );
OR2x2_ASAP7_75t_L g390 ( .A(n_344), .B(n_310), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_351), .Y(n_391) );
AND2x4_ASAP7_75t_SL g392 ( .A(n_339), .B(n_291), .Y(n_392) );
AND2x2_ASAP7_75t_L g393 ( .A(n_330), .B(n_310), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_330), .B(n_304), .Y(n_394) );
AND2x2_ASAP7_75t_L g395 ( .A(n_338), .B(n_303), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_343), .Y(n_396) );
INVx1_ASAP7_75t_L g397 ( .A(n_351), .Y(n_397) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_368), .Y(n_398) );
INVxp67_ASAP7_75t_SL g399 ( .A(n_368), .Y(n_399) );
INVx2_ASAP7_75t_L g400 ( .A(n_389), .Y(n_400) );
INVx2_ASAP7_75t_SL g401 ( .A(n_355), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_360), .B(n_340), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_383), .B(n_347), .Y(n_403) );
INVx2_ASAP7_75t_L g404 ( .A(n_389), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_389), .Y(n_406) );
AND2x4_ASAP7_75t_L g407 ( .A(n_387), .B(n_343), .Y(n_407) );
AND2x2_ASAP7_75t_L g408 ( .A(n_383), .B(n_349), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_361), .B(n_345), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_361), .Y(n_410) );
NAND2xp5_ASAP7_75t_L g411 ( .A(n_370), .B(n_348), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_370), .Y(n_412) );
NAND2xp5_ASAP7_75t_L g413 ( .A(n_377), .B(n_378), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g414 ( .A1(n_394), .A2(n_319), .B1(n_349), .B2(n_335), .Y(n_414) );
AND2x4_ASAP7_75t_L g415 ( .A(n_387), .B(n_339), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_391), .Y(n_416) );
OR2x2_ASAP7_75t_L g417 ( .A(n_385), .B(n_346), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_377), .Y(n_418) );
NAND2xp5_ASAP7_75t_L g419 ( .A(n_378), .B(n_331), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g420 ( .A1(n_394), .A2(n_306), .B1(n_331), .B2(n_316), .Y(n_420) );
INVx1_ASAP7_75t_SL g421 ( .A(n_375), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_391), .Y(n_422) );
HB1xp67_ASAP7_75t_L g423 ( .A(n_355), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_391), .Y(n_424) );
AND2x4_ASAP7_75t_L g425 ( .A(n_396), .B(n_331), .Y(n_425) );
INVx2_ASAP7_75t_L g426 ( .A(n_362), .Y(n_426) );
INVx5_ASAP7_75t_L g427 ( .A(n_375), .Y(n_427) );
INVx1_ASAP7_75t_SL g428 ( .A(n_375), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_382), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_362), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_382), .Y(n_431) );
OR2x2_ASAP7_75t_L g432 ( .A(n_385), .B(n_346), .Y(n_432) );
NOR2xp67_ASAP7_75t_L g433 ( .A(n_355), .B(n_331), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g434 ( .A(n_395), .B(n_5), .Y(n_434) );
INVx2_ASAP7_75t_L g435 ( .A(n_362), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_397), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_395), .B(n_8), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_393), .B(n_314), .Y(n_438) );
NAND2x1p5_ASAP7_75t_L g439 ( .A(n_374), .B(n_316), .Y(n_439) );
AND2x2_ASAP7_75t_L g440 ( .A(n_393), .B(n_316), .Y(n_440) );
INVx1_ASAP7_75t_L g441 ( .A(n_397), .Y(n_441) );
AND2x4_ASAP7_75t_SL g442 ( .A(n_353), .B(n_251), .Y(n_442) );
INVx1_ASAP7_75t_L g443 ( .A(n_364), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_352), .B(n_147), .Y(n_444) );
AND2x2_ASAP7_75t_L g445 ( .A(n_352), .B(n_147), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_371), .Y(n_446) );
INVx1_ASAP7_75t_L g447 ( .A(n_364), .Y(n_447) );
OR2x2_ASAP7_75t_L g448 ( .A(n_381), .B(n_174), .Y(n_448) );
AND2x2_ASAP7_75t_L g449 ( .A(n_357), .B(n_306), .Y(n_449) );
AND2x4_ASAP7_75t_L g450 ( .A(n_396), .B(n_174), .Y(n_450) );
BUFx2_ASAP7_75t_L g451 ( .A(n_379), .Y(n_451) );
INVxp67_ASAP7_75t_L g452 ( .A(n_358), .Y(n_452) );
AND2x2_ASAP7_75t_L g453 ( .A(n_357), .B(n_174), .Y(n_453) );
INVx1_ASAP7_75t_L g454 ( .A(n_364), .Y(n_454) );
BUFx2_ASAP7_75t_L g455 ( .A(n_379), .Y(n_455) );
AND2x2_ASAP7_75t_L g456 ( .A(n_359), .B(n_9), .Y(n_456) );
AND2x2_ASAP7_75t_L g457 ( .A(n_359), .B(n_9), .Y(n_457) );
AND2x2_ASAP7_75t_L g458 ( .A(n_366), .B(n_10), .Y(n_458) );
BUFx2_ASAP7_75t_L g459 ( .A(n_353), .Y(n_459) );
INVx2_ASAP7_75t_L g460 ( .A(n_371), .Y(n_460) );
AND2x4_ASAP7_75t_L g461 ( .A(n_353), .B(n_20), .Y(n_461) );
INVx2_ASAP7_75t_L g462 ( .A(n_371), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_376), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_384), .Y(n_464) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_358), .B(n_273), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_376), .Y(n_466) );
AND2x2_ASAP7_75t_L g467 ( .A(n_452), .B(n_366), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g468 ( .A(n_443), .B(n_386), .Y(n_468) );
INVx2_ASAP7_75t_SL g469 ( .A(n_427), .Y(n_469) );
INVx1_ASAP7_75t_L g470 ( .A(n_405), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_405), .Y(n_471) );
INVx2_ASAP7_75t_L g472 ( .A(n_400), .Y(n_472) );
INVx1_ASAP7_75t_SL g473 ( .A(n_421), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_408), .B(n_386), .Y(n_474) );
AND2x2_ASAP7_75t_L g475 ( .A(n_408), .B(n_373), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_403), .B(n_381), .Y(n_476) );
AND2x2_ASAP7_75t_L g477 ( .A(n_403), .B(n_373), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_410), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_410), .Y(n_479) );
AND2x2_ASAP7_75t_L g480 ( .A(n_443), .B(n_354), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_412), .Y(n_481) );
AND2x2_ASAP7_75t_L g482 ( .A(n_447), .B(n_354), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_412), .Y(n_483) );
OR2x2_ASAP7_75t_L g484 ( .A(n_402), .B(n_409), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_447), .B(n_354), .Y(n_485) );
INVx2_ASAP7_75t_L g486 ( .A(n_400), .Y(n_486) );
HB1xp67_ASAP7_75t_L g487 ( .A(n_398), .Y(n_487) );
OR2x2_ASAP7_75t_L g488 ( .A(n_454), .B(n_367), .Y(n_488) );
OR2x2_ASAP7_75t_L g489 ( .A(n_454), .B(n_367), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g490 ( .A(n_418), .B(n_363), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_418), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g492 ( .A(n_429), .B(n_363), .Y(n_492) );
INVx1_ASAP7_75t_L g493 ( .A(n_429), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_459), .B(n_354), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_459), .B(n_354), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_431), .B(n_384), .Y(n_496) );
AND2x2_ASAP7_75t_L g497 ( .A(n_456), .B(n_354), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_431), .Y(n_498) );
OR2x2_ASAP7_75t_L g499 ( .A(n_411), .B(n_390), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_436), .B(n_390), .Y(n_500) );
NAND2xp5_ASAP7_75t_L g501 ( .A(n_436), .B(n_376), .Y(n_501) );
INVx1_ASAP7_75t_L g502 ( .A(n_413), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_407), .B(n_353), .Y(n_503) );
INVx2_ASAP7_75t_L g504 ( .A(n_404), .Y(n_504) );
OR2x2_ASAP7_75t_L g505 ( .A(n_417), .B(n_380), .Y(n_505) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_441), .B(n_380), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_456), .B(n_388), .Y(n_507) );
INVx2_ASAP7_75t_SL g508 ( .A(n_427), .Y(n_508) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_441), .B(n_380), .Y(n_509) );
INVx1_ASAP7_75t_L g510 ( .A(n_464), .Y(n_510) );
OR2x2_ASAP7_75t_L g511 ( .A(n_417), .B(n_388), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_457), .B(n_388), .Y(n_512) );
INVxp67_ASAP7_75t_SL g513 ( .A(n_448), .Y(n_513) );
INVx2_ASAP7_75t_L g514 ( .A(n_404), .Y(n_514) );
INVx2_ASAP7_75t_L g515 ( .A(n_406), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_457), .B(n_369), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_432), .B(n_369), .Y(n_517) );
AND2x4_ASAP7_75t_L g518 ( .A(n_407), .B(n_369), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_464), .Y(n_519) );
HB1xp67_ASAP7_75t_L g520 ( .A(n_423), .Y(n_520) );
AND2x4_ASAP7_75t_L g521 ( .A(n_407), .B(n_372), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_432), .B(n_372), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_399), .Y(n_523) );
AND2x2_ASAP7_75t_L g524 ( .A(n_458), .B(n_372), .Y(n_524) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_433), .B(n_392), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_458), .Y(n_526) );
INVxp67_ASAP7_75t_L g527 ( .A(n_401), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_401), .B(n_392), .Y(n_528) );
OR2x2_ASAP7_75t_L g529 ( .A(n_448), .B(n_356), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_415), .B(n_356), .Y(n_530) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_444), .B(n_445), .Y(n_531) );
OR2x2_ASAP7_75t_L g532 ( .A(n_419), .B(n_356), .Y(n_532) );
INVx1_ASAP7_75t_L g533 ( .A(n_406), .Y(n_533) );
NAND2xp5_ASAP7_75t_SL g534 ( .A(n_433), .B(n_427), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_449), .B(n_392), .Y(n_535) );
AND2x2_ASAP7_75t_L g536 ( .A(n_449), .B(n_365), .Y(n_536) );
OR2x2_ASAP7_75t_SL g537 ( .A(n_434), .B(n_10), .Y(n_537) );
AND2x2_ASAP7_75t_L g538 ( .A(n_444), .B(n_365), .Y(n_538) );
INVxp67_ASAP7_75t_L g539 ( .A(n_451), .Y(n_539) );
INVxp67_ASAP7_75t_L g540 ( .A(n_451), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_416), .Y(n_541) );
NAND2x1_ASAP7_75t_L g542 ( .A(n_415), .B(n_365), .Y(n_542) );
INVx3_ASAP7_75t_L g543 ( .A(n_415), .Y(n_543) );
AND2x2_ASAP7_75t_L g544 ( .A(n_445), .B(n_11), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_425), .B(n_12), .Y(n_545) );
INVx1_ASAP7_75t_L g546 ( .A(n_416), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_422), .Y(n_547) );
AND2x2_ASAP7_75t_L g548 ( .A(n_425), .B(n_12), .Y(n_548) );
INVx1_ASAP7_75t_SL g549 ( .A(n_428), .Y(n_549) );
INVx2_ASAP7_75t_L g550 ( .A(n_422), .Y(n_550) );
INVx1_ASAP7_75t_SL g551 ( .A(n_427), .Y(n_551) );
INVx1_ASAP7_75t_L g552 ( .A(n_487), .Y(n_552) );
HB1xp67_ASAP7_75t_L g553 ( .A(n_487), .Y(n_553) );
INVx1_ASAP7_75t_SL g554 ( .A(n_473), .Y(n_554) );
AND2x2_ASAP7_75t_L g555 ( .A(n_477), .B(n_425), .Y(n_555) );
AND2x2_ASAP7_75t_L g556 ( .A(n_467), .B(n_453), .Y(n_556) );
OAI21xp33_ASAP7_75t_L g557 ( .A1(n_549), .A2(n_414), .B(n_437), .Y(n_557) );
INVx1_ASAP7_75t_L g558 ( .A(n_502), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_470), .Y(n_559) );
OR2x2_ASAP7_75t_L g560 ( .A(n_476), .B(n_453), .Y(n_560) );
AOI211xp5_ASAP7_75t_L g561 ( .A1(n_534), .A2(n_465), .B(n_461), .C(n_455), .Y(n_561) );
INVx1_ASAP7_75t_L g562 ( .A(n_471), .Y(n_562) );
INVx1_ASAP7_75t_SL g563 ( .A(n_551), .Y(n_563) );
AND2x4_ASAP7_75t_L g564 ( .A(n_503), .B(n_530), .Y(n_564) );
OR2x2_ASAP7_75t_L g565 ( .A(n_484), .B(n_424), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_475), .B(n_440), .Y(n_566) );
OR2x6_ASAP7_75t_L g567 ( .A(n_534), .B(n_455), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_520), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_511), .B(n_424), .Y(n_569) );
INVx1_ASAP7_75t_SL g570 ( .A(n_520), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g571 ( .A(n_490), .B(n_426), .Y(n_571) );
INVx2_ASAP7_75t_L g572 ( .A(n_505), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g573 ( .A(n_490), .B(n_426), .Y(n_573) );
NAND2xp5_ASAP7_75t_L g574 ( .A(n_492), .B(n_430), .Y(n_574) );
INVx1_ASAP7_75t_L g575 ( .A(n_478), .Y(n_575) );
INVxp33_ASAP7_75t_L g576 ( .A(n_525), .Y(n_576) );
NOR2xp33_ASAP7_75t_L g577 ( .A(n_537), .B(n_427), .Y(n_577) );
INVx2_ASAP7_75t_SL g578 ( .A(n_469), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_474), .B(n_440), .Y(n_579) );
AND2x4_ASAP7_75t_SL g580 ( .A(n_517), .B(n_461), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_479), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_481), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_483), .Y(n_583) );
INVx1_ASAP7_75t_L g584 ( .A(n_491), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_522), .B(n_438), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g586 ( .A(n_492), .B(n_430), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_493), .Y(n_587) );
AND2x2_ASAP7_75t_L g588 ( .A(n_507), .B(n_438), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_468), .B(n_435), .Y(n_589) );
AOI22xp5_ASAP7_75t_L g590 ( .A1(n_531), .A2(n_450), .B1(n_427), .B2(n_461), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_468), .B(n_435), .Y(n_591) );
AND2x2_ASAP7_75t_L g592 ( .A(n_512), .B(n_450), .Y(n_592) );
INVx1_ASAP7_75t_L g593 ( .A(n_498), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_510), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_519), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_523), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_472), .Y(n_597) );
NAND2xp33_ASAP7_75t_L g598 ( .A(n_508), .B(n_439), .Y(n_598) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_526), .B(n_450), .Y(n_599) );
INVx1_ASAP7_75t_L g600 ( .A(n_496), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_496), .Y(n_601) );
AND2x2_ASAP7_75t_L g602 ( .A(n_535), .B(n_439), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_497), .B(n_439), .Y(n_603) );
BUFx2_ASAP7_75t_L g604 ( .A(n_527), .Y(n_604) );
AND2x2_ASAP7_75t_L g605 ( .A(n_480), .B(n_446), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_482), .B(n_446), .Y(n_606) );
NOR2x1p5_ASAP7_75t_SL g607 ( .A(n_529), .B(n_460), .Y(n_607) );
OR2x2_ASAP7_75t_L g608 ( .A(n_499), .B(n_460), .Y(n_608) );
AND2x2_ASAP7_75t_L g609 ( .A(n_485), .B(n_462), .Y(n_609) );
INVx1_ASAP7_75t_L g610 ( .A(n_488), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_489), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_472), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_500), .Y(n_613) );
AND2x4_ASAP7_75t_L g614 ( .A(n_503), .B(n_442), .Y(n_614) );
OR2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_462), .Y(n_615) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_513), .B(n_463), .Y(n_616) );
AND2x2_ASAP7_75t_SL g617 ( .A(n_503), .B(n_442), .Y(n_617) );
NOR2xp33_ASAP7_75t_L g618 ( .A(n_545), .B(n_13), .Y(n_618) );
NAND2xp5_ASAP7_75t_L g619 ( .A(n_536), .B(n_463), .Y(n_619) );
NOR2xp33_ASAP7_75t_L g620 ( .A(n_548), .B(n_13), .Y(n_620) );
INVx3_ASAP7_75t_L g621 ( .A(n_542), .Y(n_621) );
AND2x2_ASAP7_75t_L g622 ( .A(n_494), .B(n_466), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_500), .Y(n_623) );
BUFx2_ASAP7_75t_L g624 ( .A(n_527), .Y(n_624) );
OR2x2_ASAP7_75t_L g625 ( .A(n_531), .B(n_466), .Y(n_625) );
NOR5xp2_ASAP7_75t_L g626 ( .A(n_539), .B(n_420), .C(n_15), .D(n_16), .E(n_17), .Y(n_626) );
AND2x2_ASAP7_75t_L g627 ( .A(n_495), .B(n_14), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_501), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_486), .Y(n_629) );
AND2x2_ASAP7_75t_L g630 ( .A(n_543), .B(n_16), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_613), .B(n_532), .Y(n_631) );
NAND3x2_ASAP7_75t_L g632 ( .A(n_604), .B(n_518), .C(n_521), .Y(n_632) );
AOI21xp5_ASAP7_75t_L g633 ( .A1(n_561), .A2(n_539), .B(n_540), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_552), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_553), .Y(n_635) );
INVx2_ASAP7_75t_L g636 ( .A(n_615), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_568), .Y(n_637) );
O2A1O1Ixp33_ASAP7_75t_L g638 ( .A1(n_554), .A2(n_540), .B(n_544), .C(n_543), .Y(n_638) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_557), .A2(n_530), .B1(n_538), .B2(n_524), .Y(n_639) );
AND2x2_ASAP7_75t_L g640 ( .A(n_564), .B(n_530), .Y(n_640) );
NAND3xp33_ASAP7_75t_L g641 ( .A(n_626), .B(n_533), .C(n_547), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_625), .Y(n_642) );
INVx1_ASAP7_75t_L g643 ( .A(n_628), .Y(n_643) );
INVxp67_ASAP7_75t_L g644 ( .A(n_554), .Y(n_644) );
OAI21xp5_ASAP7_75t_SL g645 ( .A1(n_577), .A2(n_518), .B(n_521), .Y(n_645) );
AND2x2_ASAP7_75t_L g646 ( .A(n_564), .B(n_518), .Y(n_646) );
INVxp67_ASAP7_75t_L g647 ( .A(n_624), .Y(n_647) );
OAI21xp33_ASAP7_75t_SL g648 ( .A1(n_617), .A2(n_528), .B(n_516), .Y(n_648) );
OAI22xp33_ASAP7_75t_L g649 ( .A1(n_576), .A2(n_521), .B1(n_501), .B2(n_506), .Y(n_649) );
AOI21xp33_ASAP7_75t_SL g650 ( .A1(n_567), .A2(n_509), .B(n_506), .Y(n_650) );
INVx2_ASAP7_75t_L g651 ( .A(n_568), .Y(n_651) );
OR2x2_ASAP7_75t_L g652 ( .A(n_619), .B(n_541), .Y(n_652) );
INVx2_ASAP7_75t_SL g653 ( .A(n_614), .Y(n_653) );
OAI22xp33_ASAP7_75t_L g654 ( .A1(n_567), .A2(n_509), .B1(n_546), .B2(n_515), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_623), .B(n_486), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_570), .Y(n_656) );
OR2x2_ASAP7_75t_L g657 ( .A(n_619), .B(n_504), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_600), .Y(n_658) );
OAI22xp33_ASAP7_75t_L g659 ( .A1(n_567), .A2(n_550), .B1(n_515), .B2(n_514), .Y(n_659) );
AOI22xp33_ASAP7_75t_L g660 ( .A1(n_557), .A2(n_550), .B1(n_514), .B2(n_504), .Y(n_660) );
INVx1_ASAP7_75t_L g661 ( .A(n_601), .Y(n_661) );
AOI21xp33_ASAP7_75t_L g662 ( .A1(n_618), .A2(n_17), .B(n_287), .Y(n_662) );
OAI322xp33_ASAP7_75t_L g663 ( .A1(n_570), .A2(n_610), .A3(n_611), .B1(n_558), .B2(n_620), .C1(n_560), .C2(n_565), .Y(n_663) );
AOI322xp5_ASAP7_75t_L g664 ( .A1(n_627), .A2(n_301), .A3(n_242), .B1(n_276), .B2(n_134), .C1(n_150), .C2(n_138), .Y(n_664) );
OR2x2_ASAP7_75t_L g665 ( .A(n_569), .B(n_238), .Y(n_665) );
OAI22xp5_ASAP7_75t_L g666 ( .A1(n_561), .A2(n_143), .B1(n_227), .B2(n_238), .Y(n_666) );
INVxp33_ASAP7_75t_L g667 ( .A(n_614), .Y(n_667) );
OR2x2_ASAP7_75t_L g668 ( .A(n_608), .B(n_220), .Y(n_668) );
AOI21xp33_ASAP7_75t_L g669 ( .A1(n_630), .A2(n_21), .B(n_26), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_589), .Y(n_670) );
AND2x2_ASAP7_75t_L g671 ( .A(n_566), .B(n_28), .Y(n_671) );
OAI21xp33_ASAP7_75t_SL g672 ( .A1(n_621), .A2(n_220), .B(n_31), .Y(n_672) );
OAI221xp5_ASAP7_75t_SL g673 ( .A1(n_590), .A2(n_241), .B1(n_230), .B2(n_35), .C(n_36), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_589), .Y(n_674) );
OAI322xp33_ASAP7_75t_L g675 ( .A1(n_591), .A2(n_30), .A3(n_33), .B1(n_37), .B2(n_39), .C1(n_41), .C2(n_46), .Y(n_675) );
OAI22xp33_ASAP7_75t_L g676 ( .A1(n_578), .A2(n_47), .B1(n_50), .B2(n_51), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_596), .B(n_53), .Y(n_677) );
OR2x2_ASAP7_75t_L g678 ( .A(n_572), .B(n_54), .Y(n_678) );
AND2x2_ASAP7_75t_L g679 ( .A(n_579), .B(n_55), .Y(n_679) );
OAI21xp33_ASAP7_75t_SL g680 ( .A1(n_621), .A2(n_60), .B(n_61), .Y(n_680) );
INVx1_ASAP7_75t_L g681 ( .A(n_591), .Y(n_681) );
NAND2xp33_ASAP7_75t_SL g682 ( .A(n_555), .B(n_64), .Y(n_682) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_607), .A2(n_65), .B(n_66), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_643), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_635), .B(n_556), .Y(n_685) );
NAND2xp5_ASAP7_75t_SL g686 ( .A(n_648), .B(n_563), .Y(n_686) );
AND2x2_ASAP7_75t_L g687 ( .A(n_640), .B(n_588), .Y(n_687) );
HB1xp67_ASAP7_75t_L g688 ( .A(n_637), .Y(n_688) );
INVx2_ASAP7_75t_L g689 ( .A(n_657), .Y(n_689) );
A2O1A1Ixp33_ASAP7_75t_L g690 ( .A1(n_645), .A2(n_580), .B(n_598), .C(n_592), .Y(n_690) );
O2A1O1Ixp33_ASAP7_75t_L g691 ( .A1(n_666), .A2(n_563), .B(n_599), .C(n_616), .Y(n_691) );
NAND2xp5_ASAP7_75t_L g692 ( .A(n_670), .B(n_571), .Y(n_692) );
OAI22xp33_ASAP7_75t_L g693 ( .A1(n_645), .A2(n_571), .B1(n_573), .B2(n_574), .Y(n_693) );
AOI321xp33_ASAP7_75t_L g694 ( .A1(n_639), .A2(n_603), .A3(n_602), .B1(n_585), .B2(n_586), .C(n_574), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_674), .B(n_573), .Y(n_695) );
AOI221xp5_ASAP7_75t_L g696 ( .A1(n_663), .A2(n_593), .B1(n_562), .B2(n_575), .C(n_581), .Y(n_696) );
OAI22xp5_ASAP7_75t_L g697 ( .A1(n_632), .A2(n_586), .B1(n_605), .B2(n_606), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_681), .Y(n_698) );
AOI21xp33_ASAP7_75t_L g699 ( .A1(n_641), .A2(n_594), .B(n_582), .Y(n_699) );
NAND3xp33_ASAP7_75t_L g700 ( .A(n_641), .B(n_595), .C(n_583), .Y(n_700) );
AOI21xp33_ASAP7_75t_SL g701 ( .A1(n_666), .A2(n_559), .B(n_584), .Y(n_701) );
AOI221xp5_ASAP7_75t_L g702 ( .A1(n_649), .A2(n_587), .B1(n_612), .B2(n_597), .C(n_629), .Y(n_702) );
AND2x2_ASAP7_75t_SL g703 ( .A(n_660), .B(n_622), .Y(n_703) );
NAND2xp5_ASAP7_75t_L g704 ( .A(n_658), .B(n_609), .Y(n_704) );
AND2x2_ASAP7_75t_L g705 ( .A(n_667), .B(n_67), .Y(n_705) );
AOI22xp5_ASAP7_75t_L g706 ( .A1(n_644), .A2(n_72), .B1(n_74), .B2(n_76), .Y(n_706) );
INVx2_ASAP7_75t_L g707 ( .A(n_652), .Y(n_707) );
INVx2_ASAP7_75t_SL g708 ( .A(n_653), .Y(n_708) );
AOI21xp5_ASAP7_75t_L g709 ( .A1(n_672), .A2(n_77), .B(n_78), .Y(n_709) );
AOI211xp5_ASAP7_75t_L g710 ( .A1(n_680), .A2(n_80), .B(n_83), .C(n_84), .Y(n_710) );
OAI22xp33_ASAP7_75t_L g711 ( .A1(n_650), .A2(n_85), .B1(n_86), .B2(n_90), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g712 ( .A(n_661), .B(n_91), .Y(n_712) );
OAI21xp5_ASAP7_75t_SL g713 ( .A1(n_696), .A2(n_638), .B(n_633), .Y(n_713) );
O2A1O1Ixp33_ASAP7_75t_L g714 ( .A1(n_699), .A2(n_662), .B(n_647), .C(n_654), .Y(n_714) );
NOR2xp33_ASAP7_75t_L g715 ( .A(n_708), .B(n_646), .Y(n_715) );
NAND4xp75_ASAP7_75t_L g716 ( .A(n_703), .B(n_679), .C(n_671), .D(n_662), .Y(n_716) );
AND2x2_ASAP7_75t_L g717 ( .A(n_687), .B(n_642), .Y(n_717) );
NAND2xp5_ASAP7_75t_SL g718 ( .A(n_696), .B(n_686), .Y(n_718) );
AOI211xp5_ASAP7_75t_L g719 ( .A1(n_700), .A2(n_682), .B(n_659), .C(n_673), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_688), .Y(n_720) );
AND2x2_ASAP7_75t_L g721 ( .A(n_690), .B(n_636), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g722 ( .A(n_698), .B(n_634), .Y(n_722) );
NOR2xp33_ASAP7_75t_SL g723 ( .A(n_711), .B(n_683), .Y(n_723) );
AOI221xp5_ASAP7_75t_L g724 ( .A1(n_693), .A2(n_631), .B1(n_656), .B2(n_651), .C(n_655), .Y(n_724) );
AOI21xp33_ASAP7_75t_SL g725 ( .A1(n_691), .A2(n_669), .B(n_676), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g726 ( .A(n_707), .B(n_665), .Y(n_726) );
AOI21xp33_ASAP7_75t_L g727 ( .A1(n_691), .A2(n_668), .B(n_677), .Y(n_727) );
AOI221x1_ASAP7_75t_L g728 ( .A1(n_720), .A2(n_701), .B1(n_705), .B2(n_709), .C(n_712), .Y(n_728) );
NAND4xp25_ASAP7_75t_L g729 ( .A(n_723), .B(n_694), .C(n_710), .D(n_709), .Y(n_729) );
NAND3xp33_ASAP7_75t_L g730 ( .A(n_718), .B(n_702), .C(n_684), .Y(n_730) );
NOR2xp33_ASAP7_75t_L g731 ( .A(n_713), .B(n_685), .Y(n_731) );
NOR2xp67_ASAP7_75t_L g732 ( .A(n_721), .B(n_697), .Y(n_732) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_723), .A2(n_702), .B(n_695), .Y(n_733) );
NAND5xp2_ASAP7_75t_L g734 ( .A(n_719), .B(n_669), .C(n_706), .D(n_664), .E(n_704), .Y(n_734) );
NAND4xp75_ASAP7_75t_L g735 ( .A(n_724), .B(n_692), .C(n_689), .D(n_675), .Y(n_735) );
OAI21xp33_ASAP7_75t_L g736 ( .A1(n_731), .A2(n_725), .B(n_714), .Y(n_736) );
NOR2x1_ASAP7_75t_SL g737 ( .A(n_735), .B(n_716), .Y(n_737) );
AOI211xp5_ASAP7_75t_L g738 ( .A1(n_734), .A2(n_727), .B(n_715), .C(n_726), .Y(n_738) );
NOR2xp67_ASAP7_75t_L g739 ( .A(n_729), .B(n_722), .Y(n_739) );
NOR3xp33_ASAP7_75t_L g740 ( .A(n_730), .B(n_717), .C(n_678), .Y(n_740) );
OR2x2_ASAP7_75t_L g741 ( .A(n_736), .B(n_733), .Y(n_741) );
NAND4xp75_ASAP7_75t_L g742 ( .A(n_739), .B(n_728), .C(n_732), .D(n_95), .Y(n_742) );
BUFx12f_ASAP7_75t_L g743 ( .A(n_737), .Y(n_743) );
INVx1_ASAP7_75t_L g744 ( .A(n_741), .Y(n_744) );
AOI31xp33_ASAP7_75t_L g745 ( .A1(n_743), .A2(n_738), .A3(n_740), .B(n_96), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_744), .Y(n_746) );
INVxp67_ASAP7_75t_SL g747 ( .A(n_745), .Y(n_747) );
AOI21xp5_ASAP7_75t_SL g748 ( .A1(n_747), .A2(n_742), .B(n_94), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_746), .B(n_93), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_748), .A2(n_746), .B(n_98), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g751 ( .A1(n_750), .A2(n_749), .B(n_99), .Y(n_751) );
OAI21xp33_ASAP7_75t_L g752 ( .A1(n_751), .A2(n_97), .B(n_100), .Y(n_752) );
OAI21xp5_ASAP7_75t_SL g753 ( .A1(n_752), .A2(n_102), .B(n_104), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g754 ( .A1(n_753), .A2(n_106), .B1(n_107), .B2(n_109), .Y(n_754) );
endmodule