module fake_jpeg_14118_n_561 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_561);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_561;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_352;
wire n_350;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx3_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_17),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

BUFx3_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

BUFx5_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_18),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_11),
.Y(n_36)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_1),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_1),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_15),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_4),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_2),
.B(n_1),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_15),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_8),
.Y(n_46)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_17),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_17),
.Y(n_49)
);

CKINVDCx14_ASAP7_75t_R g50 ( 
.A(n_10),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_10),
.Y(n_51)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_4),
.Y(n_52)
);

INVx11_ASAP7_75t_L g53 ( 
.A(n_33),
.Y(n_53)
);

BUFx10_ASAP7_75t_L g164 ( 
.A(n_53),
.Y(n_164)
);

INVx5_ASAP7_75t_L g54 ( 
.A(n_30),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g145 ( 
.A(n_54),
.Y(n_145)
);

INVx6_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_55),
.Y(n_109)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_56),
.Y(n_118)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_30),
.Y(n_57)
);

INVx3_ASAP7_75t_L g106 ( 
.A(n_57),
.Y(n_106)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_58),
.Y(n_110)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_33),
.Y(n_59)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_59),
.Y(n_126)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_26),
.Y(n_60)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_60),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_32),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g144 ( 
.A(n_61),
.Y(n_144)
);

INVx11_ASAP7_75t_L g62 ( 
.A(n_33),
.Y(n_62)
);

INVx8_ASAP7_75t_L g162 ( 
.A(n_62),
.Y(n_162)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_43),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_63),
.B(n_72),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_32),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g149 ( 
.A(n_64),
.Y(n_149)
);

BUFx12f_ASAP7_75t_L g65 ( 
.A(n_22),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g125 ( 
.A(n_65),
.Y(n_125)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_26),
.Y(n_66)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_66),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_32),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g152 ( 
.A(n_67),
.Y(n_152)
);

INVx5_ASAP7_75t_L g68 ( 
.A(n_30),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g163 ( 
.A(n_68),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_32),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_69),
.Y(n_154)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_22),
.Y(n_70)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_70),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_38),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_71),
.Y(n_169)
);

INVx2_ASAP7_75t_SL g72 ( 
.A(n_29),
.Y(n_72)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_23),
.Y(n_73)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx5_ASAP7_75t_L g117 ( 
.A(n_74),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_19),
.Y(n_75)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_75),
.Y(n_124)
);

INVx8_ASAP7_75t_L g76 ( 
.A(n_25),
.Y(n_76)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_76),
.Y(n_131)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_47),
.Y(n_77)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_78),
.Y(n_141)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_79),
.Y(n_138)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_23),
.Y(n_80)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_80),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_43),
.B(n_9),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_81),
.B(n_96),
.Y(n_107)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_82),
.Y(n_120)
);

BUFx3_ASAP7_75t_L g83 ( 
.A(n_25),
.Y(n_83)
);

INVx5_ASAP7_75t_L g150 ( 
.A(n_83),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g84 ( 
.A(n_25),
.Y(n_84)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_84),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g85 ( 
.A(n_29),
.Y(n_85)
);

INVx5_ASAP7_75t_L g153 ( 
.A(n_85),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_46),
.B(n_48),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g121 ( 
.A(n_86),
.B(n_92),
.Y(n_121)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_29),
.Y(n_87)
);

INVx3_ASAP7_75t_L g123 ( 
.A(n_87),
.Y(n_123)
);

BUFx4f_ASAP7_75t_L g88 ( 
.A(n_33),
.Y(n_88)
);

INVx3_ASAP7_75t_L g130 ( 
.A(n_88),
.Y(n_130)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_23),
.Y(n_89)
);

INVx3_ASAP7_75t_L g148 ( 
.A(n_89),
.Y(n_148)
);

INVx5_ASAP7_75t_L g90 ( 
.A(n_47),
.Y(n_90)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_90),
.Y(n_108)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_37),
.Y(n_91)
);

INVx4_ASAP7_75t_L g133 ( 
.A(n_91),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_46),
.B(n_9),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

INVx4_ASAP7_75t_L g115 ( 
.A(n_93),
.Y(n_115)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_35),
.Y(n_94)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_94),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_42),
.Y(n_95)
);

INVx4_ASAP7_75t_L g158 ( 
.A(n_95),
.Y(n_158)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_21),
.Y(n_96)
);

BUFx12f_ASAP7_75t_L g97 ( 
.A(n_37),
.Y(n_97)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_97),
.Y(n_139)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_35),
.B(n_39),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_98),
.B(n_21),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

INVx4_ASAP7_75t_L g165 ( 
.A(n_99),
.Y(n_165)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_47),
.Y(n_100)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_100),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_42),
.Y(n_101)
);

INVx3_ASAP7_75t_L g151 ( 
.A(n_101),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_42),
.Y(n_102)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_102),
.Y(n_160)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_28),
.Y(n_103)
);

INVx2_ASAP7_75t_L g129 ( 
.A(n_103),
.Y(n_129)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_28),
.Y(n_104)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_104),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_24),
.Y(n_105)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_105),
.Y(n_168)
);

AOI22xp33_ASAP7_75t_SL g112 ( 
.A1(n_72),
.A2(n_20),
.B1(n_19),
.B2(n_44),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_L g203 ( 
.A1(n_112),
.A2(n_127),
.B1(n_134),
.B2(n_147),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g127 ( 
.A1(n_87),
.A2(n_20),
.B1(n_19),
.B2(n_44),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_55),
.A2(n_24),
.B1(n_36),
.B2(n_40),
.Y(n_134)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_73),
.A2(n_50),
.B1(n_28),
.B2(n_44),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_136),
.A2(n_159),
.B1(n_70),
.B2(n_74),
.Y(n_181)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_88),
.Y(n_140)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_140),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g142 ( 
.A(n_57),
.B(n_48),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_142),
.B(n_155),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g143 ( 
.A(n_53),
.B(n_39),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_143),
.B(n_97),
.Y(n_170)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_146),
.B(n_14),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_76),
.A2(n_20),
.B1(n_31),
.B2(n_21),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_54),
.B(n_51),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g157 ( 
.A1(n_91),
.A2(n_21),
.B1(n_31),
.B2(n_40),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_83),
.B1(n_52),
.B2(n_93),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_80),
.A2(n_50),
.B1(n_36),
.B2(n_40),
.Y(n_159)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_68),
.B(n_21),
.Y(n_161)
);

AND2x2_ASAP7_75t_L g179 ( 
.A(n_161),
.B(n_85),
.Y(n_179)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_103),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_166),
.Y(n_191)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_104),
.Y(n_167)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_167),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_170),
.B(n_180),
.Y(n_240)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_107),
.B(n_59),
.C(n_62),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_171),
.B(n_212),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_118),
.B(n_41),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_172),
.B(n_0),
.Y(n_233)
);

AND2x4_ASAP7_75t_L g173 ( 
.A(n_110),
.B(n_37),
.Y(n_173)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_173),
.Y(n_274)
);

INVx13_ASAP7_75t_L g174 ( 
.A(n_164),
.Y(n_174)
);

BUFx24_ASAP7_75t_L g281 ( 
.A(n_174),
.Y(n_281)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_168),
.Y(n_175)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_175),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_114),
.A2(n_45),
.B1(n_51),
.B2(n_49),
.Y(n_176)
);

INVxp67_ASAP7_75t_L g246 ( 
.A(n_176),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_157),
.A2(n_78),
.B1(n_102),
.B2(n_101),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g254 ( 
.A1(n_177),
.A2(n_209),
.B1(n_71),
.B2(n_69),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g236 ( 
.A(n_179),
.B(n_189),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_121),
.B(n_45),
.Y(n_180)
);

CKINVDCx16_ASAP7_75t_R g276 ( 
.A(n_181),
.Y(n_276)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_129),
.Y(n_182)
);

INVx2_ASAP7_75t_L g267 ( 
.A(n_182),
.Y(n_267)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_132),
.Y(n_183)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_183),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g184 ( 
.A(n_130),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g266 ( 
.A(n_184),
.Y(n_266)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_111),
.Y(n_186)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_186),
.Y(n_237)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_122),
.Y(n_187)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_187),
.Y(n_238)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_113),
.Y(n_188)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_188),
.Y(n_247)
);

INVx4_ASAP7_75t_SL g189 ( 
.A(n_164),
.Y(n_189)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx4_ASAP7_75t_L g260 ( 
.A(n_190),
.Y(n_260)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_144),
.Y(n_192)
);

INVx6_ASAP7_75t_L g253 ( 
.A(n_192),
.Y(n_253)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_119),
.Y(n_193)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_193),
.Y(n_259)
);

INVx4_ASAP7_75t_L g194 ( 
.A(n_126),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_194),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_61),
.B1(n_99),
.B2(n_95),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_195),
.A2(n_141),
.B1(n_154),
.B2(n_169),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g196 ( 
.A(n_156),
.B(n_49),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_196),
.B(n_198),
.Y(n_251)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_143),
.Y(n_197)
);

CKINVDCx14_ASAP7_75t_R g256 ( 
.A(n_197),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_156),
.B(n_90),
.Y(n_198)
);

BUFx2_ASAP7_75t_L g199 ( 
.A(n_116),
.Y(n_199)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_124),
.Y(n_200)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_200),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_120),
.B(n_77),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_201),
.B(n_205),
.Y(n_242)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_144),
.Y(n_202)
);

INVx6_ASAP7_75t_L g271 ( 
.A(n_202),
.Y(n_271)
);

INVx1_ASAP7_75t_SL g204 ( 
.A(n_164),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g278 ( 
.A(n_204),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g205 ( 
.A(n_137),
.B(n_97),
.Y(n_205)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

INVx2_ASAP7_75t_SL g255 ( 
.A(n_207),
.Y(n_255)
);

A2O1A1Ixp33_ASAP7_75t_SL g268 ( 
.A1(n_208),
.A2(n_220),
.B(n_153),
.C(n_138),
.Y(n_268)
);

OAI22xp5_ASAP7_75t_SL g209 ( 
.A1(n_127),
.A2(n_67),
.B1(n_64),
.B2(n_79),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_133),
.A2(n_41),
.B1(n_21),
.B2(n_31),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g244 ( 
.A1(n_210),
.A2(n_231),
.B1(n_125),
.B2(n_204),
.Y(n_244)
);

INVx3_ASAP7_75t_L g211 ( 
.A(n_162),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_211),
.Y(n_232)
);

AND2x2_ASAP7_75t_L g212 ( 
.A(n_161),
.B(n_85),
.Y(n_212)
);

HB1xp67_ASAP7_75t_L g213 ( 
.A(n_145),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g234 ( 
.A(n_213),
.Y(n_234)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_128),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_214),
.B(n_216),
.Y(n_257)
);

INVx3_ASAP7_75t_L g215 ( 
.A(n_162),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_215),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_139),
.B(n_65),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_148),
.B(n_31),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_217),
.B(n_218),
.Y(n_261)
);

INVx2_ASAP7_75t_L g218 ( 
.A(n_160),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_106),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_219),
.B(n_222),
.Y(n_262)
);

O2A1O1Ixp33_ASAP7_75t_L g220 ( 
.A1(n_147),
.A2(n_52),
.B(n_65),
.C(n_31),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g221 ( 
.A(n_108),
.B(n_31),
.Y(n_221)
);

NAND2xp33_ASAP7_75t_SL g285 ( 
.A(n_221),
.B(n_34),
.Y(n_285)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_115),
.Y(n_222)
);

BUFx2_ASAP7_75t_L g223 ( 
.A(n_117),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_223),
.B(n_224),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_145),
.B(n_52),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_163),
.B(n_14),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_225),
.B(n_228),
.Y(n_243)
);

INVx2_ASAP7_75t_L g226 ( 
.A(n_115),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_226),
.B(n_227),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_163),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_108),
.B(n_14),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_229),
.B(n_230),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_125),
.B(n_24),
.Y(n_230)
);

INVx6_ASAP7_75t_L g231 ( 
.A(n_149),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_233),
.B(n_9),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_178),
.B(n_165),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_239),
.B(n_264),
.Y(n_307)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_244),
.Y(n_302)
);

AOI32xp33_ASAP7_75t_L g248 ( 
.A1(n_172),
.A2(n_112),
.A3(n_123),
.B1(n_131),
.B2(n_150),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_248),
.A2(n_279),
.B(n_285),
.Y(n_297)
);

CKINVDCx20_ASAP7_75t_R g249 ( 
.A(n_185),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_249),
.B(n_270),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_171),
.B(n_165),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_252),
.B(n_274),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_254),
.A2(n_269),
.B1(n_283),
.B2(n_34),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_258),
.A2(n_231),
.B1(n_207),
.B2(n_192),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_197),
.B(n_158),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_268),
.A2(n_199),
.B1(n_194),
.B2(n_190),
.Y(n_290)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_209),
.A2(n_177),
.B1(n_181),
.B2(n_203),
.Y(n_269)
);

OAI32xp33_ASAP7_75t_L g270 ( 
.A1(n_173),
.A2(n_158),
.A3(n_109),
.B1(n_105),
.B2(n_152),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_221),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_2),
.Y(n_330)
);

AOI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_220),
.A2(n_135),
.B1(n_141),
.B2(n_152),
.Y(n_277)
);

INVxp67_ASAP7_75t_L g308 ( 
.A(n_277),
.Y(n_308)
);

AOI32xp33_ASAP7_75t_L g279 ( 
.A1(n_173),
.A2(n_109),
.A3(n_40),
.B1(n_36),
.B2(n_34),
.Y(n_279)
);

AOI22xp33_ASAP7_75t_L g283 ( 
.A1(n_179),
.A2(n_169),
.B1(n_154),
.B2(n_36),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_173),
.B(n_0),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g310 ( 
.A(n_284),
.B(n_0),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_286),
.B(n_334),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_287),
.B(n_299),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_SL g288 ( 
.A1(n_276),
.A2(n_179),
.B1(n_212),
.B2(n_223),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g350 ( 
.A1(n_288),
.A2(n_317),
.B(n_330),
.Y(n_350)
);

INVx2_ASAP7_75t_L g289 ( 
.A(n_247),
.Y(n_289)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_289),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g339 ( 
.A1(n_290),
.A2(n_294),
.B1(n_300),
.B2(n_278),
.Y(n_339)
);

INVx2_ASAP7_75t_L g291 ( 
.A(n_247),
.Y(n_291)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_291),
.Y(n_338)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_265),
.Y(n_292)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_292),
.Y(n_372)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_281),
.Y(n_293)
);

AOI22xp33_ASAP7_75t_SL g355 ( 
.A1(n_293),
.A2(n_329),
.B1(n_331),
.B2(n_266),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g295 ( 
.A1(n_276),
.A2(n_195),
.B1(n_186),
.B2(n_187),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_295),
.A2(n_296),
.B1(n_298),
.B2(n_305),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g296 ( 
.A1(n_252),
.A2(n_218),
.B1(n_175),
.B2(n_202),
.Y(n_296)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_262),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_274),
.A2(n_212),
.B1(n_221),
.B2(n_188),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

INVx2_ASAP7_75t_SL g336 ( 
.A(n_301),
.Y(n_336)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_241),
.B(n_191),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g361 ( 
.A(n_303),
.B(n_320),
.C(n_321),
.Y(n_361)
);

CKINVDCx14_ASAP7_75t_R g304 ( 
.A(n_236),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_304),
.B(n_306),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g305 ( 
.A1(n_248),
.A2(n_200),
.B1(n_193),
.B2(n_226),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_237),
.Y(n_306)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_238),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g349 ( 
.A(n_309),
.B(n_310),
.Y(n_349)
);

INVx8_ASAP7_75t_L g311 ( 
.A(n_281),
.Y(n_311)
);

INVx4_ASAP7_75t_L g341 ( 
.A(n_311),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_233),
.B(n_183),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_312),
.B(n_315),
.Y(n_352)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_246),
.A2(n_206),
.B(n_182),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g345 ( 
.A1(n_313),
.A2(n_314),
.B(n_273),
.Y(n_345)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_246),
.A2(n_215),
.B(n_211),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g315 ( 
.A(n_281),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g316 ( 
.A(n_243),
.B(n_222),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_316),
.B(n_318),
.Y(n_363)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_236),
.B(n_189),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_259),
.Y(n_318)
);

OAI21xp5_ASAP7_75t_SL g319 ( 
.A1(n_256),
.A2(n_174),
.B(n_184),
.Y(n_319)
);

OR2x2_ASAP7_75t_L g365 ( 
.A(n_319),
.B(n_324),
.Y(n_365)
);

MAJx2_ASAP7_75t_L g320 ( 
.A(n_241),
.B(n_9),
.C(n_18),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_239),
.B(n_34),
.C(n_2),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g322 ( 
.A(n_281),
.Y(n_322)
);

CKINVDCx16_ASAP7_75t_R g368 ( 
.A(n_322),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_236),
.Y(n_323)
);

CKINVDCx16_ASAP7_75t_R g375 ( 
.A(n_323),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_240),
.B(n_8),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_263),
.Y(n_325)
);

NAND2xp5_ASAP7_75t_L g367 ( 
.A(n_325),
.B(n_333),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g326 ( 
.A1(n_284),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_326)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_326),
.A2(n_255),
.B1(n_238),
.B2(n_235),
.Y(n_356)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_243),
.B(n_11),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g369 ( 
.A(n_327),
.B(n_332),
.C(n_235),
.Y(n_369)
);

AOI22xp33_ASAP7_75t_SL g329 ( 
.A1(n_268),
.A2(n_11),
.B1(n_17),
.B2(n_16),
.Y(n_329)
);

INVx8_ASAP7_75t_L g331 ( 
.A(n_280),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_264),
.B(n_7),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_251),
.B(n_7),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_261),
.B(n_2),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_339),
.A2(n_315),
.B1(n_321),
.B2(n_299),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_328),
.A2(n_279),
.B1(n_275),
.B2(n_268),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_340),
.A2(n_346),
.B1(n_347),
.B2(n_351),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g342 ( 
.A(n_297),
.B(n_286),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_342),
.B(n_343),
.Y(n_402)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_334),
.Y(n_343)
);

INVxp67_ASAP7_75t_L g388 ( 
.A(n_345),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_SL g346 ( 
.A1(n_328),
.A2(n_268),
.B1(n_270),
.B2(n_251),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_297),
.A2(n_268),
.B1(n_272),
.B2(n_242),
.Y(n_347)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_307),
.A2(n_240),
.B1(n_258),
.B2(n_257),
.Y(n_351)
);

CKINVDCx20_ASAP7_75t_R g353 ( 
.A(n_317),
.Y(n_353)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_353),
.B(n_369),
.Y(n_404)
);

AO21x1_ASAP7_75t_L g354 ( 
.A1(n_305),
.A2(n_285),
.B(n_259),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_354),
.A2(n_355),
.B(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_SL g413 ( 
.A(n_356),
.B(n_3),
.Y(n_413)
);

OAI22xp5_ASAP7_75t_L g357 ( 
.A1(n_307),
.A2(n_249),
.B1(n_232),
.B2(n_245),
.Y(n_357)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_357),
.B(n_360),
.Y(n_389)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_304),
.A2(n_234),
.B(n_245),
.Y(n_358)
);

INVx8_ASAP7_75t_L g359 ( 
.A(n_322),
.Y(n_359)
);

INVx2_ASAP7_75t_L g408 ( 
.A(n_359),
.Y(n_408)
);

OAI22xp5_ASAP7_75t_L g360 ( 
.A1(n_308),
.A2(n_232),
.B1(n_255),
.B2(n_271),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_L g362 ( 
.A1(n_313),
.A2(n_302),
.B(n_292),
.Y(n_362)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_362),
.A2(n_366),
.B(n_377),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_L g364 ( 
.A1(n_295),
.A2(n_255),
.B1(n_280),
.B2(n_260),
.Y(n_364)
);

AOI22xp33_ASAP7_75t_L g381 ( 
.A1(n_364),
.A2(n_368),
.B1(n_296),
.B2(n_315),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_317),
.A2(n_260),
.B1(n_280),
.B2(n_273),
.Y(n_366)
);

AOI22xp5_ASAP7_75t_L g370 ( 
.A1(n_298),
.A2(n_271),
.B1(n_253),
.B2(n_234),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g384 ( 
.A1(n_370),
.A2(n_344),
.B1(n_354),
.B2(n_374),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g373 ( 
.A1(n_288),
.A2(n_282),
.B(n_267),
.Y(n_373)
);

AOI21xp5_ASAP7_75t_L g395 ( 
.A1(n_373),
.A2(n_309),
.B(n_301),
.Y(n_395)
);

AO21x2_ASAP7_75t_L g374 ( 
.A1(n_314),
.A2(n_282),
.B(n_253),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g383 ( 
.A1(n_374),
.A2(n_294),
.B1(n_300),
.B2(n_306),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_303),
.B(n_267),
.C(n_250),
.Y(n_376)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_376),
.B(n_375),
.C(n_361),
.Y(n_382)
);

OAI21xp5_ASAP7_75t_L g377 ( 
.A1(n_319),
.A2(n_266),
.B(n_250),
.Y(n_377)
);

XNOR2xp5_ASAP7_75t_L g379 ( 
.A(n_361),
.B(n_316),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_379),
.B(n_382),
.C(n_392),
.Y(n_415)
);

NAND2xp5_ASAP7_75t_L g426 ( 
.A(n_381),
.B(n_385),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g420 ( 
.A1(n_383),
.A2(n_384),
.B1(n_400),
.B2(n_405),
.Y(n_420)
);

CKINVDCx20_ASAP7_75t_R g385 ( 
.A(n_357),
.Y(n_385)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_336),
.Y(n_386)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_386),
.Y(n_428)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_336),
.Y(n_387)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_387),
.Y(n_444)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_349),
.B(n_312),
.Y(n_390)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_390),
.Y(n_416)
);

A2O1A1Ixp33_ASAP7_75t_L g391 ( 
.A1(n_365),
.A2(n_330),
.B(n_333),
.C(n_310),
.Y(n_391)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_391),
.A2(n_366),
.B(n_356),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_376),
.B(n_348),
.C(n_353),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_393),
.A2(n_413),
.B1(n_395),
.B2(n_378),
.Y(n_441)
);

CKINVDCx20_ASAP7_75t_R g394 ( 
.A(n_352),
.Y(n_394)
);

CKINVDCx14_ASAP7_75t_R g438 ( 
.A(n_394),
.Y(n_438)
);

OAI21xp5_ASAP7_75t_SL g431 ( 
.A1(n_395),
.A2(n_396),
.B(n_414),
.Y(n_431)
);

AND2x2_ASAP7_75t_L g396 ( 
.A(n_345),
.B(n_318),
.Y(n_396)
);

MAJx2_ASAP7_75t_L g397 ( 
.A(n_348),
.B(n_320),
.C(n_327),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_397),
.B(n_350),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_SL g398 ( 
.A(n_369),
.B(n_332),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_398),
.B(n_351),
.Y(n_424)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_362),
.A2(n_291),
.B(n_289),
.Y(n_399)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_399),
.A2(n_365),
.B(n_352),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_L g400 ( 
.A1(n_344),
.A2(n_253),
.B1(n_287),
.B2(n_331),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_350),
.B(n_320),
.Y(n_401)
);

MAJIxp5_ASAP7_75t_L g421 ( 
.A(n_401),
.B(n_372),
.C(n_343),
.Y(n_421)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_349),
.B(n_326),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_403),
.Y(n_425)
);

OAI22xp5_ASAP7_75t_L g405 ( 
.A1(n_354),
.A2(n_331),
.B1(n_324),
.B2(n_311),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g406 ( 
.A(n_372),
.B(n_311),
.Y(n_406)
);

NAND3xp33_ASAP7_75t_L g436 ( 
.A(n_406),
.B(n_407),
.C(n_411),
.Y(n_436)
);

NAND3xp33_ASAP7_75t_L g407 ( 
.A(n_335),
.B(n_12),
.C(n_16),
.Y(n_407)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_374),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g433 ( 
.A1(n_409),
.A2(n_360),
.B1(n_339),
.B2(n_338),
.Y(n_433)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_336),
.Y(n_410)
);

CKINVDCx20_ASAP7_75t_R g442 ( 
.A(n_410),
.Y(n_442)
);

NAND3xp33_ASAP7_75t_L g411 ( 
.A(n_335),
.B(n_13),
.C(n_5),
.Y(n_411)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_358),
.A2(n_13),
.B(n_5),
.Y(n_414)
);

AOI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_384),
.A2(n_346),
.B1(n_340),
.B2(n_347),
.Y(n_417)
);

OAI22xp5_ASAP7_75t_L g469 ( 
.A1(n_417),
.A2(n_433),
.B1(n_439),
.B2(n_414),
.Y(n_469)
);

XNOR2xp5_ASAP7_75t_SL g458 ( 
.A(n_418),
.B(n_424),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_379),
.B(n_371),
.Y(n_419)
);

XOR2xp5_ASAP7_75t_L g449 ( 
.A(n_419),
.B(n_423),
.Y(n_449)
);

MAJIxp5_ASAP7_75t_L g451 ( 
.A(n_421),
.B(n_434),
.C(n_445),
.Y(n_451)
);

AO22x1_ASAP7_75t_L g422 ( 
.A1(n_388),
.A2(n_374),
.B1(n_377),
.B2(n_342),
.Y(n_422)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_422),
.Y(n_456)
);

XNOR2xp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_371),
.Y(n_423)
);

CKINVDCx16_ASAP7_75t_R g427 ( 
.A(n_396),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_L g465 ( 
.A(n_427),
.B(n_441),
.Y(n_465)
);

AOI21x1_ASAP7_75t_L g470 ( 
.A1(n_429),
.A2(n_435),
.B(n_413),
.Y(n_470)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_382),
.B(n_363),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g461 ( 
.A(n_430),
.B(n_432),
.Y(n_461)
);

XNOR2xp5_ASAP7_75t_SL g432 ( 
.A(n_401),
.B(n_367),
.Y(n_432)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_398),
.B(n_375),
.C(n_363),
.Y(n_434)
);

OAI21xp5_ASAP7_75t_L g435 ( 
.A1(n_388),
.A2(n_365),
.B(n_373),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_385),
.A2(n_374),
.B1(n_367),
.B2(n_370),
.Y(n_437)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_437),
.A2(n_389),
.B1(n_380),
.B2(n_394),
.Y(n_450)
);

XNOR2xp5_ASAP7_75t_SL g440 ( 
.A(n_412),
.B(n_374),
.Y(n_440)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_440),
.B(n_378),
.Y(n_452)
);

OAI22xp5_ASAP7_75t_SL g443 ( 
.A1(n_412),
.A2(n_338),
.B1(n_337),
.B2(n_359),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_443),
.B(n_446),
.Y(n_460)
);

MAJIxp5_ASAP7_75t_L g445 ( 
.A(n_404),
.B(n_337),
.C(n_368),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_393),
.A2(n_359),
.B1(n_341),
.B2(n_3),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_397),
.B(n_396),
.C(n_390),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_447),
.B(n_399),
.C(n_397),
.Y(n_454)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_428),
.Y(n_448)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_448),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g476 ( 
.A1(n_450),
.A2(n_457),
.B1(n_468),
.B2(n_469),
.Y(n_476)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_452),
.B(n_470),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_429),
.Y(n_453)
);

NAND2xp5_ASAP7_75t_L g496 ( 
.A(n_453),
.B(n_459),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_454),
.B(n_425),
.C(n_431),
.Y(n_489)
);

INVx1_ASAP7_75t_L g455 ( 
.A(n_444),
.Y(n_455)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_455),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_420),
.A2(n_402),
.B1(n_380),
.B2(n_389),
.Y(n_457)
);

AND2x2_ASAP7_75t_L g459 ( 
.A(n_437),
.B(n_383),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_443),
.Y(n_462)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_462),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_442),
.B(n_387),
.Y(n_463)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_463),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g464 ( 
.A(n_415),
.B(n_403),
.C(n_410),
.Y(n_464)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_464),
.B(n_419),
.C(n_447),
.Y(n_479)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_426),
.Y(n_466)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_466),
.Y(n_498)
);

INVx1_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_L g495 ( 
.A1(n_467),
.A2(n_471),
.B1(n_341),
.B2(n_422),
.Y(n_495)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_440),
.Y(n_468)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_438),
.Y(n_471)
);

NOR2xp33_ASAP7_75t_L g472 ( 
.A(n_430),
.B(n_408),
.Y(n_472)
);

XNOR2xp5_ASAP7_75t_L g493 ( 
.A(n_472),
.B(n_473),
.Y(n_493)
);

HB1xp67_ASAP7_75t_L g473 ( 
.A(n_423),
.Y(n_473)
);

XNOR2xp5_ASAP7_75t_L g474 ( 
.A(n_415),
.B(n_405),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g494 ( 
.A(n_474),
.B(n_475),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_416),
.B(n_386),
.Y(n_475)
);

XNOR2xp5_ASAP7_75t_L g512 ( 
.A(n_479),
.B(n_487),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g480 ( 
.A1(n_457),
.A2(n_400),
.B1(n_441),
.B2(n_446),
.Y(n_480)
);

OAI22xp5_ASAP7_75t_L g506 ( 
.A1(n_480),
.A2(n_482),
.B1(n_460),
.B2(n_433),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_451),
.B(n_434),
.C(n_421),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_481),
.B(n_483),
.C(n_485),
.Y(n_501)
);

NOR3xp33_ASAP7_75t_SL g482 ( 
.A(n_456),
.B(n_391),
.C(n_436),
.Y(n_482)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_451),
.B(n_424),
.C(n_432),
.Y(n_483)
);

MAJIxp5_ASAP7_75t_L g485 ( 
.A(n_464),
.B(n_418),
.C(n_435),
.Y(n_485)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_458),
.B(n_420),
.Y(n_487)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_449),
.B(n_439),
.C(n_417),
.Y(n_488)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_488),
.B(n_491),
.C(n_492),
.Y(n_505)
);

OAI21xp5_ASAP7_75t_L g514 ( 
.A1(n_489),
.A2(n_470),
.B(n_448),
.Y(n_514)
);

BUFx24_ASAP7_75t_SL g490 ( 
.A(n_474),
.Y(n_490)
);

BUFx24_ASAP7_75t_SL g509 ( 
.A(n_490),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g491 ( 
.A(n_449),
.B(n_431),
.C(n_408),
.Y(n_491)
);

MAJIxp5_ASAP7_75t_L g492 ( 
.A(n_454),
.B(n_461),
.C(n_458),
.Y(n_492)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_495),
.Y(n_511)
);

XOR2xp5_ASAP7_75t_L g499 ( 
.A(n_491),
.B(n_452),
.Y(n_499)
);

XNOR2xp5_ASAP7_75t_L g522 ( 
.A(n_499),
.B(n_504),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_SL g500 ( 
.A1(n_496),
.A2(n_456),
.B(n_468),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_500),
.A2(n_12),
.B(n_16),
.Y(n_531)
);

BUFx6f_ASAP7_75t_L g502 ( 
.A(n_498),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_502),
.B(n_507),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g503 ( 
.A1(n_484),
.A2(n_465),
.B(n_475),
.Y(n_503)
);

OAI21xp5_ASAP7_75t_SL g519 ( 
.A1(n_503),
.A2(n_477),
.B(n_476),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g504 ( 
.A(n_494),
.B(n_461),
.Y(n_504)
);

AOI22xp5_ASAP7_75t_L g520 ( 
.A1(n_506),
.A2(n_409),
.B1(n_484),
.B2(n_482),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g507 ( 
.A(n_479),
.B(n_481),
.C(n_494),
.Y(n_507)
);

XNOR2xp5_ASAP7_75t_L g508 ( 
.A(n_493),
.B(n_422),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g526 ( 
.A(n_508),
.B(n_516),
.Y(n_526)
);

NOR2xp33_ASAP7_75t_L g510 ( 
.A(n_486),
.B(n_450),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_L g524 ( 
.A(n_510),
.B(n_515),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_SL g513 ( 
.A(n_478),
.B(n_463),
.Y(n_513)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_513),
.B(n_497),
.Y(n_517)
);

AOI21xp33_ASAP7_75t_L g530 ( 
.A1(n_514),
.A2(n_12),
.B(n_15),
.Y(n_530)
);

MAJIxp5_ASAP7_75t_L g515 ( 
.A(n_485),
.B(n_459),
.C(n_460),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_L g516 ( 
.A(n_488),
.B(n_459),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_517),
.B(n_521),
.Y(n_532)
);

AND2x2_ASAP7_75t_L g542 ( 
.A(n_519),
.B(n_520),
.Y(n_542)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_507),
.B(n_492),
.C(n_483),
.Y(n_521)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_515),
.B(n_487),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_523),
.B(n_525),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_502),
.B(n_13),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_501),
.B(n_5),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g536 ( 
.A(n_527),
.B(n_528),
.Y(n_536)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_501),
.B(n_3),
.C(n_6),
.Y(n_528)
);

XOR2xp5_ASAP7_75t_L g529 ( 
.A(n_499),
.B(n_6),
.Y(n_529)
);

XNOR2xp5_ASAP7_75t_L g537 ( 
.A(n_529),
.B(n_531),
.Y(n_537)
);

NOR2xp33_ASAP7_75t_SL g533 ( 
.A(n_530),
.B(n_18),
.Y(n_533)
);

NOR2xp33_ASAP7_75t_L g546 ( 
.A(n_533),
.B(n_535),
.Y(n_546)
);

NOR2xp33_ASAP7_75t_L g534 ( 
.A(n_518),
.B(n_511),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g545 ( 
.A(n_534),
.B(n_538),
.Y(n_545)
);

NOR2xp33_ASAP7_75t_SL g535 ( 
.A(n_521),
.B(n_509),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g538 ( 
.A(n_522),
.B(n_512),
.Y(n_538)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_524),
.B(n_505),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g547 ( 
.A(n_540),
.B(n_522),
.Y(n_547)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_519),
.B(n_500),
.Y(n_541)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_541),
.B(n_508),
.Y(n_549)
);

AOI22xp5_ASAP7_75t_SL g543 ( 
.A1(n_542),
.A2(n_505),
.B1(n_520),
.B2(n_528),
.Y(n_543)
);

NAND2xp5_ASAP7_75t_L g550 ( 
.A(n_543),
.B(n_544),
.Y(n_550)
);

OAI21xp5_ASAP7_75t_SL g544 ( 
.A1(n_532),
.A2(n_541),
.B(n_542),
.Y(n_544)
);

INVx1_ASAP7_75t_L g552 ( 
.A(n_547),
.Y(n_552)
);

AND2x2_ASAP7_75t_L g548 ( 
.A(n_539),
.B(n_516),
.Y(n_548)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_548),
.B(n_526),
.C(n_529),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g551 ( 
.A(n_549),
.Y(n_551)
);

AOI21xp5_ASAP7_75t_L g554 ( 
.A1(n_553),
.A2(n_545),
.B(n_549),
.Y(n_554)
);

AOI21x1_ASAP7_75t_L g557 ( 
.A1(n_554),
.A2(n_555),
.B(n_546),
.Y(n_557)
);

INVxp67_ASAP7_75t_L g555 ( 
.A(n_550),
.Y(n_555)
);

AO21x2_ASAP7_75t_SL g556 ( 
.A1(n_555),
.A2(n_551),
.B(n_552),
.Y(n_556)
);

OAI21xp5_ASAP7_75t_L g558 ( 
.A1(n_556),
.A2(n_557),
.B(n_531),
.Y(n_558)
);

MAJIxp5_ASAP7_75t_L g559 ( 
.A(n_558),
.B(n_537),
.C(n_536),
.Y(n_559)
);

NAND2xp5_ASAP7_75t_L g560 ( 
.A(n_559),
.B(n_526),
.Y(n_560)
);

NOR2xp33_ASAP7_75t_L g561 ( 
.A(n_560),
.B(n_504),
.Y(n_561)
);


endmodule