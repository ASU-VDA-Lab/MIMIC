module real_jpeg_23710_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_215;
wire n_176;
wire n_312;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_0),
.Y(n_65)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_1),
.A2(n_27),
.B1(n_28),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

AOI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_1),
.A2(n_35),
.B1(n_40),
.B2(n_42),
.Y(n_92)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g159 ( 
.A(n_3),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_3),
.B(n_63),
.Y(n_177)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_3),
.A2(n_67),
.B(n_83),
.C(n_219),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_3),
.A2(n_64),
.B1(n_67),
.B2(n_159),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g240 ( 
.A(n_3),
.B(n_28),
.C(n_45),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_L g243 ( 
.A1(n_3),
.A2(n_40),
.B1(n_42),
.B2(n_159),
.Y(n_243)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_3),
.A2(n_25),
.B(n_254),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_3),
.B(n_125),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_5),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_56)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_5),
.A2(n_61),
.B1(n_64),
.B2(n_67),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_5),
.A2(n_40),
.B1(n_42),
.B2(n_61),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g179 ( 
.A1(n_5),
.A2(n_27),
.B1(n_28),
.B2(n_61),
.Y(n_179)
);

INVx8_ASAP7_75t_SL g66 ( 
.A(n_6),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_7),
.A2(n_60),
.B1(n_72),
.B2(n_110),
.Y(n_109)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_7),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_7),
.A2(n_64),
.B1(n_67),
.B2(n_110),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_7),
.A2(n_40),
.B1(n_42),
.B2(n_110),
.Y(n_214)
);

AOI22xp33_ASAP7_75t_L g248 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_110),
.Y(n_248)
);

BUFx5_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

INVx13_ASAP7_75t_L g59 ( 
.A(n_9),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g71 ( 
.A1(n_10),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_10),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_10),
.A2(n_40),
.B1(n_42),
.B2(n_74),
.Y(n_155)
);

OAI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_10),
.A2(n_64),
.B1(n_67),
.B2(n_74),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_10),
.A2(n_27),
.B1(n_28),
.B2(n_74),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_11),
.A2(n_40),
.B1(n_42),
.B2(n_50),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_11),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_11),
.A2(n_27),
.B1(n_28),
.B2(n_50),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_11),
.A2(n_50),
.B1(n_64),
.B2(n_67),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_12),
.A2(n_64),
.B1(n_67),
.B2(n_87),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g87 ( 
.A(n_12),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g104 ( 
.A1(n_12),
.A2(n_40),
.B1(n_42),
.B2(n_87),
.Y(n_104)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_12),
.A2(n_60),
.B1(n_87),
.B2(n_134),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_12),
.A2(n_27),
.B1(n_28),
.B2(n_87),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_13),
.A2(n_64),
.B1(n_67),
.B2(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g149 ( 
.A(n_13),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_13),
.A2(n_59),
.B1(n_60),
.B2(n_149),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g229 ( 
.A1(n_13),
.A2(n_40),
.B1(n_42),
.B2(n_149),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_13),
.A2(n_27),
.B1(n_28),
.B2(n_149),
.Y(n_246)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_14),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_15),
.A2(n_39),
.B1(n_40),
.B2(n_42),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_15),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g88 ( 
.A1(n_15),
.A2(n_39),
.B1(n_64),
.B2(n_67),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_15),
.A2(n_27),
.B1(n_28),
.B2(n_39),
.Y(n_167)
);

INVx6_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_16),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_16),
.A2(n_26),
.B1(n_165),
.B2(n_167),
.Y(n_164)
);

INVx6_ASAP7_75t_L g182 ( 
.A(n_16),
.Y(n_182)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_16),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_16),
.A2(n_26),
.B1(n_245),
.B2(n_247),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_136),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_114),
.Y(n_20)
);

AND2x2_ASAP7_75t_L g137 ( 
.A(n_21),
.B(n_114),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_78),
.C(n_94),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g314 ( 
.A1(n_22),
.A2(n_78),
.B1(n_79),
.B2(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_22),
.Y(n_315)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_52),
.Y(n_22)
);

AOI21xp33_ASAP7_75t_L g115 ( 
.A1(n_23),
.A2(n_24),
.B(n_54),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_36),
.Y(n_23)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_24),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_24),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_24),
.A2(n_36),
.B1(n_37),
.B2(n_53),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_32),
.B(n_34),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_25),
.A2(n_34),
.B1(n_99),
.B2(n_100),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_25),
.A2(n_166),
.B1(n_179),
.B2(n_180),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_25),
.A2(n_31),
.B1(n_99),
.B2(n_196),
.Y(n_195)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_25),
.A2(n_248),
.B(n_254),
.Y(n_268)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_26),
.B(n_223),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_27),
.B(n_30),
.Y(n_26)
);

OA22x2_ASAP7_75t_L g48 ( 
.A1(n_27),
.A2(n_28),
.B1(n_45),
.B2(n_47),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_27),
.B(n_252),
.Y(n_251)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx5_ASAP7_75t_L g33 ( 
.A(n_31),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g252 ( 
.A(n_32),
.B(n_159),
.Y(n_252)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_43),
.B1(n_49),
.B2(n_51),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_38),
.A2(n_43),
.B1(n_51),
.B2(n_103),
.Y(n_102)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_40),
.Y(n_42)
);

OAI22xp33_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_42),
.B1(n_45),
.B2(n_47),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_SL g82 ( 
.A1(n_40),
.A2(n_42),
.B1(n_83),
.B2(n_84),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_40),
.B(n_240),
.Y(n_239)
);

BUFx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_42),
.A2(n_84),
.B(n_159),
.Y(n_219)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_43),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g129 ( 
.A1(n_43),
.A2(n_51),
.B(n_130),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_43),
.B(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_43),
.A2(n_51),
.B1(n_214),
.B2(n_228),
.Y(n_227)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_48),
.Y(n_43)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_45),
.Y(n_47)
);

BUFx24_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_48),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_48),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_48),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_48),
.A2(n_90),
.B1(n_104),
.B2(n_153),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_48),
.B(n_159),
.Y(n_258)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_48),
.A2(n_154),
.B(n_229),
.Y(n_267)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_51),
.B(n_155),
.Y(n_215)
);

CKINVDCx14_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_L g55 ( 
.A1(n_56),
.A2(n_62),
.B(n_69),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_56),
.A2(n_62),
.B1(n_111),
.B2(n_133),
.Y(n_132)
);

INVx8_ASAP7_75t_L g158 ( 
.A(n_57),
.Y(n_158)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

NAND3xp33_ASAP7_75t_SL g170 ( 
.A(n_58),
.B(n_66),
.C(n_67),
.Y(n_170)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g60 ( 
.A(n_59),
.Y(n_60)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_59),
.Y(n_75)
);

INVx11_ASAP7_75t_L g134 ( 
.A(n_60),
.Y(n_134)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_62),
.B(n_77),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g113 ( 
.A(n_62),
.B(n_71),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_62),
.A2(n_69),
.B(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_63),
.A2(n_76),
.B1(n_109),
.B2(n_191),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B1(n_67),
.B2(n_68),
.Y(n_63)
);

INVx5_ASAP7_75t_L g67 ( 
.A(n_64),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g85 ( 
.A1(n_64),
.A2(n_67),
.B1(n_83),
.B2(n_84),
.Y(n_85)
);

A2O1A1Ixp33_ASAP7_75t_L g169 ( 
.A1(n_64),
.A2(n_68),
.B(n_160),
.C(n_170),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_66),
.Y(n_68)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_66),
.A2(n_68),
.B1(n_72),
.B2(n_75),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_70),
.B(n_76),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

INVx8_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_73),
.B(n_159),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_76),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g156 ( 
.A1(n_76),
.A2(n_113),
.B(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_89),
.B(n_93),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_80),
.B(n_89),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_88),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_82),
.B1(n_86),
.B2(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_81),
.Y(n_124)
);

OAI21xp5_ASAP7_75t_SL g186 ( 
.A1(n_81),
.A2(n_187),
.B(n_188),
.Y(n_186)
);

OAI21xp33_ASAP7_75t_L g231 ( 
.A1(n_81),
.A2(n_188),
.B(n_232),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_85),
.Y(n_81)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_82),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_82),
.A2(n_173),
.B(n_174),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_82),
.A2(n_106),
.B(n_174),
.Y(n_298)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_83),
.Y(n_84)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_88),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_90),
.A2(n_213),
.B(n_215),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_90),
.A2(n_215),
.B(n_243),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g130 ( 
.A(n_92),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_93),
.A2(n_117),
.B1(n_118),
.B2(n_119),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g117 ( 
.A(n_93),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_94),
.A2(n_95),
.B1(n_314),
.B2(n_316),
.Y(n_313)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_105),
.C(n_107),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g307 ( 
.A1(n_96),
.A2(n_97),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g290 ( 
.A1(n_98),
.A2(n_101),
.B1(n_102),
.B2(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g291 ( 
.A(n_98),
.Y(n_291)
);

INVx3_ASAP7_75t_L g255 ( 
.A(n_100),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g257 ( 
.A1(n_100),
.A2(n_222),
.B(n_246),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_105),
.B(n_107),
.Y(n_309)
);

OAI21xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_111),
.B(n_112),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g114 ( 
.A(n_115),
.B(n_116),
.Y(n_114)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_119),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_120),
.A2(n_121),
.B1(n_132),
.B2(n_135),
.Y(n_119)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_122),
.A2(n_128),
.B1(n_129),
.B2(n_131),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_122),
.Y(n_131)
);

AOI22xp5_ASAP7_75t_L g122 ( 
.A1(n_123),
.A2(n_124),
.B1(n_125),
.B2(n_126),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_124),
.A2(n_125),
.B1(n_148),
.B2(n_150),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_124),
.B(n_175),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_125),
.B(n_175),
.Y(n_188)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_132),
.Y(n_135)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_137),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_312),
.B(n_318),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_SL g139 ( 
.A1(n_140),
.A2(n_302),
.B(n_311),
.Y(n_139)
);

O2A1O1Ixp33_ASAP7_75t_SL g140 ( 
.A1(n_141),
.A2(n_200),
.B(n_285),
.C(n_301),
.Y(n_140)
);

AND2x2_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_183),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_142),
.B(n_183),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_161),
.C(n_171),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_143),
.A2(n_144),
.B1(n_280),
.B2(n_281),
.Y(n_279)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_156),
.Y(n_144)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_146),
.A2(n_147),
.B1(n_151),
.B2(n_152),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g198 ( 
.A(n_147),
.B(n_151),
.C(n_156),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g173 ( 
.A(n_148),
.Y(n_173)
);

CKINVDCx14_ASAP7_75t_R g187 ( 
.A(n_150),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

OAI21xp33_ASAP7_75t_L g157 ( 
.A1(n_158),
.A2(n_159),
.B(n_160),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g281 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g162 ( 
.A1(n_163),
.A2(n_164),
.B1(n_168),
.B2(n_169),
.Y(n_162)
);

CKINVDCx14_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_164),
.B(n_168),
.Y(n_185)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g196 ( 
.A(n_167),
.Y(n_196)
);

CKINVDCx14_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_171),
.Y(n_282)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_172),
.B(n_208),
.Y(n_207)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_176),
.A2(n_177),
.B1(n_178),
.B2(n_209),
.Y(n_208)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_178),
.Y(n_209)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_179),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g183 ( 
.A1(n_184),
.A2(n_192),
.B1(n_193),
.B2(n_199),
.Y(n_183)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_184),
.Y(n_199)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_184),
.Y(n_319)
);

FAx1_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.CI(n_189),
.CON(n_184),
.SN(n_184)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_185),
.B(n_186),
.C(n_189),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_198),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_194),
.B(n_198),
.C(n_199),
.Y(n_300)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_197),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_195),
.B(n_197),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

AOI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_278),
.B(n_284),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_L g203 ( 
.A1(n_204),
.A2(n_233),
.B(n_277),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_SL g204 ( 
.A(n_205),
.B(n_225),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_205),
.B(n_225),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_207),
.B1(n_210),
.B2(n_224),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g283 ( 
.A(n_206),
.B(n_212),
.C(n_216),
.Y(n_283)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_210),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_211),
.A2(n_212),
.B1(n_216),
.B2(n_217),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g226 ( 
.A(n_218),
.B(n_220),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_255),
.Y(n_254)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_226),
.B(n_227),
.C(n_230),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_226),
.B(n_273),
.Y(n_272)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_227),
.A2(n_230),
.B1(n_231),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_227),
.Y(n_274)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g233 ( 
.A1(n_234),
.A2(n_271),
.B(n_276),
.Y(n_233)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_235),
.A2(n_261),
.B(n_270),
.Y(n_234)
);

AOI21xp5_ASAP7_75t_L g235 ( 
.A1(n_236),
.A2(n_249),
.B(n_260),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g236 ( 
.A(n_237),
.B(n_244),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_237),
.B(n_244),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_238),
.A2(n_239),
.B1(n_241),
.B2(n_242),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_239),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_239),
.B(n_241),
.Y(n_269)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

CKINVDCx16_ASAP7_75t_R g245 ( 
.A(n_246),
.Y(n_245)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

OAI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_256),
.B(n_259),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_257),
.B(n_258),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_257),
.B(n_258),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_269),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_262),
.B(n_269),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_268),
.Y(n_262)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_264),
.A2(n_265),
.B1(n_266),
.B2(n_267),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_264),
.B(n_267),
.C(n_268),
.Y(n_275)
);

INVx1_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_272),
.B(n_275),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g278 ( 
.A(n_279),
.B(n_283),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_279),
.B(n_283),
.Y(n_284)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_286),
.B(n_300),
.Y(n_285)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_286),
.B(n_300),
.Y(n_301)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_288),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_287),
.B(n_290),
.C(n_292),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_290),
.B1(n_292),
.B2(n_293),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_299),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_296),
.B1(n_297),
.B2(n_298),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_296),
.B(n_297),
.C(n_299),
.Y(n_310)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g311 ( 
.A(n_303),
.B(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_310),
.Y(n_304)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_306),
.B(n_307),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_306),
.B(n_307),
.C(n_310),
.Y(n_317)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_SL g312 ( 
.A(n_313),
.B(n_317),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g318 ( 
.A(n_313),
.B(n_317),
.Y(n_318)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_314),
.Y(n_316)
);


endmodule