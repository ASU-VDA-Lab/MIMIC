module real_jpeg_19533_n_9 (n_5, n_4, n_8, n_0, n_1, n_2, n_6, n_7, n_3, n_9);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_2;
input n_6;
input n_7;
input n_3;

output n_9;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_10;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_11;
wire n_47;
wire n_22;
wire n_87;
wire n_40;
wire n_105;
wire n_98;
wire n_27;
wire n_56;
wire n_48;
wire n_13;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_106;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_109;
wire n_39;
wire n_94;
wire n_26;
wire n_19;
wire n_17;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_100;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_30;
wire n_15;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_12;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_25;
wire n_53;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;
wire n_16;

INVx13_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_1),
.A2(n_16),
.B1(n_17),
.B2(n_18),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_1),
.Y(n_16)
);

AOI22xp33_ASAP7_75t_SL g32 ( 
.A1(n_1),
.A2(n_16),
.B1(n_21),
.B2(n_22),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_1),
.A2(n_16),
.B1(n_35),
.B2(n_37),
.Y(n_65)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_2),
.Y(n_51)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_2),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_3),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

AOI22xp5_ASAP7_75t_L g26 ( 
.A1(n_5),
.A2(n_17),
.B1(n_18),
.B2(n_27),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_5),
.Y(n_27)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_5),
.A2(n_21),
.B1(n_22),
.B2(n_27),
.Y(n_39)
);

AOI21xp33_ASAP7_75t_SL g44 ( 
.A1(n_5),
.A2(n_22),
.B(n_23),
.Y(n_44)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_5),
.A2(n_27),
.B1(n_35),
.B2(n_37),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_5),
.B(n_60),
.Y(n_59)
);

AOI21xp33_ASAP7_75t_L g85 ( 
.A1(n_5),
.A2(n_7),
.B(n_37),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_6),
.A2(n_17),
.B1(n_18),
.B2(n_62),
.Y(n_61)
);

INVx13_ASAP7_75t_L g62 ( 
.A(n_6),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_SL g34 ( 
.A1(n_7),
.A2(n_35),
.B1(n_36),
.B2(n_37),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g36 ( 
.A(n_7),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_L g41 ( 
.A1(n_7),
.A2(n_21),
.B1(n_22),
.B2(n_36),
.Y(n_41)
);

BUFx3_ASAP7_75t_SL g22 ( 
.A(n_8),
.Y(n_22)
);

XNOR2xp5_ASAP7_75t_L g9 ( 
.A(n_10),
.B(n_78),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g10 ( 
.A(n_11),
.B(n_77),
.Y(n_10)
);

INVxp67_ASAP7_75t_L g11 ( 
.A(n_12),
.Y(n_11)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_54),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_13),
.B(n_54),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_30),
.C(n_42),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g108 ( 
.A1(n_14),
.A2(n_30),
.B1(n_86),
.B2(n_109),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_14),
.Y(n_109)
);

AOI21xp5_ASAP7_75t_L g14 ( 
.A1(n_15),
.A2(n_19),
.B(n_25),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_15),
.Y(n_71)
);

INVx4_ASAP7_75t_SL g18 ( 
.A(n_17),
.Y(n_18)
);

A2O1A1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_17),
.A2(n_24),
.B(n_27),
.C(n_44),
.Y(n_43)
);

A2O1A1Ixp33_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_20),
.B(n_23),
.C(n_29),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_18),
.B(n_23),
.Y(n_29)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_20),
.A2(n_26),
.B1(n_28),
.B2(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_20),
.B(n_27),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_23),
.B2(n_24),
.Y(n_20)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

A2O1A1Ixp33_ASAP7_75t_L g84 ( 
.A1(n_22),
.A2(n_27),
.B(n_36),
.C(n_85),
.Y(n_84)
);

INVx11_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_28),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g90 ( 
.A(n_27),
.B(n_51),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_27),
.B(n_34),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_30),
.A2(n_83),
.B1(n_84),
.B2(n_86),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_30),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g97 ( 
.A(n_30),
.B(n_84),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_33),
.B(n_38),
.Y(n_30)
);

INVxp67_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_32),
.A2(n_34),
.B1(n_39),
.B2(n_40),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_34),
.B(n_41),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_35),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_35),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_SL g50 ( 
.A(n_37),
.B(n_51),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

XOR2xp5_ASAP7_75t_L g107 ( 
.A(n_42),
.B(n_108),
.Y(n_107)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_53),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g53 ( 
.A(n_43),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_45),
.B(n_53),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g46 ( 
.A(n_47),
.B(n_49),
.Y(n_46)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_48),
.B(n_50),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_48),
.A2(n_50),
.B1(n_51),
.B2(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_SL g49 ( 
.A(n_50),
.B(n_52),
.Y(n_49)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_51),
.Y(n_66)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_72),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_57),
.B1(n_69),
.B2(n_70),
.Y(n_55)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_57),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_58),
.A2(n_59),
.B1(n_63),
.B2(n_68),
.Y(n_57)
);

CKINVDCx16_ASAP7_75t_R g58 ( 
.A(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g68 ( 
.A(n_63),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_63),
.B(n_82),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_63),
.B(n_82),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g63 ( 
.A1(n_64),
.A2(n_66),
.B(n_67),
.Y(n_63)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_65),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_68),
.B(n_89),
.Y(n_88)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_73),
.A2(n_74),
.B1(n_75),
.B2(n_76),
.Y(n_72)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_73),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_73),
.A2(n_75),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_73),
.B(n_92),
.C(n_101),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_74),
.Y(n_76)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_105),
.B(n_110),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_SL g79 ( 
.A1(n_80),
.A2(n_96),
.B(n_104),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g80 ( 
.A1(n_81),
.A2(n_87),
.B(n_95),
.Y(n_80)
);

CKINVDCx16_ASAP7_75t_R g83 ( 
.A(n_84),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_88),
.A2(n_91),
.B(n_94),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_92),
.B(n_93),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g98 ( 
.A1(n_92),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_92),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_98),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g104 ( 
.A(n_97),
.B(n_98),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_99),
.Y(n_103)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_107),
.Y(n_110)
);


endmodule