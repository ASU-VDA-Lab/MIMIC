module real_jpeg_3135_n_17 (n_8, n_0, n_82, n_2, n_10, n_9, n_12, n_83, n_6, n_11, n_14, n_7, n_3, n_5, n_4, n_81, n_1, n_16, n_15, n_13, n_17);

input n_8;
input n_0;
input n_82;
input n_2;
input n_10;
input n_9;
input n_12;
input n_83;
input n_6;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_81;
input n_1;
input n_16;
input n_15;
input n_13;

output n_17;

wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_49;
wire n_68;
wire n_78;
wire n_64;
wire n_47;
wire n_22;
wire n_40;
wire n_27;
wire n_56;
wire n_48;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_66;
wire n_44;
wire n_28;
wire n_62;
wire n_45;
wire n_42;
wire n_18;
wire n_77;
wire n_39;
wire n_26;
wire n_19;
wire n_21;
wire n_50;
wire n_69;
wire n_31;
wire n_72;
wire n_23;
wire n_51;
wire n_71;
wire n_61;
wire n_70;
wire n_41;
wire n_74;
wire n_32;
wire n_20;
wire n_30;
wire n_43;
wire n_57;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_24;
wire n_75;
wire n_34;
wire n_60;
wire n_46;
wire n_59;
wire n_25;
wire n_53;
wire n_36;

OAI22xp5_ASAP7_75t_L g21 ( 
.A1(n_0),
.A2(n_16),
.B1(n_22),
.B2(n_23),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g18 ( 
.A1(n_1),
.A2(n_19),
.B1(n_20),
.B2(n_48),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_1),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g65 ( 
.A1(n_1),
.A2(n_48),
.B1(n_66),
.B2(n_67),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_2),
.B(n_3),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_3),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_4),
.B(n_13),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_4),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_5),
.A2(n_50),
.B1(n_53),
.B2(n_64),
.Y(n_49)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_5),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_5),
.B(n_74),
.Y(n_73)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_6),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_7),
.B(n_81),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_8),
.B(n_10),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_8),
.B(n_10),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_9),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_11),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_12),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_14),
.B(n_35),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_16),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_14),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_15),
.B(n_82),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_15),
.B(n_83),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_16),
.B(n_35),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g41 ( 
.A1(n_16),
.A2(n_22),
.B1(n_42),
.B2(n_43),
.Y(n_41)
);

AOI21xp5_ASAP7_75t_L g44 ( 
.A1(n_16),
.A2(n_45),
.B(n_47),
.Y(n_44)
);

AOI221xp5_ASAP7_75t_L g17 ( 
.A1(n_18),
.A2(n_49),
.B1(n_65),
.B2(n_73),
.C(n_78),
.Y(n_17)
);

INVxp67_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_24),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_68),
.Y(n_67)
);

NOR3xp33_ASAP7_75t_L g37 ( 
.A(n_22),
.B(n_30),
.C(n_38),
.Y(n_37)
);

OAI211xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_33),
.B(n_36),
.C(n_44),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_26),
.Y(n_25)
);

OAI21xp5_ASAP7_75t_L g26 ( 
.A1(n_27),
.A2(n_28),
.B(n_29),
.Y(n_26)
);

AOI21xp33_ASAP7_75t_L g36 ( 
.A1(n_27),
.A2(n_37),
.B(n_41),
.Y(n_36)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_28),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g70 ( 
.A(n_28),
.B(n_71),
.Y(n_70)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI21xp5_ASAP7_75t_L g72 ( 
.A1(n_30),
.A2(n_34),
.B(n_41),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_31),
.B(n_32),
.Y(n_30)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

AOI22xp33_ASAP7_75t_L g69 ( 
.A1(n_34),
.A2(n_37),
.B1(n_70),
.B2(n_71),
.Y(n_69)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_38),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_38),
.B(n_46),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_SL g38 ( 
.A(n_39),
.B(n_40),
.Y(n_38)
);

NAND3xp33_ASAP7_75t_SL g68 ( 
.A(n_44),
.B(n_69),
.C(n_72),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g77 ( 
.A(n_50),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g50 ( 
.A(n_51),
.B(n_52),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g64 ( 
.A(n_51),
.B(n_52),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_55),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_54),
.B(n_79),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g75 ( 
.A1(n_55),
.A2(n_76),
.B(n_77),
.Y(n_75)
);

AOI21xp5_ASAP7_75t_SL g55 ( 
.A1(n_56),
.A2(n_60),
.B(n_63),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g56 ( 
.A1(n_57),
.A2(n_58),
.B(n_59),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_61),
.B(n_62),
.Y(n_63)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_64),
.Y(n_76)
);

INVxp67_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);


endmodule