module fake_netlist_1_2787_n_40 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_17;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
HB1xp67_ASAP7_75t_L g15 ( .A(n_4), .Y(n_15) );
CKINVDCx20_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
INVx2_ASAP7_75t_L g17 ( .A(n_14), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_7), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_10), .Y(n_19) );
AND2x2_ASAP7_75t_L g20 ( .A(n_9), .B(n_8), .Y(n_20) );
INVx2_ASAP7_75t_L g21 ( .A(n_1), .Y(n_21) );
CKINVDCx5p33_ASAP7_75t_R g22 ( .A(n_0), .Y(n_22) );
INVx3_ASAP7_75t_L g23 ( .A(n_21), .Y(n_23) );
INVx5_ASAP7_75t_L g24 ( .A(n_20), .Y(n_24) );
INVx2_ASAP7_75t_L g25 ( .A(n_17), .Y(n_25) );
AOI22xp33_ASAP7_75t_L g26 ( .A1(n_25), .A2(n_15), .B1(n_22), .B2(n_18), .Y(n_26) );
NAND2x1_ASAP7_75t_L g27 ( .A(n_25), .B(n_17), .Y(n_27) );
AOI221xp5_ASAP7_75t_L g28 ( .A1(n_26), .A2(n_23), .B1(n_16), .B2(n_15), .C(n_19), .Y(n_28) );
AND2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_23), .Y(n_29) );
NOR4xp25_ASAP7_75t_SL g30 ( .A(n_28), .B(n_0), .C(n_2), .D(n_3), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
BUFx2_ASAP7_75t_L g32 ( .A(n_29), .Y(n_32) );
OR2x2_ASAP7_75t_L g33 ( .A(n_32), .B(n_27), .Y(n_33) );
XNOR2x1_ASAP7_75t_L g34 ( .A(n_31), .B(n_2), .Y(n_34) );
OAI322xp33_ASAP7_75t_L g35 ( .A1(n_32), .A2(n_30), .A3(n_3), .B1(n_24), .B2(n_11), .C1(n_5), .C2(n_13), .Y(n_35) );
NOR2xp33_ASAP7_75t_L g36 ( .A(n_34), .B(n_24), .Y(n_36) );
HB1xp67_ASAP7_75t_L g37 ( .A(n_33), .Y(n_37) );
CKINVDCx12_ASAP7_75t_R g38 ( .A(n_35), .Y(n_38) );
BUFx3_ASAP7_75t_L g39 ( .A(n_36), .Y(n_39) );
AOI322xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_6), .A3(n_12), .B1(n_24), .B2(n_38), .C1(n_36), .C2(n_37), .Y(n_40) );
endmodule