module real_jpeg_3887_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_498;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_366;
wire n_328;
wire n_456;
wire n_259;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_372;
wire n_219;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_515;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_494;
wire n_512;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_169;
wire n_88;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

OAI22xp33_ASAP7_75t_L g147 ( 
.A1(n_0),
.A2(n_148),
.B1(n_149),
.B2(n_152),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_0),
.Y(n_148)
);

AOI22xp33_ASAP7_75t_L g296 ( 
.A1(n_0),
.A2(n_148),
.B1(n_213),
.B2(n_231),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g376 ( 
.A1(n_0),
.A2(n_101),
.B1(n_148),
.B2(n_377),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g410 ( 
.A1(n_0),
.A2(n_93),
.B1(n_148),
.B2(n_411),
.Y(n_410)
);

INVx8_ASAP7_75t_L g220 ( 
.A(n_1),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g226 ( 
.A(n_1),
.Y(n_226)
);

BUFx6f_ASAP7_75t_L g264 ( 
.A(n_1),
.Y(n_264)
);

INVx2_ASAP7_75t_L g330 ( 
.A(n_1),
.Y(n_330)
);

BUFx6f_ASAP7_75t_L g436 ( 
.A(n_1),
.Y(n_436)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_2),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_2),
.Y(n_50)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_2),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_2),
.Y(n_151)
);

BUFx5_ASAP7_75t_L g347 ( 
.A(n_2),
.Y(n_347)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_2),
.Y(n_362)
);

BUFx6f_ASAP7_75t_L g368 ( 
.A(n_2),
.Y(n_368)
);

AOI22xp33_ASAP7_75t_SL g86 ( 
.A1(n_3),
.A2(n_87),
.B1(n_89),
.B2(n_90),
.Y(n_86)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_3),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_3),
.A2(n_90),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

OAI22xp33_ASAP7_75t_SL g386 ( 
.A1(n_3),
.A2(n_90),
.B1(n_210),
.B2(n_387),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_3),
.A2(n_90),
.B1(n_421),
.B2(n_424),
.Y(n_420)
);

OAI22xp33_ASAP7_75t_SL g207 ( 
.A1(n_4),
.A2(n_208),
.B1(n_212),
.B2(n_213),
.Y(n_207)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_4),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_SL g275 ( 
.A1(n_4),
.A2(n_182),
.B1(n_212),
.B2(n_276),
.Y(n_275)
);

AOI22xp33_ASAP7_75t_L g371 ( 
.A1(n_4),
.A2(n_212),
.B1(n_372),
.B2(n_374),
.Y(n_371)
);

AOI22xp5_ASAP7_75t_L g416 ( 
.A1(n_4),
.A2(n_212),
.B1(n_366),
.B2(n_367),
.Y(n_416)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_5),
.A2(n_182),
.B1(n_183),
.B2(n_187),
.Y(n_181)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_5),
.Y(n_187)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_5),
.B(n_197),
.C(n_200),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_5),
.B(n_78),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_5),
.B(n_226),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_5),
.B(n_123),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_282),
.Y(n_281)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_6),
.A2(n_33),
.B1(n_49),
.B2(n_51),
.Y(n_48)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_6),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_6),
.A2(n_51),
.B1(n_324),
.B2(n_325),
.Y(n_323)
);

OAI22xp33_ASAP7_75t_SL g396 ( 
.A1(n_6),
.A2(n_51),
.B1(n_397),
.B2(n_401),
.Y(n_396)
);

AOI22xp33_ASAP7_75t_SL g413 ( 
.A1(n_6),
.A2(n_51),
.B1(n_76),
.B2(n_414),
.Y(n_413)
);

AOI22xp33_ASAP7_75t_L g235 ( 
.A1(n_7),
.A2(n_182),
.B1(n_236),
.B2(n_237),
.Y(n_235)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_7),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_7),
.A2(n_208),
.B1(n_228),
.B2(n_236),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g312 ( 
.A1(n_7),
.A2(n_236),
.B1(n_313),
.B2(n_315),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g439 ( 
.A1(n_7),
.A2(n_236),
.B1(n_440),
.B2(n_442),
.Y(n_439)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_8),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_8),
.Y(n_47)
);

INVx3_ASAP7_75t_L g522 ( 
.A(n_9),
.Y(n_522)
);

BUFx3_ASAP7_75t_L g105 ( 
.A(n_10),
.Y(n_105)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_10),
.Y(n_109)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_10),
.Y(n_114)
);

INVx8_ASAP7_75t_L g81 ( 
.A(n_11),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_12),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g223 ( 
.A(n_12),
.Y(n_223)
);

BUFx3_ASAP7_75t_L g230 ( 
.A(n_12),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g525 ( 
.A(n_13),
.Y(n_525)
);

AOI22xp33_ASAP7_75t_SL g92 ( 
.A1(n_14),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_14),
.Y(n_95)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_14),
.A2(n_80),
.B1(n_95),
.B2(n_125),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_14),
.A2(n_95),
.B1(n_209),
.B2(n_392),
.Y(n_391)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_15),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_SL g54 ( 
.A1(n_16),
.A2(n_55),
.B1(n_58),
.B2(n_61),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_16),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_16),
.A2(n_61),
.B1(n_159),
.B2(n_164),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_16),
.A2(n_61),
.B1(n_228),
.B2(n_353),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_L g404 ( 
.A1(n_16),
.A2(n_61),
.B1(n_238),
.B2(n_405),
.Y(n_404)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_18),
.A2(n_126),
.B1(n_190),
.B2(n_193),
.Y(n_189)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_18),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_L g227 ( 
.A1(n_18),
.A2(n_193),
.B1(n_228),
.B2(n_231),
.Y(n_227)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_18),
.A2(n_193),
.B1(n_287),
.B2(n_290),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_L g365 ( 
.A1(n_18),
.A2(n_137),
.B1(n_193),
.B2(n_366),
.Y(n_365)
);

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_520),
.B(n_523),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_171),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_169),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_139),
.Y(n_22)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_23),
.B(n_139),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_128),
.B2(n_129),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_62),
.C(n_96),
.Y(n_25)
);

XNOR2xp5_ASAP7_75t_SL g141 ( 
.A(n_26),
.B(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_27),
.A2(n_48),
.B1(n_52),
.B2(n_54),
.Y(n_26)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_27),
.A2(n_52),
.B1(n_54),
.B2(n_134),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_27),
.A2(n_48),
.B1(n_52),
.B2(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_SL g415 ( 
.A1(n_27),
.A2(n_364),
.B(n_416),
.Y(n_415)
);

OAI22xp5_ASAP7_75t_L g438 ( 
.A1(n_27),
.A2(n_38),
.B1(n_416),
.B2(n_439),
.Y(n_438)
);

INVx2_ASAP7_75t_SL g27 ( 
.A(n_28),
.Y(n_27)
);

AOI21xp5_ASAP7_75t_L g360 ( 
.A1(n_28),
.A2(n_361),
.B(n_363),
.Y(n_360)
);

NAND2xp5_ASAP7_75t_L g465 ( 
.A(n_28),
.B(n_365),
.Y(n_465)
);

AND2x2_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_38),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_33),
.B1(n_35),
.B2(n_36),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

OAI32xp33_ASAP7_75t_L g339 ( 
.A1(n_33),
.A2(n_340),
.A3(n_341),
.B1(n_342),
.B2(n_344),
.Y(n_339)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_35),
.Y(n_152)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_36),
.Y(n_341)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g343 ( 
.A(n_37),
.Y(n_343)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_38),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_38),
.B(n_187),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_39),
.A2(n_40),
.B1(n_44),
.B2(n_46),
.Y(n_38)
);

INVx6_ASAP7_75t_L g373 ( 
.A(n_40),
.Y(n_373)
);

INVx5_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_42),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_42),
.Y(n_163)
);

BUFx6f_ASAP7_75t_L g289 ( 
.A(n_42),
.Y(n_289)
);

BUFx6f_ASAP7_75t_L g340 ( 
.A(n_42),
.Y(n_340)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_43),
.Y(n_77)
);

BUFx5_ASAP7_75t_L g168 ( 
.A(n_43),
.Y(n_168)
);

INVx3_ASAP7_75t_L g292 ( 
.A(n_43),
.Y(n_292)
);

INVx4_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

INVx6_ASAP7_75t_SL g299 ( 
.A(n_45),
.Y(n_299)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_49),
.Y(n_138)
);

INVx3_ASAP7_75t_L g443 ( 
.A(n_49),
.Y(n_443)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx2_ASAP7_75t_L g441 ( 
.A(n_50),
.Y(n_441)
);

OAI21xp5_ASAP7_75t_L g475 ( 
.A1(n_52),
.A2(n_439),
.B(n_465),
.Y(n_475)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_53),
.B(n_365),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g464 ( 
.A(n_53),
.B(n_147),
.Y(n_464)
);

INVx2_ASAP7_75t_SL g55 ( 
.A(n_56),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_60),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_62),
.A2(n_96),
.B1(n_97),
.B2(n_143),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_62),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g62 ( 
.A1(n_63),
.A2(n_86),
.B1(n_91),
.B2(n_92),
.Y(n_62)
);

INVx3_ASAP7_75t_SL g131 ( 
.A(n_63),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_63),
.A2(n_86),
.B1(n_91),
.B2(n_157),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_63),
.A2(n_91),
.B1(n_312),
.B2(n_371),
.Y(n_370)
);

OAI22xp5_ASAP7_75t_SL g409 ( 
.A1(n_63),
.A2(n_91),
.B1(n_410),
.B2(n_413),
.Y(n_409)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_64),
.B(n_78),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_70),
.B1(n_71),
.B2(n_75),
.Y(n_64)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx4_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_68),
.Y(n_85)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_69),
.Y(n_74)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_70),
.Y(n_93)
);

INVx3_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_74),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_75),
.B(n_343),
.Y(n_342)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

OAI21xp33_ASAP7_75t_SL g279 ( 
.A1(n_76),
.A2(n_187),
.B(n_280),
.Y(n_279)
);

INVx2_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx3_ASAP7_75t_L g314 ( 
.A(n_77),
.Y(n_314)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_78),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_131),
.B(n_132),
.Y(n_130)
);

AOI22x1_ASAP7_75t_L g444 ( 
.A1(n_78),
.A2(n_131),
.B1(n_319),
.B2(n_445),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_SL g452 ( 
.A1(n_78),
.A2(n_131),
.B1(n_158),
.B2(n_453),
.Y(n_452)
);

AO22x2_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_78)
);

INVx5_ASAP7_75t_L g407 ( 
.A(n_80),
.Y(n_407)
);

BUFx5_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx11_ASAP7_75t_L g83 ( 
.A(n_81),
.Y(n_83)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_81),
.Y(n_102)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_81),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_81),
.Y(n_182)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_81),
.Y(n_192)
);

BUFx3_ASAP7_75t_L g400 ( 
.A(n_81),
.Y(n_400)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx5_ASAP7_75t_L g111 ( 
.A(n_83),
.Y(n_111)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_83),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g377 ( 
.A(n_83),
.Y(n_377)
);

INVx6_ASAP7_75t_L g403 ( 
.A(n_83),
.Y(n_403)
);

AOI32xp33_ASAP7_75t_L g298 ( 
.A1(n_84),
.A2(n_182),
.A3(n_281),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVx5_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

BUFx2_ASAP7_75t_L g301 ( 
.A(n_85),
.Y(n_301)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_91),
.B(n_286),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g311 ( 
.A1(n_91),
.A2(n_312),
.B(n_318),
.Y(n_311)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_92),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_96),
.B(n_145),
.C(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g509 ( 
.A1(n_96),
.A2(n_97),
.B1(n_155),
.B2(n_156),
.Y(n_509)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_122),
.B(n_124),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_98),
.A2(n_181),
.B(n_188),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_98),
.A2(n_122),
.B1(n_235),
.B2(n_275),
.Y(n_274)
);

OAI21xp5_ASAP7_75t_SL g308 ( 
.A1(n_98),
.A2(n_188),
.B(n_275),
.Y(n_308)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_98),
.A2(n_122),
.B1(n_376),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g98 ( 
.A(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_99),
.B(n_189),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g395 ( 
.A1(n_99),
.A2(n_123),
.B1(n_396),
.B2(n_404),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_99),
.A2(n_123),
.B1(n_404),
.B2(n_420),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g455 ( 
.A1(n_99),
.A2(n_123),
.B1(n_420),
.B2(n_456),
.Y(n_455)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_100),
.B(n_112),
.Y(n_99)
);

OAI22xp33_ASAP7_75t_L g100 ( 
.A1(n_101),
.A2(n_103),
.B1(n_106),
.B2(n_110),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

BUFx5_ASAP7_75t_L g121 ( 
.A(n_109),
.Y(n_121)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_111),
.Y(n_110)
);

INVx5_ASAP7_75t_L g425 ( 
.A(n_111),
.Y(n_425)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_112),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_SL g234 ( 
.A1(n_112),
.A2(n_235),
.B(n_239),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g112 ( 
.A1(n_113),
.A2(n_115),
.B1(n_119),
.B2(n_121),
.Y(n_112)
);

INVx5_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_L g199 ( 
.A(n_114),
.Y(n_199)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx3_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g249 ( 
.A(n_117),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_118),
.Y(n_120)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_118),
.Y(n_204)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

INVx8_ASAP7_75t_L g327 ( 
.A(n_120),
.Y(n_327)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_122),
.A2(n_239),
.B(n_376),
.Y(n_375)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_123),
.B(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_124),
.Y(n_456)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_125),
.Y(n_238)
);

INVx4_ASAP7_75t_SL g125 ( 
.A(n_126),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_133),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g278 ( 
.A1(n_131),
.A2(n_279),
.B(n_285),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_131),
.B(n_319),
.Y(n_318)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_131),
.A2(n_285),
.B(n_478),
.Y(n_477)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_144),
.C(n_153),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g515 ( 
.A1(n_140),
.A2(n_141),
.B1(n_144),
.B2(n_145),
.Y(n_515)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_144),
.A2(n_145),
.B1(n_509),
.B2(n_510),
.Y(n_508)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVxp67_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

INVx8_ASAP7_75t_L g150 ( 
.A(n_151),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_L g513 ( 
.A1(n_153),
.A2(n_154),
.B1(n_514),
.B2(n_515),
.Y(n_513)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx4_ASAP7_75t_SL g161 ( 
.A(n_162),
.Y(n_161)
);

INVx5_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_165),
.Y(n_164)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

INVx6_ASAP7_75t_L g284 ( 
.A(n_168),
.Y(n_284)
);

INVx2_ASAP7_75t_L g317 ( 
.A(n_168),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_173),
.A2(n_504),
.B(n_517),
.Y(n_172)
);

OAI311xp33_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_380),
.A3(n_480),
.B1(n_498),
.C1(n_499),
.Y(n_173)
);

AOI21x1_ASAP7_75t_L g174 ( 
.A1(n_175),
.A2(n_333),
.B(n_379),
.Y(n_174)
);

AO21x1_ASAP7_75t_L g175 ( 
.A1(n_176),
.A2(n_303),
.B(n_332),
.Y(n_175)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_269),
.B(n_302),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_242),
.B(n_268),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_179),
.B(n_205),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_179),
.B(n_205),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g179 ( 
.A(n_180),
.B(n_194),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_180),
.A2(n_194),
.B1(n_195),
.B2(n_266),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_180),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_183),
.B(n_196),
.Y(n_195)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx6_ASAP7_75t_L g423 ( 
.A(n_186),
.Y(n_423)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_187),
.A2(n_217),
.B(n_224),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_187),
.B(n_345),
.Y(n_344)
);

OAI21xp33_ASAP7_75t_SL g361 ( 
.A1(n_187),
.A2(n_344),
.B(n_362),
.Y(n_361)
);

INVx4_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_191),
.Y(n_276)
);

INVx4_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

BUFx6f_ASAP7_75t_L g231 ( 
.A(n_203),
.Y(n_231)
);

INVx5_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_204),
.Y(n_211)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_204),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_206),
.B(n_232),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_206),
.B(n_233),
.C(n_241),
.Y(n_270)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_217),
.B(n_224),
.Y(n_206)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_207),
.Y(n_262)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_210),
.Y(n_209)
);

INVx6_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx4_ASAP7_75t_SL g214 ( 
.A(n_215),
.Y(n_214)
);

INVx4_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI22xp5_ASAP7_75t_L g349 ( 
.A1(n_217),
.A2(n_297),
.B1(n_350),
.B2(n_351),
.Y(n_349)
);

AOI22xp5_ASAP7_75t_L g385 ( 
.A1(n_217),
.A2(n_386),
.B1(n_389),
.B2(n_391),
.Y(n_385)
);

OAI21xp5_ASAP7_75t_SL g426 ( 
.A1(n_217),
.A2(n_391),
.B(n_427),
.Y(n_426)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_218),
.B(n_227),
.Y(n_256)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_218),
.A2(n_261),
.B1(n_262),
.B2(n_263),
.Y(n_260)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_218),
.A2(n_296),
.B1(n_323),
.B2(n_328),
.Y(n_322)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_218),
.A2(n_352),
.B1(n_434),
.B2(n_435),
.Y(n_433)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_219),
.B(n_221),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

INVx2_ASAP7_75t_L g427 ( 
.A(n_220),
.Y(n_427)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g222 ( 
.A(n_223),
.Y(n_222)
);

BUFx5_ASAP7_75t_L g388 ( 
.A(n_223),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_227),
.Y(n_224)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_225),
.Y(n_255)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_226),
.Y(n_390)
);

INVx8_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

BUFx8_ASAP7_75t_L g229 ( 
.A(n_230),
.Y(n_229)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_230),
.Y(n_354)
);

BUFx5_ASAP7_75t_L g394 ( 
.A(n_230),
.Y(n_394)
);

INVx3_ASAP7_75t_L g324 ( 
.A(n_231),
.Y(n_324)
);

AOI22xp5_ASAP7_75t_SL g232 ( 
.A1(n_233),
.A2(n_234),
.B1(n_240),
.B2(n_241),
.Y(n_232)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp33_ASAP7_75t_SL g300 ( 
.A(n_237),
.B(n_301),
.Y(n_300)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_243),
.A2(n_259),
.B(n_267),
.Y(n_242)
);

AOI21xp5_ASAP7_75t_L g243 ( 
.A1(n_244),
.A2(n_252),
.B(n_258),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_251),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_250),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_248),
.Y(n_247)
);

INVx4_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_257),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_253),
.B(n_257),
.Y(n_258)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_254),
.A2(n_255),
.B(n_256),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_254),
.Y(n_261)
);

AOI21xp5_ASAP7_75t_L g294 ( 
.A1(n_256),
.A2(n_295),
.B(n_297),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_265),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_260),
.B(n_265),
.Y(n_267)
);

INVx4_ASAP7_75t_L g297 ( 
.A(n_263),
.Y(n_297)
);

INVx4_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_271),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_270),
.B(n_271),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_293),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_274),
.B1(n_277),
.B2(n_278),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_277),
.C(n_293),
.Y(n_304)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

INVxp33_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx3_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx2_ASAP7_75t_L g283 ( 
.A(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_286),
.Y(n_319)
);

INVx3_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx12f_ASAP7_75t_L g288 ( 
.A(n_289),
.Y(n_288)
);

INVx2_ASAP7_75t_L g412 ( 
.A(n_289),
.Y(n_412)
);

INVx8_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_292),
.Y(n_291)
);

INVx4_ASAP7_75t_L g414 ( 
.A(n_292),
.Y(n_414)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_298),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_294),
.B(n_298),
.Y(n_309)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_296),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

NOR2xp33_ASAP7_75t_SL g332 ( 
.A(n_304),
.B(n_305),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_310),
.B2(n_331),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_309),
.Y(n_307)
);

MAJIxp5_ASAP7_75t_L g334 ( 
.A(n_308),
.B(n_309),
.C(n_331),
.Y(n_334)
);

INVx1_ASAP7_75t_L g331 ( 
.A(n_310),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_320),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g355 ( 
.A(n_311),
.B(n_321),
.C(n_322),
.Y(n_355)
);

INVx5_ASAP7_75t_L g374 ( 
.A(n_313),
.Y(n_374)
);

INVx4_ASAP7_75t_L g313 ( 
.A(n_314),
.Y(n_313)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_317),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_322),
.Y(n_320)
);

INVxp67_ASAP7_75t_L g350 ( 
.A(n_323),
.Y(n_350)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

INVx5_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx2_ASAP7_75t_L g329 ( 
.A(n_330),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_335),
.Y(n_333)
);

NOR2xp33_ASAP7_75t_SL g379 ( 
.A(n_334),
.B(n_335),
.Y(n_379)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_358),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_355),
.B1(n_356),
.B2(n_357),
.Y(n_336)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_337),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_348),
.B2(n_349),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_339),
.B(n_348),
.Y(n_476)
);

INVx4_ASAP7_75t_L g345 ( 
.A(n_346),
.Y(n_345)
);

INVx3_ASAP7_75t_L g346 ( 
.A(n_347),
.Y(n_346)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_349),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g351 ( 
.A(n_352),
.Y(n_351)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_354),
.Y(n_353)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_355),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g494 ( 
.A(n_355),
.B(n_356),
.C(n_358),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_359),
.A2(n_360),
.B1(n_369),
.B2(n_378),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g489 ( 
.A(n_359),
.B(n_370),
.C(n_375),
.Y(n_489)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_364),
.Y(n_363)
);

INVx3_ASAP7_75t_L g366 ( 
.A(n_367),
.Y(n_366)
);

INVx4_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

INVx1_ASAP7_75t_L g378 ( 
.A(n_369),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_SL g369 ( 
.A(n_370),
.B(n_375),
.Y(n_369)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_371),
.Y(n_478)
);

INVx3_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp33_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_466),
.Y(n_380)
);

A2O1A1Ixp33_ASAP7_75t_SL g499 ( 
.A1(n_381),
.A2(n_466),
.B(n_500),
.C(n_503),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_446),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g498 ( 
.A(n_382),
.B(n_446),
.Y(n_498)
);

MAJIxp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_417),
.C(n_429),
.Y(n_382)
);

FAx1_ASAP7_75t_SL g479 ( 
.A(n_383),
.B(n_417),
.CI(n_429),
.CON(n_479),
.SN(n_479)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_408),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_384),
.B(n_409),
.C(n_415),
.Y(n_447)
);

NOR2xp33_ASAP7_75t_L g384 ( 
.A(n_385),
.B(n_395),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g472 ( 
.A(n_385),
.B(n_395),
.Y(n_472)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_386),
.Y(n_434)
);

INVx5_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

BUFx3_ASAP7_75t_L g389 ( 
.A(n_390),
.Y(n_389)
);

CKINVDCx14_ASAP7_75t_R g392 ( 
.A(n_393),
.Y(n_392)
);

INVx2_ASAP7_75t_L g393 ( 
.A(n_394),
.Y(n_393)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_396),
.Y(n_432)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx2_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

INVx3_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

INVx3_ASAP7_75t_SL g401 ( 
.A(n_402),
.Y(n_401)
);

INVx8_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_406),
.Y(n_405)
);

INVx2_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_409),
.B(n_415),
.Y(n_408)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_410),
.Y(n_445)
);

INVx2_ASAP7_75t_L g411 ( 
.A(n_412),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_413),
.Y(n_453)
);

OAI22xp5_ASAP7_75t_SL g417 ( 
.A1(n_418),
.A2(n_419),
.B1(n_426),
.B2(n_428),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g460 ( 
.A(n_419),
.B(n_426),
.Y(n_460)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_422),
.Y(n_421)
);

INVx3_ASAP7_75t_L g422 ( 
.A(n_423),
.Y(n_422)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_425),
.Y(n_424)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_426),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g461 ( 
.A1(n_426),
.A2(n_428),
.B1(n_462),
.B2(n_463),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_L g507 ( 
.A1(n_426),
.A2(n_460),
.B(n_463),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_430),
.B(n_437),
.C(n_444),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g469 ( 
.A(n_430),
.B(n_470),
.Y(n_469)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_433),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g488 ( 
.A(n_431),
.B(n_433),
.Y(n_488)
);

INVx3_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

AOI22xp5_ASAP7_75t_SL g470 ( 
.A1(n_437),
.A2(n_438),
.B1(n_444),
.B2(n_471),
.Y(n_470)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_438),
.Y(n_437)
);

INVx4_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_443),
.Y(n_442)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_444),
.Y(n_471)
);

XNOR2xp5_ASAP7_75t_L g446 ( 
.A(n_447),
.B(n_448),
.Y(n_446)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_447),
.B(n_450),
.C(n_458),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g448 ( 
.A1(n_449),
.A2(n_450),
.B1(n_458),
.B2(n_459),
.Y(n_448)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_450),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_L g450 ( 
.A1(n_451),
.A2(n_454),
.B(n_457),
.Y(n_450)
);

INVxp67_ASAP7_75t_L g451 ( 
.A(n_452),
.Y(n_451)
);

AND2x2_ASAP7_75t_L g457 ( 
.A(n_452),
.B(n_455),
.Y(n_457)
);

INVxp67_ASAP7_75t_L g454 ( 
.A(n_455),
.Y(n_454)
);

FAx1_ASAP7_75t_SL g506 ( 
.A(n_457),
.B(n_507),
.CI(n_508),
.CON(n_506),
.SN(n_506)
);

MAJIxp5_ASAP7_75t_L g516 ( 
.A(n_457),
.B(n_507),
.C(n_508),
.Y(n_516)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_459),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

NAND2xp5_ASAP7_75t_L g463 ( 
.A(n_464),
.B(n_465),
.Y(n_463)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_467),
.B(n_479),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g503 ( 
.A(n_467),
.B(n_479),
.Y(n_503)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_468),
.B(n_472),
.C(n_473),
.Y(n_467)
);

AOI22xp5_ASAP7_75t_SL g491 ( 
.A1(n_468),
.A2(n_469),
.B1(n_472),
.B2(n_492),
.Y(n_491)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_469),
.Y(n_468)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_472),
.Y(n_492)
);

XNOR2xp5_ASAP7_75t_L g490 ( 
.A(n_473),
.B(n_491),
.Y(n_490)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_474),
.B(n_476),
.C(n_477),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_474),
.A2(n_475),
.B1(n_477),
.B2(n_486),
.Y(n_485)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_475),
.Y(n_474)
);

XOR2xp5_ASAP7_75t_L g484 ( 
.A(n_476),
.B(n_485),
.Y(n_484)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_477),
.Y(n_486)
);

BUFx24_ASAP7_75t_SL g527 ( 
.A(n_479),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g480 ( 
.A(n_481),
.B(n_493),
.Y(n_480)
);

INVx1_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

OAI21xp5_ASAP7_75t_L g500 ( 
.A1(n_482),
.A2(n_501),
.B(n_502),
.Y(n_500)
);

NOR2x1_ASAP7_75t_L g482 ( 
.A(n_483),
.B(n_490),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_483),
.B(n_490),
.Y(n_502)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_484),
.B(n_487),
.C(n_489),
.Y(n_483)
);

XOR2xp5_ASAP7_75t_L g495 ( 
.A(n_484),
.B(n_496),
.Y(n_495)
);

AOI22xp5_ASAP7_75t_L g496 ( 
.A1(n_487),
.A2(n_488),
.B1(n_489),
.B2(n_497),
.Y(n_496)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g497 ( 
.A(n_489),
.Y(n_497)
);

OR2x2_ASAP7_75t_L g493 ( 
.A(n_494),
.B(n_495),
.Y(n_493)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_495),
.Y(n_501)
);

NOR2xp33_ASAP7_75t_L g504 ( 
.A(n_505),
.B(n_512),
.Y(n_504)
);

NOR2xp33_ASAP7_75t_SL g505 ( 
.A(n_506),
.B(n_511),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g518 ( 
.A(n_506),
.B(n_511),
.Y(n_518)
);

BUFx24_ASAP7_75t_SL g526 ( 
.A(n_506),
.Y(n_526)
);

INVx1_ASAP7_75t_L g510 ( 
.A(n_509),
.Y(n_510)
);

OAI21xp5_ASAP7_75t_L g517 ( 
.A1(n_512),
.A2(n_518),
.B(n_519),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_513),
.B(n_516),
.Y(n_512)
);

NAND2xp5_ASAP7_75t_L g519 ( 
.A(n_513),
.B(n_516),
.Y(n_519)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

BUFx4f_ASAP7_75t_SL g520 ( 
.A(n_521),
.Y(n_520)
);

INVx13_ASAP7_75t_L g521 ( 
.A(n_522),
.Y(n_521)
);

INVx6_ASAP7_75t_L g524 ( 
.A(n_522),
.Y(n_524)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_524),
.B(n_525),
.Y(n_523)
);


endmodule