module fake_jpeg_22965_n_135 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_135);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_135;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

HB1xp67_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx6_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

BUFx16f_ASAP7_75t_L g15 ( 
.A(n_3),
.Y(n_15)
);

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

INVx2_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_0),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_11),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_12),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_16),
.B(n_0),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_26),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_14),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g37 ( 
.A1(n_29),
.A2(n_14),
.B1(n_21),
.B2(n_27),
.Y(n_37)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_31),
.Y(n_46)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_17),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_32),
.B(n_35),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_33),
.Y(n_39)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

CKINVDCx14_ASAP7_75t_R g35 ( 
.A(n_15),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

AOI21xp5_ASAP7_75t_L g55 ( 
.A1(n_37),
.A2(n_50),
.B(n_25),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_SL g56 ( 
.A(n_40),
.B(n_29),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_33),
.Y(n_43)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_44),
.B(n_47),
.Y(n_53)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_49),
.B(n_20),
.Y(n_54)
);

AOI22xp33_ASAP7_75t_SL g50 ( 
.A1(n_31),
.A2(n_14),
.B1(n_25),
.B2(n_20),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g51 ( 
.A1(n_46),
.A2(n_36),
.B1(n_34),
.B2(n_31),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g76 ( 
.A1(n_51),
.A2(n_57),
.B1(n_65),
.B2(n_47),
.Y(n_76)
);

HAxp5_ASAP7_75t_SL g73 ( 
.A(n_54),
.B(n_55),
.CON(n_73),
.SN(n_73)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_56),
.B(n_57),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g57 ( 
.A1(n_40),
.A2(n_34),
.B1(n_32),
.B2(n_29),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_30),
.C(n_33),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_58),
.B(n_59),
.Y(n_71)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_49),
.B(n_30),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_41),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_46),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_38),
.B(n_24),
.Y(n_61)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_61),
.Y(n_66)
);

HB1xp67_ASAP7_75t_L g62 ( 
.A(n_44),
.Y(n_62)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_62),
.Y(n_74)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_44),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_64),
.B(n_15),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_45),
.A2(n_24),
.B1(n_27),
.B2(n_23),
.Y(n_65)
);

INVx1_ASAP7_75t_SL g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_68),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_60),
.B(n_46),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_70),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_65),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_72),
.B(n_75),
.Y(n_93)
);

INVxp67_ASAP7_75t_L g75 ( 
.A(n_53),
.Y(n_75)
);

AO21x1_ASAP7_75t_L g88 ( 
.A1(n_76),
.A2(n_63),
.B(n_43),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_54),
.B(n_38),
.Y(n_77)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_77),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_39),
.Y(n_78)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_78),
.Y(n_89)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_64),
.Y(n_79)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_56),
.A2(n_48),
.B1(n_45),
.B2(n_42),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g84 ( 
.A1(n_80),
.A2(n_39),
.B1(n_42),
.B2(n_52),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_81),
.A2(n_44),
.B(n_74),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_71),
.B(n_58),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_91),
.Y(n_97)
);

CKINVDCx14_ASAP7_75t_R g96 ( 
.A(n_84),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_87),
.B(n_80),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_88),
.B(n_76),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_71),
.B(n_63),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_43),
.C(n_52),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g102 ( 
.A(n_92),
.B(n_94),
.Y(n_102)
);

XNOR2xp5_ASAP7_75t_L g94 ( 
.A(n_72),
.B(n_15),
.Y(n_94)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_90),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_95),
.B(n_100),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_91),
.B(n_93),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_89),
.B(n_68),
.Y(n_99)
);

AOI322xp5_ASAP7_75t_SL g100 ( 
.A1(n_85),
.A2(n_73),
.A3(n_66),
.B1(n_67),
.B2(n_77),
.C1(n_69),
.C2(n_70),
.Y(n_100)
);

INVx2_ASAP7_75t_SL g101 ( 
.A(n_86),
.Y(n_101)
);

CKINVDCx14_ASAP7_75t_R g112 ( 
.A(n_101),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g103 ( 
.A(n_82),
.B(n_66),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_103),
.A2(n_92),
.B1(n_84),
.B2(n_88),
.Y(n_108)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_104),
.A2(n_105),
.B(n_106),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g105 ( 
.A1(n_83),
.A2(n_74),
.B(n_79),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_97),
.B(n_94),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g122 ( 
.A(n_107),
.B(n_111),
.Y(n_122)
);

OAI21xp5_ASAP7_75t_SL g117 ( 
.A1(n_108),
.A2(n_113),
.B(n_115),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_97),
.B(n_87),
.C(n_86),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_109),
.B(n_99),
.C(n_98),
.Y(n_118)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_105),
.A2(n_23),
.B(n_19),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_106),
.A2(n_52),
.B1(n_19),
.B2(n_18),
.Y(n_115)
);

BUFx24_ASAP7_75t_SL g116 ( 
.A(n_107),
.Y(n_116)
);

BUFx24_ASAP7_75t_SL g123 ( 
.A(n_116),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_118),
.B(n_119),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_109),
.B(n_102),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_114),
.B(n_102),
.C(n_96),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_121),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_108),
.B(n_101),
.C(n_18),
.Y(n_121)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_122),
.A2(n_111),
.B(n_117),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_124),
.B(n_110),
.C(n_112),
.Y(n_128)
);

OR2x6_ASAP7_75t_L g127 ( 
.A(n_117),
.B(n_113),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_128),
.B(n_129),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_127),
.A2(n_110),
.B1(n_115),
.B2(n_101),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_126),
.B(n_9),
.Y(n_130)
);

AOI322xp5_ASAP7_75t_L g132 ( 
.A1(n_130),
.A2(n_125),
.A3(n_123),
.B1(n_16),
.B2(n_8),
.C1(n_10),
.C2(n_7),
.Y(n_132)
);

AOI21xp5_ASAP7_75t_SL g133 ( 
.A1(n_132),
.A2(n_2),
.B(n_4),
.Y(n_133)
);

AOI21x1_ASAP7_75t_L g134 ( 
.A1(n_133),
.A2(n_131),
.B(n_22),
.Y(n_134)
);

BUFx24_ASAP7_75t_SL g135 ( 
.A(n_134),
.Y(n_135)
);


endmodule