module fake_jpeg_10989_n_525 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_525);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_525;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_524;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_12),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_0),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_2),
.Y(n_22)
);

BUFx4f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_0),
.Y(n_25)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_4),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_18),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g31 ( 
.A(n_1),
.B(n_7),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_6),
.B(n_3),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx8_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_3),
.B(n_10),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_5),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_5),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_16),
.Y(n_42)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_4),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_17),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_4),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_10),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_6),
.Y(n_47)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_13),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_51),
.Y(n_151)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_23),
.Y(n_52)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_20),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g157 ( 
.A(n_53),
.Y(n_157)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

CKINVDCx16_ASAP7_75t_R g108 ( 
.A(n_54),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_32),
.B(n_18),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_55),
.B(n_83),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g56 ( 
.A(n_37),
.B(n_18),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_56),
.B(n_58),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_57),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_37),
.B(n_30),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_20),
.Y(n_59)
);

INVx6_ASAP7_75t_L g119 ( 
.A(n_59),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g60 ( 
.A(n_34),
.Y(n_60)
);

INVx1_ASAP7_75t_SL g139 ( 
.A(n_60),
.Y(n_139)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_46),
.Y(n_61)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_61),
.Y(n_107)
);

BUFx12f_ASAP7_75t_L g62 ( 
.A(n_34),
.Y(n_62)
);

INVx5_ASAP7_75t_L g161 ( 
.A(n_62),
.Y(n_161)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_34),
.Y(n_63)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx12_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

BUFx2_ASAP7_75t_L g144 ( 
.A(n_64),
.Y(n_144)
);

INVx4_ASAP7_75t_SL g65 ( 
.A(n_22),
.Y(n_65)
);

INVx4_ASAP7_75t_L g122 ( 
.A(n_65),
.Y(n_122)
);

INVx4_ASAP7_75t_SL g66 ( 
.A(n_22),
.Y(n_66)
);

INVx4_ASAP7_75t_L g140 ( 
.A(n_66),
.Y(n_140)
);

INVx3_ASAP7_75t_L g67 ( 
.A(n_34),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g145 ( 
.A(n_67),
.Y(n_145)
);

INVx4_ASAP7_75t_L g68 ( 
.A(n_43),
.Y(n_68)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_68),
.Y(n_104)
);

INVx11_ASAP7_75t_L g69 ( 
.A(n_34),
.Y(n_69)
);

BUFx2_ASAP7_75t_SL g142 ( 
.A(n_69),
.Y(n_142)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_70),
.Y(n_106)
);

BUFx5_ASAP7_75t_L g71 ( 
.A(n_22),
.Y(n_71)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_71),
.Y(n_150)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_43),
.Y(n_72)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_72),
.Y(n_133)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_22),
.Y(n_73)
);

INVx6_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx8_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_74),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_31),
.B(n_0),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_76),
.Y(n_115)
);

INVx8_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

INVx6_ASAP7_75t_L g135 ( 
.A(n_77),
.Y(n_135)
);

INVx8_ASAP7_75t_L g78 ( 
.A(n_38),
.Y(n_78)
);

INVx6_ASAP7_75t_L g154 ( 
.A(n_78),
.Y(n_154)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_38),
.Y(n_79)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_79),
.Y(n_111)
);

INVx8_ASAP7_75t_L g80 ( 
.A(n_38),
.Y(n_80)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_80),
.Y(n_153)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_23),
.Y(n_81)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_81),
.Y(n_114)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_82),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_32),
.B(n_30),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_23),
.Y(n_84)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_84),
.Y(n_137)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_26),
.Y(n_85)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_85),
.Y(n_148)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_43),
.Y(n_86)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_86),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_23),
.Y(n_87)
);

INVx2_ASAP7_75t_L g159 ( 
.A(n_87),
.Y(n_159)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_23),
.Y(n_88)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_88),
.Y(n_162)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_43),
.Y(n_89)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_89),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_26),
.Y(n_90)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_90),
.Y(n_117)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_43),
.Y(n_91)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_91),
.Y(n_120)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_43),
.Y(n_92)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_21),
.B(n_45),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_93),
.B(n_94),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_21),
.B(n_1),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_95),
.Y(n_131)
);

BUFx3_ASAP7_75t_L g96 ( 
.A(n_24),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_50),
.Y(n_97)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_97),
.Y(n_149)
);

BUFx5_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_98),
.B(n_99),
.Y(n_110)
);

BUFx12f_ASAP7_75t_L g99 ( 
.A(n_19),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g100 ( 
.A(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_101),
.Y(n_121)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_31),
.B(n_1),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_54),
.A2(n_31),
.B1(n_50),
.B2(n_27),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g178 ( 
.A1(n_113),
.A2(n_132),
.B1(n_141),
.B2(n_147),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_101),
.B(n_48),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g200 ( 
.A(n_123),
.B(n_126),
.Y(n_200)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_69),
.A2(n_33),
.B1(n_19),
.B2(n_49),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_124),
.A2(n_60),
.B1(n_62),
.B2(n_47),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_64),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_75),
.B(n_48),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_129),
.B(n_136),
.Y(n_180)
);

AOI22xp33_ASAP7_75t_L g132 ( 
.A1(n_51),
.A2(n_31),
.B1(n_19),
.B2(n_33),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_99),
.B(n_36),
.Y(n_136)
);

AOI21xp33_ASAP7_75t_SL g138 ( 
.A1(n_64),
.A2(n_2),
.B(n_3),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g216 ( 
.A(n_138),
.B(n_2),
.Y(n_216)
);

OAI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_53),
.A2(n_25),
.B1(n_47),
.B2(n_41),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_99),
.B(n_45),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_143),
.B(n_146),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_68),
.B(n_36),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_L g147 ( 
.A1(n_57),
.A2(n_33),
.B1(n_40),
.B2(n_44),
.Y(n_147)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_96),
.Y(n_155)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_155),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_156),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_61),
.B(n_40),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_158),
.B(n_74),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_59),
.A2(n_42),
.B1(n_44),
.B2(n_47),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g183 ( 
.A1(n_160),
.A2(n_27),
.B1(n_49),
.B2(n_41),
.Y(n_183)
);

INVx1_ASAP7_75t_SL g163 ( 
.A(n_139),
.Y(n_163)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_163),
.Y(n_223)
);

INVx4_ASAP7_75t_L g164 ( 
.A(n_161),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g267 ( 
.A(n_164),
.Y(n_267)
);

INVxp67_ASAP7_75t_L g261 ( 
.A(n_166),
.Y(n_261)
);

INVx13_ASAP7_75t_L g167 ( 
.A(n_144),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g246 ( 
.A(n_167),
.Y(n_246)
);

BUFx4f_ASAP7_75t_L g168 ( 
.A(n_111),
.Y(n_168)
);

INVx3_ASAP7_75t_L g254 ( 
.A(n_168),
.Y(n_254)
);

INVx3_ASAP7_75t_L g169 ( 
.A(n_153),
.Y(n_169)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_169),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_109),
.B(n_42),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_170),
.B(n_172),
.Y(n_247)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_102),
.Y(n_171)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_171),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_134),
.B(n_86),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_112),
.B(n_72),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_182),
.Y(n_226)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

INVx3_ASAP7_75t_SL g250 ( 
.A(n_174),
.Y(n_250)
);

OAI22xp33_ASAP7_75t_SL g176 ( 
.A1(n_138),
.A2(n_90),
.B1(n_79),
.B2(n_97),
.Y(n_176)
);

AOI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_176),
.A2(n_214),
.B1(n_215),
.B2(n_150),
.Y(n_262)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_152),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_177),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_112),
.A2(n_73),
.B1(n_80),
.B2(n_78),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_179),
.A2(n_183),
.B1(n_187),
.B2(n_192),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g181 ( 
.A1(n_160),
.A2(n_60),
.B1(n_62),
.B2(n_41),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_181),
.A2(n_139),
.B1(n_140),
.B2(n_122),
.Y(n_229)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_125),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g184 ( 
.A(n_146),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_184),
.B(n_185),
.Y(n_233)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

INVx2_ASAP7_75t_L g257 ( 
.A(n_186),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_L g187 ( 
.A1(n_121),
.A2(n_77),
.B1(n_87),
.B2(n_84),
.Y(n_187)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_103),
.Y(n_188)
);

BUFx3_ASAP7_75t_L g248 ( 
.A(n_188),
.Y(n_248)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

INVx3_ASAP7_75t_L g258 ( 
.A(n_189),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_105),
.B(n_49),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_190),
.B(n_198),
.Y(n_236)
);

BUFx2_ASAP7_75t_SL g191 ( 
.A(n_103),
.Y(n_191)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_191),
.Y(n_224)
);

OAI22xp33_ASAP7_75t_L g192 ( 
.A1(n_131),
.A2(n_91),
.B1(n_81),
.B2(n_95),
.Y(n_192)
);

INVx8_ASAP7_75t_L g193 ( 
.A(n_130),
.Y(n_193)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_193),
.Y(n_265)
);

INVx2_ASAP7_75t_L g194 ( 
.A(n_162),
.Y(n_194)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_194),
.Y(n_227)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_162),
.Y(n_195)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_195),
.Y(n_228)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_120),
.Y(n_196)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_196),
.Y(n_230)
);

INVx5_ASAP7_75t_L g197 ( 
.A(n_107),
.Y(n_197)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_197),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_145),
.Y(n_198)
);

INVx3_ASAP7_75t_SL g199 ( 
.A(n_111),
.Y(n_199)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_199),
.Y(n_243)
);

INVx6_ASAP7_75t_L g201 ( 
.A(n_151),
.Y(n_201)
);

BUFx3_ASAP7_75t_L g272 ( 
.A(n_201),
.Y(n_272)
);

INVx2_ASAP7_75t_SL g202 ( 
.A(n_107),
.Y(n_202)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_202),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_117),
.A2(n_35),
.B1(n_27),
.B2(n_28),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_204),
.A2(n_219),
.B1(n_133),
.B2(n_104),
.Y(n_268)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_130),
.Y(n_205)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_205),
.Y(n_266)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_152),
.Y(n_206)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_206),
.Y(n_270)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_114),
.Y(n_207)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_207),
.Y(n_271)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_135),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_208),
.B(n_209),
.Y(n_263)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_114),
.Y(n_209)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_159),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g269 ( 
.A(n_210),
.B(n_211),
.Y(n_269)
);

BUFx6f_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_106),
.B(n_39),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_212),
.B(n_217),
.Y(n_225)
);

OR2x2_ASAP7_75t_L g213 ( 
.A(n_122),
.B(n_39),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_213),
.A2(n_25),
.B(n_35),
.Y(n_245)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_157),
.Y(n_214)
);

INVx11_ASAP7_75t_L g215 ( 
.A(n_142),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_SL g264 ( 
.A1(n_216),
.A2(n_4),
.B(n_5),
.Y(n_264)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_137),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g218 ( 
.A(n_115),
.B(n_39),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_218),
.B(n_220),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g219 ( 
.A1(n_149),
.A2(n_35),
.B1(n_28),
.B2(n_25),
.Y(n_219)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_116),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_128),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_221),
.B(n_148),
.Y(n_238)
);

AO22x2_ASAP7_75t_L g222 ( 
.A1(n_153),
.A2(n_66),
.B1(n_65),
.B2(n_74),
.Y(n_222)
);

O2A1O1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_222),
.A2(n_28),
.B(n_144),
.C(n_133),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g317 ( 
.A(n_229),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_183),
.A2(n_140),
.B1(n_148),
.B2(n_127),
.Y(n_232)
);

OAI22xp5_ASAP7_75t_L g291 ( 
.A1(n_232),
.A2(n_217),
.B1(n_207),
.B2(n_210),
.Y(n_291)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_213),
.A2(n_135),
.B1(n_154),
.B2(n_118),
.Y(n_237)
);

AOI22xp5_ASAP7_75t_L g292 ( 
.A1(n_237),
.A2(n_249),
.B1(n_260),
.B2(n_215),
.Y(n_292)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_238),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_165),
.B(n_110),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_239),
.B(n_242),
.Y(n_280)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_216),
.A2(n_200),
.B(n_180),
.Y(n_241)
);

OAI21xp5_ASAP7_75t_SL g295 ( 
.A1(n_241),
.A2(n_222),
.B(n_196),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_216),
.B(n_104),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_194),
.B(n_178),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_244),
.B(n_259),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g277 ( 
.A(n_245),
.B(n_163),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_193),
.A2(n_118),
.B1(n_119),
.B2(n_154),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_175),
.B(n_127),
.C(n_108),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_251),
.B(n_264),
.Y(n_302)
);

OA21x2_ASAP7_75t_L g290 ( 
.A1(n_255),
.A2(n_262),
.B(n_222),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g259 ( 
.A(n_171),
.B(n_186),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_205),
.A2(n_119),
.B1(n_137),
.B2(n_159),
.Y(n_260)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_268),
.Y(n_286)
);

BUFx2_ASAP7_75t_L g273 ( 
.A(n_265),
.Y(n_273)
);

INVx1_ASAP7_75t_SL g321 ( 
.A(n_273),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g274 ( 
.A1(n_244),
.A2(n_192),
.B1(n_208),
.B2(n_201),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_L g318 ( 
.A1(n_274),
.A2(n_278),
.B1(n_306),
.B2(n_243),
.Y(n_318)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_259),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_275),
.B(n_281),
.Y(n_330)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_271),
.Y(n_276)
);

HB1xp67_ASAP7_75t_L g325 ( 
.A(n_276),
.Y(n_325)
);

NOR3xp33_ASAP7_75t_L g329 ( 
.A(n_277),
.B(n_224),
.C(n_264),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_240),
.A2(n_262),
.B1(n_261),
.B2(n_268),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_238),
.Y(n_281)
);

XOR2xp5_ASAP7_75t_L g283 ( 
.A(n_239),
.B(n_203),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_283),
.B(n_228),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g284 ( 
.A(n_263),
.Y(n_284)
);

NOR2xp33_ASAP7_75t_L g339 ( 
.A(n_284),
.B(n_313),
.Y(n_339)
);

AOI22xp33_ASAP7_75t_SL g285 ( 
.A1(n_261),
.A2(n_199),
.B1(n_188),
.B2(n_202),
.Y(n_285)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_285),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g287 ( 
.A(n_235),
.B(n_182),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_287),
.B(n_293),
.Y(n_334)
);

INVx1_ASAP7_75t_SL g288 ( 
.A(n_223),
.Y(n_288)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_288),
.B(n_291),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_255),
.A2(n_219),
.B(n_204),
.Y(n_289)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_289),
.A2(n_307),
.B(n_248),
.Y(n_338)
);

OAI21xp5_ASAP7_75t_SL g348 ( 
.A1(n_290),
.A2(n_230),
.B(n_270),
.Y(n_348)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_292),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_235),
.B(n_236),
.Y(n_293)
);

INVx3_ASAP7_75t_L g294 ( 
.A(n_272),
.Y(n_294)
);

INVx4_ASAP7_75t_L g322 ( 
.A(n_294),
.Y(n_322)
);

INVxp67_ASAP7_75t_L g355 ( 
.A(n_295),
.Y(n_355)
);

INVx3_ASAP7_75t_L g296 ( 
.A(n_272),
.Y(n_296)
);

INVx4_ASAP7_75t_L g349 ( 
.A(n_296),
.Y(n_349)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_271),
.Y(n_297)
);

HB1xp67_ASAP7_75t_L g340 ( 
.A(n_297),
.Y(n_340)
);

OAI21xp5_ASAP7_75t_SL g298 ( 
.A1(n_242),
.A2(n_222),
.B(n_206),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g357 ( 
.A1(n_298),
.A2(n_300),
.B(n_308),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_237),
.A2(n_174),
.B1(n_169),
.B2(n_209),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_SL g324 ( 
.A1(n_299),
.A2(n_309),
.B1(n_310),
.B2(n_316),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g300 ( 
.A1(n_226),
.A2(n_167),
.B(n_197),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_227),
.Y(n_301)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_301),
.Y(n_336)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_253),
.Y(n_303)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_303),
.Y(n_341)
);

INVx1_ASAP7_75t_SL g304 ( 
.A(n_223),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_L g346 ( 
.A(n_305),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_240),
.A2(n_214),
.B1(n_211),
.B2(n_150),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_L g307 ( 
.A1(n_245),
.A2(n_189),
.B(n_164),
.Y(n_307)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_224),
.A2(n_168),
.B(n_8),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_225),
.A2(n_168),
.B1(n_8),
.B2(n_9),
.Y(n_309)
);

AOI22xp5_ASAP7_75t_L g310 ( 
.A1(n_225),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_SL g311 ( 
.A1(n_243),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_311)
);

AOI22xp33_ASAP7_75t_SL g332 ( 
.A1(n_311),
.A2(n_250),
.B1(n_267),
.B2(n_254),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_247),
.B(n_9),
.Y(n_312)
);

INVxp33_ASAP7_75t_L g353 ( 
.A(n_312),
.Y(n_353)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_269),
.Y(n_313)
);

BUFx8_ASAP7_75t_L g314 ( 
.A(n_246),
.Y(n_314)
);

BUFx12_ASAP7_75t_L g326 ( 
.A(n_314),
.Y(n_326)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_230),
.Y(n_315)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_315),
.Y(n_347)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_251),
.A2(n_266),
.B1(n_233),
.B2(n_252),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g388 ( 
.A(n_318),
.B(n_348),
.Y(n_388)
);

BUFx24_ASAP7_75t_SL g319 ( 
.A(n_283),
.Y(n_319)
);

INVxp67_ASAP7_75t_L g367 ( 
.A(n_319),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g320 ( 
.A1(n_278),
.A2(n_266),
.B1(n_234),
.B2(n_265),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g381 ( 
.A1(n_320),
.A2(n_331),
.B1(n_354),
.B2(n_305),
.Y(n_381)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_282),
.A2(n_241),
.B1(n_250),
.B2(n_252),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g369 ( 
.A1(n_327),
.A2(n_289),
.B1(n_306),
.B2(n_307),
.Y(n_369)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_329),
.Y(n_374)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_286),
.A2(n_234),
.B1(n_250),
.B2(n_231),
.Y(n_331)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_332),
.A2(n_317),
.B1(n_288),
.B2(n_304),
.Y(n_366)
);

XNOR2xp5_ASAP7_75t_SL g391 ( 
.A(n_333),
.B(n_327),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_275),
.B(n_281),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_335),
.B(n_337),
.Y(n_359)
);

INVx2_ASAP7_75t_SL g337 ( 
.A(n_315),
.Y(n_337)
);

OAI21xp5_ASAP7_75t_L g364 ( 
.A1(n_338),
.A2(n_351),
.B(n_356),
.Y(n_364)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_291),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_343),
.B(n_301),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_279),
.B(n_231),
.Y(n_344)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_344),
.B(n_282),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_SL g345 ( 
.A(n_280),
.B(n_228),
.Y(n_345)
);

NOR2xp33_ASAP7_75t_SL g371 ( 
.A(n_345),
.B(n_313),
.Y(n_371)
);

INVx1_ASAP7_75t_L g350 ( 
.A(n_276),
.Y(n_350)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_350),
.Y(n_358)
);

OAI21xp5_ASAP7_75t_SL g351 ( 
.A1(n_290),
.A2(n_270),
.B(n_257),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g354 ( 
.A1(n_286),
.A2(n_256),
.B1(n_258),
.B2(n_254),
.Y(n_354)
);

OAI21xp5_ASAP7_75t_SL g356 ( 
.A1(n_290),
.A2(n_317),
.B(n_280),
.Y(n_356)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_336),
.Y(n_360)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_360),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g361 ( 
.A(n_330),
.B(n_279),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g406 ( 
.A(n_361),
.B(n_362),
.Y(n_406)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_336),
.Y(n_363)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_363),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g365 ( 
.A(n_345),
.B(n_284),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_365),
.B(n_368),
.Y(n_410)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_366),
.A2(n_369),
.B1(n_373),
.B2(n_378),
.Y(n_401)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_325),
.Y(n_368)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_346),
.Y(n_370)
);

INVx1_ASAP7_75t_L g405 ( 
.A(n_370),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g400 ( 
.A(n_371),
.B(n_386),
.Y(n_400)
);

XNOR2xp5_ASAP7_75t_L g372 ( 
.A(n_333),
.B(n_302),
.Y(n_372)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_372),
.B(n_382),
.C(n_334),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g373 ( 
.A1(n_352),
.A2(n_274),
.B1(n_298),
.B2(n_295),
.Y(n_373)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_346),
.Y(n_375)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_375),
.Y(n_414)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_347),
.Y(n_376)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_376),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g377 ( 
.A(n_339),
.B(n_316),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g393 ( 
.A(n_377),
.B(n_379),
.Y(n_393)
);

AOI22xp33_ASAP7_75t_L g378 ( 
.A1(n_352),
.A2(n_292),
.B1(n_273),
.B2(n_299),
.Y(n_378)
);

CKINVDCx16_ASAP7_75t_R g379 ( 
.A(n_340),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_335),
.A2(n_308),
.B1(n_309),
.B2(n_310),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g415 ( 
.A1(n_380),
.A2(n_381),
.B1(n_385),
.B2(n_328),
.Y(n_415)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_344),
.B(n_302),
.Y(n_382)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_383),
.Y(n_403)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_357),
.A2(n_300),
.B(n_297),
.Y(n_384)
);

OAI21xp5_ASAP7_75t_SL g394 ( 
.A1(n_384),
.A2(n_390),
.B(n_355),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_SL g385 ( 
.A1(n_355),
.A2(n_273),
.B1(n_296),
.B2(n_294),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g386 ( 
.A(n_356),
.B(n_303),
.Y(n_386)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_326),
.Y(n_387)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_387),
.B(n_342),
.Y(n_411)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_347),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g420 ( 
.A(n_389),
.Y(n_420)
);

OAI21xp5_ASAP7_75t_SL g390 ( 
.A1(n_357),
.A2(n_314),
.B(n_248),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g398 ( 
.A(n_391),
.B(n_348),
.Y(n_398)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_372),
.B(n_382),
.Y(n_392)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_392),
.B(n_402),
.Y(n_423)
);

OAI21xp5_ASAP7_75t_SL g427 ( 
.A1(n_394),
.A2(n_418),
.B(n_386),
.Y(n_427)
);

INVx3_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_395),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g397 ( 
.A1(n_373),
.A2(n_318),
.B1(n_338),
.B2(n_320),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_397),
.A2(n_407),
.B1(n_363),
.B2(n_360),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g446 ( 
.A(n_398),
.B(n_326),
.Y(n_446)
);

XOR2xp5_ASAP7_75t_L g402 ( 
.A(n_391),
.B(n_351),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_404),
.B(n_359),
.C(n_384),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g407 ( 
.A1(n_369),
.A2(n_343),
.B1(n_323),
.B2(n_331),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_365),
.B(n_353),
.Y(n_408)
);

CKINVDCx14_ASAP7_75t_R g425 ( 
.A(n_408),
.Y(n_425)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_362),
.B(n_342),
.Y(n_409)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_409),
.B(n_412),
.Y(n_440)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_411),
.Y(n_429)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_361),
.B(n_324),
.Y(n_412)
);

XOR2xp5_ASAP7_75t_L g413 ( 
.A(n_364),
.B(n_324),
.Y(n_413)
);

XOR2xp5_ASAP7_75t_L g445 ( 
.A(n_413),
.B(n_341),
.Y(n_445)
);

OAI22xp5_ASAP7_75t_L g430 ( 
.A1(n_415),
.A2(n_364),
.B1(n_383),
.B2(n_388),
.Y(n_430)
);

NAND2xp5_ASAP7_75t_SL g416 ( 
.A(n_371),
.B(n_314),
.Y(n_416)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_416),
.Y(n_436)
);

AOI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_388),
.A2(n_323),
.B1(n_328),
.B2(n_337),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_SL g419 ( 
.A(n_377),
.B(n_314),
.Y(n_419)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_419),
.Y(n_438)
);

OAI22xp5_ASAP7_75t_L g421 ( 
.A1(n_374),
.A2(n_354),
.B1(n_337),
.B2(n_350),
.Y(n_421)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_421),
.Y(n_443)
);

XNOR2xp5_ASAP7_75t_L g450 ( 
.A(n_422),
.B(n_428),
.Y(n_450)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_392),
.B(n_359),
.C(n_390),
.Y(n_426)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_426),
.B(n_432),
.C(n_439),
.Y(n_447)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_427),
.B(n_433),
.Y(n_459)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_404),
.B(n_388),
.Y(n_428)
);

AND2x2_ASAP7_75t_L g452 ( 
.A(n_430),
.B(n_407),
.Y(n_452)
);

OAI21xp33_ASAP7_75t_SL g431 ( 
.A1(n_403),
.A2(n_387),
.B(n_368),
.Y(n_431)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_431),
.B(n_434),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_402),
.B(n_398),
.C(n_413),
.Y(n_432)
);

XNOR2xp5_ASAP7_75t_L g433 ( 
.A(n_393),
.B(n_385),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_SL g434 ( 
.A1(n_400),
.A2(n_379),
.B(n_389),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_401),
.A2(n_381),
.B1(n_380),
.B2(n_328),
.Y(n_435)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_435),
.A2(n_417),
.B1(n_414),
.B2(n_405),
.Y(n_462)
);

CKINVDCx16_ASAP7_75t_R g437 ( 
.A(n_410),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_437),
.B(n_406),
.Y(n_456)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_409),
.B(n_358),
.C(n_375),
.Y(n_439)
);

OA21x2_ASAP7_75t_L g441 ( 
.A1(n_397),
.A2(n_376),
.B(n_370),
.Y(n_441)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_441),
.A2(n_444),
.B(n_414),
.C(n_405),
.Y(n_465)
);

OAI22xp5_ASAP7_75t_SL g451 ( 
.A1(n_442),
.A2(n_415),
.B1(n_418),
.B2(n_403),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_SL g444 ( 
.A1(n_394),
.A2(n_326),
.B(n_341),
.C(n_321),
.Y(n_444)
);

XNOR2xp5_ASAP7_75t_SL g461 ( 
.A(n_445),
.B(n_446),
.Y(n_461)
);

BUFx24_ASAP7_75t_SL g449 ( 
.A(n_425),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_449),
.B(n_458),
.Y(n_477)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_451),
.A2(n_452),
.B1(n_462),
.B2(n_441),
.Y(n_471)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_429),
.Y(n_453)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_453),
.Y(n_474)
);

INVx1_ASAP7_75t_L g454 ( 
.A(n_436),
.Y(n_454)
);

NOR2xp33_ASAP7_75t_L g469 ( 
.A(n_454),
.B(n_463),
.Y(n_469)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_428),
.B(n_412),
.C(n_410),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g473 ( 
.A(n_455),
.B(n_457),
.C(n_460),
.Y(n_473)
);

OAI21x1_ASAP7_75t_L g479 ( 
.A1(n_456),
.A2(n_452),
.B(n_466),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_422),
.B(n_406),
.C(n_420),
.Y(n_457)
);

NOR2xp33_ASAP7_75t_SL g458 ( 
.A(n_438),
.B(n_367),
.Y(n_458)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_426),
.B(n_420),
.C(n_417),
.Y(n_460)
);

INVx1_ASAP7_75t_L g463 ( 
.A(n_424),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g464 ( 
.A1(n_435),
.A2(n_442),
.B1(n_443),
.B2(n_439),
.Y(n_464)
);

NOR2xp33_ASAP7_75t_L g476 ( 
.A(n_464),
.B(n_466),
.Y(n_476)
);

OAI21xp5_ASAP7_75t_L g468 ( 
.A1(n_465),
.A2(n_427),
.B(n_444),
.Y(n_468)
);

INVxp33_ASAP7_75t_L g466 ( 
.A(n_433),
.Y(n_466)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_423),
.B(n_399),
.C(n_396),
.Y(n_467)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_467),
.B(n_440),
.C(n_444),
.Y(n_475)
);

AOI21xp5_ASAP7_75t_L g491 ( 
.A1(n_468),
.A2(n_479),
.B(n_349),
.Y(n_491)
);

AOI21xp5_ASAP7_75t_L g470 ( 
.A1(n_448),
.A2(n_445),
.B(n_432),
.Y(n_470)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_470),
.A2(n_461),
.B(n_326),
.Y(n_489)
);

XOR2xp5_ASAP7_75t_L g493 ( 
.A(n_471),
.B(n_322),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_452),
.A2(n_441),
.B1(n_440),
.B2(n_423),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g486 ( 
.A(n_472),
.B(n_475),
.Y(n_486)
);

MAJIxp5_ASAP7_75t_L g478 ( 
.A(n_450),
.B(n_446),
.C(n_444),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g488 ( 
.A(n_478),
.B(n_481),
.C(n_482),
.Y(n_488)
);

OAI22xp5_ASAP7_75t_SL g480 ( 
.A1(n_457),
.A2(n_399),
.B1(n_396),
.B2(n_395),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g484 ( 
.A1(n_480),
.A2(n_451),
.B1(n_459),
.B2(n_465),
.Y(n_484)
);

MAJIxp5_ASAP7_75t_L g481 ( 
.A(n_450),
.B(n_321),
.C(n_258),
.Y(n_481)
);

MAJIxp5_ASAP7_75t_L g482 ( 
.A(n_467),
.B(n_447),
.C(n_460),
.Y(n_482)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_447),
.B(n_256),
.Y(n_483)
);

NOR2xp33_ASAP7_75t_L g490 ( 
.A(n_483),
.B(n_461),
.Y(n_490)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_484),
.Y(n_507)
);

NOR2xp33_ASAP7_75t_SL g485 ( 
.A(n_477),
.B(n_455),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_485),
.B(n_469),
.Y(n_503)
);

AOI22xp33_ASAP7_75t_SL g487 ( 
.A1(n_474),
.A2(n_349),
.B1(n_322),
.B2(n_459),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_487),
.B(n_490),
.Y(n_498)
);

AND2x2_ASAP7_75t_L g500 ( 
.A(n_489),
.B(n_492),
.Y(n_500)
);

OAI21xp5_ASAP7_75t_L g502 ( 
.A1(n_491),
.A2(n_495),
.B(n_496),
.Y(n_502)
);

AOI22xp5_ASAP7_75t_L g492 ( 
.A1(n_480),
.A2(n_468),
.B1(n_475),
.B2(n_473),
.Y(n_492)
);

AOI22xp5_ASAP7_75t_L g506 ( 
.A1(n_493),
.A2(n_11),
.B1(n_13),
.B2(n_14),
.Y(n_506)
);

AOI22xp5_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_267),
.B1(n_257),
.B2(n_253),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g501 ( 
.A(n_494),
.B(n_497),
.Y(n_501)
);

AOI21xp5_ASAP7_75t_L g495 ( 
.A1(n_471),
.A2(n_267),
.B(n_12),
.Y(n_495)
);

AOI21xp5_ASAP7_75t_L g496 ( 
.A1(n_478),
.A2(n_17),
.B(n_12),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_482),
.B(n_17),
.C(n_12),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_488),
.B(n_483),
.C(n_476),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g509 ( 
.A(n_499),
.B(n_503),
.Y(n_509)
);

MAJIxp5_ASAP7_75t_L g504 ( 
.A(n_488),
.B(n_481),
.C(n_472),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g513 ( 
.A1(n_504),
.A2(n_506),
.B(n_13),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_492),
.B(n_11),
.Y(n_505)
);

NOR3xp33_ASAP7_75t_L g512 ( 
.A(n_505),
.B(n_497),
.C(n_494),
.Y(n_512)
);

MAJx2_ASAP7_75t_L g508 ( 
.A(n_500),
.B(n_486),
.C(n_491),
.Y(n_508)
);

OR2x2_ASAP7_75t_L g514 ( 
.A(n_508),
.B(n_512),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g510 ( 
.A1(n_500),
.A2(n_484),
.B(n_496),
.Y(n_510)
);

AOI21xp5_ASAP7_75t_L g516 ( 
.A1(n_510),
.A2(n_513),
.B(n_502),
.Y(n_516)
);

AOI21x1_ASAP7_75t_SL g511 ( 
.A1(n_507),
.A2(n_495),
.B(n_493),
.Y(n_511)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_511),
.B(n_498),
.C(n_501),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_L g515 ( 
.A(n_509),
.B(n_499),
.Y(n_515)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_515),
.A2(n_516),
.B(n_14),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_504),
.Y(n_518)
);

AOI21xp5_ASAP7_75t_L g520 ( 
.A1(n_518),
.A2(n_519),
.B(n_514),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_520),
.B(n_521),
.C(n_14),
.Y(n_522)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_518),
.B(n_14),
.C(n_15),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_15),
.B(n_16),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_15),
.C(n_16),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g525 ( 
.A(n_524),
.B(n_15),
.Y(n_525)
);


endmodule