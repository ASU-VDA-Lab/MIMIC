module real_jpeg_26257_n_18 (n_17, n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_18);

input n_17;
input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

INVxp67_ASAP7_75t_L g63 ( 
.A(n_0),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_0),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_0),
.B(n_89),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_0),
.B(n_116),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_0),
.B(n_185),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_0),
.B(n_32),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_0),
.B(n_51),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_1),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_1),
.B(n_46),
.Y(n_86)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_1),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_1),
.B(n_51),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_1),
.B(n_66),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_1),
.B(n_185),
.Y(n_274)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_SL g115 ( 
.A(n_3),
.B(n_116),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_3),
.B(n_48),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_3),
.B(n_46),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_3),
.B(n_51),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g214 ( 
.A(n_3),
.B(n_32),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_3),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_3),
.B(n_66),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_3),
.B(n_89),
.Y(n_264)
);

CKINVDCx14_ASAP7_75t_R g25 ( 
.A(n_4),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_4),
.B(n_73),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_4),
.B(n_46),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_4),
.B(n_66),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_4),
.B(n_17),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_4),
.B(n_32),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_4),
.B(n_51),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_4),
.B(n_48),
.Y(n_280)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

INVx8_ASAP7_75t_SL g27 ( 
.A(n_7),
.Y(n_27)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_8),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_8),
.B(n_51),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_9),
.B(n_32),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_9),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_9),
.B(n_48),
.Y(n_87)
);

CKINVDCx14_ASAP7_75t_R g111 ( 
.A(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_9),
.B(n_46),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_10),
.B(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_10),
.B(n_89),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_10),
.B(n_51),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g169 ( 
.A(n_10),
.B(n_48),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_10),
.B(n_32),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_10),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_10),
.B(n_46),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_10),
.B(n_66),
.Y(n_275)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

INVx13_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

CKINVDCx14_ASAP7_75t_R g58 ( 
.A(n_13),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_13),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_13),
.B(n_32),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_13),
.B(n_51),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_13),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_13),
.B(n_48),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_SL g262 ( 
.A(n_13),
.B(n_46),
.Y(n_262)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_13),
.B(n_66),
.Y(n_296)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

INVxp67_ASAP7_75t_L g60 ( 
.A(n_14),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_14),
.B(n_66),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_14),
.B(n_185),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g263 ( 
.A(n_14),
.B(n_32),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_14),
.B(n_51),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_16),
.B(n_46),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_16),
.B(n_66),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_16),
.B(n_48),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_16),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_16),
.B(n_32),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_16),
.B(n_89),
.Y(n_247)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_17),
.Y(n_114)
);

INVx6_ASAP7_75t_L g186 ( 
.A(n_17),
.Y(n_186)
);

XNOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_152),
.Y(n_18)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_123),
.Y(n_19)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_77),
.C(n_90),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g333 ( 
.A(n_21),
.B(n_77),
.Y(n_333)
);

XNOR2xp5_ASAP7_75t_SL g21 ( 
.A(n_22),
.B(n_53),
.Y(n_21)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_22),
.B(n_54),
.C(n_70),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_38),
.C(n_44),
.Y(n_22)
);

XOR2xp5_ASAP7_75t_L g326 ( 
.A(n_23),
.B(n_327),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_28),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g76 ( 
.A(n_24),
.B(n_29),
.C(n_36),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_25),
.B(n_26),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_26),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_26),
.B(n_60),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g28 ( 
.A1(n_29),
.A2(n_34),
.B1(n_36),
.B2(n_37),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_29),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_29),
.A2(n_37),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_SL g137 ( 
.A(n_29),
.B(n_79),
.C(n_82),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_31),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_SL g34 ( 
.A(n_30),
.B(n_35),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_30),
.B(n_61),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_31),
.B(n_120),
.Y(n_119)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_34),
.A2(n_36),
.B1(n_39),
.B2(n_103),
.Y(n_102)
);

INVx5_ASAP7_75t_L g198 ( 
.A(n_35),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_36),
.B(n_39),
.C(n_40),
.Y(n_38)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_38),
.B(n_44),
.Y(n_327)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_39),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_40),
.A2(n_41),
.B1(n_101),
.B2(n_102),
.Y(n_100)
);

CKINVDCx16_ASAP7_75t_R g40 ( 
.A(n_41),
.Y(n_40)
);

INVx11_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

INVx6_ASAP7_75t_L g118 ( 
.A(n_43),
.Y(n_118)
);

BUFx24_ASAP7_75t_SL g337 ( 
.A(n_44),
.Y(n_337)
);

FAx1_ASAP7_75t_SL g44 ( 
.A(n_45),
.B(n_47),
.CI(n_50),
.CON(n_44),
.SN(n_44)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_45),
.B(n_47),
.C(n_50),
.Y(n_84)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_46),
.Y(n_64)
);

INVx8_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx13_ASAP7_75t_L g219 ( 
.A(n_51),
.Y(n_219)
);

BUFx24_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_54),
.B(n_70),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_65),
.C(n_69),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_55),
.A2(n_56),
.B1(n_105),
.B2(n_107),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_56),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_57),
.B(n_59),
.C(n_62),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g93 ( 
.A(n_57),
.B(n_62),
.Y(n_93)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_59),
.B(n_93),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_61),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_63),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_64),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_65),
.A2(n_72),
.B1(n_74),
.B2(n_75),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_65),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g105 ( 
.A1(n_65),
.A2(n_69),
.B1(n_75),
.B2(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_65),
.B(n_74),
.C(n_76),
.Y(n_143)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_69),
.Y(n_106)
);

XOR2xp5_ASAP7_75t_L g70 ( 
.A(n_71),
.B(n_76),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_72),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_78),
.B(n_83),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_78),
.B(n_84),
.C(n_85),
.Y(n_140)
);

XOR2xp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_80),
.Y(n_78)
);

AOI22xp33_ASAP7_75t_L g131 ( 
.A1(n_81),
.A2(n_82),
.B1(n_132),
.B2(n_133),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_82),
.Y(n_81)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_85),
.Y(n_83)
);

BUFx24_ASAP7_75t_SL g334 ( 
.A(n_85),
.Y(n_334)
);

FAx1_ASAP7_75t_SL g85 ( 
.A(n_86),
.B(n_87),
.CI(n_88),
.CON(n_85),
.SN(n_85)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_86),
.B(n_87),
.C(n_88),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_90),
.B(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_104),
.C(n_108),
.Y(n_90)
);

XOR2xp5_ASAP7_75t_L g328 ( 
.A(n_91),
.B(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_92),
.B(n_94),
.C(n_100),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_92),
.B(n_312),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_94),
.B(n_100),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_97),
.C(n_98),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_95),
.A2(n_96),
.B1(n_98),
.B2(n_99),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_97),
.B(n_291),
.Y(n_290)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g329 ( 
.A(n_104),
.B(n_108),
.Y(n_329)
);

INVx1_ASAP7_75t_L g107 ( 
.A(n_105),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_109),
.B(n_121),
.C(n_122),
.Y(n_108)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_109),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_115),
.C(n_119),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g305 ( 
.A(n_110),
.B(n_119),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_112),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_SL g304 ( 
.A(n_115),
.B(n_305),
.Y(n_304)
);

INVx8_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_117),
.B(n_218),
.Y(n_278)
);

INVx8_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_121),
.B(n_122),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_125),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_138),
.B2(n_139),
.Y(n_125)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_129),
.B1(n_134),
.B2(n_135),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_131),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_132),
.Y(n_133)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_135),
.Y(n_134)
);

XOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_137),
.Y(n_135)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_142),
.A2(n_143),
.B1(n_144),
.B2(n_145),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_143),
.Y(n_142)
);

CKINVDCx16_ASAP7_75t_R g144 ( 
.A(n_145),
.Y(n_144)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_146),
.B(n_147),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g147 ( 
.A1(n_148),
.A2(n_149),
.B1(n_150),
.B2(n_151),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g148 ( 
.A(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g151 ( 
.A(n_150),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_331),
.C(n_332),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_321),
.C(n_322),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_307),
.C(n_308),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_284),
.C(n_285),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_254),
.C(n_255),
.Y(n_156)
);

MAJIxp5_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_229),
.C(n_230),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_188),
.C(n_200),
.Y(n_158)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_160),
.B(n_173),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_168),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_161),
.B(n_168),
.C(n_173),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.C(n_166),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g189 ( 
.A1(n_162),
.A2(n_163),
.B1(n_190),
.B2(n_191),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g162 ( 
.A(n_163),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_164),
.A2(n_165),
.B1(n_166),
.B2(n_167),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_165),
.Y(n_164)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_169),
.B(n_170),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_169),
.B(n_171),
.C(n_172),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_172),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_179),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_174),
.B(n_180),
.C(n_181),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_SL g199 ( 
.A1(n_175),
.A2(n_176),
.B1(n_177),
.B2(n_178),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_176),
.Y(n_175)
);

CKINVDCx16_ASAP7_75t_R g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_182),
.A2(n_183),
.B1(n_184),
.B2(n_187),
.Y(n_181)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_182),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_183),
.B(n_187),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g183 ( 
.A(n_184),
.Y(n_183)
);

INVx5_ASAP7_75t_L g224 ( 
.A(n_185),
.Y(n_224)
);

INVx8_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

INVx5_ASAP7_75t_L g212 ( 
.A(n_186),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_189),
.B(n_192),
.C(n_199),
.Y(n_188)
);

XNOR2xp5_ASAP7_75t_L g226 ( 
.A(n_189),
.B(n_227),
.Y(n_226)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_191),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_L g227 ( 
.A1(n_192),
.A2(n_193),
.B1(n_199),
.B2(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_196),
.Y(n_193)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_197),
.Y(n_204)
);

CKINVDCx16_ASAP7_75t_R g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_199),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_225),
.C(n_226),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_209),
.C(n_215),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_SL g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g225 ( 
.A(n_203),
.B(n_207),
.C(n_208),
.Y(n_225)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_210),
.B(n_213),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_210),
.A2(n_211),
.B1(n_213),
.B2(n_214),
.Y(n_216)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_211),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g213 ( 
.A(n_214),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_216),
.B(n_217),
.C(n_220),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_219),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_L g220 ( 
.A(n_221),
.B(n_222),
.Y(n_220)
);

INVx3_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_243),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_244),
.C(n_253),
.Y(n_254)
);

XNOR2xp5_ASAP7_75t_SL g231 ( 
.A(n_232),
.B(n_239),
.Y(n_231)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_238),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g258 ( 
.A(n_233),
.B(n_238),
.C(n_239),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_SL g233 ( 
.A1(n_234),
.A2(n_235),
.B1(n_236),
.B2(n_237),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_234),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_235),
.B(n_237),
.Y(n_267)
);

CKINVDCx16_ASAP7_75t_R g235 ( 
.A(n_236),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g336 ( 
.A(n_239),
.Y(n_336)
);

FAx1_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_241),
.CI(n_242),
.CON(n_239),
.SN(n_239)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_240),
.B(n_241),
.C(n_242),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_244),
.B(n_253),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g244 ( 
.A1(n_245),
.A2(n_246),
.B1(n_251),
.B2(n_252),
.Y(n_244)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_246),
.Y(n_245)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_247),
.A2(n_248),
.B1(n_249),
.B2(n_250),
.Y(n_246)
);

CKINVDCx16_ASAP7_75t_R g250 ( 
.A(n_247),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_248),
.B(n_250),
.C(n_252),
.Y(n_271)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_251),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g255 ( 
.A(n_256),
.B(n_270),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_258),
.B1(n_259),
.B2(n_260),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_258),
.B(n_259),
.C(n_270),
.Y(n_284)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_265),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_261),
.B(n_266),
.C(n_269),
.Y(n_288)
);

BUFx24_ASAP7_75t_SL g338 ( 
.A(n_261),
.Y(n_338)
);

FAx1_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_263),
.CI(n_264),
.CON(n_261),
.SN(n_261)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_262),
.B(n_263),
.C(n_264),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_266),
.A2(n_267),
.B1(n_268),
.B2(n_269),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

CKINVDCx16_ASAP7_75t_R g268 ( 
.A(n_269),
.Y(n_268)
);

XNOR2xp5_ASAP7_75t_SL g270 ( 
.A(n_271),
.B(n_272),
.Y(n_270)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_271),
.B(n_277),
.C(n_282),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g272 ( 
.A1(n_273),
.A2(n_277),
.B1(n_282),
.B2(n_283),
.Y(n_272)
);

CKINVDCx20_ASAP7_75t_R g282 ( 
.A(n_273),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_274),
.A2(n_275),
.B(n_276),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_274),
.B(n_275),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_303),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_276),
.B(n_303),
.C(n_304),
.Y(n_314)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_277),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_278),
.B(n_280),
.C(n_281),
.Y(n_298)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_280),
.B(n_281),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_299),
.B2(n_306),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_286),
.B(n_300),
.C(n_301),
.Y(n_307)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

XNOR2xp5_ASAP7_75t_SL g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_288),
.B(n_290),
.C(n_292),
.Y(n_309)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_292),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_298),
.Y(n_292)
);

AOI22xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_295),
.B1(n_296),
.B2(n_297),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_294),
.B(n_297),
.C(n_298),
.Y(n_316)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_295),
.Y(n_294)
);

CKINVDCx20_ASAP7_75t_R g297 ( 
.A(n_296),
.Y(n_297)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_299),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_SL g299 ( 
.A(n_300),
.B(n_301),
.Y(n_299)
);

XNOR2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_304),
.Y(n_301)
);

AOI22xp5_ASAP7_75t_L g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_319),
.B2(n_320),
.Y(n_308)
);

CKINVDCx14_ASAP7_75t_R g319 ( 
.A(n_309),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_310),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g310 ( 
.A(n_311),
.B(n_313),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_311),
.B(n_313),
.C(n_319),
.Y(n_321)
);

XNOR2xp5_ASAP7_75t_L g313 ( 
.A(n_314),
.B(n_315),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_314),
.B(n_316),
.C(n_317),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_L g322 ( 
.A(n_323),
.B(n_324),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_325),
.C(n_330),
.Y(n_331)
);

AOI22xp5_ASAP7_75t_L g324 ( 
.A1(n_325),
.A2(n_326),
.B1(n_328),
.B2(n_330),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_326),
.Y(n_325)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_328),
.Y(n_330)
);


endmodule