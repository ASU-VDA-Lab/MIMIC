module fake_jpeg_13058_n_69 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_69);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_69;

wire n_13;
wire n_21;
wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_55;
wire n_64;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_62;
wire n_25;
wire n_17;
wire n_31;
wire n_56;
wire n_67;
wire n_37;
wire n_29;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_15;
wire n_66;

INVx1_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_2),
.Y(n_10)
);

INVx13_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

BUFx12f_ASAP7_75t_L g12 ( 
.A(n_6),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_8),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_6),
.Y(n_14)
);

INVx4_ASAP7_75t_SL g15 ( 
.A(n_2),
.Y(n_15)
);

NOR2xp33_ASAP7_75t_L g16 ( 
.A(n_2),
.B(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_7),
.Y(n_17)
);

CKINVDCx5p33_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_18),
.B(n_19),
.Y(n_27)
);

OR2x4_ASAP7_75t_L g19 ( 
.A(n_15),
.B(n_0),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_L g20 ( 
.A(n_16),
.B(n_0),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_20),
.B(n_10),
.Y(n_25)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_15),
.Y(n_21)
);

INVx6_ASAP7_75t_L g26 ( 
.A(n_21),
.Y(n_26)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_22),
.Y(n_30)
);

INVx5_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_23),
.B(n_24),
.Y(n_29)
);

INVx11_ASAP7_75t_L g24 ( 
.A(n_15),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g35 ( 
.A(n_25),
.B(n_17),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_20),
.B(n_9),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_28),
.B(n_10),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g31 ( 
.A(n_19),
.B(n_17),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_31),
.B(n_18),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_32),
.B(n_33),
.Y(n_43)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_30),
.Y(n_34)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_35),
.B(n_13),
.Y(n_45)
);

CKINVDCx14_ASAP7_75t_R g36 ( 
.A(n_27),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g41 ( 
.A(n_36),
.B(n_37),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g37 ( 
.A(n_30),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_21),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_38),
.B(n_39),
.Y(n_44)
);

AND2x2_ASAP7_75t_L g39 ( 
.A(n_25),
.B(n_21),
.Y(n_39)
);

AOI21xp5_ASAP7_75t_L g42 ( 
.A1(n_38),
.A2(n_29),
.B(n_24),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_42),
.B(n_26),
.C(n_11),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_47),
.Y(n_52)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_33),
.B(n_22),
.Y(n_46)
);

XNOR2xp5_ASAP7_75t_SL g50 ( 
.A(n_46),
.B(n_24),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_37),
.Y(n_47)
);

AOI22xp5_ASAP7_75t_L g48 ( 
.A1(n_40),
.A2(n_14),
.B1(n_13),
.B2(n_23),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_48),
.B(n_49),
.Y(n_55)
);

INVxp33_ASAP7_75t_SL g49 ( 
.A(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_50),
.B(n_51),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_44),
.A2(n_12),
.B1(n_14),
.B2(n_21),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_53),
.B(n_42),
.C(n_26),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_52),
.B(n_43),
.Y(n_54)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_54),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_49),
.C(n_46),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_56),
.B(n_57),
.C(n_12),
.Y(n_60)
);

A2O1A1Ixp33_ASAP7_75t_SL g59 ( 
.A1(n_58),
.A2(n_0),
.B(n_1),
.C(n_12),
.Y(n_59)
);

AOI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_59),
.A2(n_3),
.B(n_5),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_60),
.B(n_1),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_61),
.B(n_55),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_62),
.Y(n_66)
);

AOI31xp67_ASAP7_75t_L g65 ( 
.A1(n_63),
.A2(n_64),
.A3(n_3),
.B(n_5),
.Y(n_65)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_65),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_66),
.B(n_7),
.Y(n_68)
);

XNOR2xp5_ASAP7_75t_L g69 ( 
.A(n_68),
.B(n_8),
.Y(n_69)
);


endmodule