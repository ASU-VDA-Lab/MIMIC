module fake_jpeg_12186_n_93 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_93);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_93;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_22;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

INVx1_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_9),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

BUFx3_ASAP7_75t_L g14 ( 
.A(n_5),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

BUFx2_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx8_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

INVxp67_ASAP7_75t_L g21 ( 
.A(n_1),
.Y(n_21)
);

INVx2_ASAP7_75t_R g22 ( 
.A(n_8),
.Y(n_22)
);

AOI22xp33_ASAP7_75t_SL g23 ( 
.A1(n_16),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_23)
);

AOI22xp33_ASAP7_75t_SL g41 ( 
.A1(n_23),
.A2(n_29),
.B1(n_13),
.B2(n_14),
.Y(n_41)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_24),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_19),
.Y(n_25)
);

INVx5_ASAP7_75t_L g39 ( 
.A(n_25),
.Y(n_39)
);

INVx5_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_27),
.Y(n_32)
);

AOI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g37 ( 
.A(n_28),
.B(n_22),
.Y(n_37)
);

AOI22xp33_ASAP7_75t_L g29 ( 
.A1(n_16),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_20),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_30),
.B(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_21),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_31),
.B(n_22),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_SL g51 ( 
.A(n_33),
.B(n_38),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_41),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_18),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_27),
.B(n_18),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g43 ( 
.A(n_40),
.B(n_12),
.Y(n_43)
);

INVx1_ASAP7_75t_SL g42 ( 
.A(n_34),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_50),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g60 ( 
.A(n_43),
.B(n_52),
.Y(n_60)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_39),
.Y(n_44)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_44),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_38),
.A2(n_37),
.B1(n_25),
.B2(n_39),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_46),
.B(n_30),
.Y(n_59)
);

AOI32xp33_ASAP7_75t_L g47 ( 
.A1(n_33),
.A2(n_13),
.A3(n_30),
.B1(n_12),
.B2(n_11),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_47),
.B(n_53),
.Y(n_58)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_32),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g49 ( 
.A1(n_36),
.A2(n_25),
.B1(n_26),
.B2(n_19),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_49),
.A2(n_30),
.B1(n_26),
.B2(n_34),
.Y(n_55)
);

OAI21xp5_ASAP7_75t_L g50 ( 
.A1(n_36),
.A2(n_24),
.B(n_11),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_40),
.B(n_15),
.Y(n_52)
);

INVxp67_ASAP7_75t_SL g53 ( 
.A(n_39),
.Y(n_53)
);

INVxp67_ASAP7_75t_L g67 ( 
.A(n_55),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_32),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_56),
.B(n_61),
.Y(n_69)
);

INVxp67_ASAP7_75t_L g71 ( 
.A(n_59),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_51),
.B(n_14),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_6),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_62),
.B(n_7),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_64),
.B(n_66),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g65 ( 
.A(n_60),
.B(n_57),
.Y(n_65)
);

XNOR2xp5_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_69),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_57),
.B(n_46),
.Y(n_66)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_54),
.Y(n_68)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_68),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g70 ( 
.A(n_63),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_70),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_72),
.B(n_77),
.C(n_74),
.Y(n_80)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_67),
.A2(n_58),
.B(n_45),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_73),
.B(n_76),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g77 ( 
.A(n_71),
.B(n_59),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_71),
.A2(n_55),
.B1(n_49),
.B2(n_42),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_67),
.B1(n_44),
.B2(n_68),
.Y(n_82)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_79),
.B(n_80),
.Y(n_84)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_75),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_72),
.B(n_8),
.Y(n_83)
);

OAI21xp5_ASAP7_75t_L g85 ( 
.A1(n_83),
.A2(n_35),
.B(n_78),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_SL g89 ( 
.A(n_85),
.B(n_17),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_84),
.B(n_80),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_87),
.B(n_88),
.Y(n_90)
);

NAND2xp33_ASAP7_75t_L g88 ( 
.A(n_86),
.B(n_77),
.Y(n_88)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_89),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g92 ( 
.A1(n_90),
.A2(n_91),
.B(n_35),
.Y(n_92)
);

XOR2xp5_ASAP7_75t_L g93 ( 
.A(n_92),
.B(n_17),
.Y(n_93)
);


endmodule