module fake_netlist_1_1645_n_8 (n_3, n_1, n_2, n_0, n_8);
input n_3;
input n_1;
input n_2;
input n_0;
output n_8;
wire n_6;
wire n_4;
wire n_5;
wire n_7;
NOR2xp33_ASAP7_75t_R g4 ( .A(n_0), .B(n_2), .Y(n_4) );
CKINVDCx5p33_ASAP7_75t_R g5 ( .A(n_2), .Y(n_5) );
NAND2xp5_ASAP7_75t_L g6 ( .A(n_5), .B(n_3), .Y(n_6) );
OAI211xp5_ASAP7_75t_SL g7 ( .A1(n_6), .A2(n_4), .B(n_1), .C(n_3), .Y(n_7) );
AOI22xp5_ASAP7_75t_L g8 ( .A1(n_7), .A2(n_4), .B1(n_0), .B2(n_1), .Y(n_8) );
endmodule