module real_jpeg_6275_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_425;
wire n_50;
wire n_409;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_339;
wire n_326;
wire n_80;
wire n_30;
wire n_332;
wire n_149;
wire n_328;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_423;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_378;
wire n_98;
wire n_200;
wire n_432;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_383;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_18;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_450;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AND2x2_ASAP7_75t_SL g24 ( 
.A(n_0),
.B(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_0),
.B(n_45),
.Y(n_44)
);

AND2x2_ASAP7_75t_SL g62 ( 
.A(n_0),
.B(n_63),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_0),
.B(n_81),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_0),
.B(n_51),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_0),
.B(n_122),
.Y(n_121)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_0),
.Y(n_150)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_2),
.B(n_220),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_246),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_2),
.B(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g265 ( 
.A(n_2),
.B(n_266),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_2),
.B(n_301),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_2),
.B(n_114),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g386 ( 
.A(n_2),
.Y(n_386)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_3),
.B(n_51),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_3),
.B(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g225 ( 
.A(n_3),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_3),
.B(n_258),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g326 ( 
.A(n_3),
.B(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_3),
.B(n_360),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_3),
.B(n_163),
.Y(n_404)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_4),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g138 ( 
.A(n_4),
.Y(n_138)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_4),
.Y(n_256)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_5),
.Y(n_72)
);

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_6),
.B(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_6),
.Y(n_55)
);

AND2x2_ASAP7_75t_L g70 ( 
.A(n_6),
.B(n_71),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_6),
.B(n_74),
.Y(n_73)
);

AND2x2_ASAP7_75t_SL g106 ( 
.A(n_6),
.B(n_107),
.Y(n_106)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_6),
.B(n_114),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_6),
.B(n_145),
.Y(n_144)
);

AND2x2_ASAP7_75t_L g180 ( 
.A(n_6),
.B(n_181),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_7),
.Y(n_63)
);

INVx8_ASAP7_75t_L g148 ( 
.A(n_7),
.Y(n_148)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_7),
.Y(n_233)
);

BUFx6f_ASAP7_75t_L g260 ( 
.A(n_7),
.Y(n_260)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_7),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g376 ( 
.A(n_7),
.Y(n_376)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_8),
.Y(n_83)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_8),
.Y(n_115)
);

BUFx5_ASAP7_75t_L g163 ( 
.A(n_8),
.Y(n_163)
);

BUFx5_ASAP7_75t_L g378 ( 
.A(n_8),
.Y(n_378)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_9),
.Y(n_41)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_10),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g60 ( 
.A(n_10),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_10),
.Y(n_154)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_10),
.Y(n_182)
);

AND2x2_ASAP7_75t_L g153 ( 
.A(n_11),
.B(n_154),
.Y(n_153)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_11),
.B(n_211),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_11),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_11),
.B(n_253),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_11),
.B(n_270),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_11),
.B(n_299),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_11),
.B(n_318),
.Y(n_317)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_11),
.A2(n_373),
.B(n_378),
.Y(n_377)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_12),
.Y(n_49)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

BUFx5_ASAP7_75t_L g122 ( 
.A(n_12),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g287 ( 
.A(n_12),
.Y(n_287)
);

AND2x2_ASAP7_75t_L g59 ( 
.A(n_13),
.B(n_60),
.Y(n_59)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_13),
.B(n_88),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_13),
.B(n_161),
.Y(n_160)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_13),
.Y(n_230)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_13),
.B(n_227),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_13),
.B(n_287),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_13),
.B(n_332),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_13),
.B(n_383),
.Y(n_382)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_14),
.B(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_14),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_14),
.B(n_103),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_14),
.B(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_14),
.B(n_196),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g374 ( 
.A(n_14),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_15),
.B(n_77),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_15),
.B(n_88),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_15),
.B(n_156),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_15),
.B(n_192),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_15),
.B(n_316),
.Y(n_315)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_15),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g403 ( 
.A(n_15),
.B(n_287),
.Y(n_403)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_201),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_199),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_167),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_19),
.B(n_167),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_96),
.C(n_124),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_20),
.B(n_96),
.Y(n_428)
);

XOR2xp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_67),
.Y(n_20)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_21),
.B(n_68),
.C(n_84),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_43),
.C(n_53),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_L g422 ( 
.A(n_22),
.B(n_43),
.Y(n_422)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_24),
.B1(n_29),
.B2(n_30),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_23),
.B(n_32),
.C(n_37),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_23),
.A2(n_24),
.B1(n_119),
.B2(n_120),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_23),
.B(n_119),
.C(n_123),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g288 ( 
.A1(n_23),
.A2(n_24),
.B1(n_143),
.B2(n_144),
.Y(n_288)
);

INVx1_ASAP7_75t_SL g23 ( 
.A(n_24),
.Y(n_23)
);

NAND2xp5_ASAP7_75t_SL g321 ( 
.A(n_24),
.B(n_144),
.Y(n_321)
);

BUFx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_27),
.Y(n_75)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g228 ( 
.A(n_28),
.Y(n_228)
);

BUFx3_ASAP7_75t_L g357 ( 
.A(n_28),
.Y(n_357)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_32),
.B1(n_37),
.B2(n_42),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_36),
.Y(n_35)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_36),
.Y(n_109)
);

INVx11_ASAP7_75t_L g158 ( 
.A(n_36),
.Y(n_158)
);

INVx3_ASAP7_75t_L g247 ( 
.A(n_36),
.Y(n_247)
);

BUFx3_ASAP7_75t_L g335 ( 
.A(n_36),
.Y(n_335)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_37),
.Y(n_42)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx3_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_41),
.Y(n_46)
);

INVx6_ASAP7_75t_L g91 ( 
.A(n_41),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g197 ( 
.A(n_41),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_44),
.B(n_47),
.C(n_50),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_44),
.B(n_140),
.Y(n_139)
);

INVx4_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx6_ASAP7_75t_SL g318 ( 
.A(n_46),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_47),
.B(n_50),
.Y(n_140)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_49),
.Y(n_218)
);

INVx8_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g421 ( 
.A(n_53),
.B(n_422),
.Y(n_421)
);

OAI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_65),
.B2(n_66),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g65 ( 
.A(n_54),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_54),
.B(n_59),
.C(n_62),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_54),
.A2(n_65),
.B1(n_381),
.B2(n_382),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_54),
.B(n_382),
.C(n_385),
.Y(n_400)
);

OR2x2_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_56),
.Y(n_54)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_56),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g243 ( 
.A(n_57),
.Y(n_243)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_58),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g58 ( 
.A1(n_59),
.A2(n_61),
.B1(n_62),
.B2(n_64),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_59),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_61),
.A2(n_62),
.B1(n_73),
.B2(n_130),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_61),
.A2(n_62),
.B1(n_235),
.B2(n_236),
.Y(n_234)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_70),
.C(n_73),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g289 ( 
.A(n_62),
.B(n_236),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_68),
.B(n_84),
.Y(n_67)
);

MAJx2_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_76),
.C(n_80),
.Y(n_68)
);

XOR2xp5_ASAP7_75t_L g164 ( 
.A(n_69),
.B(n_165),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_70),
.A2(n_127),
.B1(n_128),
.B2(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_70),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_70),
.A2(n_127),
.B1(n_195),
.B2(n_198),
.Y(n_194)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_72),
.Y(n_79)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_72),
.Y(n_105)
);

INVx3_ASAP7_75t_L g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx3_ASAP7_75t_L g384 ( 
.A(n_72),
.Y(n_384)
);

CKINVDCx16_ASAP7_75t_R g130 ( 
.A(n_73),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g337 ( 
.A1(n_73),
.A2(n_130),
.B1(n_338),
.B2(n_339),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_73),
.B(n_338),
.Y(n_366)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_75),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_76),
.A2(n_80),
.B1(n_92),
.B2(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_76),
.Y(n_166)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_80),
.A2(n_86),
.B1(n_87),
.B2(n_92),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_80),
.Y(n_92)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_82),
.Y(n_81)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

INVx4_ASAP7_75t_L g193 ( 
.A(n_83),
.Y(n_193)
);

OA22x2_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_93),
.B1(n_94),
.B2(n_95),
.Y(n_84)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_87),
.B(n_92),
.C(n_95),
.Y(n_188)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx5_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g362 ( 
.A(n_91),
.Y(n_362)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_93),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g96 ( 
.A(n_97),
.B(n_116),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_99),
.Y(n_97)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_98),
.B(n_99),
.C(n_116),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_100),
.A2(n_101),
.B1(n_112),
.B2(n_113),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_102),
.A2(n_106),
.B1(n_110),
.B2(n_111),
.Y(n_101)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_102),
.Y(n_110)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_104),
.Y(n_221)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_105),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g111 ( 
.A(n_106),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_106),
.B(n_110),
.C(n_113),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g397 ( 
.A(n_106),
.B(n_133),
.Y(n_397)
);

INVx4_ASAP7_75t_SL g107 ( 
.A(n_108),
.Y(n_107)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_111),
.B(n_132),
.C(n_134),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx6_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g116 ( 
.A1(n_117),
.A2(n_118),
.B1(n_121),
.B2(n_123),
.Y(n_116)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

CKINVDCx14_ASAP7_75t_R g120 ( 
.A(n_119),
.Y(n_120)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_121),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_121),
.A2(n_123),
.B1(n_180),
.B2(n_183),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_121),
.A2(n_123),
.B1(n_326),
.B2(n_330),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g368 ( 
.A(n_121),
.B(n_326),
.C(n_331),
.Y(n_368)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_124),
.B(n_428),
.Y(n_427)
);

MAJIxp5_ASAP7_75t_L g124 ( 
.A(n_125),
.B(n_141),
.C(n_164),
.Y(n_124)
);

XNOR2x1_ASAP7_75t_L g423 ( 
.A(n_125),
.B(n_424),
.Y(n_423)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_126),
.B(n_131),
.C(n_139),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_126),
.B(n_409),
.Y(n_408)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XNOR2xp5_ASAP7_75t_L g409 ( 
.A(n_131),
.B(n_139),
.Y(n_409)
);

INVxp67_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XOR2xp5_ASAP7_75t_L g396 ( 
.A(n_134),
.B(n_397),
.Y(n_396)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx3_ASAP7_75t_SL g136 ( 
.A(n_137),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

XNOR2x1_ASAP7_75t_L g424 ( 
.A(n_141),
.B(n_164),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_155),
.C(n_159),
.Y(n_141)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_142),
.B(n_406),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_149),
.C(n_153),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_SL g415 ( 
.A1(n_143),
.A2(n_144),
.B1(n_153),
.B2(n_416),
.Y(n_415)
);

INVx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx3_ASAP7_75t_L g146 ( 
.A(n_147),
.Y(n_146)
);

INVx3_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx4_ASAP7_75t_L g316 ( 
.A(n_148),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g412 ( 
.A1(n_149),
.A2(n_413),
.B1(n_414),
.B2(n_415),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_149),
.Y(n_413)
);

OR2x2_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_151),
.Y(n_149)
);

OR2x2_ASAP7_75t_L g175 ( 
.A(n_150),
.B(n_176),
.Y(n_175)
);

INVx8_ASAP7_75t_L g329 ( 
.A(n_151),
.Y(n_329)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g416 ( 
.A(n_153),
.Y(n_416)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_154),
.Y(n_387)
);

AOI22xp5_ASAP7_75t_SL g406 ( 
.A1(n_155),
.A2(n_159),
.B1(n_160),
.B2(n_407),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_155),
.Y(n_407)
);

INVx4_ASAP7_75t_L g156 ( 
.A(n_157),
.Y(n_156)
);

INVx5_ASAP7_75t_L g157 ( 
.A(n_158),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_158),
.Y(n_177)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_158),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g295 ( 
.A(n_158),
.Y(n_295)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx6_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

XOR2xp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_169),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_184),
.Y(n_169)
);

BUFx24_ASAP7_75t_SL g451 ( 
.A(n_170),
.Y(n_451)
);

FAx1_ASAP7_75t_SL g170 ( 
.A(n_171),
.B(n_172),
.CI(n_173),
.CON(n_170),
.SN(n_170)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_174),
.A2(n_175),
.B1(n_178),
.B2(n_179),
.Y(n_173)
);

AOI22xp5_ASAP7_75t_L g358 ( 
.A1(n_174),
.A2(n_175),
.B1(n_359),
.B2(n_363),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_174),
.B(n_352),
.C(n_363),
.Y(n_398)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

INVx11_ASAP7_75t_L g176 ( 
.A(n_177),
.Y(n_176)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_180),
.Y(n_183)
);

INVx3_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_SL g184 ( 
.A(n_185),
.B(n_186),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_190),
.Y(n_186)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

XNOR2xp5_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_194),
.Y(n_190)
);

INVx6_ASAP7_75t_L g192 ( 
.A(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_193),
.B(n_240),
.Y(n_372)
);

CKINVDCx14_ASAP7_75t_R g198 ( 
.A(n_195),
.Y(n_198)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_197),
.Y(n_196)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_197),
.Y(n_303)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

AOI221xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_390),
.B1(n_444),
.B2(n_449),
.C(n_450),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g203 ( 
.A1(n_204),
.A2(n_345),
.B(n_389),
.Y(n_203)
);

AOI21xp5_ASAP7_75t_L g204 ( 
.A1(n_205),
.A2(n_306),
.B(n_344),
.Y(n_204)
);

OAI21xp5_ASAP7_75t_L g205 ( 
.A1(n_206),
.A2(n_281),
.B(n_305),
.Y(n_205)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_207),
.A2(n_248),
.B(n_280),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_SL g207 ( 
.A(n_208),
.B(n_237),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_208),
.B(n_237),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_209),
.B(n_222),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_209),
.B(n_223),
.C(n_234),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_214),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_210),
.B(n_215),
.C(n_219),
.Y(n_291)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_212),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_219),
.Y(n_214)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g217 ( 
.A(n_218),
.Y(n_217)
);

INVx3_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_234),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_229),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_224),
.B(n_229),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_225),
.B(n_226),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g293 ( 
.A(n_225),
.B(n_294),
.Y(n_293)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

INVx4_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx8_ASAP7_75t_L g268 ( 
.A(n_228),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_231),
.Y(n_229)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

INVx3_ASAP7_75t_L g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_235),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g237 ( 
.A(n_238),
.B(n_239),
.C(n_244),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g276 ( 
.A(n_238),
.B(n_277),
.Y(n_276)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_239),
.A2(n_244),
.B1(n_245),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_239),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

INVx2_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_245),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g246 ( 
.A(n_247),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_249),
.A2(n_274),
.B(n_279),
.Y(n_248)
);

AOI21xp5_ASAP7_75t_L g249 ( 
.A1(n_250),
.A2(n_264),
.B(n_273),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g250 ( 
.A(n_251),
.B(n_261),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_261),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_252),
.B(n_257),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_252),
.B(n_257),
.Y(n_275)
);

INVx2_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx2_ASAP7_75t_L g254 ( 
.A(n_255),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_259),
.Y(n_258)
);

INVx3_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_269),
.Y(n_264)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_267),
.Y(n_266)
);

INVx4_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx2_ASAP7_75t_L g270 ( 
.A(n_271),
.Y(n_270)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_275),
.B(n_276),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_282),
.B(n_283),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_282),
.B(n_283),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_290),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_284),
.B(n_291),
.C(n_292),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_289),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_286),
.B(n_288),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_286),
.B(n_288),
.C(n_289),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_293),
.B(n_296),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_293),
.B(n_297),
.C(n_304),
.Y(n_340)
);

INVx4_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g296 ( 
.A1(n_297),
.A2(n_298),
.B1(n_300),
.B2(n_304),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_300),
.Y(n_304)
);

INVx4_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

INVx3_ASAP7_75t_L g302 ( 
.A(n_303),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_343),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g344 ( 
.A(n_307),
.B(n_343),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_323),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g308 ( 
.A1(n_309),
.A2(n_310),
.B1(n_311),
.B2(n_312),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_309),
.B(n_312),
.C(n_323),
.Y(n_346)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_312),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_313),
.A2(n_320),
.B1(n_321),
.B2(n_322),
.Y(n_312)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_313),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_314),
.A2(n_315),
.B1(n_317),
.B2(n_319),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_314),
.B(n_319),
.C(n_320),
.Y(n_388)
);

CKINVDCx14_ASAP7_75t_R g314 ( 
.A(n_315),
.Y(n_314)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_317),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_336),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_324),
.B(n_340),
.C(n_342),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g324 ( 
.A(n_325),
.B(n_331),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_326),
.Y(n_330)
);

INVx2_ASAP7_75t_L g327 ( 
.A(n_328),
.Y(n_327)
);

INVx4_ASAP7_75t_L g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

INVx2_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

INVx3_ASAP7_75t_L g334 ( 
.A(n_335),
.Y(n_334)
);

AOI22xp5_ASAP7_75t_L g336 ( 
.A1(n_337),
.A2(n_340),
.B1(n_341),
.B2(n_342),
.Y(n_336)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_337),
.Y(n_342)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_346),
.B(n_347),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g347 ( 
.A(n_348),
.B(n_369),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g348 ( 
.A(n_349),
.B(n_350),
.Y(n_348)
);

MAJIxp5_ASAP7_75t_L g441 ( 
.A(n_349),
.B(n_350),
.C(n_369),
.Y(n_441)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_364),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_351),
.B(n_365),
.C(n_368),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g351 ( 
.A(n_352),
.B(n_358),
.Y(n_351)
);

NOR2xp33_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_354),
.Y(n_352)
);

INVx2_ASAP7_75t_L g354 ( 
.A(n_355),
.Y(n_354)
);

INVx4_ASAP7_75t_L g355 ( 
.A(n_356),
.Y(n_355)
);

BUFx6f_ASAP7_75t_L g356 ( 
.A(n_357),
.Y(n_356)
);

INVx1_ASAP7_75t_L g363 ( 
.A(n_359),
.Y(n_363)
);

INVx6_ASAP7_75t_L g360 ( 
.A(n_361),
.Y(n_360)
);

INVx5_ASAP7_75t_L g361 ( 
.A(n_362),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g364 ( 
.A1(n_365),
.A2(n_366),
.B1(n_367),
.B2(n_368),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_366),
.Y(n_365)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_368),
.Y(n_367)
);

XOR2xp5_ASAP7_75t_L g369 ( 
.A(n_370),
.B(n_388),
.Y(n_369)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_371),
.B(n_379),
.Y(n_370)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_371),
.B(n_379),
.C(n_388),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g371 ( 
.A1(n_372),
.A2(n_373),
.B(n_377),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_374),
.B(n_375),
.Y(n_373)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_376),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g402 ( 
.A(n_377),
.B(n_403),
.C(n_404),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g417 ( 
.A(n_377),
.B(n_418),
.Y(n_417)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_380),
.B(n_385),
.Y(n_379)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_382),
.Y(n_381)
);

INVx6_ASAP7_75t_L g383 ( 
.A(n_384),
.Y(n_383)
);

NOR2xp33_ASAP7_75t_L g385 ( 
.A(n_386),
.B(n_387),
.Y(n_385)
);

NOR3xp33_ASAP7_75t_SL g390 ( 
.A(n_391),
.B(n_426),
.C(n_430),
.Y(n_390)
);

OAI21xp5_ASAP7_75t_SL g444 ( 
.A1(n_391),
.A2(n_445),
.B(n_448),
.Y(n_444)
);

AND2x2_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_419),
.Y(n_391)
);

OR2x2_ASAP7_75t_L g448 ( 
.A(n_392),
.B(n_419),
.Y(n_448)
);

MAJIxp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_408),
.C(n_410),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g439 ( 
.A(n_393),
.B(n_408),
.Y(n_439)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_394),
.B(n_401),
.Y(n_393)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_394),
.B(n_402),
.C(n_405),
.Y(n_425)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.C(n_399),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_396),
.Y(n_395)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_396),
.B(n_400),
.Y(n_437)
);

XOR2xp5_ASAP7_75t_L g436 ( 
.A(n_398),
.B(n_437),
.Y(n_436)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_400),
.Y(n_399)
);

XNOR2xp5_ASAP7_75t_L g401 ( 
.A(n_402),
.B(n_405),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_403),
.B(n_404),
.Y(n_418)
);

XOR2xp5_ASAP7_75t_L g438 ( 
.A(n_410),
.B(n_439),
.Y(n_438)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.C(n_417),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g433 ( 
.A(n_411),
.B(n_434),
.Y(n_433)
);

XNOR2xp5_ASAP7_75t_L g434 ( 
.A(n_412),
.B(n_417),
.Y(n_434)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_415),
.Y(n_414)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_420),
.B(n_425),
.Y(n_419)
);

XNOR2xp5_ASAP7_75t_L g420 ( 
.A(n_421),
.B(n_423),
.Y(n_420)
);

MAJIxp5_ASAP7_75t_L g429 ( 
.A(n_421),
.B(n_423),
.C(n_425),
.Y(n_429)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_426),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_429),
.Y(n_426)
);

AND2x2_ASAP7_75t_L g450 ( 
.A(n_427),
.B(n_429),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g430 ( 
.A(n_431),
.B(n_440),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g445 ( 
.A1(n_431),
.A2(n_446),
.B(n_447),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_L g431 ( 
.A(n_432),
.B(n_438),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_L g447 ( 
.A(n_432),
.B(n_438),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_433),
.B(n_435),
.C(n_436),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g442 ( 
.A(n_433),
.B(n_443),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_L g443 ( 
.A(n_435),
.B(n_436),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_442),
.Y(n_440)
);

NOR2xp33_ASAP7_75t_L g446 ( 
.A(n_441),
.B(n_442),
.Y(n_446)
);


endmodule