module fake_aes_7411_n_22 (n_1, n_2, n_4, n_3, n_5, n_0, n_22);
input n_1;
input n_2;
input n_4;
input n_3;
input n_5;
input n_0;
output n_22;
wire n_20;
wire n_8;
wire n_11;
wire n_16;
wire n_13;
wire n_18;
wire n_12;
wire n_9;
wire n_17;
wire n_14;
wire n_10;
wire n_15;
wire n_19;
wire n_21;
wire n_6;
wire n_7;
INVx1_ASAP7_75t_L g6 ( .A(n_1), .Y(n_6) );
NAND2xp5_ASAP7_75t_L g7 ( .A(n_5), .B(n_4), .Y(n_7) );
CKINVDCx5p33_ASAP7_75t_R g8 ( .A(n_0), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_3), .B(n_0), .Y(n_9) );
BUFx6f_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
NAND2xp5_ASAP7_75t_L g11 ( .A(n_6), .B(n_1), .Y(n_11) );
BUFx6f_ASAP7_75t_L g12 ( .A(n_9), .Y(n_12) );
AO31x2_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_7), .A3(n_9), .B(n_8), .Y(n_13) );
INVx1_ASAP7_75t_L g14 ( .A(n_12), .Y(n_14) );
AND2x2_ASAP7_75t_L g15 ( .A(n_13), .B(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_14), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_16), .Y(n_17) );
OR2x2_ASAP7_75t_L g18 ( .A(n_17), .B(n_15), .Y(n_18) );
BUFx2_ASAP7_75t_L g19 ( .A(n_18), .Y(n_19) );
INVx1_ASAP7_75t_SL g20 ( .A(n_18), .Y(n_20) );
XOR2xp5_ASAP7_75t_L g21 ( .A(n_20), .B(n_2), .Y(n_21) );
AOI22xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_19), .B1(n_10), .B2(n_13), .Y(n_22) );
endmodule