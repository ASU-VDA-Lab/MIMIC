module fake_aes_6252_n_723 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_79, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_723);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_79;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_723;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_490;
wire n_613;
wire n_247;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_191;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_446;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_621;
wire n_285;
wire n_666;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_653;
wire n_716;
wire n_260;
wire n_539;
wire n_197;
wire n_201;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_200;
wire n_208;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_717;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_722;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_132;
wire n_109;
wire n_99;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g80 ( .A(n_16), .Y(n_80) );
INVx1_ASAP7_75t_L g81 ( .A(n_22), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_27), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_6), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
CKINVDCx20_ASAP7_75t_R g86 ( .A(n_40), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_71), .Y(n_87) );
BUFx10_ASAP7_75t_L g88 ( .A(n_39), .Y(n_88) );
INVxp67_ASAP7_75t_SL g89 ( .A(n_41), .Y(n_89) );
INVxp33_ASAP7_75t_L g90 ( .A(n_59), .Y(n_90) );
INVx2_ASAP7_75t_L g91 ( .A(n_77), .Y(n_91) );
CKINVDCx5p33_ASAP7_75t_R g92 ( .A(n_45), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_69), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_47), .Y(n_94) );
CKINVDCx5p33_ASAP7_75t_R g95 ( .A(n_10), .Y(n_95) );
CKINVDCx16_ASAP7_75t_R g96 ( .A(n_7), .Y(n_96) );
INVx1_ASAP7_75t_L g97 ( .A(n_46), .Y(n_97) );
CKINVDCx20_ASAP7_75t_R g98 ( .A(n_60), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_21), .Y(n_99) );
CKINVDCx16_ASAP7_75t_R g100 ( .A(n_34), .Y(n_100) );
INVxp67_ASAP7_75t_L g101 ( .A(n_29), .Y(n_101) );
INVxp33_ASAP7_75t_SL g102 ( .A(n_0), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_72), .Y(n_103) );
CKINVDCx5p33_ASAP7_75t_R g104 ( .A(n_26), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_28), .Y(n_105) );
INVx1_ASAP7_75t_L g106 ( .A(n_20), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_32), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_48), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_68), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_20), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_51), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_44), .Y(n_112) );
INVx2_ASAP7_75t_L g113 ( .A(n_33), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_19), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_53), .Y(n_115) );
BUFx5_ASAP7_75t_L g116 ( .A(n_25), .Y(n_116) );
INVxp67_ASAP7_75t_SL g117 ( .A(n_11), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_14), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_58), .Y(n_119) );
BUFx2_ASAP7_75t_L g120 ( .A(n_52), .Y(n_120) );
INVxp67_ASAP7_75t_SL g121 ( .A(n_57), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_62), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_2), .Y(n_123) );
CKINVDCx5p33_ASAP7_75t_R g124 ( .A(n_7), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_17), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_12), .Y(n_126) );
CKINVDCx16_ASAP7_75t_R g127 ( .A(n_42), .Y(n_127) );
INVx1_ASAP7_75t_L g128 ( .A(n_37), .Y(n_128) );
BUFx6f_ASAP7_75t_L g129 ( .A(n_91), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_116), .Y(n_130) );
HB1xp67_ASAP7_75t_L g131 ( .A(n_95), .Y(n_131) );
AND2x4_ASAP7_75t_L g132 ( .A(n_120), .B(n_0), .Y(n_132) );
INVx1_ASAP7_75t_L g133 ( .A(n_81), .Y(n_133) );
AND2x4_ASAP7_75t_L g134 ( .A(n_120), .B(n_1), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_83), .Y(n_135) );
AND2x2_ASAP7_75t_L g136 ( .A(n_96), .B(n_1), .Y(n_136) );
AND2x4_ASAP7_75t_L g137 ( .A(n_91), .B(n_2), .Y(n_137) );
INVx1_ASAP7_75t_L g138 ( .A(n_87), .Y(n_138) );
BUFx2_ASAP7_75t_L g139 ( .A(n_95), .Y(n_139) );
BUFx3_ASAP7_75t_L g140 ( .A(n_116), .Y(n_140) );
CKINVDCx11_ASAP7_75t_R g141 ( .A(n_88), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_93), .Y(n_142) );
INVx2_ASAP7_75t_L g143 ( .A(n_116), .Y(n_143) );
NAND2xp5_ASAP7_75t_SL g144 ( .A(n_116), .B(n_3), .Y(n_144) );
AND2x4_ASAP7_75t_L g145 ( .A(n_113), .B(n_3), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_114), .B(n_4), .Y(n_146) );
INVx1_ASAP7_75t_L g147 ( .A(n_94), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_116), .Y(n_148) );
INVx2_ASAP7_75t_L g149 ( .A(n_116), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_97), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_116), .Y(n_151) );
INVx2_ASAP7_75t_L g152 ( .A(n_116), .Y(n_152) );
INVx2_ASAP7_75t_L g153 ( .A(n_113), .Y(n_153) );
BUFx2_ASAP7_75t_L g154 ( .A(n_114), .Y(n_154) );
INVx1_ASAP7_75t_L g155 ( .A(n_103), .Y(n_155) );
NOR2xp33_ASAP7_75t_L g156 ( .A(n_108), .B(n_4), .Y(n_156) );
INVxp67_ASAP7_75t_L g157 ( .A(n_80), .Y(n_157) );
INVx3_ASAP7_75t_L g158 ( .A(n_88), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_109), .Y(n_159) );
INVx2_ASAP7_75t_L g160 ( .A(n_111), .Y(n_160) );
BUFx8_ASAP7_75t_L g161 ( .A(n_112), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_124), .B(n_5), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_124), .B(n_5), .Y(n_163) );
BUFx6f_ASAP7_75t_L g164 ( .A(n_115), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_119), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_122), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_128), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_82), .Y(n_168) );
INVx1_ASAP7_75t_L g169 ( .A(n_84), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_88), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g171 ( .A(n_102), .B(n_6), .Y(n_171) );
INVx2_ASAP7_75t_L g172 ( .A(n_85), .Y(n_172) );
INVx4_ASAP7_75t_L g173 ( .A(n_132), .Y(n_173) );
AND2x4_ASAP7_75t_L g174 ( .A(n_132), .B(n_123), .Y(n_174) );
AND2x6_ASAP7_75t_L g175 ( .A(n_132), .B(n_126), .Y(n_175) );
INVx1_ASAP7_75t_L g176 ( .A(n_130), .Y(n_176) );
AND2x6_ASAP7_75t_L g177 ( .A(n_132), .B(n_125), .Y(n_177) );
BUFx3_ASAP7_75t_L g178 ( .A(n_170), .Y(n_178) );
INVx1_ASAP7_75t_L g179 ( .A(n_137), .Y(n_179) );
BUFx4f_ASAP7_75t_L g180 ( .A(n_137), .Y(n_180) );
AND2x4_ASAP7_75t_L g181 ( .A(n_134), .B(n_118), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_158), .B(n_90), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g183 ( .A1(n_134), .A2(n_102), .B1(n_127), .B2(n_100), .Y(n_183) );
BUFx3_ASAP7_75t_L g184 ( .A(n_170), .Y(n_184) );
AOI22xp5_ASAP7_75t_L g185 ( .A1(n_134), .A2(n_86), .B1(n_98), .B2(n_105), .Y(n_185) );
AND2x4_ASAP7_75t_L g186 ( .A(n_134), .B(n_110), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_129), .Y(n_187) );
INVx2_ASAP7_75t_L g188 ( .A(n_129), .Y(n_188) );
AND2x2_ASAP7_75t_L g189 ( .A(n_139), .B(n_99), .Y(n_189) );
INVx2_ASAP7_75t_L g190 ( .A(n_129), .Y(n_190) );
BUFx3_ASAP7_75t_L g191 ( .A(n_170), .Y(n_191) );
INVx1_ASAP7_75t_L g192 ( .A(n_137), .Y(n_192) );
AOI22xp33_ASAP7_75t_L g193 ( .A1(n_137), .A2(n_106), .B1(n_117), .B2(n_107), .Y(n_193) );
NOR3xp33_ASAP7_75t_L g194 ( .A(n_146), .B(n_101), .C(n_121), .Y(n_194) );
AND2x4_ASAP7_75t_L g195 ( .A(n_158), .B(n_89), .Y(n_195) );
INVx4_ASAP7_75t_L g196 ( .A(n_170), .Y(n_196) );
INVx1_ASAP7_75t_L g197 ( .A(n_145), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_129), .Y(n_198) );
CKINVDCx14_ASAP7_75t_R g199 ( .A(n_139), .Y(n_199) );
AND2x4_ASAP7_75t_L g200 ( .A(n_158), .B(n_107), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_129), .Y(n_201) );
INVxp67_ASAP7_75t_L g202 ( .A(n_154), .Y(n_202) );
INVx1_ASAP7_75t_L g203 ( .A(n_145), .Y(n_203) );
BUFx2_ASAP7_75t_L g204 ( .A(n_154), .Y(n_204) );
AND2x4_ASAP7_75t_L g205 ( .A(n_158), .B(n_104), .Y(n_205) );
AND2x6_ASAP7_75t_L g206 ( .A(n_145), .B(n_105), .Y(n_206) );
OAI22xp33_ASAP7_75t_L g207 ( .A1(n_162), .A2(n_98), .B1(n_86), .B2(n_104), .Y(n_207) );
AOI22xp33_ASAP7_75t_L g208 ( .A1(n_145), .A2(n_92), .B1(n_99), .B2(n_10), .Y(n_208) );
AO22x2_ASAP7_75t_L g209 ( .A1(n_136), .A2(n_8), .B1(n_9), .B2(n_11), .Y(n_209) );
AO22x2_ASAP7_75t_L g210 ( .A1(n_136), .A2(n_8), .B1(n_9), .B2(n_12), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_168), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_129), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_168), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g214 ( .A1(n_157), .A2(n_92), .B1(n_14), .B2(n_15), .Y(n_214) );
BUFx6f_ASAP7_75t_L g215 ( .A(n_140), .Y(n_215) );
INVx4_ASAP7_75t_L g216 ( .A(n_170), .Y(n_216) );
INVx1_ASAP7_75t_L g217 ( .A(n_169), .Y(n_217) );
BUFx4f_ASAP7_75t_L g218 ( .A(n_170), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_130), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_169), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_172), .Y(n_221) );
AND2x4_ASAP7_75t_L g222 ( .A(n_133), .B(n_13), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_140), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_141), .Y(n_224) );
INVx4_ASAP7_75t_L g225 ( .A(n_140), .Y(n_225) );
INVx2_ASAP7_75t_L g226 ( .A(n_130), .Y(n_226) );
AND2x6_ASAP7_75t_L g227 ( .A(n_133), .B(n_55), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_143), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_172), .Y(n_229) );
INVx3_ASAP7_75t_L g230 ( .A(n_164), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_131), .B(n_13), .Y(n_231) );
BUFx6f_ASAP7_75t_L g232 ( .A(n_164), .Y(n_232) );
BUFx3_ASAP7_75t_L g233 ( .A(n_161), .Y(n_233) );
INVx1_ASAP7_75t_L g234 ( .A(n_172), .Y(n_234) );
AND2x2_ASAP7_75t_L g235 ( .A(n_135), .B(n_16), .Y(n_235) );
OAI22xp5_ASAP7_75t_L g236 ( .A1(n_163), .A2(n_17), .B1(n_18), .B2(n_23), .Y(n_236) );
INVx2_ASAP7_75t_SL g237 ( .A(n_161), .Y(n_237) );
NOR2xp33_ASAP7_75t_L g238 ( .A(n_202), .B(n_161), .Y(n_238) );
AOI22xp33_ASAP7_75t_L g239 ( .A1(n_222), .A2(n_161), .B1(n_167), .B2(n_166), .Y(n_239) );
AND2x2_ASAP7_75t_L g240 ( .A(n_189), .B(n_135), .Y(n_240) );
NAND2xp5_ASAP7_75t_L g241 ( .A(n_195), .B(n_138), .Y(n_241) );
BUFx3_ASAP7_75t_L g242 ( .A(n_233), .Y(n_242) );
INVx3_ASAP7_75t_SL g243 ( .A(n_224), .Y(n_243) );
INVx2_ASAP7_75t_L g244 ( .A(n_232), .Y(n_244) );
AOI22xp5_ASAP7_75t_L g245 ( .A1(n_183), .A2(n_171), .B1(n_156), .B2(n_166), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_222), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_232), .Y(n_247) );
INVx3_ASAP7_75t_L g248 ( .A(n_196), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_221), .Y(n_249) );
NAND2xp5_ASAP7_75t_L g250 ( .A(n_195), .B(n_167), .Y(n_250) );
BUFx3_ASAP7_75t_L g251 ( .A(n_233), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_229), .Y(n_252) );
BUFx2_ASAP7_75t_L g253 ( .A(n_199), .Y(n_253) );
INVx2_ASAP7_75t_SL g254 ( .A(n_180), .Y(n_254) );
OR2x6_ASAP7_75t_L g255 ( .A(n_237), .B(n_165), .Y(n_255) );
AOI22xp5_ASAP7_75t_L g256 ( .A1(n_175), .A2(n_150), .B1(n_142), .B2(n_147), .Y(n_256) );
BUFx3_ASAP7_75t_L g257 ( .A(n_178), .Y(n_257) );
O2A1O1Ixp33_ASAP7_75t_L g258 ( .A1(n_179), .A2(n_165), .B(n_138), .C(n_142), .Y(n_258) );
BUFx2_ASAP7_75t_L g259 ( .A(n_199), .Y(n_259) );
NOR2xp33_ASAP7_75t_L g260 ( .A(n_189), .B(n_150), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_234), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_195), .B(n_147), .Y(n_262) );
INVx3_ASAP7_75t_L g263 ( .A(n_196), .Y(n_263) );
AND2x4_ASAP7_75t_L g264 ( .A(n_200), .B(n_159), .Y(n_264) );
AND2x4_ASAP7_75t_L g265 ( .A(n_200), .B(n_159), .Y(n_265) );
INVx2_ASAP7_75t_L g266 ( .A(n_232), .Y(n_266) );
BUFx3_ASAP7_75t_L g267 ( .A(n_178), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_182), .B(n_155), .Y(n_268) );
INVx1_ASAP7_75t_L g269 ( .A(n_222), .Y(n_269) );
NAND2xp5_ASAP7_75t_L g270 ( .A(n_200), .B(n_155), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_235), .Y(n_271) );
INVx6_ASAP7_75t_L g272 ( .A(n_196), .Y(n_272) );
BUFx6f_ASAP7_75t_L g273 ( .A(n_227), .Y(n_273) );
AND2x4_ASAP7_75t_L g274 ( .A(n_205), .B(n_160), .Y(n_274) );
BUFx6f_ASAP7_75t_SL g275 ( .A(n_206), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_205), .B(n_160), .Y(n_276) );
INVx3_ASAP7_75t_L g277 ( .A(n_216), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_235), .Y(n_278) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_205), .B(n_160), .Y(n_279) );
CKINVDCx8_ASAP7_75t_R g280 ( .A(n_224), .Y(n_280) );
AOI22xp5_ASAP7_75t_L g281 ( .A1(n_175), .A2(n_144), .B1(n_153), .B2(n_164), .Y(n_281) );
OR2x2_ASAP7_75t_L g282 ( .A(n_204), .B(n_153), .Y(n_282) );
AO22x1_ASAP7_75t_L g283 ( .A1(n_206), .A2(n_153), .B1(n_164), .B2(n_152), .Y(n_283) );
INVx5_ASAP7_75t_L g284 ( .A(n_227), .Y(n_284) );
INVx2_ASAP7_75t_L g285 ( .A(n_232), .Y(n_285) );
AND2x2_ASAP7_75t_L g286 ( .A(n_204), .B(n_152), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_232), .Y(n_287) );
INVx3_ASAP7_75t_L g288 ( .A(n_216), .Y(n_288) );
CKINVDCx5p33_ASAP7_75t_R g289 ( .A(n_185), .Y(n_289) );
BUFx3_ASAP7_75t_L g290 ( .A(n_184), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_187), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_237), .Y(n_292) );
AND2x2_ASAP7_75t_L g293 ( .A(n_180), .B(n_152), .Y(n_293) );
OAI22xp5_ASAP7_75t_SL g294 ( .A1(n_208), .A2(n_164), .B1(n_151), .B2(n_149), .Y(n_294) );
NAND2xp5_ASAP7_75t_SL g295 ( .A(n_180), .B(n_164), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_192), .Y(n_296) );
INVx3_ASAP7_75t_L g297 ( .A(n_216), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_206), .Y(n_298) );
INVx4_ASAP7_75t_L g299 ( .A(n_175), .Y(n_299) );
INVx2_ASAP7_75t_SL g300 ( .A(n_175), .Y(n_300) );
AND2x4_ASAP7_75t_L g301 ( .A(n_174), .B(n_151), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_197), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_203), .Y(n_303) );
AND2x2_ASAP7_75t_L g304 ( .A(n_173), .B(n_151), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_211), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_174), .B(n_149), .Y(n_306) );
INVx2_ASAP7_75t_SL g307 ( .A(n_255), .Y(n_307) );
INVx2_ASAP7_75t_L g308 ( .A(n_249), .Y(n_308) );
BUFx6f_ASAP7_75t_L g309 ( .A(n_255), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g310 ( .A(n_286), .B(n_174), .Y(n_310) );
INVx2_ASAP7_75t_SL g311 ( .A(n_255), .Y(n_311) );
BUFx6f_ASAP7_75t_L g312 ( .A(n_255), .Y(n_312) );
BUFx2_ASAP7_75t_L g313 ( .A(n_253), .Y(n_313) );
BUFx2_ASAP7_75t_L g314 ( .A(n_253), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_286), .B(n_186), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g316 ( .A1(n_268), .A2(n_223), .B(n_225), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_260), .B(n_186), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_238), .B(n_207), .Y(n_318) );
INVx1_ASAP7_75t_L g319 ( .A(n_249), .Y(n_319) );
INVxp67_ASAP7_75t_SL g320 ( .A(n_242), .Y(n_320) );
BUFx2_ASAP7_75t_L g321 ( .A(n_259), .Y(n_321) );
INVx2_ASAP7_75t_L g322 ( .A(n_252), .Y(n_322) );
INVx1_ASAP7_75t_L g323 ( .A(n_252), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_261), .Y(n_324) );
INVx1_ASAP7_75t_L g325 ( .A(n_261), .Y(n_325) );
INVx2_ASAP7_75t_L g326 ( .A(n_248), .Y(n_326) );
INVx6_ASAP7_75t_L g327 ( .A(n_299), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_305), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_259), .Y(n_329) );
INVx3_ASAP7_75t_L g330 ( .A(n_299), .Y(n_330) );
NOR2xp33_ASAP7_75t_L g331 ( .A(n_240), .B(n_231), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_304), .Y(n_332) );
INVx2_ASAP7_75t_L g333 ( .A(n_248), .Y(n_333) );
INVx2_ASAP7_75t_L g334 ( .A(n_248), .Y(n_334) );
INVx1_ASAP7_75t_L g335 ( .A(n_304), .Y(n_335) );
INVx2_ASAP7_75t_L g336 ( .A(n_263), .Y(n_336) );
BUFx6f_ASAP7_75t_SL g337 ( .A(n_299), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_L g338 ( .A1(n_258), .A2(n_181), .B(n_186), .C(n_213), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_296), .Y(n_339) );
BUFx2_ASAP7_75t_L g340 ( .A(n_242), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_263), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_243), .Y(n_342) );
INVx2_ASAP7_75t_L g343 ( .A(n_263), .Y(n_343) );
INVx2_ASAP7_75t_L g344 ( .A(n_277), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_282), .B(n_231), .Y(n_345) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_240), .B(n_181), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_243), .Y(n_347) );
OAI22xp33_ASAP7_75t_L g348 ( .A1(n_289), .A2(n_173), .B1(n_220), .B2(n_217), .Y(n_348) );
NAND2xp5_ASAP7_75t_SL g349 ( .A(n_251), .B(n_173), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_282), .Y(n_350) );
BUFx6f_ASAP7_75t_L g351 ( .A(n_251), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_277), .Y(n_352) );
INVx2_ASAP7_75t_L g353 ( .A(n_277), .Y(n_353) );
NOR2xp33_ASAP7_75t_L g354 ( .A(n_245), .B(n_181), .Y(n_354) );
INVx1_ASAP7_75t_SL g355 ( .A(n_264), .Y(n_355) );
INVx2_ASAP7_75t_L g356 ( .A(n_288), .Y(n_356) );
BUFx12f_ASAP7_75t_L g357 ( .A(n_289), .Y(n_357) );
AOI22xp33_ASAP7_75t_L g358 ( .A1(n_294), .A2(n_206), .B1(n_175), .B2(n_177), .Y(n_358) );
INVx3_ASAP7_75t_L g359 ( .A(n_288), .Y(n_359) );
INVx5_ASAP7_75t_L g360 ( .A(n_273), .Y(n_360) );
NOR2xp67_ASAP7_75t_SL g361 ( .A(n_309), .B(n_284), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_308), .Y(n_362) );
CKINVDCx5p33_ASAP7_75t_R g363 ( .A(n_342), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_308), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_354), .A2(n_206), .B1(n_177), .B2(n_175), .Y(n_365) );
NOR2xp33_ASAP7_75t_L g366 ( .A(n_329), .B(n_271), .Y(n_366) );
NAND3x1_ASAP7_75t_L g367 ( .A(n_318), .B(n_209), .C(n_210), .Y(n_367) );
OR2x2_ASAP7_75t_L g368 ( .A(n_350), .B(n_270), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_308), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_338), .A2(n_269), .B(n_246), .C(n_239), .Y(n_370) );
CKINVDCx8_ASAP7_75t_R g371 ( .A(n_347), .Y(n_371) );
AND2x2_ASAP7_75t_L g372 ( .A(n_322), .B(n_264), .Y(n_372) );
AOI221xp5_ASAP7_75t_L g373 ( .A1(n_331), .A2(n_278), .B1(n_193), .B2(n_264), .C(n_265), .Y(n_373) );
INVxp67_ASAP7_75t_L g374 ( .A(n_313), .Y(n_374) );
BUFx2_ASAP7_75t_L g375 ( .A(n_309), .Y(n_375) );
BUFx2_ASAP7_75t_L g376 ( .A(n_309), .Y(n_376) );
AND2x2_ASAP7_75t_L g377 ( .A(n_322), .B(n_265), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_322), .B(n_265), .Y(n_378) );
AOI22xp33_ASAP7_75t_L g379 ( .A1(n_346), .A2(n_206), .B1(n_177), .B2(n_194), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g380 ( .A1(n_313), .A2(n_177), .B1(n_209), .B2(n_210), .Y(n_380) );
INVx8_ASAP7_75t_L g381 ( .A(n_337), .Y(n_381) );
BUFx2_ASAP7_75t_R g382 ( .A(n_314), .Y(n_382) );
BUFx6f_ASAP7_75t_L g383 ( .A(n_309), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_319), .Y(n_384) );
INVx3_ASAP7_75t_L g385 ( .A(n_309), .Y(n_385) );
A2O1A1Ixp33_ASAP7_75t_L g386 ( .A1(n_328), .A2(n_339), .B(n_325), .C(n_319), .Y(n_386) );
AOI22xp33_ASAP7_75t_L g387 ( .A1(n_314), .A2(n_177), .B1(n_209), .B2(n_210), .Y(n_387) );
INVx2_ASAP7_75t_L g388 ( .A(n_323), .Y(n_388) );
OAI22xp5_ASAP7_75t_L g389 ( .A1(n_309), .A2(n_256), .B1(n_210), .B2(n_209), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_357), .Y(n_390) );
A2O1A1Ixp33_ASAP7_75t_L g391 ( .A1(n_328), .A2(n_303), .B(n_302), .C(n_276), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_323), .Y(n_392) );
OAI221xp5_ASAP7_75t_L g393 ( .A1(n_345), .A2(n_280), .B1(n_241), .B2(n_250), .C(n_262), .Y(n_393) );
OAI221xp5_ASAP7_75t_L g394 ( .A1(n_345), .A2(n_317), .B1(n_280), .B2(n_355), .C(n_310), .Y(n_394) );
BUFx3_ASAP7_75t_L g395 ( .A(n_381), .Y(n_395) );
AND2x4_ASAP7_75t_SL g396 ( .A(n_372), .B(n_312), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_372), .B(n_377), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_362), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_364), .Y(n_399) );
AOI21x1_ASAP7_75t_L g400 ( .A1(n_361), .A2(n_283), .B(n_324), .Y(n_400) );
AOI22xp33_ASAP7_75t_L g401 ( .A1(n_393), .A2(n_357), .B1(n_348), .B2(n_177), .Y(n_401) );
INVx2_ASAP7_75t_L g402 ( .A(n_362), .Y(n_402) );
AOI22xp5_ASAP7_75t_L g403 ( .A1(n_367), .A2(n_274), .B1(n_339), .B2(n_311), .Y(n_403) );
NOR2x1p5_ASAP7_75t_L g404 ( .A(n_390), .B(n_312), .Y(n_404) );
HB1xp67_ASAP7_75t_L g405 ( .A(n_374), .Y(n_405) );
OAI22xp33_ASAP7_75t_L g406 ( .A1(n_389), .A2(n_312), .B1(n_307), .B2(n_311), .Y(n_406) );
OAI221xp5_ASAP7_75t_L g407 ( .A1(n_380), .A2(n_321), .B1(n_358), .B2(n_315), .C(n_214), .Y(n_407) );
OAI22xp5_ASAP7_75t_L g408 ( .A1(n_387), .A2(n_312), .B1(n_307), .B2(n_324), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_373), .B(n_332), .Y(n_409) );
AOI21xp5_ASAP7_75t_L g410 ( .A1(n_370), .A2(n_312), .B(n_325), .Y(n_410) );
AOI31xp33_ASAP7_75t_L g411 ( .A1(n_389), .A2(n_292), .A3(n_298), .B(n_236), .Y(n_411) );
INVx2_ASAP7_75t_L g412 ( .A(n_362), .Y(n_412) );
INVx4_ASAP7_75t_L g413 ( .A(n_381), .Y(n_413) );
OAI22xp5_ASAP7_75t_L g414 ( .A1(n_367), .A2(n_312), .B1(n_292), .B2(n_298), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_364), .Y(n_415) );
AOI22xp33_ASAP7_75t_L g416 ( .A1(n_394), .A2(n_274), .B1(n_321), .B2(n_275), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_369), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g418 ( .A1(n_369), .A2(n_386), .B(n_391), .Y(n_418) );
HB1xp67_ASAP7_75t_L g419 ( .A(n_368), .Y(n_419) );
AOI221xp5_ASAP7_75t_L g420 ( .A1(n_366), .A2(n_274), .B1(n_335), .B2(n_332), .C(n_279), .Y(n_420) );
AOI22xp33_ASAP7_75t_SL g421 ( .A1(n_381), .A2(n_275), .B1(n_273), .B2(n_337), .Y(n_421) );
AOI221xp5_ASAP7_75t_L g422 ( .A1(n_368), .A2(n_335), .B1(n_283), .B2(n_301), .C(n_306), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g423 ( .A1(n_379), .A2(n_275), .B1(n_254), .B2(n_340), .Y(n_423) );
AND2x2_ASAP7_75t_L g424 ( .A(n_399), .B(n_369), .Y(n_424) );
OA21x2_ASAP7_75t_L g425 ( .A1(n_418), .A2(n_388), .B(n_384), .Y(n_425) );
OAI22xp5_ASAP7_75t_L g426 ( .A1(n_403), .A2(n_388), .B1(n_384), .B2(n_392), .Y(n_426) );
AOI222xp33_ASAP7_75t_L g427 ( .A1(n_420), .A2(n_392), .B1(n_377), .B2(n_378), .C1(n_384), .C2(n_388), .Y(n_427) );
AOI221xp5_ASAP7_75t_L g428 ( .A1(n_419), .A2(n_378), .B1(n_363), .B2(n_365), .C(n_301), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_399), .B(n_375), .Y(n_429) );
AND2x2_ASAP7_75t_L g430 ( .A(n_415), .B(n_375), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_415), .Y(n_431) );
AOI33xp33_ASAP7_75t_L g432 ( .A1(n_401), .A2(n_143), .A3(n_148), .B1(n_149), .B2(n_188), .B3(n_201), .Y(n_432) );
INVxp67_ASAP7_75t_SL g433 ( .A(n_398), .Y(n_433) );
BUFx2_ASAP7_75t_L g434 ( .A(n_398), .Y(n_434) );
OAI221xp5_ASAP7_75t_L g435 ( .A1(n_416), .A2(n_371), .B1(n_254), .B2(n_281), .C(n_340), .Y(n_435) );
AND2x4_ASAP7_75t_L g436 ( .A(n_413), .B(n_385), .Y(n_436) );
OR2x2_ASAP7_75t_L g437 ( .A(n_417), .B(n_376), .Y(n_437) );
OAI211xp5_ASAP7_75t_SL g438 ( .A1(n_405), .A2(n_371), .B(n_382), .C(n_295), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_398), .Y(n_439) );
NOR2xp33_ASAP7_75t_L g440 ( .A(n_407), .B(n_385), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_397), .B(n_376), .Y(n_441) );
OAI22xp5_ASAP7_75t_L g442 ( .A1(n_403), .A2(n_381), .B1(n_383), .B2(n_385), .Y(n_442) );
BUFx2_ASAP7_75t_L g443 ( .A(n_402), .Y(n_443) );
INVx2_ASAP7_75t_L g444 ( .A(n_402), .Y(n_444) );
NAND5xp2_ASAP7_75t_L g445 ( .A(n_422), .B(n_381), .C(n_293), .D(n_316), .E(n_320), .Y(n_445) );
INVx1_ASAP7_75t_L g446 ( .A(n_417), .Y(n_446) );
OA21x2_ASAP7_75t_L g447 ( .A1(n_410), .A2(n_198), .B(n_201), .Y(n_447) );
BUFx3_ASAP7_75t_L g448 ( .A(n_395), .Y(n_448) );
OAI22xp5_ASAP7_75t_L g449 ( .A1(n_411), .A2(n_383), .B1(n_385), .B2(n_273), .Y(n_449) );
OA21x2_ASAP7_75t_L g450 ( .A1(n_400), .A2(n_187), .B(n_198), .Y(n_450) );
OA211x2_ASAP7_75t_L g451 ( .A1(n_411), .A2(n_361), .B(n_227), .C(n_383), .Y(n_451) );
AOI221xp5_ASAP7_75t_L g452 ( .A1(n_409), .A2(n_301), .B1(n_143), .B2(n_148), .C(n_293), .Y(n_452) );
INVx2_ASAP7_75t_L g453 ( .A(n_402), .Y(n_453) );
AOI221xp5_ASAP7_75t_L g454 ( .A1(n_406), .A2(n_148), .B1(n_184), .B2(n_191), .C(n_359), .Y(n_454) );
OR2x2_ASAP7_75t_L g455 ( .A(n_412), .B(n_383), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_412), .Y(n_456) );
OAI211xp5_ASAP7_75t_L g457 ( .A1(n_413), .A2(n_191), .B(n_349), .C(n_359), .Y(n_457) );
NAND2xp5_ASAP7_75t_L g458 ( .A(n_397), .B(n_326), .Y(n_458) );
OR2x6_ASAP7_75t_L g459 ( .A(n_413), .B(n_383), .Y(n_459) );
AOI221x1_ASAP7_75t_L g460 ( .A1(n_445), .A2(n_414), .B1(n_408), .B2(n_412), .C(n_413), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_SL g461 ( .A1(n_449), .A2(n_404), .B(n_395), .C(n_421), .Y(n_461) );
OAI221xp5_ASAP7_75t_SL g462 ( .A1(n_428), .A2(n_395), .B1(n_423), .B2(n_343), .C(n_336), .Y(n_462) );
INVx2_ASAP7_75t_L g463 ( .A(n_439), .Y(n_463) );
NAND4xp25_ASAP7_75t_L g464 ( .A(n_427), .B(n_18), .C(n_230), .D(n_188), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g465 ( .A(n_431), .B(n_404), .Y(n_465) );
NAND2xp5_ASAP7_75t_L g466 ( .A(n_431), .B(n_396), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_427), .B(n_396), .Y(n_467) );
BUFx2_ASAP7_75t_L g468 ( .A(n_434), .Y(n_468) );
INVx2_ASAP7_75t_L g469 ( .A(n_439), .Y(n_469) );
NAND2xp5_ASAP7_75t_SL g470 ( .A(n_448), .B(n_396), .Y(n_470) );
NOR2xp33_ASAP7_75t_R g471 ( .A(n_448), .B(n_337), .Y(n_471) );
INVx3_ASAP7_75t_L g472 ( .A(n_459), .Y(n_472) );
INVx2_ASAP7_75t_L g473 ( .A(n_439), .Y(n_473) );
OR2x2_ASAP7_75t_L g474 ( .A(n_434), .B(n_326), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_446), .Y(n_475) );
INVx1_ASAP7_75t_L g476 ( .A(n_446), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_443), .Y(n_477) );
HB1xp67_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_424), .B(n_326), .Y(n_479) );
OR2x2_ASAP7_75t_L g480 ( .A(n_437), .B(n_333), .Y(n_480) );
OAI31xp33_ASAP7_75t_L g481 ( .A1(n_426), .A2(n_359), .A3(n_333), .B(n_334), .Y(n_481) );
CKINVDCx16_ASAP7_75t_R g482 ( .A(n_448), .Y(n_482) );
INVx1_ASAP7_75t_L g483 ( .A(n_444), .Y(n_483) );
INVx2_ASAP7_75t_L g484 ( .A(n_444), .Y(n_484) );
NAND2xp5_ASAP7_75t_L g485 ( .A(n_441), .B(n_333), .Y(n_485) );
AND2x2_ASAP7_75t_L g486 ( .A(n_424), .B(n_334), .Y(n_486) );
INVxp67_ASAP7_75t_L g487 ( .A(n_437), .Y(n_487) );
INVx1_ASAP7_75t_L g488 ( .A(n_444), .Y(n_488) );
OAI22xp33_ASAP7_75t_L g489 ( .A1(n_449), .A2(n_273), .B1(n_400), .B2(n_284), .Y(n_489) );
OAI211xp5_ASAP7_75t_SL g490 ( .A1(n_435), .A2(n_230), .B(n_190), .C(n_212), .Y(n_490) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_441), .B(n_334), .Y(n_491) );
OR2x2_ASAP7_75t_L g492 ( .A(n_453), .B(n_341), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_458), .B(n_341), .Y(n_493) );
INVx1_ASAP7_75t_L g494 ( .A(n_453), .Y(n_494) );
AND2x2_ASAP7_75t_L g495 ( .A(n_453), .B(n_341), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g496 ( .A(n_429), .B(n_344), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_456), .Y(n_497) );
AOI22xp33_ASAP7_75t_L g498 ( .A1(n_440), .A2(n_227), .B1(n_273), .B2(n_351), .Y(n_498) );
INVx4_ASAP7_75t_L g499 ( .A(n_459), .Y(n_499) );
AND2x2_ASAP7_75t_L g500 ( .A(n_456), .B(n_344), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_456), .Y(n_501) );
AND2x2_ASAP7_75t_L g502 ( .A(n_433), .B(n_344), .Y(n_502) );
INVx2_ASAP7_75t_L g503 ( .A(n_425), .Y(n_503) );
AND2x2_ASAP7_75t_L g504 ( .A(n_429), .B(n_352), .Y(n_504) );
OAI21xp5_ASAP7_75t_SL g505 ( .A1(n_442), .A2(n_330), .B(n_351), .Y(n_505) );
INVx2_ASAP7_75t_L g506 ( .A(n_425), .Y(n_506) );
HB1xp67_ASAP7_75t_L g507 ( .A(n_430), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_430), .B(n_352), .Y(n_508) );
INVx1_ASAP7_75t_SL g509 ( .A(n_455), .Y(n_509) );
OAI221xp5_ASAP7_75t_L g510 ( .A1(n_438), .A2(n_218), .B1(n_359), .B2(n_356), .C(n_343), .Y(n_510) );
NAND2x1p5_ASAP7_75t_L g511 ( .A(n_499), .B(n_436), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_475), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_475), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g514 ( .A1(n_464), .A2(n_442), .B1(n_426), .B2(n_451), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_476), .Y(n_515) );
INVx2_ASAP7_75t_L g516 ( .A(n_503), .Y(n_516) );
AND2x2_ASAP7_75t_SL g517 ( .A(n_482), .B(n_436), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_476), .B(n_425), .Y(n_518) );
INVx1_ASAP7_75t_L g519 ( .A(n_465), .Y(n_519) );
AND2x2_ASAP7_75t_L g520 ( .A(n_482), .B(n_436), .Y(n_520) );
OAI31xp33_ASAP7_75t_L g521 ( .A1(n_464), .A2(n_436), .A3(n_457), .B(n_455), .Y(n_521) );
AOI22xp33_ASAP7_75t_SL g522 ( .A1(n_499), .A2(n_459), .B1(n_425), .B2(n_451), .Y(n_522) );
INVx1_ASAP7_75t_L g523 ( .A(n_507), .Y(n_523) );
NOR2xp33_ASAP7_75t_L g524 ( .A(n_487), .B(n_459), .Y(n_524) );
INVx2_ASAP7_75t_L g525 ( .A(n_503), .Y(n_525) );
INVxp67_ASAP7_75t_L g526 ( .A(n_478), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_483), .B(n_459), .Y(n_527) );
INVx1_ASAP7_75t_SL g528 ( .A(n_471), .Y(n_528) );
NAND2xp5_ASAP7_75t_L g529 ( .A(n_504), .B(n_432), .Y(n_529) );
NOR2xp67_ASAP7_75t_L g530 ( .A(n_505), .B(n_24), .Y(n_530) );
OAI221xp5_ASAP7_75t_L g531 ( .A1(n_462), .A2(n_452), .B1(n_454), .B2(n_218), .C(n_447), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_504), .B(n_447), .Y(n_532) );
NOR2x1p5_ASAP7_75t_SL g533 ( .A(n_506), .B(n_447), .Y(n_533) );
INVx2_ASAP7_75t_L g534 ( .A(n_506), .Y(n_534) );
AND2x2_ASAP7_75t_L g535 ( .A(n_479), .B(n_447), .Y(n_535) );
HB1xp67_ASAP7_75t_L g536 ( .A(n_468), .Y(n_536) );
INVx2_ASAP7_75t_L g537 ( .A(n_463), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_477), .Y(n_538) );
AND2x2_ASAP7_75t_L g539 ( .A(n_479), .B(n_450), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_483), .B(n_450), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_488), .B(n_450), .Y(n_541) );
OAI211xp5_ASAP7_75t_L g542 ( .A1(n_460), .A2(n_284), .B(n_450), .C(n_212), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_477), .Y(n_543) );
OR2x2_ASAP7_75t_L g544 ( .A(n_509), .B(n_352), .Y(n_544) );
INVxp67_ASAP7_75t_L g545 ( .A(n_468), .Y(n_545) );
CKINVDCx16_ASAP7_75t_R g546 ( .A(n_499), .Y(n_546) );
OR2x2_ASAP7_75t_L g547 ( .A(n_509), .B(n_353), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_488), .Y(n_548) );
OR2x2_ASAP7_75t_L g549 ( .A(n_494), .B(n_353), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_494), .B(n_190), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_497), .Y(n_551) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_486), .B(n_227), .Y(n_552) );
INVx1_ASAP7_75t_L g553 ( .A(n_497), .Y(n_553) );
AND2x4_ASAP7_75t_L g554 ( .A(n_472), .B(n_30), .Y(n_554) );
OR2x2_ASAP7_75t_L g555 ( .A(n_501), .B(n_353), .Y(n_555) );
NAND3xp33_ASAP7_75t_L g556 ( .A(n_460), .B(n_351), .C(n_230), .Y(n_556) );
AOI221xp5_ASAP7_75t_L g557 ( .A1(n_467), .A2(n_218), .B1(n_356), .B2(n_336), .C(n_176), .Y(n_557) );
INVx2_ASAP7_75t_L g558 ( .A(n_463), .Y(n_558) );
INVx1_ASAP7_75t_L g559 ( .A(n_501), .Y(n_559) );
AOI221xp5_ASAP7_75t_L g560 ( .A1(n_461), .A2(n_176), .B1(n_288), .B2(n_297), .C(n_219), .Y(n_560) );
OR2x2_ASAP7_75t_L g561 ( .A(n_474), .B(n_351), .Y(n_561) );
OR2x2_ASAP7_75t_L g562 ( .A(n_474), .B(n_351), .Y(n_562) );
OR2x2_ASAP7_75t_L g563 ( .A(n_466), .B(n_351), .Y(n_563) );
OAI33xp33_ASAP7_75t_L g564 ( .A1(n_485), .A2(n_31), .A3(n_35), .B1(n_36), .B2(n_38), .B3(n_43), .Y(n_564) );
AND2x2_ASAP7_75t_SL g565 ( .A(n_499), .B(n_337), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_469), .Y(n_566) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_486), .B(n_227), .Y(n_567) );
OR2x2_ASAP7_75t_L g568 ( .A(n_469), .B(n_49), .Y(n_568) );
OR2x2_ASAP7_75t_L g569 ( .A(n_473), .B(n_50), .Y(n_569) );
AND2x2_ASAP7_75t_L g570 ( .A(n_473), .B(n_54), .Y(n_570) );
NAND2x1p5_ASAP7_75t_L g571 ( .A(n_517), .B(n_470), .Y(n_571) );
NOR2xp33_ASAP7_75t_L g572 ( .A(n_528), .B(n_472), .Y(n_572) );
OR2x2_ASAP7_75t_L g573 ( .A(n_523), .B(n_484), .Y(n_573) );
INVxp67_ASAP7_75t_L g574 ( .A(n_536), .Y(n_574) );
HB1xp67_ASAP7_75t_L g575 ( .A(n_536), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_520), .B(n_472), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_512), .Y(n_577) );
INVxp67_ASAP7_75t_L g578 ( .A(n_519), .Y(n_578) );
AND2x2_ASAP7_75t_L g579 ( .A(n_517), .B(n_484), .Y(n_579) );
INVx1_ASAP7_75t_SL g580 ( .A(n_546), .Y(n_580) );
OAI21xp33_ASAP7_75t_L g581 ( .A1(n_514), .A2(n_505), .B(n_498), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_513), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_515), .Y(n_583) );
INVx1_ASAP7_75t_SL g584 ( .A(n_527), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_538), .Y(n_585) );
NOR3xp33_ASAP7_75t_L g586 ( .A(n_542), .B(n_510), .C(n_490), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_543), .Y(n_587) );
INVx1_ASAP7_75t_L g588 ( .A(n_526), .Y(n_588) );
OR2x2_ASAP7_75t_L g589 ( .A(n_526), .B(n_480), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_548), .Y(n_590) );
AND2x4_ASAP7_75t_L g591 ( .A(n_527), .B(n_502), .Y(n_591) );
OAI22xp5_ASAP7_75t_L g592 ( .A1(n_530), .A2(n_565), .B1(n_522), .B2(n_511), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_524), .B(n_502), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g594 ( .A(n_518), .B(n_481), .Y(n_594) );
INVx1_ASAP7_75t_L g595 ( .A(n_551), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_564), .A2(n_481), .B(n_489), .Y(n_596) );
INVx1_ASAP7_75t_L g597 ( .A(n_553), .Y(n_597) );
AND2x2_ASAP7_75t_L g598 ( .A(n_524), .B(n_500), .Y(n_598) );
OAI21xp5_ASAP7_75t_L g599 ( .A1(n_531), .A2(n_480), .B(n_500), .Y(n_599) );
AND2x2_ASAP7_75t_L g600 ( .A(n_545), .B(n_495), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g601 ( .A(n_518), .B(n_495), .Y(n_601) );
INVxp67_ASAP7_75t_L g602 ( .A(n_561), .Y(n_602) );
AND2x4_ASAP7_75t_L g603 ( .A(n_545), .B(n_492), .Y(n_603) );
INVx2_ASAP7_75t_L g604 ( .A(n_516), .Y(n_604) );
OR2x2_ASAP7_75t_L g605 ( .A(n_559), .B(n_491), .Y(n_605) );
INVxp67_ASAP7_75t_L g606 ( .A(n_562), .Y(n_606) );
AND2x2_ASAP7_75t_L g607 ( .A(n_511), .B(n_508), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_532), .B(n_496), .Y(n_608) );
OR2x2_ASAP7_75t_L g609 ( .A(n_537), .B(n_492), .Y(n_609) );
OAI21xp5_ASAP7_75t_L g610 ( .A1(n_556), .A2(n_493), .B(n_284), .Y(n_610) );
NAND4xp25_ASAP7_75t_SL g611 ( .A(n_521), .B(n_56), .C(n_61), .D(n_63), .Y(n_611) );
INVxp67_ASAP7_75t_L g612 ( .A(n_544), .Y(n_612) );
INVx2_ASAP7_75t_L g613 ( .A(n_516), .Y(n_613) );
OAI22xp33_ASAP7_75t_SL g614 ( .A1(n_554), .A2(n_360), .B1(n_284), .B2(n_327), .Y(n_614) );
INVx2_ASAP7_75t_L g615 ( .A(n_525), .Y(n_615) );
OR2x2_ASAP7_75t_L g616 ( .A(n_537), .B(n_64), .Y(n_616) );
NOR2x1_ASAP7_75t_L g617 ( .A(n_554), .B(n_330), .Y(n_617) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_525), .B(n_65), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_535), .B(n_539), .Y(n_619) );
OR2x2_ASAP7_75t_L g620 ( .A(n_558), .B(n_66), .Y(n_620) );
INVxp67_ASAP7_75t_L g621 ( .A(n_547), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_558), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g623 ( .A(n_534), .B(n_67), .Y(n_623) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_565), .B(n_360), .Y(n_624) );
NAND4xp25_ASAP7_75t_SL g625 ( .A(n_580), .B(n_522), .C(n_560), .D(n_557), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_580), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_578), .B(n_534), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g628 ( .A(n_612), .B(n_540), .Y(n_628) );
AND2x2_ASAP7_75t_L g629 ( .A(n_619), .B(n_566), .Y(n_629) );
NAND2xp5_ASAP7_75t_SL g630 ( .A(n_592), .B(n_554), .Y(n_630) );
AOI221xp5_ASAP7_75t_L g631 ( .A1(n_588), .A2(n_564), .B1(n_529), .B2(n_540), .C(n_541), .Y(n_631) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_621), .B(n_541), .Y(n_632) );
A2O1A1Ixp33_ASAP7_75t_L g633 ( .A1(n_592), .A2(n_533), .B(n_570), .C(n_568), .Y(n_633) );
INVx1_ASAP7_75t_L g634 ( .A(n_585), .Y(n_634) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_611), .A2(n_570), .B(n_569), .Y(n_635) );
XNOR2xp5_ASAP7_75t_L g636 ( .A(n_576), .B(n_563), .Y(n_636) );
OAI22xp33_ASAP7_75t_L g637 ( .A1(n_571), .A2(n_549), .B1(n_555), .B2(n_566), .Y(n_637) );
INVx1_ASAP7_75t_L g638 ( .A(n_587), .Y(n_638) );
OAI22xp5_ASAP7_75t_L g639 ( .A1(n_571), .A2(n_567), .B1(n_552), .B2(n_550), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_574), .B(n_550), .Y(n_640) );
NAND2xp5_ASAP7_75t_L g641 ( .A(n_575), .B(n_70), .Y(n_641) );
NOR2xp33_ASAP7_75t_L g642 ( .A(n_581), .B(n_73), .Y(n_642) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_617), .B(n_327), .Y(n_643) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_602), .B(n_74), .Y(n_644) );
AND2x2_ASAP7_75t_L g645 ( .A(n_584), .B(n_591), .Y(n_645) );
OR2x2_ASAP7_75t_L g646 ( .A(n_601), .B(n_75), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_577), .Y(n_647) );
OAI211xp5_ASAP7_75t_SL g648 ( .A1(n_599), .A2(n_297), .B(n_330), .C(n_228), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_582), .Y(n_649) );
NAND2xp5_ASAP7_75t_SL g650 ( .A(n_614), .B(n_360), .Y(n_650) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_624), .B(n_603), .Y(n_651) );
OA21x2_ASAP7_75t_L g652 ( .A1(n_594), .A2(n_266), .B(n_287), .Y(n_652) );
INVx2_ASAP7_75t_L g653 ( .A(n_604), .Y(n_653) );
NAND3xp33_ASAP7_75t_L g654 ( .A(n_599), .B(n_360), .C(n_330), .Y(n_654) );
INVxp67_ASAP7_75t_L g655 ( .A(n_572), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_613), .Y(n_656) );
INVx2_ASAP7_75t_L g657 ( .A(n_615), .Y(n_657) );
NOR2xp67_ASAP7_75t_SL g658 ( .A(n_616), .B(n_360), .Y(n_658) );
NAND2xp5_ASAP7_75t_SL g659 ( .A(n_624), .B(n_360), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_603), .Y(n_660) );
NAND2x1_ASAP7_75t_L g661 ( .A(n_579), .B(n_327), .Y(n_661) );
AOI21x1_ASAP7_75t_SL g662 ( .A1(n_594), .A2(n_76), .B(n_78), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g663 ( .A1(n_583), .A2(n_297), .B1(n_219), .B2(n_226), .C(n_228), .Y(n_663) );
AO22x2_ASAP7_75t_L g664 ( .A1(n_584), .A2(n_79), .B1(n_300), .B2(n_266), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g665 ( .A(n_606), .B(n_226), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_607), .A2(n_327), .B1(n_300), .B2(n_272), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_590), .B(n_267), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_573), .Y(n_668) );
XNOR2xp5_ASAP7_75t_L g669 ( .A(n_598), .B(n_267), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_595), .Y(n_670) );
INVx1_ASAP7_75t_SL g671 ( .A(n_589), .Y(n_671) );
NOR2xp33_ASAP7_75t_L g672 ( .A(n_605), .B(n_257), .Y(n_672) );
XNOR2xp5_ASAP7_75t_L g673 ( .A(n_593), .B(n_257), .Y(n_673) );
AOI222xp33_ASAP7_75t_L g674 ( .A1(n_600), .A2(n_290), .B1(n_272), .B2(n_291), .C1(n_244), .C2(n_247), .Y(n_674) );
OAI21xp5_ASAP7_75t_L g675 ( .A1(n_596), .A2(n_290), .B(n_287), .Y(n_675) );
OAI31xp33_ASAP7_75t_L g676 ( .A1(n_586), .A2(n_247), .A3(n_285), .B(n_244), .Y(n_676) );
NAND4xp75_ASAP7_75t_L g677 ( .A(n_608), .B(n_285), .C(n_291), .D(n_272), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_597), .Y(n_678) );
OAI22xp33_ASAP7_75t_SL g679 ( .A1(n_601), .A2(n_272), .B1(n_223), .B2(n_225), .Y(n_679) );
XNOR2x1_ASAP7_75t_L g680 ( .A(n_591), .B(n_215), .Y(n_680) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_622), .B(n_215), .Y(n_681) );
XOR2xp5_ASAP7_75t_L g682 ( .A(n_609), .B(n_215), .Y(n_682) );
AO22x2_ASAP7_75t_L g683 ( .A1(n_610), .A2(n_223), .B1(n_225), .B2(n_215), .Y(n_683) );
XNOR2xp5_ASAP7_75t_L g684 ( .A(n_618), .B(n_215), .Y(n_684) );
NAND2xp5_ASAP7_75t_L g685 ( .A(n_618), .B(n_623), .Y(n_685) );
INVx1_ASAP7_75t_L g686 ( .A(n_623), .Y(n_686) );
OAI221xp5_ASAP7_75t_SL g687 ( .A1(n_626), .A2(n_633), .B1(n_655), .B2(n_637), .C(n_631), .Y(n_687) );
OAI22xp5_ASAP7_75t_L g688 ( .A1(n_630), .A2(n_633), .B1(n_680), .B2(n_651), .Y(n_688) );
OAI21xp5_ASAP7_75t_SL g689 ( .A1(n_630), .A2(n_651), .B(n_648), .Y(n_689) );
NAND5xp2_ASAP7_75t_L g690 ( .A(n_642), .B(n_675), .C(n_635), .D(n_674), .E(n_676), .Y(n_690) );
AOI22xp33_ASAP7_75t_L g691 ( .A1(n_625), .A2(n_682), .B1(n_642), .B2(n_654), .Y(n_691) );
AOI22xp33_ASAP7_75t_SL g692 ( .A1(n_664), .A2(n_671), .B1(n_645), .B2(n_639), .Y(n_692) );
INVx1_ASAP7_75t_L g693 ( .A(n_627), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_638), .Y(n_694) );
INVx1_ASAP7_75t_L g695 ( .A(n_634), .Y(n_695) );
INVx1_ASAP7_75t_SL g696 ( .A(n_629), .Y(n_696) );
INVx1_ASAP7_75t_L g697 ( .A(n_649), .Y(n_697) );
AOI21xp5_ASAP7_75t_SL g698 ( .A1(n_650), .A2(n_659), .B(n_679), .Y(n_698) );
AO22x2_ASAP7_75t_L g699 ( .A1(n_678), .A2(n_670), .B1(n_647), .B2(n_660), .Y(n_699) );
AOI221xp5_ASAP7_75t_L g700 ( .A1(n_668), .A2(n_637), .B1(n_628), .B2(n_632), .C(n_686), .Y(n_700) );
OAI221xp5_ASAP7_75t_L g701 ( .A1(n_692), .A2(n_661), .B1(n_636), .B2(n_650), .C(n_640), .Y(n_701) );
OAI211xp5_ASAP7_75t_SL g702 ( .A1(n_689), .A2(n_646), .B(n_665), .C(n_644), .Y(n_702) );
OAI21xp5_ASAP7_75t_L g703 ( .A1(n_688), .A2(n_659), .B(n_677), .Y(n_703) );
INVx1_ASAP7_75t_SL g704 ( .A(n_696), .Y(n_704) );
INVx1_ASAP7_75t_L g705 ( .A(n_694), .Y(n_705) );
OAI21xp5_ASAP7_75t_SL g706 ( .A1(n_691), .A2(n_684), .B(n_673), .Y(n_706) );
AOI22xp5_ASAP7_75t_L g707 ( .A1(n_700), .A2(n_672), .B1(n_669), .B2(n_664), .Y(n_707) );
AOI211xp5_ASAP7_75t_L g708 ( .A1(n_687), .A2(n_685), .B(n_641), .C(n_658), .Y(n_708) );
NOR2x1_ASAP7_75t_L g709 ( .A(n_703), .B(n_698), .Y(n_709) );
AOI221xp5_ASAP7_75t_L g710 ( .A1(n_701), .A2(n_699), .B1(n_690), .B2(n_693), .C(n_695), .Y(n_710) );
NAND3xp33_ASAP7_75t_SL g711 ( .A(n_708), .B(n_643), .C(n_666), .Y(n_711) );
AOI222xp33_ASAP7_75t_L g712 ( .A1(n_704), .A2(n_699), .B1(n_697), .B2(n_653), .C1(n_656), .C2(n_657), .Y(n_712) );
OA22x2_ASAP7_75t_L g713 ( .A1(n_707), .A2(n_706), .B1(n_705), .B2(n_699), .Y(n_713) );
NOR2xp33_ASAP7_75t_L g714 ( .A(n_709), .B(n_702), .Y(n_714) );
BUFx2_ASAP7_75t_L g715 ( .A(n_713), .Y(n_715) );
NOR4xp25_ASAP7_75t_L g716 ( .A(n_710), .B(n_681), .C(n_667), .D(n_663), .Y(n_716) );
AOI22xp5_ASAP7_75t_L g717 ( .A1(n_715), .A2(n_711), .B1(n_712), .B2(n_683), .Y(n_717) );
OAI222xp33_ASAP7_75t_L g718 ( .A1(n_714), .A2(n_666), .B1(n_653), .B2(n_620), .C1(n_662), .C2(n_683), .Y(n_718) );
INVx1_ASAP7_75t_L g719 ( .A(n_717), .Y(n_719) );
INVx1_ASAP7_75t_L g720 ( .A(n_718), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_719), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g722 ( .A1(n_721), .A2(n_720), .B(n_716), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g723 ( .A1(n_722), .A2(n_610), .B1(n_652), .B2(n_716), .C(n_715), .Y(n_723) );
endmodule