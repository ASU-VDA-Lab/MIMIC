module real_jpeg_6496_n_20 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_19, n_16, n_15, n_13, n_20);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_19;
input n_16;
input n_15;
input n_13;

output n_20;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_446;
wire n_199;
wire n_95;
wire n_441;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_456;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_466;
wire n_353;
wire n_453;
wire n_230;
wire n_417;
wire n_428;
wire n_216;
wire n_128;
wire n_202;
wire n_483;
wire n_367;
wire n_127;
wire n_365;
wire n_356;
wire n_464;
wire n_423;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_422;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_393;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_131;
wire n_439;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_469;
wire n_378;
wire n_200;
wire n_432;
wire n_465;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_459;
wire n_139;
wire n_33;
wire n_338;
wire n_175;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_470;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_21;
wire n_476;
wire n_69;
wire n_31;
wire n_426;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_411;
wire n_382;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_448;
wire n_212;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_25;
wire n_480;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_412;
wire n_405;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_427;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_152;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_201;
wire n_484;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_472;
wire n_343;
wire n_292;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_444;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_143;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_368;
wire n_100;
wire n_51;
wire n_205;
wire n_361;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_438;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_257;
wire n_447;
wire n_344;
wire n_210;
wire n_206;
wire n_408;
wire n_85;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

NAND2xp5_ASAP7_75t_L g37 ( 
.A(n_0),
.B(n_38),
.Y(n_37)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_0),
.B(n_42),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_0),
.B(n_98),
.Y(n_97)
);

AND2x2_ASAP7_75t_SL g114 ( 
.A(n_0),
.B(n_115),
.Y(n_114)
);

AND2x2_ASAP7_75t_SL g143 ( 
.A(n_0),
.B(n_64),
.Y(n_143)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_1),
.Y(n_99)
);

INVx8_ASAP7_75t_L g221 ( 
.A(n_1),
.Y(n_221)
);

BUFx6f_ASAP7_75t_L g303 ( 
.A(n_1),
.Y(n_303)
);

BUFx6f_ASAP7_75t_L g310 ( 
.A(n_1),
.Y(n_310)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_2),
.Y(n_78)
);

BUFx6f_ASAP7_75t_L g104 ( 
.A(n_2),
.Y(n_104)
);

BUFx5_ASAP7_75t_L g139 ( 
.A(n_2),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_2),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g276 ( 
.A(n_2),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_3),
.B(n_213),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_3),
.B(n_255),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g298 ( 
.A(n_3),
.B(n_299),
.Y(n_298)
);

AND2x2_ASAP7_75t_L g323 ( 
.A(n_3),
.B(n_324),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_3),
.B(n_338),
.Y(n_337)
);

AND2x2_ASAP7_75t_L g375 ( 
.A(n_3),
.B(n_64),
.Y(n_375)
);

AND2x2_ASAP7_75t_L g384 ( 
.A(n_3),
.B(n_249),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_4),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_4),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_4),
.B(n_107),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_4),
.B(n_179),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_4),
.B(n_200),
.Y(n_199)
);

AND2x2_ASAP7_75t_SL g277 ( 
.A(n_4),
.B(n_278),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_4),
.B(n_303),
.Y(n_356)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_4),
.B(n_404),
.Y(n_403)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_5),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_5),
.B(n_102),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_5),
.B(n_204),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_5),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_5),
.B(n_115),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g334 ( 
.A(n_5),
.B(n_219),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g358 ( 
.A(n_5),
.B(n_359),
.Y(n_358)
);

AND2x2_ASAP7_75t_L g398 ( 
.A(n_5),
.B(n_53),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_SL g160 ( 
.A(n_6),
.B(n_104),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_6),
.B(n_198),
.Y(n_197)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_6),
.B(n_249),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_6),
.B(n_303),
.Y(n_302)
);

AND2x2_ASAP7_75t_L g317 ( 
.A(n_6),
.B(n_216),
.Y(n_317)
);

AND2x2_ASAP7_75t_L g342 ( 
.A(n_6),
.B(n_343),
.Y(n_342)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_6),
.B(n_368),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g395 ( 
.A(n_6),
.B(n_396),
.Y(n_395)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_7),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g95 ( 
.A(n_7),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_7),
.Y(n_127)
);

INVx3_ASAP7_75t_L g389 ( 
.A(n_7),
.Y(n_389)
);

INVx3_ASAP7_75t_L g484 ( 
.A(n_8),
.Y(n_484)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_9),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g182 ( 
.A(n_9),
.B(n_183),
.Y(n_182)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_9),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_9),
.B(n_285),
.Y(n_284)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_9),
.B(n_319),
.Y(n_318)
);

AND2x2_ASAP7_75t_L g333 ( 
.A(n_9),
.B(n_216),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g399 ( 
.A(n_9),
.B(n_115),
.Y(n_399)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_10),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g279 ( 
.A(n_10),
.Y(n_279)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_10),
.Y(n_283)
);

INVx8_ASAP7_75t_L g58 ( 
.A(n_11),
.Y(n_58)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g217 ( 
.A(n_12),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g261 ( 
.A(n_12),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_13),
.B(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_13),
.B(n_49),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g116 ( 
.A(n_13),
.B(n_117),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_13),
.B(n_137),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g176 ( 
.A(n_13),
.B(n_177),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_13),
.B(n_259),
.Y(n_258)
);

AND2x2_ASAP7_75t_L g282 ( 
.A(n_13),
.B(n_283),
.Y(n_282)
);

AND2x2_ASAP7_75t_L g406 ( 
.A(n_13),
.B(n_407),
.Y(n_406)
);

INVx6_ASAP7_75t_L g51 ( 
.A(n_14),
.Y(n_51)
);

INVxp33_ASAP7_75t_L g486 ( 
.A(n_15),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_16),
.B(n_56),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_16),
.B(n_62),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_16),
.B(n_86),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_16),
.B(n_125),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_16),
.B(n_216),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_16),
.B(n_223),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_16),
.B(n_247),
.Y(n_246)
);

INVx8_ASAP7_75t_L g34 ( 
.A(n_17),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_18),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_18),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_18),
.B(n_82),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_18),
.B(n_129),
.Y(n_128)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_18),
.B(n_162),
.Y(n_161)
);

AND2x2_ASAP7_75t_SL g218 ( 
.A(n_18),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_19),
.B(n_274),
.Y(n_273)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_19),
.B(n_305),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_19),
.B(n_310),
.Y(n_309)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_19),
.B(n_115),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g341 ( 
.A(n_19),
.B(n_179),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_19),
.B(n_373),
.Y(n_372)
);

AND2x2_ASAP7_75t_L g385 ( 
.A(n_19),
.B(n_386),
.Y(n_385)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_482),
.B(n_485),
.Y(n_20)
);

XNOR2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_186),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_185),
.Y(n_22)
);

INVxp67_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_149),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_25),
.B(n_149),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_27),
.B1(n_109),
.B2(n_148),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

MAJIxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_73),
.C(n_89),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_28),
.B(n_151),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g28 ( 
.A(n_29),
.B(n_47),
.C(n_59),
.Y(n_28)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_29),
.B(n_229),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_35),
.Y(n_29)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_30),
.B(n_37),
.C(n_41),
.Y(n_118)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_32),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

BUFx5_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx6_ASAP7_75t_L g87 ( 
.A(n_34),
.Y(n_87)
);

INVx3_ASAP7_75t_L g227 ( 
.A(n_34),
.Y(n_227)
);

BUFx6f_ASAP7_75t_L g374 ( 
.A(n_34),
.Y(n_374)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_36),
.A2(n_37),
.B1(n_41),
.B2(n_46),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g112 ( 
.A1(n_36),
.A2(n_37),
.B1(n_113),
.B2(n_114),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_36),
.B(n_113),
.C(n_116),
.Y(n_134)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g223 ( 
.A(n_39),
.Y(n_223)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g307 ( 
.A(n_40),
.Y(n_307)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_41),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_41),
.B(n_92),
.C(n_96),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_41),
.A2(n_46),
.B1(n_96),
.B2(n_97),
.Y(n_158)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

INVx2_ASAP7_75t_L g301 ( 
.A(n_44),
.Y(n_301)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_45),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_47),
.B(n_59),
.Y(n_229)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_55),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_48),
.B(n_55),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_50),
.Y(n_204)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

BUFx3_ASAP7_75t_L g180 ( 
.A(n_51),
.Y(n_180)
);

INVx3_ASAP7_75t_L g266 ( 
.A(n_51),
.Y(n_266)
);

XNOR2xp5_ASAP7_75t_L g165 ( 
.A(n_52),
.B(n_166),
.Y(n_165)
);

INVx4_ASAP7_75t_L g354 ( 
.A(n_53),
.Y(n_354)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

INVx11_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx3_ASAP7_75t_L g370 ( 
.A(n_58),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_L g59 ( 
.A(n_60),
.B(n_70),
.Y(n_59)
);

XNOR2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_65),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g119 ( 
.A(n_61),
.B(n_65),
.C(n_70),
.Y(n_119)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_67),
.Y(n_177)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_68),
.Y(n_67)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_69),
.Y(n_68)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_69),
.Y(n_115)
);

INVx3_ASAP7_75t_L g202 ( 
.A(n_69),
.Y(n_202)
);

INVx5_ASAP7_75t_L g339 ( 
.A(n_69),
.Y(n_339)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_72),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_73),
.A2(n_89),
.B1(n_90),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_73),
.Y(n_152)
);

XOR2xp5_ASAP7_75t_L g73 ( 
.A(n_74),
.B(n_79),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_74),
.B(n_80),
.C(n_88),
.Y(n_132)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_78),
.Y(n_77)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_78),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_80),
.A2(n_81),
.B1(n_85),
.B2(n_88),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

INVx3_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_85),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_87),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g251 ( 
.A(n_87),
.Y(n_251)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_100),
.C(n_105),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_91),
.B(n_168),
.Y(n_167)
);

XNOR2xp5_ASAP7_75t_SL g157 ( 
.A(n_92),
.B(n_158),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_94),
.Y(n_92)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_94),
.Y(n_198)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g206 ( 
.A1(n_96),
.A2(n_97),
.B1(n_161),
.B2(n_207),
.Y(n_206)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_97),
.B(n_160),
.C(n_161),
.Y(n_159)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_100),
.A2(n_101),
.B1(n_105),
.B2(n_106),
.Y(n_168)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx8_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

INVx8_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_105),
.A2(n_106),
.B1(n_181),
.B2(n_182),
.Y(n_209)
);

INVx1_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_106),
.B(n_170),
.C(n_181),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_109),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_120),
.Y(n_109)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_118),
.C(n_119),
.Y(n_110)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_111),
.B(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_SL g111 ( 
.A(n_112),
.B(n_116),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_L g141 ( 
.A1(n_113),
.A2(n_114),
.B1(n_142),
.B2(n_143),
.Y(n_141)
);

CKINVDCx16_ASAP7_75t_R g113 ( 
.A(n_114),
.Y(n_113)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_118),
.B(n_119),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_121),
.A2(n_122),
.B1(n_133),
.B2(n_147),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_122),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_132),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_128),
.Y(n_123)
);

INVx6_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_127),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_127),
.Y(n_175)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_127),
.Y(n_256)
);

INVx4_ASAP7_75t_SL g129 ( 
.A(n_130),
.Y(n_129)
);

INVx5_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_133),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g133 ( 
.A1(n_134),
.A2(n_135),
.B1(n_145),
.B2(n_146),
.Y(n_133)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_134),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_135),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_136),
.A2(n_140),
.B1(n_141),
.B2(n_144),
.Y(n_135)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_136),
.Y(n_144)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVx8_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_141),
.Y(n_140)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_143),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_153),
.C(n_155),
.Y(n_149)
);

FAx1_ASAP7_75t_L g478 ( 
.A(n_150),
.B(n_153),
.CI(n_155),
.CON(n_478),
.SN(n_478)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_167),
.C(n_169),
.Y(n_155)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_156),
.B(n_231),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_157),
.B(n_159),
.C(n_165),
.Y(n_156)
);

XOR2xp5_ASAP7_75t_L g237 ( 
.A(n_157),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_159),
.B(n_165),
.Y(n_238)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_160),
.B(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_161),
.Y(n_207)
);

INVx4_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

BUFx6f_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_167),
.B(n_169),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_171),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g208 ( 
.A(n_171),
.B(n_209),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_176),
.C(n_178),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_L g194 ( 
.A(n_172),
.B(n_178),
.Y(n_194)
);

INVx3_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx8_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

XNOR2xp5_ASAP7_75t_SL g193 ( 
.A(n_176),
.B(n_194),
.Y(n_193)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

BUFx6f_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

AO21x1_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_476),
.B(n_480),
.Y(n_186)
);

HB1xp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_287),
.B(n_475),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_SL g189 ( 
.A(n_190),
.B(n_232),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_190),
.B(n_232),
.Y(n_475)
);

BUFx24_ASAP7_75t_SL g489 ( 
.A(n_190),
.Y(n_489)
);

FAx1_ASAP7_75t_L g190 ( 
.A(n_191),
.B(n_228),
.CI(n_230),
.CON(n_190),
.SN(n_190)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_191),
.B(n_228),
.C(n_230),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g191 ( 
.A(n_192),
.B(n_208),
.C(n_210),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_192),
.B(n_235),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_195),
.C(n_205),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g460 ( 
.A(n_193),
.B(n_461),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_L g461 ( 
.A1(n_195),
.A2(n_196),
.B1(n_205),
.B2(n_462),
.Y(n_461)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.C(n_203),
.Y(n_196)
);

XNOR2xp5_ASAP7_75t_L g451 ( 
.A(n_197),
.B(n_203),
.Y(n_451)
);

XOR2xp5_ASAP7_75t_L g450 ( 
.A(n_199),
.B(n_451),
.Y(n_450)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_205),
.Y(n_462)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_208),
.B(n_210),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g210 ( 
.A(n_211),
.B(n_222),
.C(n_224),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_211),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_212),
.B(n_214),
.C(n_218),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g243 ( 
.A(n_212),
.B(n_244),
.Y(n_243)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_215),
.B(n_218),
.Y(n_244)
);

BUFx5_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx2_ASAP7_75t_L g405 ( 
.A(n_217),
.Y(n_405)
);

INVx8_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_221),
.Y(n_319)
);

INVx4_ASAP7_75t_L g407 ( 
.A(n_221),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g269 ( 
.A(n_222),
.B(n_224),
.Y(n_269)
);

INVx6_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx4_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

MAJIxp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_236),
.C(n_239),
.Y(n_232)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

XNOR2xp5_ASAP7_75t_L g471 ( 
.A(n_234),
.B(n_237),
.Y(n_471)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_237),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g470 ( 
.A(n_239),
.B(n_471),
.Y(n_470)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_267),
.C(n_270),
.Y(n_239)
);

INVxp67_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_241),
.B(n_464),
.Y(n_463)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_245),
.C(n_252),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_242),
.A2(n_243),
.B1(n_442),
.B2(n_443),
.Y(n_441)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_243),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g429 ( 
.A1(n_245),
.A2(n_246),
.B(n_248),
.Y(n_429)
);

XNOR2xp5_ASAP7_75t_L g442 ( 
.A(n_245),
.B(n_252),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

INVx5_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

INVx3_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx4_ASAP7_75t_L g286 ( 
.A(n_251),
.Y(n_286)
);

MAJx2_ASAP7_75t_L g252 ( 
.A(n_253),
.B(n_257),
.C(n_262),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_L g419 ( 
.A1(n_253),
.A2(n_254),
.B1(n_257),
.B2(n_258),
.Y(n_419)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_258),
.Y(n_257)
);

INVx6_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_261),
.Y(n_260)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_261),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g418 ( 
.A(n_262),
.B(n_419),
.Y(n_418)
);

NOR2xp33_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_L g353 ( 
.A(n_263),
.B(n_354),
.Y(n_353)
);

INVx5_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_266),
.Y(n_265)
);

INVx3_ASAP7_75t_L g397 ( 
.A(n_266),
.Y(n_397)
);

AOI22xp33_ASAP7_75t_L g464 ( 
.A1(n_267),
.A2(n_268),
.B1(n_270),
.B2(n_465),
.Y(n_464)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_268),
.Y(n_267)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_270),
.Y(n_465)
);

MAJx2_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_282),
.C(n_284),
.Y(n_270)
);

INVx1_ASAP7_75t_SL g271 ( 
.A(n_272),
.Y(n_271)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_272),
.B(n_453),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_273),
.B(n_277),
.C(n_280),
.Y(n_272)
);

XOR2xp5_ASAP7_75t_L g430 ( 
.A(n_273),
.B(n_431),
.Y(n_430)
);

INVx4_ASAP7_75t_L g274 ( 
.A(n_275),
.Y(n_274)
);

INVx8_ASAP7_75t_L g275 ( 
.A(n_276),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g431 ( 
.A1(n_277),
.A2(n_280),
.B1(n_281),
.B2(n_432),
.Y(n_431)
);

INVx1_ASAP7_75t_SL g432 ( 
.A(n_277),
.Y(n_432)
);

BUFx6f_ASAP7_75t_L g278 ( 
.A(n_279),
.Y(n_278)
);

INVx3_ASAP7_75t_L g325 ( 
.A(n_279),
.Y(n_325)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g453 ( 
.A(n_282),
.B(n_284),
.Y(n_453)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_286),
.Y(n_285)
);

AOI21xp5_ASAP7_75t_SL g287 ( 
.A1(n_288),
.A2(n_469),
.B(n_474),
.Y(n_287)
);

OAI21x1_ASAP7_75t_L g288 ( 
.A1(n_289),
.A2(n_456),
.B(n_468),
.Y(n_288)
);

AOI21x1_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_438),
.B(n_455),
.Y(n_289)
);

OAI21x1_ASAP7_75t_L g290 ( 
.A1(n_291),
.A2(n_412),
.B(n_437),
.Y(n_290)
);

AOI21x1_ASAP7_75t_L g291 ( 
.A1(n_292),
.A2(n_379),
.B(n_411),
.Y(n_291)
);

OAI21xp5_ASAP7_75t_L g292 ( 
.A1(n_293),
.A2(n_346),
.B(n_378),
.Y(n_292)
);

AOI21xp5_ASAP7_75t_L g293 ( 
.A1(n_294),
.A2(n_329),
.B(n_345),
.Y(n_293)
);

OAI21xp5_ASAP7_75t_L g294 ( 
.A1(n_295),
.A2(n_312),
.B(n_328),
.Y(n_294)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_296),
.A2(n_308),
.B(n_311),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_304),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_297),
.B(n_304),
.Y(n_311)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_298),
.B(n_302),
.Y(n_297)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_298),
.B(n_309),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_298),
.B(n_302),
.Y(n_313)
);

INVx4_ASAP7_75t_SL g299 ( 
.A(n_300),
.Y(n_299)
);

INVx4_ASAP7_75t_L g300 ( 
.A(n_301),
.Y(n_300)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_306),
.Y(n_305)
);

HB1xp67_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_313),
.B(n_314),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_314),
.Y(n_328)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_315),
.A2(n_316),
.B1(n_320),
.B2(n_321),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_315),
.B(n_323),
.C(n_326),
.Y(n_344)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_316),
.Y(n_315)
);

XNOR2xp5_ASAP7_75t_SL g316 ( 
.A(n_317),
.B(n_318),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_317),
.B(n_318),
.Y(n_335)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

OAI22xp5_ASAP7_75t_SL g321 ( 
.A1(n_322),
.A2(n_323),
.B1(n_326),
.B2(n_327),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_325),
.Y(n_324)
);

INVx2_ASAP7_75t_L g343 ( 
.A(n_325),
.Y(n_343)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_SL g329 ( 
.A(n_330),
.B(n_344),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_330),
.B(n_344),
.Y(n_345)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_336),
.Y(n_330)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_335),
.Y(n_331)
);

MAJIxp5_ASAP7_75t_L g347 ( 
.A(n_332),
.B(n_335),
.C(n_348),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_333),
.B(n_334),
.Y(n_332)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_333),
.B(n_334),
.Y(n_351)
);

INVxp67_ASAP7_75t_L g348 ( 
.A(n_336),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_340),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_364),
.C(n_365),
.Y(n_363)
);

HB1xp67_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

XNOR2xp5_ASAP7_75t_L g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g364 ( 
.A(n_341),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_342),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_347),
.B(n_349),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_347),
.B(n_349),
.Y(n_378)
);

XNOR2xp5_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_362),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g410 ( 
.A(n_350),
.B(n_363),
.C(n_366),
.Y(n_410)
);

XOR2xp5_ASAP7_75t_L g350 ( 
.A(n_351),
.B(n_352),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_351),
.B(n_353),
.C(n_355),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g352 ( 
.A(n_353),
.B(n_355),
.Y(n_352)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_356),
.A2(n_357),
.B1(n_358),
.B2(n_361),
.Y(n_355)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_356),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g390 ( 
.A(n_357),
.B(n_361),
.Y(n_390)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_358),
.Y(n_357)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_360),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_366),
.Y(n_362)
);

XNOR2xp5_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_371),
.Y(n_366)
);

MAJx2_ASAP7_75t_L g409 ( 
.A(n_367),
.B(n_375),
.C(n_376),
.Y(n_409)
);

INVx5_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

INVx3_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

AOI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_372),
.A2(n_375),
.B1(n_376),
.B2(n_377),
.Y(n_371)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_372),
.Y(n_376)
);

INVx4_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_375),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_SL g379 ( 
.A(n_380),
.B(n_410),
.Y(n_379)
);

NOR2xp33_ASAP7_75t_L g411 ( 
.A(n_380),
.B(n_410),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g380 ( 
.A(n_381),
.B(n_392),
.Y(n_380)
);

XOR2xp5_ASAP7_75t_L g381 ( 
.A(n_382),
.B(n_391),
.Y(n_381)
);

MAJIxp5_ASAP7_75t_L g435 ( 
.A(n_382),
.B(n_391),
.C(n_436),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_390),
.Y(n_382)
);

XNOR2xp5_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_385),
.Y(n_383)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_384),
.Y(n_426)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_385),
.Y(n_427)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_387),
.Y(n_386)
);

INVx6_ASAP7_75t_L g387 ( 
.A(n_388),
.Y(n_387)
);

INVx5_ASAP7_75t_L g388 ( 
.A(n_389),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g425 ( 
.A(n_390),
.B(n_426),
.C(n_427),
.Y(n_425)
);

INVxp67_ASAP7_75t_L g436 ( 
.A(n_392),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_393),
.B(n_400),
.Y(n_392)
);

MAJIxp5_ASAP7_75t_L g415 ( 
.A(n_393),
.B(n_402),
.C(n_408),
.Y(n_415)
);

XOR2xp5_ASAP7_75t_L g393 ( 
.A(n_394),
.B(n_399),
.Y(n_393)
);

XNOR2xp5_ASAP7_75t_L g394 ( 
.A(n_395),
.B(n_398),
.Y(n_394)
);

MAJx2_ASAP7_75t_L g423 ( 
.A(n_395),
.B(n_398),
.C(n_399),
.Y(n_423)
);

INVx6_ASAP7_75t_L g396 ( 
.A(n_397),
.Y(n_396)
);

AOI22xp5_ASAP7_75t_L g400 ( 
.A1(n_401),
.A2(n_402),
.B1(n_408),
.B2(n_409),
.Y(n_400)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_403),
.B(n_406),
.Y(n_402)
);

AND2x2_ASAP7_75t_L g422 ( 
.A(n_403),
.B(n_406),
.Y(n_422)
);

INVx2_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

INVx1_ASAP7_75t_SL g408 ( 
.A(n_409),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_413),
.B(n_435),
.Y(n_412)
);

NAND2xp5_ASAP7_75t_L g437 ( 
.A(n_413),
.B(n_435),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g413 ( 
.A(n_414),
.B(n_424),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g414 ( 
.A(n_415),
.B(n_416),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g454 ( 
.A(n_415),
.B(n_416),
.C(n_424),
.Y(n_454)
);

OAI22xp5_ASAP7_75t_SL g416 ( 
.A1(n_417),
.A2(n_418),
.B1(n_420),
.B2(n_421),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g446 ( 
.A(n_417),
.B(n_447),
.C(n_448),
.Y(n_446)
);

INVx1_ASAP7_75t_SL g417 ( 
.A(n_418),
.Y(n_417)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_421),
.Y(n_420)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_422),
.B(n_423),
.Y(n_421)
);

CKINVDCx16_ASAP7_75t_R g447 ( 
.A(n_422),
.Y(n_447)
);

INVx1_ASAP7_75t_L g448 ( 
.A(n_423),
.Y(n_448)
);

XNOR2xp5_ASAP7_75t_SL g424 ( 
.A(n_425),
.B(n_428),
.Y(n_424)
);

MAJIxp5_ASAP7_75t_L g444 ( 
.A(n_425),
.B(n_429),
.C(n_434),
.Y(n_444)
);

AOI22xp5_ASAP7_75t_L g428 ( 
.A1(n_429),
.A2(n_430),
.B1(n_433),
.B2(n_434),
.Y(n_428)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_430),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_439),
.B(n_454),
.Y(n_438)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_439),
.B(n_454),
.Y(n_455)
);

XNOR2xp5_ASAP7_75t_SL g439 ( 
.A(n_440),
.B(n_445),
.Y(n_439)
);

XOR2xp5_ASAP7_75t_L g440 ( 
.A(n_441),
.B(n_444),
.Y(n_440)
);

MAJIxp5_ASAP7_75t_L g466 ( 
.A(n_441),
.B(n_444),
.C(n_467),
.Y(n_466)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_442),
.Y(n_443)
);

INVxp67_ASAP7_75t_L g467 ( 
.A(n_445),
.Y(n_467)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_446),
.B(n_449),
.Y(n_445)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_446),
.B(n_450),
.C(n_452),
.Y(n_458)
);

XNOR2xp5_ASAP7_75t_L g449 ( 
.A(n_450),
.B(n_452),
.Y(n_449)
);

NOR2xp33_ASAP7_75t_SL g456 ( 
.A(n_457),
.B(n_466),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_457),
.B(n_466),
.Y(n_468)
);

XNOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

INVx1_ASAP7_75t_L g473 ( 
.A(n_458),
.Y(n_473)
);

XOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_463),
.Y(n_459)
);

MAJIxp5_ASAP7_75t_L g472 ( 
.A(n_460),
.B(n_463),
.C(n_473),
.Y(n_472)
);

NAND2xp5_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_472),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g474 ( 
.A(n_470),
.B(n_472),
.Y(n_474)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

NOR2xp33_ASAP7_75t_SL g477 ( 
.A(n_478),
.B(n_479),
.Y(n_477)
);

NAND2xp5_ASAP7_75t_L g481 ( 
.A(n_478),
.B(n_479),
.Y(n_481)
);

BUFx24_ASAP7_75t_SL g488 ( 
.A(n_478),
.Y(n_488)
);

INVxp67_ASAP7_75t_L g480 ( 
.A(n_481),
.Y(n_480)
);

NOR2xp33_ASAP7_75t_L g485 ( 
.A(n_482),
.B(n_486),
.Y(n_485)
);

BUFx12f_ASAP7_75t_L g482 ( 
.A(n_483),
.Y(n_482)
);

INVx5_ASAP7_75t_L g483 ( 
.A(n_484),
.Y(n_483)
);


endmodule