module fake_jpeg_26118_n_137 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_137);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_137;

wire n_117;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_44;
wire n_24;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_12;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_3),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_11),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_7),
.Y(n_16)
);

INVx3_ASAP7_75t_L g17 ( 
.A(n_11),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_0),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_4),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

INVx3_ASAP7_75t_SL g27 ( 
.A(n_25),
.Y(n_27)
);

BUFx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_16),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_29),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_16),
.B(n_25),
.Y(n_30)
);

AND2x2_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_16),
.Y(n_43)
);

AOI21xp5_ASAP7_75t_L g31 ( 
.A1(n_13),
.A2(n_0),
.B(n_1),
.Y(n_31)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_31),
.B(n_18),
.C(n_21),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g32 ( 
.A(n_25),
.Y(n_32)
);

BUFx10_ASAP7_75t_L g35 ( 
.A(n_32),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_16),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_33),
.Y(n_47)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_34),
.B(n_15),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_36),
.B(n_39),
.Y(n_60)
);

INVxp67_ASAP7_75t_L g39 ( 
.A(n_30),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_29),
.Y(n_42)
);

INVx3_ASAP7_75t_SL g53 ( 
.A(n_42),
.Y(n_53)
);

INVx1_ASAP7_75t_SL g57 ( 
.A(n_43),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_34),
.B(n_14),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g59 ( 
.A(n_44),
.Y(n_59)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_45),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g56 ( 
.A(n_46),
.Y(n_56)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_39),
.A2(n_27),
.B1(n_32),
.B2(n_17),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_48),
.A2(n_52),
.B1(n_61),
.B2(n_19),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_50),
.Y(n_65)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_38),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_51),
.B(n_54),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g52 ( 
.A1(n_43),
.A2(n_27),
.B1(n_32),
.B2(n_17),
.Y(n_52)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_38),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_35),
.Y(n_55)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_55),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_40),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_58),
.B(n_40),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_SL g61 ( 
.A1(n_46),
.A2(n_17),
.B1(n_19),
.B2(n_20),
.Y(n_61)
);

AND2x4_ASAP7_75t_L g62 ( 
.A(n_49),
.B(n_35),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_SL g83 ( 
.A1(n_62),
.A2(n_67),
.B(n_69),
.Y(n_83)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_63),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_64),
.A2(n_54),
.B1(n_51),
.B2(n_48),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_66),
.Y(n_89)
);

O2A1O1Ixp33_ASAP7_75t_L g67 ( 
.A1(n_49),
.A2(n_35),
.B(n_20),
.C(n_22),
.Y(n_67)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_53),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g78 ( 
.A(n_68),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_28),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_70),
.B(n_72),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_56),
.B(n_60),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_50),
.Y(n_73)
);

AOI22xp33_ASAP7_75t_SL g81 ( 
.A1(n_73),
.A2(n_53),
.B1(n_42),
.B2(n_47),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_14),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_74),
.B(n_75),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_59),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_28),
.Y(n_76)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_76),
.B(n_33),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_L g92 ( 
.A1(n_77),
.A2(n_81),
.B1(n_65),
.B2(n_62),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g79 ( 
.A1(n_70),
.A2(n_57),
.B(n_55),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_79),
.B(n_80),
.Y(n_95)
);

NOR2x1_ASAP7_75t_L g80 ( 
.A(n_62),
.B(n_22),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_82),
.B(n_83),
.Y(n_94)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_76),
.B(n_33),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_SL g96 ( 
.A(n_84),
.B(n_33),
.Y(n_96)
);

OAI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_62),
.A2(n_12),
.B1(n_26),
.B2(n_29),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g100 ( 
.A1(n_85),
.A2(n_13),
.B1(n_24),
.B2(n_23),
.Y(n_100)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_90),
.B(n_91),
.Y(n_105)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_78),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g104 ( 
.A1(n_92),
.A2(n_93),
.B1(n_100),
.B2(n_80),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_72),
.B1(n_67),
.B2(n_71),
.Y(n_93)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_96),
.A2(n_79),
.B(n_84),
.Y(n_103)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_86),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_97),
.B(n_98),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g99 ( 
.A(n_82),
.B(n_71),
.C(n_29),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_99),
.B(n_87),
.C(n_89),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_88),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_SL g117 ( 
.A(n_101),
.B(n_24),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_103),
.B(n_106),
.Y(n_114)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_104),
.A2(n_107),
.B(n_100),
.Y(n_112)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_83),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_99),
.B(n_94),
.C(n_84),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g113 ( 
.A(n_108),
.B(n_110),
.C(n_41),
.Y(n_113)
);

INVxp33_ASAP7_75t_SL g109 ( 
.A(n_93),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_66),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_110),
.B(n_97),
.C(n_89),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_111),
.B(n_113),
.C(n_118),
.Y(n_121)
);

XOR2xp5_ASAP7_75t_L g119 ( 
.A(n_112),
.B(n_109),
.Y(n_119)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_115),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_102),
.B(n_105),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_116),
.B(n_117),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_107),
.B(n_41),
.C(n_47),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_119),
.B(n_120),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_114),
.A2(n_23),
.B1(n_21),
.B2(n_18),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_111),
.A2(n_8),
.B1(n_10),
.B2(n_9),
.Y(n_124)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_124),
.A2(n_6),
.B1(n_2),
.B2(n_5),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_41),
.C(n_8),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_125),
.B(n_126),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_121),
.B(n_9),
.C(n_10),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g127 ( 
.A1(n_123),
.A2(n_2),
.B(n_4),
.Y(n_127)
);

AOI21xp5_ASAP7_75t_L g131 ( 
.A1(n_127),
.A2(n_5),
.B(n_6),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_128),
.A2(n_122),
.B(n_124),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_130),
.A2(n_131),
.B1(n_129),
.B2(n_132),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_133),
.B(n_134),
.Y(n_135)
);

NAND3xp33_ASAP7_75t_SL g134 ( 
.A(n_130),
.B(n_123),
.C(n_119),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g136 ( 
.A(n_135),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_136),
.B(n_5),
.Y(n_137)
);


endmodule