module fake_aes_3146_n_32 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
CKINVDCx20_ASAP7_75t_R g12 ( .A(n_3), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_7), .Y(n_13) );
INVxp67_ASAP7_75t_L g14 ( .A(n_4), .Y(n_14) );
CKINVDCx5p33_ASAP7_75t_R g15 ( .A(n_8), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_0), .Y(n_16) );
INVx3_ASAP7_75t_L g17 ( .A(n_11), .Y(n_17) );
NAND2xp5_ASAP7_75t_L g18 ( .A(n_17), .B(n_1), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_12), .Y(n_19) );
INVx1_ASAP7_75t_L g20 ( .A(n_16), .Y(n_20) );
NOR2x1_ASAP7_75t_L g21 ( .A(n_20), .B(n_13), .Y(n_21) );
AOI22xp33_ASAP7_75t_L g22 ( .A1(n_18), .A2(n_14), .B1(n_15), .B2(n_6), .Y(n_22) );
OAI21xp5_ASAP7_75t_L g23 ( .A1(n_22), .A2(n_19), .B(n_5), .Y(n_23) );
OR2x4_ASAP7_75t_L g24 ( .A(n_23), .B(n_21), .Y(n_24) );
INVx1_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
CKINVDCx20_ASAP7_75t_R g27 ( .A(n_25), .Y(n_27) );
INVx2_ASAP7_75t_SL g28 ( .A(n_26), .Y(n_28) );
OR2x2_ASAP7_75t_L g29 ( .A(n_28), .B(n_2), .Y(n_29) );
HB1xp67_ASAP7_75t_L g30 ( .A(n_27), .Y(n_30) );
INVxp67_ASAP7_75t_L g31 ( .A(n_30), .Y(n_31) );
AOI22xp5_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_29), .B1(n_9), .B2(n_10), .Y(n_32) );
endmodule