module fake_aes_3391_n_1027 (n_117, n_219, n_44, n_133, n_149, n_289, n_220, n_81, n_69, n_214, n_267, n_204, n_221, n_249, n_185, n_22, n_203, n_57, n_88, n_52, n_244, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_284, n_107, n_158, n_278, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_240, n_254, n_9, n_161, n_262, n_10, n_177, n_130, n_189, n_103, n_239, n_19, n_87, n_137, n_180, n_104, n_277, n_160, n_98, n_74, n_206, n_276, n_154, n_272, n_7, n_29, n_285, n_195, n_165, n_146, n_45, n_85, n_250, n_237, n_181, n_101, n_62, n_255, n_36, n_47, n_215, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_217, n_139, n_229, n_230, n_274, n_16, n_13, n_198, n_169, n_193, n_273, n_282, n_252, n_152, n_113, n_241, n_95, n_124, n_156, n_238, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_247, n_197, n_201, n_242, n_260, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_210, n_38, n_64, n_142, n_184, n_245, n_265, n_191, n_264, n_281, n_232, n_200, n_46, n_31, n_208, n_211, n_58, n_122, n_187, n_138, n_126, n_275, n_178, n_118, n_258, n_253, n_32, n_0, n_179, n_84, n_131, n_112, n_266, n_55, n_205, n_12, n_86, n_143, n_213, n_235, n_243, n_182, n_263, n_166, n_162, n_186, n_75, n_163, n_226, n_105, n_159, n_174, n_227, n_248, n_268, n_231, n_72, n_136, n_283, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_256, n_67, n_77, n_216, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_212, n_228, n_92, n_11, n_223, n_251, n_25, n_30, n_59, n_236, n_150, n_218, n_168, n_194, n_3, n_287, n_18, n_110, n_261, n_66, n_134, n_222, n_234, n_1, n_164, n_233, n_271, n_82, n_106, n_175, n_15, n_173, n_190, n_286, n_145, n_270, n_246, n_153, n_61, n_259, n_280, n_21, n_99, n_109, n_93, n_132, n_288, n_151, n_51, n_140, n_207, n_257, n_224, n_96, n_269, n_225, n_39, n_279, n_1027);
input n_117;
input n_219;
input n_44;
input n_133;
input n_149;
input n_289;
input n_220;
input n_81;
input n_69;
input n_214;
input n_267;
input n_204;
input n_221;
input n_249;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_244;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_284;
input n_107;
input n_158;
input n_278;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_240;
input n_254;
input n_9;
input n_161;
input n_262;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_239;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_277;
input n_160;
input n_98;
input n_74;
input n_206;
input n_276;
input n_154;
input n_272;
input n_7;
input n_29;
input n_285;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_250;
input n_237;
input n_181;
input n_101;
input n_62;
input n_255;
input n_36;
input n_47;
input n_215;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_217;
input n_139;
input n_229;
input n_230;
input n_274;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_273;
input n_282;
input n_252;
input n_152;
input n_113;
input n_241;
input n_95;
input n_124;
input n_156;
input n_238;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_247;
input n_197;
input n_201;
input n_242;
input n_260;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_210;
input n_38;
input n_64;
input n_142;
input n_184;
input n_245;
input n_265;
input n_191;
input n_264;
input n_281;
input n_232;
input n_200;
input n_46;
input n_31;
input n_208;
input n_211;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_275;
input n_178;
input n_118;
input n_258;
input n_253;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_266;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_213;
input n_235;
input n_243;
input n_182;
input n_263;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_226;
input n_105;
input n_159;
input n_174;
input n_227;
input n_248;
input n_268;
input n_231;
input n_72;
input n_136;
input n_283;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_256;
input n_67;
input n_77;
input n_216;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_212;
input n_228;
input n_92;
input n_11;
input n_223;
input n_251;
input n_25;
input n_30;
input n_59;
input n_236;
input n_150;
input n_218;
input n_168;
input n_194;
input n_3;
input n_287;
input n_18;
input n_110;
input n_261;
input n_66;
input n_134;
input n_222;
input n_234;
input n_1;
input n_164;
input n_233;
input n_271;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_286;
input n_145;
input n_270;
input n_246;
input n_153;
input n_61;
input n_259;
input n_280;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_288;
input n_151;
input n_51;
input n_140;
input n_207;
input n_257;
input n_224;
input n_96;
input n_269;
input n_225;
input n_39;
input n_279;
output n_1027;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_963;
wire n_838;
wire n_705;
wire n_949;
wire n_998;
wire n_603;
wire n_604;
wire n_858;
wire n_964;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_500;
wire n_925;
wire n_848;
wire n_607;
wire n_957;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_988;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_958;
wire n_328;
wire n_655;
wire n_468;
wire n_917;
wire n_743;
wire n_523;
wire n_903;
wire n_920;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_965;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_918;
wire n_1022;
wire n_878;
wire n_814;
wire n_911;
wire n_980;
wire n_637;
wire n_999;
wire n_817;
wire n_985;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_993;
wire n_779;
wire n_528;
wire n_383;
wire n_971;
wire n_904;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_981;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_987;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_462;
wire n_1015;
wire n_316;
wire n_545;
wire n_896;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_1019;
wire n_940;
wire n_715;
wire n_463;
wire n_789;
wire n_973;
wire n_330;
wire n_1003;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_476;
wire n_434;
wire n_384;
wire n_617;
wire n_452;
wire n_518;
wire n_978;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_752;
wire n_732;
wire n_1012;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_786;
wire n_724;
wire n_857;
wire n_360;
wire n_345;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_922;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_914;
wire n_909;
wire n_366;
wire n_927;
wire n_596;
wire n_1005;
wire n_951;
wire n_321;
wire n_702;
wire n_1016;
wire n_1024;
wire n_572;
wire n_1017;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_968;
wire n_303;
wire n_975;
wire n_437;
wire n_512;
wire n_326;
wire n_333;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_540;
wire n_563;
wire n_638;
wire n_937;
wire n_517;
wire n_560;
wire n_945;
wire n_479;
wire n_623;
wire n_593;
wire n_955;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_897;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_1009;
wire n_502;
wire n_921;
wire n_543;
wire n_1010;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_1011;
wire n_1025;
wire n_880;
wire n_630;
wire n_511;
wire n_1002;
wire n_467;
wire n_692;
wire n_865;
wire n_915;
wire n_647;
wire n_367;
wire n_644;
wire n_764;
wire n_314;
wire n_426;
wire n_624;
wire n_725;
wire n_818;
wire n_769;
wire n_844;
wire n_1018;
wire n_738;
wire n_979;
wire n_319;
wire n_969;
wire n_499;
wire n_895;
wire n_417;
wire n_798;
wire n_575;
wire n_711;
wire n_977;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_1014;
wire n_828;
wire n_767;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_863;
wire n_322;
wire n_310;
wire n_907;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_696;
wire n_735;
wire n_771;
wire n_784;
wire n_1013;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_1000;
wire n_939;
wire n_953;
wire n_413;
wire n_676;
wire n_391;
wire n_910;
wire n_427;
wire n_935;
wire n_950;
wire n_460;
wire n_478;
wire n_482;
wire n_415;
wire n_394;
wire n_703;
wire n_442;
wire n_331;
wire n_485;
wire n_938;
wire n_928;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_501;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_729;
wire n_699;
wire n_805;
wire n_693;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_961;
wire n_995;
wire n_1020;
wire n_982;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_905;
wire n_902;
wire n_525;
wire n_876;
wire n_886;
wire n_986;
wire n_959;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_760;
wire n_941;
wire n_751;
wire n_800;
wire n_626;
wire n_990;
wire n_302;
wire n_466;
wire n_900;
wire n_952;
wire n_710;
wire n_685;
wire n_362;
wire n_931;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_788;
wire n_475;
wire n_926;
wire n_578;
wire n_542;
wire n_537;
wire n_660;
wire n_430;
wire n_839;
wire n_1001;
wire n_943;
wire n_450;
wire n_936;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_549;
wire n_622;
wire n_832;
wire n_556;
wire n_439;
wire n_601;
wire n_996;
wire n_379;
wire n_641;
wire n_966;
wire n_614;
wire n_527;
wire n_526;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_420;
wire n_446;
wire n_666;
wire n_423;
wire n_342;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_954;
wire n_643;
wire n_574;
wire n_874;
wire n_388;
wire n_454;
wire n_687;
wire n_505;
wire n_706;
wire n_970;
wire n_822;
wire n_823;
wire n_984;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_906;
wire n_720;
wire n_568;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_899;
wire n_806;
wire n_539;
wire n_974;
wire n_591;
wire n_933;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_956;
wire n_522;
wire n_883;
wire n_573;
wire n_948;
wire n_898;
wire n_989;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_315;
wire n_363;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_1023;
wire n_503;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_577;
wire n_870;
wire n_942;
wire n_790;
wire n_761;
wire n_615;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_445;
wire n_398;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_908;
wire n_429;
wire n_488;
wire n_763;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_944;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_972;
wire n_1021;
wire n_811;
wire n_749;
wire n_835;
wire n_535;
wire n_1006;
wire n_530;
wire n_737;
wire n_778;
wire n_358;
wire n_795;
wire n_456;
wire n_962;
wire n_782;
wire n_449;
wire n_997;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_919;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_912;
wire n_620;
wire n_841;
wire n_924;
wire n_947;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_923;
wire n_561;
wire n_335;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_1008;
wire n_1026;
wire n_306;
wire n_766;
wire n_602;
wire n_831;
wire n_1007;
wire n_859;
wire n_930;
wire n_994;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_932;
wire n_837;
wire n_946;
wire n_960;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_830;
wire n_510;
wire n_343;
wire n_675;
wire n_967;
wire n_291;
wire n_504;
wire n_458;
wire n_581;
wire n_493;
wire n_418;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_901;
wire n_727;
wire n_690;
wire n_356;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_991;
wire n_558;
wire n_515;
wire n_670;
wire n_843;
wire n_820;
wire n_1004;
wire n_683;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_929;
wire n_753;
wire n_368;
wire n_355;
wire n_976;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_913;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_494;
wire n_559;
wire n_480;
wire n_453;
wire n_372;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_934;
wire n_350;
wire n_433;
wire n_983;
wire n_781;
wire n_916;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_992;
INVx1_ASAP7_75t_SL g290 ( .A(n_125), .Y(n_290) );
CKINVDCx20_ASAP7_75t_R g291 ( .A(n_262), .Y(n_291) );
CKINVDCx5p33_ASAP7_75t_R g292 ( .A(n_245), .Y(n_292) );
BUFx6f_ASAP7_75t_L g293 ( .A(n_231), .Y(n_293) );
CKINVDCx5p33_ASAP7_75t_R g294 ( .A(n_191), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_209), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_100), .Y(n_296) );
CKINVDCx5p33_ASAP7_75t_R g297 ( .A(n_244), .Y(n_297) );
CKINVDCx5p33_ASAP7_75t_R g298 ( .A(n_180), .Y(n_298) );
BUFx2_ASAP7_75t_L g299 ( .A(n_230), .Y(n_299) );
INVx2_ASAP7_75t_L g300 ( .A(n_264), .Y(n_300) );
CKINVDCx5p33_ASAP7_75t_R g301 ( .A(n_253), .Y(n_301) );
INVx1_ASAP7_75t_L g302 ( .A(n_252), .Y(n_302) );
CKINVDCx16_ASAP7_75t_R g303 ( .A(n_5), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_10), .Y(n_304) );
CKINVDCx5p33_ASAP7_75t_R g305 ( .A(n_223), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_65), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_256), .Y(n_307) );
CKINVDCx5p33_ASAP7_75t_R g308 ( .A(n_257), .Y(n_308) );
CKINVDCx5p33_ASAP7_75t_R g309 ( .A(n_172), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_61), .Y(n_310) );
INVx1_ASAP7_75t_L g311 ( .A(n_50), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_242), .Y(n_312) );
CKINVDCx5p33_ASAP7_75t_R g313 ( .A(n_73), .Y(n_313) );
CKINVDCx5p33_ASAP7_75t_R g314 ( .A(n_203), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_200), .Y(n_315) );
INVx1_ASAP7_75t_L g316 ( .A(n_77), .Y(n_316) );
CKINVDCx20_ASAP7_75t_R g317 ( .A(n_259), .Y(n_317) );
NOR2xp67_ASAP7_75t_L g318 ( .A(n_101), .B(n_123), .Y(n_318) );
BUFx5_ASAP7_75t_L g319 ( .A(n_277), .Y(n_319) );
CKINVDCx5p33_ASAP7_75t_R g320 ( .A(n_281), .Y(n_320) );
BUFx6f_ASAP7_75t_L g321 ( .A(n_267), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_127), .Y(n_322) );
CKINVDCx5p33_ASAP7_75t_R g323 ( .A(n_16), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_250), .Y(n_324) );
CKINVDCx5p33_ASAP7_75t_R g325 ( .A(n_30), .Y(n_325) );
BUFx3_ASAP7_75t_L g326 ( .A(n_278), .Y(n_326) );
CKINVDCx5p33_ASAP7_75t_R g327 ( .A(n_121), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_33), .Y(n_328) );
CKINVDCx5p33_ASAP7_75t_R g329 ( .A(n_67), .Y(n_329) );
CKINVDCx5p33_ASAP7_75t_R g330 ( .A(n_232), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_110), .Y(n_331) );
CKINVDCx5p33_ASAP7_75t_R g332 ( .A(n_43), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_246), .Y(n_333) );
BUFx10_ASAP7_75t_L g334 ( .A(n_219), .Y(n_334) );
BUFx6f_ASAP7_75t_L g335 ( .A(n_3), .Y(n_335) );
INVx1_ASAP7_75t_SL g336 ( .A(n_62), .Y(n_336) );
BUFx10_ASAP7_75t_L g337 ( .A(n_40), .Y(n_337) );
CKINVDCx5p33_ASAP7_75t_R g338 ( .A(n_42), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_270), .Y(n_339) );
INVx1_ASAP7_75t_L g340 ( .A(n_265), .Y(n_340) );
CKINVDCx5p33_ASAP7_75t_R g341 ( .A(n_161), .Y(n_341) );
CKINVDCx5p33_ASAP7_75t_R g342 ( .A(n_38), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_156), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_248), .Y(n_344) );
NOR2xp67_ASAP7_75t_L g345 ( .A(n_105), .B(n_22), .Y(n_345) );
INVx1_ASAP7_75t_L g346 ( .A(n_44), .Y(n_346) );
CKINVDCx5p33_ASAP7_75t_R g347 ( .A(n_107), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_60), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_120), .Y(n_349) );
HB1xp67_ASAP7_75t_L g350 ( .A(n_141), .Y(n_350) );
INVx2_ASAP7_75t_L g351 ( .A(n_279), .Y(n_351) );
CKINVDCx20_ASAP7_75t_R g352 ( .A(n_34), .Y(n_352) );
INVx1_ASAP7_75t_SL g353 ( .A(n_192), .Y(n_353) );
CKINVDCx5p33_ASAP7_75t_R g354 ( .A(n_261), .Y(n_354) );
CKINVDCx5p33_ASAP7_75t_R g355 ( .A(n_12), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_21), .Y(n_356) );
INVx1_ASAP7_75t_L g357 ( .A(n_226), .Y(n_357) );
CKINVDCx5p33_ASAP7_75t_R g358 ( .A(n_216), .Y(n_358) );
BUFx6f_ASAP7_75t_L g359 ( .A(n_108), .Y(n_359) );
CKINVDCx20_ASAP7_75t_R g360 ( .A(n_237), .Y(n_360) );
CKINVDCx16_ASAP7_75t_R g361 ( .A(n_51), .Y(n_361) );
CKINVDCx20_ASAP7_75t_R g362 ( .A(n_243), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_234), .Y(n_363) );
BUFx10_ASAP7_75t_L g364 ( .A(n_251), .Y(n_364) );
INVx2_ASAP7_75t_SL g365 ( .A(n_136), .Y(n_365) );
INVxp67_ASAP7_75t_SL g366 ( .A(n_186), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_89), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_233), .Y(n_368) );
INVx2_ASAP7_75t_L g369 ( .A(n_88), .Y(n_369) );
CKINVDCx20_ASAP7_75t_R g370 ( .A(n_193), .Y(n_370) );
CKINVDCx5p33_ASAP7_75t_R g371 ( .A(n_205), .Y(n_371) );
CKINVDCx5p33_ASAP7_75t_R g372 ( .A(n_249), .Y(n_372) );
CKINVDCx5p33_ASAP7_75t_R g373 ( .A(n_84), .Y(n_373) );
CKINVDCx16_ASAP7_75t_R g374 ( .A(n_240), .Y(n_374) );
INVx1_ASAP7_75t_L g375 ( .A(n_159), .Y(n_375) );
INVx1_ASAP7_75t_SL g376 ( .A(n_27), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_112), .Y(n_377) );
INVx1_ASAP7_75t_L g378 ( .A(n_285), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_266), .Y(n_379) );
CKINVDCx5p33_ASAP7_75t_R g380 ( .A(n_228), .Y(n_380) );
INVx1_ASAP7_75t_L g381 ( .A(n_206), .Y(n_381) );
CKINVDCx5p33_ASAP7_75t_R g382 ( .A(n_196), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_124), .Y(n_383) );
CKINVDCx20_ASAP7_75t_R g384 ( .A(n_260), .Y(n_384) );
NOR2xp67_ASAP7_75t_L g385 ( .A(n_163), .B(n_241), .Y(n_385) );
BUFx3_ASAP7_75t_L g386 ( .A(n_268), .Y(n_386) );
BUFx10_ASAP7_75t_L g387 ( .A(n_82), .Y(n_387) );
INVx1_ASAP7_75t_L g388 ( .A(n_214), .Y(n_388) );
BUFx6f_ASAP7_75t_L g389 ( .A(n_23), .Y(n_389) );
CKINVDCx5p33_ASAP7_75t_R g390 ( .A(n_258), .Y(n_390) );
INVx1_ASAP7_75t_L g391 ( .A(n_272), .Y(n_391) );
CKINVDCx5p33_ASAP7_75t_R g392 ( .A(n_276), .Y(n_392) );
CKINVDCx5p33_ASAP7_75t_R g393 ( .A(n_102), .Y(n_393) );
OR2x2_ASAP7_75t_L g394 ( .A(n_151), .B(n_176), .Y(n_394) );
INVx1_ASAP7_75t_L g395 ( .A(n_75), .Y(n_395) );
BUFx6f_ASAP7_75t_L g396 ( .A(n_239), .Y(n_396) );
CKINVDCx5p33_ASAP7_75t_R g397 ( .A(n_255), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_254), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_263), .Y(n_399) );
INVx1_ASAP7_75t_SL g400 ( .A(n_273), .Y(n_400) );
INVx2_ASAP7_75t_L g401 ( .A(n_170), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_145), .Y(n_402) );
BUFx6f_ASAP7_75t_L g403 ( .A(n_280), .Y(n_403) );
CKINVDCx20_ASAP7_75t_R g404 ( .A(n_71), .Y(n_404) );
INVx1_ASAP7_75t_L g405 ( .A(n_45), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_194), .Y(n_406) );
INVx1_ASAP7_75t_L g407 ( .A(n_247), .Y(n_407) );
INVx1_ASAP7_75t_L g408 ( .A(n_148), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_269), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_17), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_41), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_204), .Y(n_412) );
CKINVDCx5p33_ASAP7_75t_R g413 ( .A(n_275), .Y(n_413) );
CKINVDCx5p33_ASAP7_75t_R g414 ( .A(n_271), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_18), .Y(n_415) );
CKINVDCx5p33_ASAP7_75t_R g416 ( .A(n_111), .Y(n_416) );
INVx1_ASAP7_75t_L g417 ( .A(n_274), .Y(n_417) );
INVx1_ASAP7_75t_L g418 ( .A(n_90), .Y(n_418) );
INVxp67_ASAP7_75t_L g419 ( .A(n_87), .Y(n_419) );
CKINVDCx6p67_ASAP7_75t_R g420 ( .A(n_334), .Y(n_420) );
INVx2_ASAP7_75t_L g421 ( .A(n_319), .Y(n_421) );
AND2x4_ASAP7_75t_L g422 ( .A(n_299), .B(n_0), .Y(n_422) );
INVx2_ASAP7_75t_L g423 ( .A(n_319), .Y(n_423) );
BUFx8_ASAP7_75t_L g424 ( .A(n_335), .Y(n_424) );
INVx1_ASAP7_75t_L g425 ( .A(n_350), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_302), .Y(n_426) );
BUFx6f_ASAP7_75t_L g427 ( .A(n_293), .Y(n_427) );
OAI21x1_ASAP7_75t_L g428 ( .A1(n_300), .A2(n_20), .B(n_19), .Y(n_428) );
INVx1_ASAP7_75t_L g429 ( .A(n_306), .Y(n_429) );
AND2x4_ASAP7_75t_L g430 ( .A(n_365), .B(n_0), .Y(n_430) );
INVx5_ASAP7_75t_L g431 ( .A(n_337), .Y(n_431) );
AND2x4_ASAP7_75t_L g432 ( .A(n_304), .B(n_1), .Y(n_432) );
INVx2_ASAP7_75t_L g433 ( .A(n_319), .Y(n_433) );
INVxp33_ASAP7_75t_SL g434 ( .A(n_323), .Y(n_434) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_293), .Y(n_435) );
INVx5_ASAP7_75t_L g436 ( .A(n_364), .Y(n_436) );
INVx6_ASAP7_75t_L g437 ( .A(n_387), .Y(n_437) );
INVx2_ASAP7_75t_L g438 ( .A(n_319), .Y(n_438) );
INVx1_ASAP7_75t_L g439 ( .A(n_307), .Y(n_439) );
INVx2_ASAP7_75t_L g440 ( .A(n_351), .Y(n_440) );
INVx2_ASAP7_75t_L g441 ( .A(n_369), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_421), .Y(n_442) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_426), .B(n_401), .Y(n_443) );
NAND2xp5_ASAP7_75t_SL g444 ( .A(n_431), .B(n_361), .Y(n_444) );
INVx1_ASAP7_75t_L g445 ( .A(n_423), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_426), .B(n_406), .Y(n_446) );
INVx2_ASAP7_75t_SL g447 ( .A(n_437), .Y(n_447) );
INVx2_ASAP7_75t_L g448 ( .A(n_433), .Y(n_448) );
INVxp33_ASAP7_75t_L g449 ( .A(n_425), .Y(n_449) );
INVx2_ASAP7_75t_L g450 ( .A(n_438), .Y(n_450) );
NAND3xp33_ASAP7_75t_L g451 ( .A(n_422), .B(n_355), .C(n_335), .Y(n_451) );
NAND2xp5_ASAP7_75t_SL g452 ( .A(n_431), .B(n_374), .Y(n_452) );
NAND2xp33_ASAP7_75t_L g453 ( .A(n_429), .B(n_292), .Y(n_453) );
INVxp67_ASAP7_75t_L g454 ( .A(n_429), .Y(n_454) );
AND2x2_ASAP7_75t_L g455 ( .A(n_420), .B(n_303), .Y(n_455) );
INVx1_ASAP7_75t_L g456 ( .A(n_432), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_440), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_430), .Y(n_458) );
AOI21x1_ASAP7_75t_L g459 ( .A1(n_428), .A2(n_311), .B(n_310), .Y(n_459) );
NAND2xp5_ASAP7_75t_SL g460 ( .A(n_431), .B(n_419), .Y(n_460) );
INVx2_ASAP7_75t_L g461 ( .A(n_442), .Y(n_461) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_454), .B(n_439), .Y(n_462) );
A2O1A1Ixp33_ASAP7_75t_L g463 ( .A1(n_454), .A2(n_439), .B(n_441), .C(n_312), .Y(n_463) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_449), .B(n_434), .Y(n_464) );
INVx2_ASAP7_75t_L g465 ( .A(n_448), .Y(n_465) );
AND2x4_ASAP7_75t_L g466 ( .A(n_458), .B(n_436), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_450), .Y(n_467) );
BUFx3_ASAP7_75t_L g468 ( .A(n_447), .Y(n_468) );
AO221x1_ASAP7_75t_L g469 ( .A1(n_456), .A2(n_317), .B1(n_352), .B2(n_315), .C(n_291), .Y(n_469) );
NOR2xp67_ASAP7_75t_L g470 ( .A(n_451), .B(n_394), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g471 ( .A(n_443), .B(n_436), .Y(n_471) );
AND2x6_ASAP7_75t_SL g472 ( .A(n_455), .B(n_424), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_443), .B(n_436), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g474 ( .A(n_444), .B(n_294), .Y(n_474) );
NAND2xp5_ASAP7_75t_SL g475 ( .A(n_452), .B(n_295), .Y(n_475) );
OR2x6_ASAP7_75t_L g476 ( .A(n_460), .B(n_437), .Y(n_476) );
AND2x6_ASAP7_75t_SL g477 ( .A(n_446), .B(n_316), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_446), .Y(n_478) );
INVx1_ASAP7_75t_L g479 ( .A(n_457), .Y(n_479) );
NOR2xp33_ASAP7_75t_L g480 ( .A(n_453), .B(n_290), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g481 ( .A(n_445), .B(n_296), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_459), .B(n_336), .Y(n_482) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_454), .A2(n_324), .B(n_331), .C(n_328), .Y(n_483) );
NAND2xp33_ASAP7_75t_L g484 ( .A(n_458), .B(n_297), .Y(n_484) );
NAND2xp5_ASAP7_75t_SL g485 ( .A(n_454), .B(n_298), .Y(n_485) );
NAND2xp5_ASAP7_75t_SL g486 ( .A(n_454), .B(n_301), .Y(n_486) );
AOI22xp5_ASAP7_75t_L g487 ( .A1(n_478), .A2(n_362), .B1(n_370), .B2(n_360), .Y(n_487) );
BUFx12f_ASAP7_75t_L g488 ( .A(n_472), .Y(n_488) );
CKINVDCx8_ASAP7_75t_R g489 ( .A(n_477), .Y(n_489) );
BUFx4f_ASAP7_75t_L g490 ( .A(n_476), .Y(n_490) );
BUFx3_ASAP7_75t_L g491 ( .A(n_468), .Y(n_491) );
A2O1A1Ixp33_ASAP7_75t_L g492 ( .A1(n_462), .A2(n_333), .B(n_340), .C(n_339), .Y(n_492) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_464), .B(n_384), .Y(n_493) );
INVx2_ASAP7_75t_L g494 ( .A(n_479), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_482), .A2(n_366), .B(n_346), .Y(n_495) );
NOR2x1_ASAP7_75t_L g496 ( .A(n_476), .B(n_404), .Y(n_496) );
NOR2x1_ASAP7_75t_L g497 ( .A(n_470), .B(n_344), .Y(n_497) );
INVx1_ASAP7_75t_L g498 ( .A(n_461), .Y(n_498) );
AOI21xp5_ASAP7_75t_L g499 ( .A1(n_481), .A2(n_349), .B(n_348), .Y(n_499) );
CKINVDCx5p33_ASAP7_75t_R g500 ( .A(n_466), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g501 ( .A(n_474), .Y(n_501) );
NOR3xp33_ASAP7_75t_L g502 ( .A(n_484), .B(n_376), .C(n_353), .Y(n_502) );
OAI21xp5_ASAP7_75t_L g503 ( .A1(n_463), .A2(n_357), .B(n_356), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_483), .B(n_305), .Y(n_504) );
INVx2_ASAP7_75t_L g505 ( .A(n_465), .Y(n_505) );
OAI21xp5_ASAP7_75t_L g506 ( .A1(n_467), .A2(n_367), .B(n_363), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_470), .A2(n_375), .B(n_377), .C(n_368), .Y(n_507) );
AOI21xp5_ASAP7_75t_L g508 ( .A1(n_485), .A2(n_486), .B(n_473), .Y(n_508) );
AOI22xp5_ASAP7_75t_L g509 ( .A1(n_466), .A2(n_379), .B1(n_381), .B2(n_378), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_475), .B(n_400), .Y(n_510) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_471), .A2(n_388), .B(n_383), .Y(n_511) );
INVx1_ASAP7_75t_L g512 ( .A(n_480), .Y(n_512) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_469), .B(n_308), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_478), .B(n_309), .Y(n_514) );
AOI22xp5_ASAP7_75t_L g515 ( .A1(n_478), .A2(n_395), .B1(n_398), .B2(n_391), .Y(n_515) );
AOI22xp33_ASAP7_75t_L g516 ( .A1(n_493), .A2(n_402), .B1(n_405), .B2(n_399), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_512), .B(n_407), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g518 ( .A(n_492), .B(n_408), .Y(n_518) );
OAI22xp5_ASAP7_75t_L g519 ( .A1(n_487), .A2(n_314), .B1(n_320), .B2(n_313), .Y(n_519) );
BUFx8_ASAP7_75t_L g520 ( .A(n_488), .Y(n_520) );
OAI21x1_ASAP7_75t_L g521 ( .A1(n_508), .A2(n_410), .B(n_409), .Y(n_521) );
INVx4_ASAP7_75t_L g522 ( .A(n_491), .Y(n_522) );
AND2x6_ASAP7_75t_L g523 ( .A(n_496), .B(n_411), .Y(n_523) );
OAI22xp5_ASAP7_75t_L g524 ( .A1(n_487), .A2(n_322), .B1(n_327), .B2(n_325), .Y(n_524) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_495), .A2(n_415), .B(n_412), .Y(n_525) );
OAI21xp5_ASAP7_75t_L g526 ( .A1(n_499), .A2(n_418), .B(n_417), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_515), .B(n_329), .Y(n_527) );
OAI21x1_ASAP7_75t_L g528 ( .A1(n_506), .A2(n_345), .B(n_318), .Y(n_528) );
NAND2xp5_ASAP7_75t_SL g529 ( .A(n_514), .B(n_330), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g530 ( .A(n_507), .B(n_332), .Y(n_530) );
INVx1_ASAP7_75t_L g531 ( .A(n_494), .Y(n_531) );
A2O1A1Ixp33_ASAP7_75t_L g532 ( .A1(n_511), .A2(n_385), .B(n_326), .C(n_343), .Y(n_532) );
OAI21x1_ASAP7_75t_L g533 ( .A1(n_497), .A2(n_359), .B(n_321), .Y(n_533) );
OAI21x1_ASAP7_75t_L g534 ( .A1(n_503), .A2(n_359), .B(n_321), .Y(n_534) );
AO31x2_ASAP7_75t_L g535 ( .A1(n_498), .A2(n_389), .A3(n_403), .B(n_396), .Y(n_535) );
OAI21x1_ASAP7_75t_L g536 ( .A1(n_505), .A2(n_396), .B(n_389), .Y(n_536) );
AOI21xp5_ASAP7_75t_L g537 ( .A1(n_504), .A2(n_341), .B(n_338), .Y(n_537) );
HB1xp67_ASAP7_75t_L g538 ( .A(n_500), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_509), .Y(n_539) );
INVx3_ASAP7_75t_L g540 ( .A(n_489), .Y(n_540) );
AND2x4_ASAP7_75t_L g541 ( .A(n_502), .B(n_386), .Y(n_541) );
AO31x2_ASAP7_75t_L g542 ( .A1(n_510), .A2(n_403), .A3(n_435), .B(n_427), .Y(n_542) );
OA22x2_ASAP7_75t_L g543 ( .A1(n_513), .A2(n_347), .B1(n_354), .B2(n_342), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_490), .B(n_358), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g545 ( .A1(n_490), .A2(n_372), .B(n_371), .Y(n_545) );
AND2x2_ASAP7_75t_L g546 ( .A(n_501), .B(n_1), .Y(n_546) );
INVx2_ASAP7_75t_L g547 ( .A(n_494), .Y(n_547) );
NAND2xp5_ASAP7_75t_L g548 ( .A(n_512), .B(n_373), .Y(n_548) );
AOI21xp5_ASAP7_75t_L g549 ( .A1(n_495), .A2(n_382), .B(n_380), .Y(n_549) );
OAI21x1_ASAP7_75t_L g550 ( .A1(n_508), .A2(n_25), .B(n_24), .Y(n_550) );
OAI21x1_ASAP7_75t_L g551 ( .A1(n_534), .A2(n_28), .B(n_26), .Y(n_551) );
INVx2_ASAP7_75t_L g552 ( .A(n_547), .Y(n_552) );
AOI21xp5_ASAP7_75t_SL g553 ( .A1(n_532), .A2(n_392), .B(n_390), .Y(n_553) );
AOI22xp33_ASAP7_75t_L g554 ( .A1(n_539), .A2(n_523), .B1(n_541), .B2(n_543), .Y(n_554) );
INVx3_ASAP7_75t_L g555 ( .A(n_522), .Y(n_555) );
INVx6_ASAP7_75t_L g556 ( .A(n_520), .Y(n_556) );
AOI21xp5_ASAP7_75t_L g557 ( .A1(n_517), .A2(n_397), .B(n_393), .Y(n_557) );
HB1xp67_ASAP7_75t_L g558 ( .A(n_531), .Y(n_558) );
INVx2_ASAP7_75t_L g559 ( .A(n_521), .Y(n_559) );
BUFx12f_ASAP7_75t_L g560 ( .A(n_523), .Y(n_560) );
INVx1_ASAP7_75t_SL g561 ( .A(n_538), .Y(n_561) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_527), .A2(n_414), .B1(n_416), .B2(n_413), .Y(n_562) );
AOI22xp33_ASAP7_75t_L g563 ( .A1(n_523), .A2(n_435), .B1(n_427), .B2(n_4), .Y(n_563) );
OAI21x1_ASAP7_75t_L g564 ( .A1(n_536), .A2(n_31), .B(n_29), .Y(n_564) );
OAI22xp5_ASAP7_75t_SL g565 ( .A1(n_540), .A2(n_4), .B1(n_2), .B2(n_3), .Y(n_565) );
INVx5_ASAP7_75t_L g566 ( .A(n_546), .Y(n_566) );
AO21x2_ASAP7_75t_L g567 ( .A1(n_528), .A2(n_35), .B(n_32), .Y(n_567) );
BUFx4_ASAP7_75t_R g568 ( .A(n_545), .Y(n_568) );
INVx1_ASAP7_75t_L g569 ( .A(n_518), .Y(n_569) );
INVx1_ASAP7_75t_L g570 ( .A(n_533), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_526), .A2(n_37), .B(n_36), .Y(n_571) );
INVx1_ASAP7_75t_L g572 ( .A(n_548), .Y(n_572) );
OAI221xp5_ASAP7_75t_L g573 ( .A1(n_516), .A2(n_2), .B1(n_5), .B2(n_6), .C(n_7), .Y(n_573) );
NOR2xp67_ASAP7_75t_L g574 ( .A(n_544), .B(n_6), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_541), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_542), .Y(n_576) );
OA21x2_ASAP7_75t_L g577 ( .A1(n_550), .A2(n_46), .B(n_39), .Y(n_577) );
O2A1O1Ixp33_ASAP7_75t_SL g578 ( .A1(n_529), .A2(n_48), .B(n_49), .C(n_47), .Y(n_578) );
INVxp67_ASAP7_75t_L g579 ( .A(n_519), .Y(n_579) );
INVx1_ASAP7_75t_L g580 ( .A(n_525), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_542), .Y(n_581) );
INVx1_ASAP7_75t_L g582 ( .A(n_535), .Y(n_582) );
INVx1_ASAP7_75t_L g583 ( .A(n_535), .Y(n_583) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_530), .B(n_7), .Y(n_584) );
INVx1_ASAP7_75t_L g585 ( .A(n_537), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_549), .Y(n_586) );
AND2x4_ASAP7_75t_L g587 ( .A(n_524), .B(n_8), .Y(n_587) );
OAI21x1_ASAP7_75t_L g588 ( .A1(n_534), .A2(n_53), .B(n_52), .Y(n_588) );
OAI21x1_ASAP7_75t_L g589 ( .A1(n_534), .A2(n_55), .B(n_54), .Y(n_589) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_522), .B(n_8), .Y(n_590) );
CKINVDCx5p33_ASAP7_75t_R g591 ( .A(n_520), .Y(n_591) );
INVx2_ASAP7_75t_L g592 ( .A(n_547), .Y(n_592) );
OAI21x1_ASAP7_75t_SL g593 ( .A1(n_547), .A2(n_9), .B(n_10), .Y(n_593) );
OAI21x1_ASAP7_75t_L g594 ( .A1(n_534), .A2(n_57), .B(n_56), .Y(n_594) );
OAI21x1_ASAP7_75t_L g595 ( .A1(n_534), .A2(n_59), .B(n_58), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_547), .Y(n_596) );
INVx2_ASAP7_75t_L g597 ( .A(n_547), .Y(n_597) );
AO21x2_ASAP7_75t_L g598 ( .A1(n_534), .A2(n_64), .B(n_63), .Y(n_598) );
OAI21x1_ASAP7_75t_L g599 ( .A1(n_534), .A2(n_68), .B(n_66), .Y(n_599) );
INVx2_ASAP7_75t_L g600 ( .A(n_547), .Y(n_600) );
O2A1O1Ixp33_ASAP7_75t_SL g601 ( .A1(n_532), .A2(n_70), .B(n_72), .C(n_69), .Y(n_601) );
OAI21x1_ASAP7_75t_L g602 ( .A1(n_534), .A2(n_76), .B(n_74), .Y(n_602) );
AND2x2_ASAP7_75t_L g603 ( .A(n_558), .B(n_9), .Y(n_603) );
AND2x2_ASAP7_75t_L g604 ( .A(n_572), .B(n_11), .Y(n_604) );
AO21x2_ASAP7_75t_L g605 ( .A1(n_582), .A2(n_583), .B(n_581), .Y(n_605) );
OAI21x1_ASAP7_75t_SL g606 ( .A1(n_593), .A2(n_11), .B(n_12), .Y(n_606) );
INVx2_ASAP7_75t_L g607 ( .A(n_596), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_596), .Y(n_608) );
INVx2_ASAP7_75t_L g609 ( .A(n_552), .Y(n_609) );
INVx2_ASAP7_75t_SL g610 ( .A(n_556), .Y(n_610) );
AND2x2_ASAP7_75t_L g611 ( .A(n_587), .B(n_13), .Y(n_611) );
NOR2xp33_ASAP7_75t_L g612 ( .A(n_575), .B(n_13), .Y(n_612) );
BUFx2_ASAP7_75t_L g613 ( .A(n_555), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_592), .Y(n_614) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_579), .B(n_14), .Y(n_615) );
BUFx2_ASAP7_75t_L g616 ( .A(n_555), .Y(n_616) );
NAND2xp33_ASAP7_75t_R g617 ( .A(n_587), .B(n_14), .Y(n_617) );
INVx1_ASAP7_75t_L g618 ( .A(n_597), .Y(n_618) );
INVx2_ASAP7_75t_L g619 ( .A(n_600), .Y(n_619) );
INVx2_ASAP7_75t_L g620 ( .A(n_569), .Y(n_620) );
OAI211xp5_ASAP7_75t_L g621 ( .A1(n_554), .A2(n_15), .B(n_16), .C(n_78), .Y(n_621) );
INVx1_ASAP7_75t_L g622 ( .A(n_590), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_574), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_584), .Y(n_624) );
OAI21x1_ASAP7_75t_L g625 ( .A1(n_559), .A2(n_80), .B(n_79), .Y(n_625) );
BUFx2_ASAP7_75t_SL g626 ( .A(n_566), .Y(n_626) );
INVx1_ASAP7_75t_L g627 ( .A(n_580), .Y(n_627) );
OAI21x1_ASAP7_75t_L g628 ( .A1(n_570), .A2(n_83), .B(n_81), .Y(n_628) );
INVx1_ASAP7_75t_L g629 ( .A(n_573), .Y(n_629) );
INVx1_ASAP7_75t_L g630 ( .A(n_565), .Y(n_630) );
INVx2_ASAP7_75t_L g631 ( .A(n_586), .Y(n_631) );
INVx1_ASAP7_75t_L g632 ( .A(n_586), .Y(n_632) );
AND2x2_ASAP7_75t_L g633 ( .A(n_566), .B(n_561), .Y(n_633) );
INVx2_ASAP7_75t_L g634 ( .A(n_585), .Y(n_634) );
INVx1_ASAP7_75t_L g635 ( .A(n_566), .Y(n_635) );
INVx1_ASAP7_75t_L g636 ( .A(n_568), .Y(n_636) );
INVx1_ASAP7_75t_L g637 ( .A(n_560), .Y(n_637) );
BUFx2_ASAP7_75t_SL g638 ( .A(n_576), .Y(n_638) );
INVx1_ASAP7_75t_L g639 ( .A(n_567), .Y(n_639) );
INVx2_ASAP7_75t_L g640 ( .A(n_570), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_578), .Y(n_641) );
HB1xp67_ASAP7_75t_SL g642 ( .A(n_591), .Y(n_642) );
INVxp67_ASAP7_75t_L g643 ( .A(n_557), .Y(n_643) );
INVx2_ASAP7_75t_L g644 ( .A(n_564), .Y(n_644) );
OAI21x1_ASAP7_75t_L g645 ( .A1(n_551), .A2(n_86), .B(n_85), .Y(n_645) );
INVx1_ASAP7_75t_L g646 ( .A(n_563), .Y(n_646) );
INVx1_ASAP7_75t_L g647 ( .A(n_601), .Y(n_647) );
INVx1_ASAP7_75t_L g648 ( .A(n_588), .Y(n_648) );
INVx1_ASAP7_75t_L g649 ( .A(n_589), .Y(n_649) );
INVx2_ASAP7_75t_L g650 ( .A(n_594), .Y(n_650) );
INVx1_ASAP7_75t_SL g651 ( .A(n_556), .Y(n_651) );
INVx2_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
INVx3_ASAP7_75t_L g653 ( .A(n_599), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_602), .Y(n_654) );
INVx3_ASAP7_75t_L g655 ( .A(n_598), .Y(n_655) );
INVx2_ASAP7_75t_L g656 ( .A(n_577), .Y(n_656) );
INVx1_ASAP7_75t_L g657 ( .A(n_577), .Y(n_657) );
BUFx6f_ASAP7_75t_L g658 ( .A(n_553), .Y(n_658) );
INVx3_ASAP7_75t_L g659 ( .A(n_562), .Y(n_659) );
INVx1_ASAP7_75t_SL g660 ( .A(n_571), .Y(n_660) );
INVx2_ASAP7_75t_SL g661 ( .A(n_556), .Y(n_661) );
INVx1_ASAP7_75t_L g662 ( .A(n_558), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_596), .Y(n_663) );
INVx3_ASAP7_75t_L g664 ( .A(n_555), .Y(n_664) );
OA21x2_ASAP7_75t_L g665 ( .A1(n_582), .A2(n_92), .B(n_91), .Y(n_665) );
INVx2_ASAP7_75t_L g666 ( .A(n_596), .Y(n_666) );
INVx1_ASAP7_75t_L g667 ( .A(n_558), .Y(n_667) );
INVxp67_ASAP7_75t_L g668 ( .A(n_558), .Y(n_668) );
INVx2_ASAP7_75t_SL g669 ( .A(n_556), .Y(n_669) );
INVx1_ASAP7_75t_L g670 ( .A(n_596), .Y(n_670) );
HB1xp67_ASAP7_75t_L g671 ( .A(n_558), .Y(n_671) );
AND2x4_ASAP7_75t_L g672 ( .A(n_596), .B(n_15), .Y(n_672) );
INVx1_ASAP7_75t_SL g673 ( .A(n_555), .Y(n_673) );
INVx1_ASAP7_75t_L g674 ( .A(n_558), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_558), .Y(n_675) );
INVx1_ASAP7_75t_L g676 ( .A(n_558), .Y(n_676) );
NAND2x1p5_ASAP7_75t_L g677 ( .A(n_555), .B(n_93), .Y(n_677) );
INVx1_ASAP7_75t_L g678 ( .A(n_558), .Y(n_678) );
INVx1_ASAP7_75t_L g679 ( .A(n_558), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_596), .Y(n_680) );
INVx2_ASAP7_75t_L g681 ( .A(n_596), .Y(n_681) );
INVxp67_ASAP7_75t_SL g682 ( .A(n_558), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g683 ( .A(n_575), .B(n_94), .Y(n_683) );
OAI22xp5_ASAP7_75t_L g684 ( .A1(n_587), .A2(n_95), .B1(n_96), .B2(n_97), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_558), .Y(n_685) );
INVx3_ASAP7_75t_L g686 ( .A(n_664), .Y(n_686) );
INVx2_ASAP7_75t_L g687 ( .A(n_607), .Y(n_687) );
AND2x2_ASAP7_75t_L g688 ( .A(n_611), .B(n_98), .Y(n_688) );
BUFx3_ASAP7_75t_L g689 ( .A(n_613), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g690 ( .A(n_630), .B(n_289), .Y(n_690) );
INVx2_ASAP7_75t_L g691 ( .A(n_608), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_627), .Y(n_692) );
AND2x2_ASAP7_75t_L g693 ( .A(n_671), .B(n_99), .Y(n_693) );
INVx1_ASAP7_75t_L g694 ( .A(n_627), .Y(n_694) );
AOI22xp33_ASAP7_75t_SL g695 ( .A1(n_626), .A2(n_103), .B1(n_104), .B2(n_106), .Y(n_695) );
INVx1_ASAP7_75t_L g696 ( .A(n_670), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_663), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_670), .Y(n_698) );
INVx1_ASAP7_75t_L g699 ( .A(n_680), .Y(n_699) );
INVx2_ASAP7_75t_L g700 ( .A(n_666), .Y(n_700) );
INVx2_ASAP7_75t_L g701 ( .A(n_681), .Y(n_701) );
AND2x2_ASAP7_75t_L g702 ( .A(n_603), .B(n_109), .Y(n_702) );
INVx1_ASAP7_75t_L g703 ( .A(n_680), .Y(n_703) );
INVx1_ASAP7_75t_L g704 ( .A(n_662), .Y(n_704) );
INVx2_ASAP7_75t_SL g705 ( .A(n_616), .Y(n_705) );
AND2x2_ASAP7_75t_L g706 ( .A(n_682), .B(n_113), .Y(n_706) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_668), .Y(n_707) );
INVx2_ASAP7_75t_L g708 ( .A(n_609), .Y(n_708) );
INVx1_ASAP7_75t_L g709 ( .A(n_667), .Y(n_709) );
OR2x2_ASAP7_75t_L g710 ( .A(n_674), .B(n_114), .Y(n_710) );
NAND2xp5_ASAP7_75t_L g711 ( .A(n_620), .B(n_288), .Y(n_711) );
INVx2_ASAP7_75t_L g712 ( .A(n_619), .Y(n_712) );
INVx1_ASAP7_75t_L g713 ( .A(n_632), .Y(n_713) );
AND2x2_ASAP7_75t_L g714 ( .A(n_673), .B(n_115), .Y(n_714) );
INVx2_ASAP7_75t_SL g715 ( .A(n_610), .Y(n_715) );
INVx2_ASAP7_75t_L g716 ( .A(n_614), .Y(n_716) );
INVx1_ASAP7_75t_L g717 ( .A(n_675), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_676), .Y(n_718) );
INVx2_ASAP7_75t_L g719 ( .A(n_618), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g720 ( .A(n_624), .B(n_287), .Y(n_720) );
INVx1_ASAP7_75t_L g721 ( .A(n_678), .Y(n_721) );
HB1xp67_ASAP7_75t_L g722 ( .A(n_679), .Y(n_722) );
AND2x4_ASAP7_75t_SL g723 ( .A(n_661), .B(n_116), .Y(n_723) );
INVx2_ASAP7_75t_L g724 ( .A(n_634), .Y(n_724) );
INVx1_ASAP7_75t_L g725 ( .A(n_685), .Y(n_725) );
INVx1_ASAP7_75t_L g726 ( .A(n_672), .Y(n_726) );
BUFx3_ASAP7_75t_L g727 ( .A(n_669), .Y(n_727) );
INVx1_ASAP7_75t_L g728 ( .A(n_672), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_604), .Y(n_729) );
AND2x2_ASAP7_75t_L g730 ( .A(n_633), .B(n_117), .Y(n_730) );
AO31x2_ASAP7_75t_L g731 ( .A1(n_639), .A2(n_118), .A3(n_119), .B(n_122), .Y(n_731) );
AND2x2_ASAP7_75t_L g732 ( .A(n_664), .B(n_126), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_646), .B(n_128), .Y(n_733) );
INVx4_ASAP7_75t_R g734 ( .A(n_642), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_631), .Y(n_735) );
BUFx6f_ASAP7_75t_L g736 ( .A(n_658), .Y(n_736) );
INVx1_ASAP7_75t_L g737 ( .A(n_640), .Y(n_737) );
AND2x2_ASAP7_75t_L g738 ( .A(n_615), .B(n_129), .Y(n_738) );
BUFx3_ASAP7_75t_L g739 ( .A(n_651), .Y(n_739) );
OA21x2_ASAP7_75t_L g740 ( .A1(n_657), .A2(n_130), .B(n_131), .Y(n_740) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_629), .B(n_132), .Y(n_741) );
INVx2_ASAP7_75t_SL g742 ( .A(n_637), .Y(n_742) );
AND2x2_ASAP7_75t_L g743 ( .A(n_622), .B(n_133), .Y(n_743) );
AND2x2_ASAP7_75t_L g744 ( .A(n_612), .B(n_134), .Y(n_744) );
INVxp67_ASAP7_75t_SL g745 ( .A(n_617), .Y(n_745) );
INVxp67_ASAP7_75t_SL g746 ( .A(n_636), .Y(n_746) );
INVx1_ASAP7_75t_L g747 ( .A(n_605), .Y(n_747) );
HB1xp67_ASAP7_75t_L g748 ( .A(n_635), .Y(n_748) );
AND2x4_ASAP7_75t_L g749 ( .A(n_658), .B(n_135), .Y(n_749) );
AND2x2_ASAP7_75t_L g750 ( .A(n_626), .B(n_137), .Y(n_750) );
AND2x2_ASAP7_75t_L g751 ( .A(n_623), .B(n_138), .Y(n_751) );
INVx1_ASAP7_75t_L g752 ( .A(n_606), .Y(n_752) );
INVx2_ASAP7_75t_L g753 ( .A(n_677), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_659), .B(n_643), .Y(n_754) );
AND2x2_ASAP7_75t_L g755 ( .A(n_659), .B(n_139), .Y(n_755) );
INVx2_ASAP7_75t_L g756 ( .A(n_628), .Y(n_756) );
INVx5_ASAP7_75t_L g757 ( .A(n_658), .Y(n_757) );
INVx2_ASAP7_75t_L g758 ( .A(n_638), .Y(n_758) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_649), .Y(n_759) );
INVx1_ASAP7_75t_L g760 ( .A(n_638), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_621), .Y(n_761) );
BUFx3_ASAP7_75t_L g762 ( .A(n_683), .Y(n_762) );
OR2x2_ASAP7_75t_L g763 ( .A(n_684), .B(n_286), .Y(n_763) );
INVx1_ASAP7_75t_L g764 ( .A(n_649), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g765 ( .A(n_641), .B(n_140), .Y(n_765) );
INVxp67_ASAP7_75t_SL g766 ( .A(n_656), .Y(n_766) );
INVx6_ASAP7_75t_L g767 ( .A(n_625), .Y(n_767) );
AND2x2_ASAP7_75t_L g768 ( .A(n_665), .B(n_142), .Y(n_768) );
NAND2xp5_ASAP7_75t_L g769 ( .A(n_660), .B(n_143), .Y(n_769) );
BUFx2_ASAP7_75t_L g770 ( .A(n_665), .Y(n_770) );
NAND2xp5_ASAP7_75t_L g771 ( .A(n_647), .B(n_284), .Y(n_771) );
HB1xp67_ASAP7_75t_L g772 ( .A(n_648), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_654), .B(n_144), .Y(n_773) );
OR2x2_ASAP7_75t_L g774 ( .A(n_655), .B(n_283), .Y(n_774) );
AND2x2_ASAP7_75t_L g775 ( .A(n_645), .B(n_146), .Y(n_775) );
INVx3_ASAP7_75t_L g776 ( .A(n_653), .Y(n_776) );
AND2x4_ASAP7_75t_SL g777 ( .A(n_653), .B(n_147), .Y(n_777) );
AND2x2_ASAP7_75t_L g778 ( .A(n_655), .B(n_149), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_644), .Y(n_779) );
INVx2_ASAP7_75t_L g780 ( .A(n_650), .Y(n_780) );
OR2x2_ASAP7_75t_L g781 ( .A(n_652), .B(n_282), .Y(n_781) );
INVx1_ASAP7_75t_L g782 ( .A(n_670), .Y(n_782) );
INVx2_ASAP7_75t_L g783 ( .A(n_607), .Y(n_783) );
INVx1_ASAP7_75t_L g784 ( .A(n_627), .Y(n_784) );
BUFx2_ASAP7_75t_L g785 ( .A(n_613), .Y(n_785) );
INVxp67_ASAP7_75t_SL g786 ( .A(n_682), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_607), .Y(n_787) );
INVx1_ASAP7_75t_L g788 ( .A(n_670), .Y(n_788) );
INVx3_ASAP7_75t_L g789 ( .A(n_664), .Y(n_789) );
INVx2_ASAP7_75t_L g790 ( .A(n_607), .Y(n_790) );
INVx1_ASAP7_75t_L g791 ( .A(n_722), .Y(n_791) );
INVx1_ASAP7_75t_L g792 ( .A(n_704), .Y(n_792) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_786), .B(n_150), .Y(n_793) );
NOR2xp33_ASAP7_75t_L g794 ( .A(n_727), .B(n_152), .Y(n_794) );
INVx3_ASAP7_75t_L g795 ( .A(n_758), .Y(n_795) );
INVx2_ASAP7_75t_L g796 ( .A(n_687), .Y(n_796) );
NAND2xp5_ASAP7_75t_L g797 ( .A(n_709), .B(n_153), .Y(n_797) );
AND2x2_ASAP7_75t_L g798 ( .A(n_717), .B(n_154), .Y(n_798) );
INVxp67_ASAP7_75t_L g799 ( .A(n_785), .Y(n_799) );
NAND2xp5_ASAP7_75t_L g800 ( .A(n_718), .B(n_155), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_721), .Y(n_801) );
NOR2x1_ASAP7_75t_L g802 ( .A(n_689), .B(n_157), .Y(n_802) );
AND2x2_ASAP7_75t_L g803 ( .A(n_725), .B(n_748), .Y(n_803) );
OR2x2_ASAP7_75t_L g804 ( .A(n_707), .B(n_158), .Y(n_804) );
INVx2_ASAP7_75t_L g805 ( .A(n_691), .Y(n_805) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_716), .B(n_160), .Y(n_806) );
INVxp67_ASAP7_75t_L g807 ( .A(n_705), .Y(n_807) );
OR2x2_ASAP7_75t_L g808 ( .A(n_719), .B(n_162), .Y(n_808) );
INVx4_ASAP7_75t_L g809 ( .A(n_757), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_729), .B(n_164), .Y(n_810) );
INVx2_ASAP7_75t_L g811 ( .A(n_790), .Y(n_811) );
INVx1_ASAP7_75t_L g812 ( .A(n_696), .Y(n_812) );
NAND2xp5_ASAP7_75t_L g813 ( .A(n_698), .B(n_165), .Y(n_813) );
AOI22xp5_ASAP7_75t_L g814 ( .A1(n_745), .A2(n_166), .B1(n_167), .B2(n_168), .Y(n_814) );
AND2x2_ASAP7_75t_L g815 ( .A(n_754), .B(n_169), .Y(n_815) );
INVx2_ASAP7_75t_L g816 ( .A(n_697), .Y(n_816) );
NOR2xp33_ASAP7_75t_L g817 ( .A(n_739), .B(n_171), .Y(n_817) );
INVx3_ASAP7_75t_L g818 ( .A(n_686), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_699), .Y(n_819) );
AND2x2_ASAP7_75t_L g820 ( .A(n_708), .B(n_173), .Y(n_820) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_715), .Y(n_821) );
OR2x2_ASAP7_75t_L g822 ( .A(n_700), .B(n_174), .Y(n_822) );
AND2x2_ASAP7_75t_L g823 ( .A(n_712), .B(n_175), .Y(n_823) );
AND2x2_ASAP7_75t_L g824 ( .A(n_701), .B(n_177), .Y(n_824) );
AND2x4_ASAP7_75t_SL g825 ( .A(n_760), .B(n_178), .Y(n_825) );
INVx1_ASAP7_75t_L g826 ( .A(n_703), .Y(n_826) );
AND2x2_ASAP7_75t_L g827 ( .A(n_783), .B(n_179), .Y(n_827) );
INVx1_ASAP7_75t_L g828 ( .A(n_692), .Y(n_828) );
INVx1_ASAP7_75t_SL g829 ( .A(n_723), .Y(n_829) );
AND2x2_ASAP7_75t_L g830 ( .A(n_787), .B(n_181), .Y(n_830) );
INVxp67_ASAP7_75t_SL g831 ( .A(n_759), .Y(n_831) );
INVx2_ASAP7_75t_L g832 ( .A(n_724), .Y(n_832) );
OR2x2_ASAP7_75t_L g833 ( .A(n_782), .B(n_182), .Y(n_833) );
INVx1_ASAP7_75t_L g834 ( .A(n_788), .Y(n_834) );
AND2x2_ASAP7_75t_L g835 ( .A(n_746), .B(n_183), .Y(n_835) );
AND2x2_ASAP7_75t_L g836 ( .A(n_726), .B(n_184), .Y(n_836) );
OR2x2_ASAP7_75t_L g837 ( .A(n_735), .B(n_185), .Y(n_837) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_713), .B(n_187), .Y(n_838) );
INVx1_ASAP7_75t_L g839 ( .A(n_692), .Y(n_839) );
INVxp67_ASAP7_75t_L g840 ( .A(n_742), .Y(n_840) );
INVx1_ASAP7_75t_L g841 ( .A(n_694), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_713), .B(n_188), .Y(n_842) );
NAND2xp5_ASAP7_75t_L g843 ( .A(n_694), .B(n_189), .Y(n_843) );
INVx3_ASAP7_75t_L g844 ( .A(n_686), .Y(n_844) );
INVx2_ASAP7_75t_L g845 ( .A(n_784), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_784), .Y(n_846) );
AND2x2_ASAP7_75t_L g847 ( .A(n_728), .B(n_190), .Y(n_847) );
AND2x2_ASAP7_75t_L g848 ( .A(n_789), .B(n_195), .Y(n_848) );
INVx2_ASAP7_75t_L g849 ( .A(n_737), .Y(n_849) );
AND2x2_ASAP7_75t_L g850 ( .A(n_789), .B(n_197), .Y(n_850) );
AND2x4_ASAP7_75t_SL g851 ( .A(n_734), .B(n_198), .Y(n_851) );
INVx3_ASAP7_75t_L g852 ( .A(n_757), .Y(n_852) );
OR2x2_ASAP7_75t_L g853 ( .A(n_737), .B(n_199), .Y(n_853) );
INVx1_ASAP7_75t_L g854 ( .A(n_764), .Y(n_854) );
AND2x2_ASAP7_75t_L g855 ( .A(n_706), .B(n_201), .Y(n_855) );
INVx1_ASAP7_75t_L g856 ( .A(n_764), .Y(n_856) );
BUFx2_ASAP7_75t_L g857 ( .A(n_757), .Y(n_857) );
INVx1_ASAP7_75t_L g858 ( .A(n_772), .Y(n_858) );
OR2x2_ASAP7_75t_L g859 ( .A(n_710), .B(n_202), .Y(n_859) );
INVx1_ASAP7_75t_L g860 ( .A(n_747), .Y(n_860) );
AND2x2_ASAP7_75t_L g861 ( .A(n_693), .B(n_207), .Y(n_861) );
AND2x2_ASAP7_75t_L g862 ( .A(n_730), .B(n_208), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_747), .Y(n_863) );
NOR2xp33_ASAP7_75t_L g864 ( .A(n_762), .B(n_210), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_779), .Y(n_865) );
AND2x2_ASAP7_75t_L g866 ( .A(n_688), .B(n_211), .Y(n_866) );
AND2x2_ASAP7_75t_L g867 ( .A(n_752), .B(n_212), .Y(n_867) );
OR2x2_ASAP7_75t_L g868 ( .A(n_773), .B(n_213), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_766), .Y(n_869) );
AND2x2_ASAP7_75t_L g870 ( .A(n_702), .B(n_215), .Y(n_870) );
NAND2xp5_ASAP7_75t_L g871 ( .A(n_791), .B(n_761), .Y(n_871) );
AND2x2_ASAP7_75t_L g872 ( .A(n_803), .B(n_755), .Y(n_872) );
INVx1_ASAP7_75t_L g873 ( .A(n_828), .Y(n_873) );
INVx2_ASAP7_75t_L g874 ( .A(n_869), .Y(n_874) );
INVx2_ASAP7_75t_L g875 ( .A(n_869), .Y(n_875) );
INVx1_ASAP7_75t_L g876 ( .A(n_792), .Y(n_876) );
AND2x2_ASAP7_75t_L g877 ( .A(n_799), .B(n_776), .Y(n_877) );
INVx2_ASAP7_75t_L g878 ( .A(n_849), .Y(n_878) );
NAND5xp2_ASAP7_75t_L g879 ( .A(n_864), .B(n_695), .C(n_690), .D(n_750), .E(n_744), .Y(n_879) );
AND2x2_ASAP7_75t_L g880 ( .A(n_807), .B(n_776), .Y(n_880) );
OR2x2_ASAP7_75t_L g881 ( .A(n_858), .B(n_780), .Y(n_881) );
INVx1_ASAP7_75t_L g882 ( .A(n_828), .Y(n_882) );
OR2x2_ASAP7_75t_L g883 ( .A(n_832), .B(n_774), .Y(n_883) );
NAND2xp5_ASAP7_75t_L g884 ( .A(n_801), .B(n_733), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g885 ( .A(n_812), .B(n_819), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_796), .Y(n_886) );
INVxp67_ASAP7_75t_SL g887 ( .A(n_831), .Y(n_887) );
OR2x2_ASAP7_75t_L g888 ( .A(n_805), .B(n_781), .Y(n_888) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_826), .B(n_753), .Y(n_889) );
OR2x2_ASAP7_75t_L g890 ( .A(n_811), .B(n_736), .Y(n_890) );
INVxp67_ASAP7_75t_SL g891 ( .A(n_795), .Y(n_891) );
OR2x2_ASAP7_75t_L g892 ( .A(n_816), .B(n_736), .Y(n_892) );
INVx1_ASAP7_75t_L g893 ( .A(n_839), .Y(n_893) );
AND2x2_ASAP7_75t_L g894 ( .A(n_795), .B(n_778), .Y(n_894) );
INVx2_ASAP7_75t_L g895 ( .A(n_845), .Y(n_895) );
OR2x2_ASAP7_75t_L g896 ( .A(n_834), .B(n_736), .Y(n_896) );
INVx1_ASAP7_75t_L g897 ( .A(n_841), .Y(n_897) );
NAND2xp5_ASAP7_75t_L g898 ( .A(n_846), .B(n_741), .Y(n_898) );
INVx1_ASAP7_75t_L g899 ( .A(n_854), .Y(n_899) );
OR2x2_ASAP7_75t_L g900 ( .A(n_865), .B(n_770), .Y(n_900) );
INVxp67_ASAP7_75t_L g901 ( .A(n_840), .Y(n_901) );
AND2x2_ASAP7_75t_L g902 ( .A(n_818), .B(n_751), .Y(n_902) );
OR2x2_ASAP7_75t_L g903 ( .A(n_865), .B(n_769), .Y(n_903) );
INVx1_ASAP7_75t_L g904 ( .A(n_856), .Y(n_904) );
INVx2_ASAP7_75t_L g905 ( .A(n_860), .Y(n_905) );
INVx1_ASAP7_75t_L g906 ( .A(n_863), .Y(n_906) );
INVxp67_ASAP7_75t_SL g907 ( .A(n_818), .Y(n_907) );
AND2x4_ASAP7_75t_L g908 ( .A(n_844), .B(n_749), .Y(n_908) );
AND2x2_ASAP7_75t_L g909 ( .A(n_844), .B(n_714), .Y(n_909) );
NOR2xp33_ASAP7_75t_L g910 ( .A(n_829), .B(n_738), .Y(n_910) );
INVx1_ASAP7_75t_L g911 ( .A(n_804), .Y(n_911) );
NAND2xp5_ASAP7_75t_L g912 ( .A(n_815), .B(n_720), .Y(n_912) );
AND2x2_ASAP7_75t_L g913 ( .A(n_857), .B(n_777), .Y(n_913) );
OR2x2_ASAP7_75t_L g914 ( .A(n_853), .B(n_711), .Y(n_914) );
INVx2_ASAP7_75t_L g915 ( .A(n_852), .Y(n_915) );
INVx1_ASAP7_75t_L g916 ( .A(n_843), .Y(n_916) );
INVx1_ASAP7_75t_L g917 ( .A(n_838), .Y(n_917) );
AND2x4_ASAP7_75t_L g918 ( .A(n_852), .B(n_749), .Y(n_918) );
INVx2_ASAP7_75t_L g919 ( .A(n_809), .Y(n_919) );
INVx2_ASAP7_75t_L g920 ( .A(n_874), .Y(n_920) );
NAND2xp5_ASAP7_75t_L g921 ( .A(n_887), .B(n_867), .Y(n_921) );
HB1xp67_ASAP7_75t_L g922 ( .A(n_891), .Y(n_922) );
AND2x2_ASAP7_75t_L g923 ( .A(n_880), .B(n_872), .Y(n_923) );
INVx1_ASAP7_75t_L g924 ( .A(n_876), .Y(n_924) );
AND2x2_ASAP7_75t_L g925 ( .A(n_877), .B(n_821), .Y(n_925) );
NAND2xp5_ASAP7_75t_L g926 ( .A(n_871), .B(n_798), .Y(n_926) );
OR2x2_ASAP7_75t_L g927 ( .A(n_881), .B(n_886), .Y(n_927) );
INVx1_ASAP7_75t_L g928 ( .A(n_885), .Y(n_928) );
INVx1_ASAP7_75t_L g929 ( .A(n_906), .Y(n_929) );
BUFx2_ASAP7_75t_L g930 ( .A(n_919), .Y(n_930) );
INVx2_ASAP7_75t_L g931 ( .A(n_875), .Y(n_931) );
BUFx2_ASAP7_75t_L g932 ( .A(n_915), .Y(n_932) );
INVx2_ASAP7_75t_L g933 ( .A(n_905), .Y(n_933) );
NAND2xp5_ASAP7_75t_L g934 ( .A(n_873), .B(n_835), .Y(n_934) );
NAND2xp5_ASAP7_75t_L g935 ( .A(n_873), .B(n_793), .Y(n_935) );
NAND2xp5_ASAP7_75t_L g936 ( .A(n_893), .B(n_842), .Y(n_936) );
INVx1_ASAP7_75t_L g937 ( .A(n_882), .Y(n_937) );
INVxp67_ASAP7_75t_L g938 ( .A(n_910), .Y(n_938) );
INVx1_ASAP7_75t_L g939 ( .A(n_882), .Y(n_939) );
INVx1_ASAP7_75t_L g940 ( .A(n_897), .Y(n_940) );
INVx2_ASAP7_75t_L g941 ( .A(n_878), .Y(n_941) );
AND2x2_ASAP7_75t_L g942 ( .A(n_901), .B(n_809), .Y(n_942) );
INVxp67_ASAP7_75t_SL g943 ( .A(n_907), .Y(n_943) );
OR2x2_ASAP7_75t_L g944 ( .A(n_900), .B(n_808), .Y(n_944) );
OAI21xp33_ASAP7_75t_L g945 ( .A1(n_879), .A2(n_851), .B(n_802), .Y(n_945) );
AND2x4_ASAP7_75t_L g946 ( .A(n_908), .B(n_825), .Y(n_946) );
AND2x2_ASAP7_75t_L g947 ( .A(n_894), .B(n_848), .Y(n_947) );
AND2x2_ASAP7_75t_L g948 ( .A(n_909), .B(n_902), .Y(n_948) );
AND2x2_ASAP7_75t_L g949 ( .A(n_913), .B(n_850), .Y(n_949) );
INVx2_ASAP7_75t_L g950 ( .A(n_922), .Y(n_950) );
AOI32xp33_ASAP7_75t_L g951 ( .A1(n_945), .A2(n_918), .A3(n_911), .B1(n_817), .B2(n_908), .Y(n_951) );
NOR2xp33_ASAP7_75t_L g952 ( .A(n_938), .B(n_889), .Y(n_952) );
INVx1_ASAP7_75t_L g953 ( .A(n_924), .Y(n_953) );
INVx1_ASAP7_75t_L g954 ( .A(n_929), .Y(n_954) );
INVx2_ASAP7_75t_SL g955 ( .A(n_927), .Y(n_955) );
CKINVDCx16_ASAP7_75t_R g956 ( .A(n_925), .Y(n_956) );
INVxp67_ASAP7_75t_L g957 ( .A(n_930), .Y(n_957) );
NOR2xp67_ASAP7_75t_L g958 ( .A(n_945), .B(n_918), .Y(n_958) );
NAND2xp5_ASAP7_75t_L g959 ( .A(n_928), .B(n_899), .Y(n_959) );
INVx1_ASAP7_75t_SL g960 ( .A(n_932), .Y(n_960) );
INVx1_ASAP7_75t_L g961 ( .A(n_940), .Y(n_961) );
NAND2xp5_ASAP7_75t_L g962 ( .A(n_935), .B(n_904), .Y(n_962) );
AOI22xp5_ASAP7_75t_L g963 ( .A1(n_921), .A2(n_917), .B1(n_916), .B2(n_912), .Y(n_963) );
INVx1_ASAP7_75t_L g964 ( .A(n_937), .Y(n_964) );
OAI31xp33_ASAP7_75t_L g965 ( .A1(n_946), .A2(n_794), .A3(n_859), .B(n_870), .Y(n_965) );
INVxp67_ASAP7_75t_L g966 ( .A(n_942), .Y(n_966) );
INVx1_ASAP7_75t_L g967 ( .A(n_939), .Y(n_967) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_935), .B(n_917), .Y(n_968) );
INVx1_ASAP7_75t_L g969 ( .A(n_933), .Y(n_969) );
OAI22xp33_ASAP7_75t_L g970 ( .A1(n_958), .A2(n_943), .B1(n_921), .B2(n_944), .Y(n_970) );
O2A1O1Ixp33_ASAP7_75t_SL g971 ( .A1(n_957), .A2(n_926), .B(n_934), .C(n_868), .Y(n_971) );
AOI31xp33_ASAP7_75t_L g972 ( .A1(n_960), .A2(n_946), .A3(n_949), .B(n_866), .Y(n_972) );
OAI221xp5_ASAP7_75t_L g973 ( .A1(n_951), .A2(n_934), .B1(n_936), .B2(n_916), .C(n_884), .Y(n_973) );
NOR2xp33_ASAP7_75t_L g974 ( .A(n_956), .B(n_923), .Y(n_974) );
AOI22xp5_ASAP7_75t_L g975 ( .A1(n_966), .A2(n_947), .B1(n_948), .B2(n_941), .Y(n_975) );
INVxp67_ASAP7_75t_L g976 ( .A(n_968), .Y(n_976) );
INVx1_ASAP7_75t_L g977 ( .A(n_964), .Y(n_977) );
OR2x2_ASAP7_75t_L g978 ( .A(n_955), .B(n_920), .Y(n_978) );
INVx1_ASAP7_75t_L g979 ( .A(n_967), .Y(n_979) );
OAI22xp5_ASAP7_75t_L g980 ( .A1(n_963), .A2(n_931), .B1(n_896), .B2(n_903), .Y(n_980) );
OAI321xp33_ASAP7_75t_L g981 ( .A1(n_950), .A2(n_814), .A3(n_898), .B1(n_892), .B2(n_890), .C(n_883), .Y(n_981) );
INVxp67_ASAP7_75t_SL g982 ( .A(n_969), .Y(n_982) );
NOR4xp25_ASAP7_75t_L g983 ( .A(n_973), .B(n_952), .C(n_959), .D(n_961), .Y(n_983) );
OAI221xp5_ASAP7_75t_L g984 ( .A1(n_972), .A2(n_965), .B1(n_962), .B2(n_954), .C(n_953), .Y(n_984) );
NAND2xp5_ASAP7_75t_L g985 ( .A(n_976), .B(n_965), .Y(n_985) );
AOI22xp5_ASAP7_75t_L g986 ( .A1(n_970), .A2(n_855), .B1(n_862), .B2(n_861), .Y(n_986) );
OAI21xp5_ASAP7_75t_SL g987 ( .A1(n_974), .A2(n_914), .B(n_836), .Y(n_987) );
BUFx3_ASAP7_75t_L g988 ( .A(n_978), .Y(n_988) );
AOI21xp5_ASAP7_75t_L g989 ( .A1(n_971), .A2(n_810), .B(n_895), .Y(n_989) );
O2A1O1Ixp33_ASAP7_75t_SL g990 ( .A1(n_982), .A2(n_833), .B(n_763), .C(n_797), .Y(n_990) );
AOI221xp5_ASAP7_75t_L g991 ( .A1(n_980), .A2(n_800), .B1(n_847), .B2(n_743), .C(n_813), .Y(n_991) );
NOR2xp33_ASAP7_75t_L g992 ( .A(n_984), .B(n_977), .Y(n_992) );
AND2x2_ASAP7_75t_L g993 ( .A(n_988), .B(n_975), .Y(n_993) );
NAND2xp5_ASAP7_75t_L g994 ( .A(n_983), .B(n_979), .Y(n_994) );
INVx1_ASAP7_75t_SL g995 ( .A(n_985), .Y(n_995) );
NAND2xp5_ASAP7_75t_L g996 ( .A(n_987), .B(n_888), .Y(n_996) );
INVx1_ASAP7_75t_L g997 ( .A(n_986), .Y(n_997) );
NOR2xp33_ASAP7_75t_SL g998 ( .A(n_995), .B(n_993), .Y(n_998) );
NOR3xp33_ASAP7_75t_L g999 ( .A(n_994), .B(n_981), .C(n_990), .Y(n_999) );
NOR3xp33_ASAP7_75t_L g1000 ( .A(n_992), .B(n_997), .C(n_996), .Y(n_1000) );
A2O1A1Ixp33_ASAP7_75t_L g1001 ( .A1(n_992), .A2(n_989), .B(n_991), .C(n_768), .Y(n_1001) );
AOI22xp5_ASAP7_75t_L g1002 ( .A1(n_995), .A2(n_732), .B1(n_775), .B2(n_806), .Y(n_1002) );
NAND2xp5_ASAP7_75t_L g1003 ( .A(n_1000), .B(n_824), .Y(n_1003) );
INVx1_ASAP7_75t_L g1004 ( .A(n_1002), .Y(n_1004) );
NOR2x1_ASAP7_75t_L g1005 ( .A(n_1001), .B(n_740), .Y(n_1005) );
INVx1_ASAP7_75t_L g1006 ( .A(n_998), .Y(n_1006) );
OA21x2_ASAP7_75t_L g1007 ( .A1(n_1006), .A2(n_999), .B(n_765), .Y(n_1007) );
XNOR2x1_ASAP7_75t_L g1008 ( .A(n_1004), .B(n_837), .Y(n_1008) );
INVx1_ASAP7_75t_L g1009 ( .A(n_1003), .Y(n_1009) );
OAI22xp5_ASAP7_75t_L g1010 ( .A1(n_1007), .A2(n_1005), .B1(n_822), .B2(n_771), .Y(n_1010) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_1009), .B(n_827), .Y(n_1011) );
INVx2_ASAP7_75t_L g1012 ( .A(n_1008), .Y(n_1012) );
AOI22xp5_ASAP7_75t_L g1013 ( .A1(n_1012), .A2(n_830), .B1(n_823), .B2(n_820), .Y(n_1013) );
HB1xp67_ASAP7_75t_L g1014 ( .A(n_1011), .Y(n_1014) );
INVx1_ASAP7_75t_L g1015 ( .A(n_1010), .Y(n_1015) );
NAND2xp5_ASAP7_75t_L g1016 ( .A(n_1014), .B(n_731), .Y(n_1016) );
INVx1_ASAP7_75t_L g1017 ( .A(n_1015), .Y(n_1017) );
OAI22x1_ASAP7_75t_L g1018 ( .A1(n_1013), .A2(n_740), .B1(n_756), .B2(n_731), .Y(n_1018) );
HB1xp67_ASAP7_75t_L g1019 ( .A(n_1017), .Y(n_1019) );
NAND2xp5_ASAP7_75t_L g1020 ( .A(n_1016), .B(n_731), .Y(n_1020) );
OAI21xp5_ASAP7_75t_L g1021 ( .A1(n_1018), .A2(n_217), .B(n_218), .Y(n_1021) );
OAI21x1_ASAP7_75t_L g1022 ( .A1(n_1019), .A2(n_767), .B(n_221), .Y(n_1022) );
NAND2xp5_ASAP7_75t_L g1023 ( .A(n_1021), .B(n_220), .Y(n_1023) );
AOI221xp5_ASAP7_75t_SL g1024 ( .A1(n_1020), .A2(n_222), .B1(n_224), .B2(n_225), .C(n_227), .Y(n_1024) );
AO21x2_ASAP7_75t_L g1025 ( .A1(n_1023), .A2(n_1022), .B(n_1024), .Y(n_1025) );
OR2x2_ASAP7_75t_L g1026 ( .A(n_1025), .B(n_229), .Y(n_1026) );
AOI22xp33_ASAP7_75t_SL g1027 ( .A1(n_1026), .A2(n_235), .B1(n_236), .B2(n_238), .Y(n_1027) );
endmodule