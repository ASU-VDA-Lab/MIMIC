module fake_ariane_2054_n_1901 (n_83, n_8, n_56, n_60, n_170, n_160, n_64, n_179, n_180, n_119, n_124, n_167, n_90, n_38, n_47, n_110, n_153, n_18, n_86, n_75, n_89, n_67, n_176, n_149, n_34, n_158, n_172, n_69, n_95, n_175, n_92, n_143, n_183, n_150, n_98, n_74, n_113, n_114, n_33, n_19, n_40, n_181, n_152, n_120, n_169, n_106, n_12, n_53, n_173, n_111, n_21, n_115, n_133, n_66, n_71, n_24, n_7, n_109, n_96, n_156, n_49, n_20, n_174, n_100, n_17, n_50, n_132, n_62, n_147, n_51, n_166, n_76, n_103, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_91, n_159, n_107, n_72, n_105, n_128, n_44, n_30, n_82, n_178, n_31, n_42, n_57, n_131, n_70, n_10, n_117, n_139, n_165, n_85, n_130, n_144, n_6, n_48, n_94, n_101, n_4, n_134, n_185, n_2, n_32, n_37, n_58, n_65, n_123, n_9, n_138, n_112, n_45, n_162, n_11, n_129, n_126, n_137, n_122, n_148, n_164, n_52, n_157, n_184, n_177, n_135, n_73, n_77, n_171, n_15, n_118, n_93, n_121, n_23, n_61, n_108, n_102, n_182, n_125, n_22, n_168, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_140, n_55, n_151, n_136, n_28, n_80, n_146, n_97, n_154, n_142, n_161, n_14, n_163, n_88, n_141, n_68, n_116, n_104, n_145, n_78, n_39, n_59, n_63, n_99, n_16, n_5, n_155, n_127, n_35, n_54, n_25, n_1901);

input n_83;
input n_8;
input n_56;
input n_60;
input n_170;
input n_160;
input n_64;
input n_179;
input n_180;
input n_119;
input n_124;
input n_167;
input n_90;
input n_38;
input n_47;
input n_110;
input n_153;
input n_18;
input n_86;
input n_75;
input n_89;
input n_67;
input n_176;
input n_149;
input n_34;
input n_158;
input n_172;
input n_69;
input n_95;
input n_175;
input n_92;
input n_143;
input n_183;
input n_150;
input n_98;
input n_74;
input n_113;
input n_114;
input n_33;
input n_19;
input n_40;
input n_181;
input n_152;
input n_120;
input n_169;
input n_106;
input n_12;
input n_53;
input n_173;
input n_111;
input n_21;
input n_115;
input n_133;
input n_66;
input n_71;
input n_24;
input n_7;
input n_109;
input n_96;
input n_156;
input n_49;
input n_20;
input n_174;
input n_100;
input n_17;
input n_50;
input n_132;
input n_62;
input n_147;
input n_51;
input n_166;
input n_76;
input n_103;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_91;
input n_159;
input n_107;
input n_72;
input n_105;
input n_128;
input n_44;
input n_30;
input n_82;
input n_178;
input n_31;
input n_42;
input n_57;
input n_131;
input n_70;
input n_10;
input n_117;
input n_139;
input n_165;
input n_85;
input n_130;
input n_144;
input n_6;
input n_48;
input n_94;
input n_101;
input n_4;
input n_134;
input n_185;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_123;
input n_9;
input n_138;
input n_112;
input n_45;
input n_162;
input n_11;
input n_129;
input n_126;
input n_137;
input n_122;
input n_148;
input n_164;
input n_52;
input n_157;
input n_184;
input n_177;
input n_135;
input n_73;
input n_77;
input n_171;
input n_15;
input n_118;
input n_93;
input n_121;
input n_23;
input n_61;
input n_108;
input n_102;
input n_182;
input n_125;
input n_22;
input n_168;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_140;
input n_55;
input n_151;
input n_136;
input n_28;
input n_80;
input n_146;
input n_97;
input n_154;
input n_142;
input n_161;
input n_14;
input n_163;
input n_88;
input n_141;
input n_68;
input n_116;
input n_104;
input n_145;
input n_78;
input n_39;
input n_59;
input n_63;
input n_99;
input n_16;
input n_5;
input n_155;
input n_127;
input n_35;
input n_54;
input n_25;

output n_1901;

wire n_913;
wire n_1681;
wire n_1486;
wire n_1507;
wire n_589;
wire n_1174;
wire n_1469;
wire n_691;
wire n_1353;
wire n_1355;
wire n_423;
wire n_1383;
wire n_603;
wire n_373;
wire n_1250;
wire n_1169;
wire n_789;
wire n_850;
wire n_610;
wire n_245;
wire n_1713;
wire n_319;
wire n_1436;
wire n_690;
wire n_416;
wire n_1109;
wire n_1430;
wire n_525;
wire n_187;
wire n_1463;
wire n_1238;
wire n_1515;
wire n_817;
wire n_1837;
wire n_924;
wire n_781;
wire n_1566;
wire n_189;
wire n_717;
wire n_952;
wire n_864;
wire n_1096;
wire n_1379;
wire n_1706;
wire n_524;
wire n_634;
wire n_1214;
wire n_1839;
wire n_1246;
wire n_1138;
wire n_214;
wire n_1853;
wire n_764;
wire n_1503;
wire n_462;
wire n_1196;
wire n_1181;
wire n_410;
wire n_1187;
wire n_1131;
wire n_1225;
wire n_737;
wire n_1298;
wire n_1745;
wire n_1366;
wire n_232;
wire n_568;
wire n_1088;
wire n_1424;
wire n_766;
wire n_1835;
wire n_1457;
wire n_377;
wire n_1682;
wire n_1836;
wire n_520;
wire n_870;
wire n_1453;
wire n_279;
wire n_958;
wire n_945;
wire n_813;
wire n_419;
wire n_270;
wire n_338;
wire n_995;
wire n_285;
wire n_1184;
wire n_202;
wire n_1535;
wire n_500;
wire n_665;
wire n_754;
wire n_903;
wire n_871;
wire n_1073;
wire n_239;
wire n_402;
wire n_1277;
wire n_1746;
wire n_829;
wire n_1761;
wire n_1062;
wire n_339;
wire n_738;
wire n_1690;
wire n_672;
wire n_740;
wire n_1283;
wire n_1736;
wire n_1018;
wire n_259;
wire n_953;
wire n_1364;
wire n_1888;
wire n_1224;
wire n_1425;
wire n_625;
wire n_557;
wire n_1107;
wire n_1688;
wire n_989;
wire n_242;
wire n_645;
wire n_331;
wire n_559;
wire n_495;
wire n_267;
wire n_350;
wire n_381;
wire n_795;
wire n_721;
wire n_1084;
wire n_1718;
wire n_1276;
wire n_200;
wire n_1428;
wire n_1284;
wire n_1241;
wire n_821;
wire n_561;
wire n_770;
wire n_1514;
wire n_1528;
wire n_507;
wire n_486;
wire n_901;
wire n_569;
wire n_1145;
wire n_971;
wire n_787;
wire n_1650;
wire n_1519;
wire n_1195;
wire n_1522;
wire n_518;
wire n_1207;
wire n_222;
wire n_786;
wire n_1404;
wire n_868;
wire n_1847;
wire n_1542;
wire n_1314;
wire n_1512;
wire n_1539;
wire n_884;
wire n_1851;
wire n_1415;
wire n_1034;
wire n_1652;
wire n_1676;
wire n_1085;
wire n_277;
wire n_1636;
wire n_432;
wire n_293;
wire n_823;
wire n_1900;
wire n_620;
wire n_1074;
wire n_859;
wire n_1765;
wire n_1889;
wire n_587;
wire n_693;
wire n_863;
wire n_303;
wire n_1254;
wire n_929;
wire n_206;
wire n_352;
wire n_899;
wire n_1703;
wire n_611;
wire n_1295;
wire n_1850;
wire n_365;
wire n_238;
wire n_1013;
wire n_1495;
wire n_1637;
wire n_334;
wire n_192;
wire n_661;
wire n_1751;
wire n_300;
wire n_533;
wire n_438;
wire n_1560;
wire n_1654;
wire n_1548;
wire n_1811;
wire n_440;
wire n_273;
wire n_1396;
wire n_1230;
wire n_612;
wire n_333;
wire n_1840;
wire n_376;
wire n_512;
wire n_1597;
wire n_1771;
wire n_1544;
wire n_579;
wire n_844;
wire n_1012;
wire n_1267;
wire n_1354;
wire n_1790;
wire n_1213;
wire n_237;
wire n_780;
wire n_1021;
wire n_1443;
wire n_491;
wire n_1465;
wire n_1595;
wire n_1142;
wire n_1140;
wire n_705;
wire n_570;
wire n_260;
wire n_942;
wire n_1437;
wire n_1378;
wire n_461;
wire n_1121;
wire n_1416;
wire n_209;
wire n_490;
wire n_1461;
wire n_1391;
wire n_225;
wire n_1599;
wire n_1876;
wire n_1006;
wire n_1830;
wire n_575;
wire n_546;
wire n_503;
wire n_1112;
wire n_700;
wire n_1159;
wire n_772;
wire n_1216;
wire n_1245;
wire n_1669;
wire n_1675;
wire n_676;
wire n_1838;
wire n_1594;
wire n_680;
wire n_287;
wire n_1716;
wire n_302;
wire n_1872;
wire n_380;
wire n_1585;
wire n_1432;
wire n_249;
wire n_1108;
wire n_355;
wire n_212;
wire n_444;
wire n_851;
wire n_1590;
wire n_1351;
wire n_1274;
wire n_257;
wire n_652;
wire n_1819;
wire n_475;
wire n_947;
wire n_930;
wire n_1260;
wire n_1179;
wire n_468;
wire n_696;
wire n_1442;
wire n_482;
wire n_798;
wire n_577;
wire n_1833;
wire n_407;
wire n_1691;
wire n_916;
wire n_1386;
wire n_912;
wire n_1884;
wire n_460;
wire n_1555;
wire n_1842;
wire n_366;
wire n_762;
wire n_1253;
wire n_1468;
wire n_1661;
wire n_555;
wire n_804;
wire n_1656;
wire n_1382;
wire n_966;
wire n_992;
wire n_955;
wire n_1182;
wire n_794;
wire n_1692;
wire n_1562;
wire n_514;
wire n_418;
wire n_1376;
wire n_513;
wire n_288;
wire n_1292;
wire n_1178;
wire n_1435;
wire n_1750;
wire n_1026;
wire n_1506;
wire n_1610;
wire n_306;
wire n_203;
wire n_436;
wire n_324;
wire n_669;
wire n_931;
wire n_1491;
wire n_619;
wire n_437;
wire n_337;
wire n_274;
wire n_967;
wire n_1083;
wire n_1418;
wire n_746;
wire n_1357;
wire n_292;
wire n_1079;
wire n_1787;
wire n_1389;
wire n_615;
wire n_1139;
wire n_517;
wire n_1312;
wire n_1717;
wire n_1812;
wire n_824;
wire n_428;
wire n_892;
wire n_1880;
wire n_959;
wire n_1399;
wire n_1101;
wire n_1567;
wire n_1343;
wire n_563;
wire n_1855;
wire n_990;
wire n_1623;
wire n_867;
wire n_1226;
wire n_944;
wire n_749;
wire n_1780;
wire n_815;
wire n_542;
wire n_1340;
wire n_470;
wire n_1240;
wire n_1087;
wire n_632;
wire n_477;
wire n_650;
wire n_425;
wire n_1433;
wire n_1825;
wire n_1155;
wire n_1071;
wire n_712;
wire n_976;
wire n_909;
wire n_1392;
wire n_767;
wire n_1832;
wire n_1841;
wire n_1680;
wire n_964;
wire n_1627;
wire n_382;
wire n_489;
wire n_251;
wire n_974;
wire n_506;
wire n_1731;
wire n_799;
wire n_1147;
wire n_397;
wire n_471;
wire n_351;
wire n_965;
wire n_934;
wire n_1447;
wire n_1220;
wire n_356;
wire n_698;
wire n_1674;
wire n_307;
wire n_1209;
wire n_1020;
wire n_1563;
wire n_646;
wire n_1633;
wire n_404;
wire n_1058;
wire n_347;
wire n_1042;
wire n_1234;
wire n_479;
wire n_1578;
wire n_1455;
wire n_299;
wire n_836;
wire n_1279;
wire n_564;
wire n_205;
wire n_1029;
wire n_1247;
wire n_760;
wire n_522;
wire n_1568;
wire n_1483;
wire n_1363;
wire n_367;
wire n_1111;
wire n_970;
wire n_1689;
wire n_713;
wire n_1255;
wire n_1646;
wire n_598;
wire n_345;
wire n_1237;
wire n_927;
wire n_261;
wire n_1095;
wire n_1728;
wire n_370;
wire n_706;
wire n_286;
wire n_1401;
wire n_1419;
wire n_1531;
wire n_776;
wire n_424;
wire n_1651;
wire n_1387;
wire n_466;
wire n_1263;
wire n_346;
wire n_1817;
wire n_552;
wire n_348;
wire n_670;
wire n_1826;
wire n_379;
wire n_264;
wire n_441;
wire n_1032;
wire n_1217;
wire n_1496;
wire n_637;
wire n_1592;
wire n_327;
wire n_1259;
wire n_1177;
wire n_1231;
wire n_980;
wire n_1618;
wire n_1869;
wire n_1743;
wire n_905;
wire n_207;
wire n_720;
wire n_926;
wire n_194;
wire n_1802;
wire n_1163;
wire n_186;
wire n_1795;
wire n_1384;
wire n_1868;
wire n_1501;
wire n_1173;
wire n_1068;
wire n_1198;
wire n_1570;
wire n_487;
wire n_1518;
wire n_1456;
wire n_1879;
wire n_1886;
wire n_1648;
wire n_1413;
wire n_855;
wire n_808;
wire n_1365;
wire n_553;
wire n_1439;
wire n_814;
wire n_578;
wire n_1665;
wire n_1287;
wire n_405;
wire n_1611;
wire n_320;
wire n_1414;
wire n_1134;
wire n_1484;
wire n_647;
wire n_1423;
wire n_481;
wire n_600;
wire n_1053;
wire n_1609;
wire n_529;
wire n_1899;
wire n_502;
wire n_218;
wire n_1467;
wire n_247;
wire n_1828;
wire n_1798;
wire n_1304;
wire n_1608;
wire n_1744;
wire n_1105;
wire n_547;
wire n_439;
wire n_604;
wire n_677;
wire n_478;
wire n_703;
wire n_1349;
wire n_1709;
wire n_1061;
wire n_326;
wire n_681;
wire n_227;
wire n_874;
wire n_1278;
wire n_707;
wire n_983;
wire n_590;
wire n_699;
wire n_727;
wire n_301;
wire n_1726;
wire n_545;
wire n_1015;
wire n_1377;
wire n_1162;
wire n_536;
wire n_1614;
wire n_325;
wire n_1740;
wire n_1602;
wire n_688;
wire n_636;
wire n_427;
wire n_1098;
wire n_1490;
wire n_442;
wire n_777;
wire n_1553;
wire n_1080;
wire n_920;
wire n_1760;
wire n_1086;
wire n_1092;
wire n_986;
wire n_1104;
wire n_729;
wire n_887;
wire n_1122;
wire n_1205;
wire n_1408;
wire n_1693;
wire n_1132;
wire n_390;
wire n_1156;
wire n_501;
wire n_314;
wire n_1823;
wire n_1120;
wire n_1202;
wire n_627;
wire n_1188;
wire n_1498;
wire n_1371;
wire n_233;
wire n_957;
wire n_388;
wire n_1402;
wire n_1242;
wire n_1607;
wire n_1489;
wire n_1218;
wire n_321;
wire n_221;
wire n_1586;
wire n_861;
wire n_1543;
wire n_1431;
wire n_877;
wire n_1119;
wire n_1863;
wire n_1763;
wire n_1666;
wire n_1500;
wire n_616;
wire n_1055;
wire n_1395;
wire n_1346;
wire n_1189;
wire n_1089;
wire n_281;
wire n_1859;
wire n_262;
wire n_1502;
wire n_1523;
wire n_1478;
wire n_1883;
wire n_735;
wire n_297;
wire n_1005;
wire n_527;
wire n_1294;
wire n_1667;
wire n_845;
wire n_888;
wire n_1649;
wire n_1677;
wire n_1297;
wire n_551;
wire n_417;
wire n_1708;
wire n_343;
wire n_1222;
wire n_1844;
wire n_582;
wire n_755;
wire n_1097;
wire n_1219;
wire n_1711;
wire n_710;
wire n_534;
wire n_1791;
wire n_1894;
wire n_1460;
wire n_1239;
wire n_278;
wire n_560;
wire n_890;
wire n_842;
wire n_1898;
wire n_451;
wire n_745;
wire n_1741;
wire n_1572;
wire n_1793;
wire n_742;
wire n_1081;
wire n_1373;
wire n_1388;
wire n_1266;
wire n_1540;
wire n_1719;
wire n_769;
wire n_1797;
wire n_1753;
wire n_1372;
wire n_476;
wire n_832;
wire n_535;
wire n_744;
wire n_1895;
wire n_982;
wire n_1800;
wire n_915;
wire n_215;
wire n_1075;
wire n_454;
wire n_298;
wire n_1331;
wire n_1890;
wire n_1529;
wire n_1227;
wire n_655;
wire n_1734;
wire n_1860;
wire n_403;
wire n_1007;
wire n_1580;
wire n_1319;
wire n_657;
wire n_837;
wire n_812;
wire n_606;
wire n_951;
wire n_862;
wire n_1700;
wire n_659;
wire n_1332;
wire n_509;
wire n_1854;
wire n_666;
wire n_1747;
wire n_430;
wire n_1206;
wire n_1729;
wire n_722;
wire n_1508;
wire n_1532;
wire n_1171;
wire n_1030;
wire n_785;
wire n_1309;
wire n_999;
wire n_1766;
wire n_1338;
wire n_1342;
wire n_456;
wire n_1867;
wire n_852;
wire n_1394;
wire n_704;
wire n_1060;
wire n_1044;
wire n_1714;
wire n_521;
wire n_873;
wire n_1301;
wire n_1748;
wire n_1243;
wire n_1400;
wire n_342;
wire n_1466;
wire n_1513;
wire n_1527;
wire n_358;
wire n_1783;
wire n_608;
wire n_1538;
wire n_1037;
wire n_1329;
wire n_317;
wire n_1545;
wire n_1257;
wire n_1480;
wire n_1668;
wire n_1878;
wire n_1605;
wire n_1078;
wire n_266;
wire n_1897;
wire n_1161;
wire n_811;
wire n_624;
wire n_791;
wire n_876;
wire n_618;
wire n_1191;
wire n_736;
wire n_1025;
wire n_1215;
wire n_241;
wire n_1449;
wire n_687;
wire n_797;
wire n_1786;
wire n_480;
wire n_1327;
wire n_1475;
wire n_211;
wire n_642;
wire n_1804;
wire n_408;
wire n_1406;
wire n_595;
wire n_1405;
wire n_602;
wire n_1757;
wire n_592;
wire n_1499;
wire n_854;
wire n_1318;
wire n_393;
wire n_1632;
wire n_1769;
wire n_474;
wire n_805;
wire n_295;
wire n_1658;
wire n_190;
wire n_1072;
wire n_695;
wire n_1526;
wire n_1305;
wire n_730;
wire n_386;
wire n_1596;
wire n_1281;
wire n_516;
wire n_1137;
wire n_1873;
wire n_1258;
wire n_197;
wire n_640;
wire n_463;
wire n_1476;
wire n_1524;
wire n_1733;
wire n_1856;
wire n_943;
wire n_1118;
wire n_678;
wire n_651;
wire n_1874;
wire n_1293;
wire n_961;
wire n_469;
wire n_1046;
wire n_1807;
wire n_726;
wire n_1123;
wire n_1657;
wire n_878;
wire n_1784;
wire n_771;
wire n_1321;
wire n_752;
wire n_1488;
wire n_985;
wire n_421;
wire n_1330;
wire n_906;
wire n_1180;
wire n_1697;
wire n_283;
wire n_806;
wire n_1350;
wire n_1556;
wire n_649;
wire n_1561;
wire n_374;
wire n_1352;
wire n_1824;
wire n_643;
wire n_1492;
wire n_226;
wire n_1441;
wire n_1822;
wire n_682;
wire n_1616;
wire n_819;
wire n_586;
wire n_1324;
wire n_1429;
wire n_1778;
wire n_1776;
wire n_686;
wire n_605;
wire n_1154;
wire n_584;
wire n_1557;
wire n_1759;
wire n_1829;
wire n_1130;
wire n_1450;
wire n_349;
wire n_756;
wire n_1016;
wire n_1149;
wire n_1505;
wire n_979;
wire n_1642;
wire n_1815;
wire n_897;
wire n_949;
wire n_1493;
wire n_515;
wire n_807;
wire n_891;
wire n_885;
wire n_1659;
wire n_198;
wire n_1864;
wire n_1887;
wire n_1208;
wire n_396;
wire n_802;
wire n_1151;
wire n_554;
wire n_960;
wire n_1256;
wire n_714;
wire n_790;
wire n_354;
wire n_725;
wire n_1577;
wire n_1448;
wire n_1009;
wire n_230;
wire n_1133;
wire n_883;
wire n_473;
wire n_1852;
wire n_801;
wire n_1286;
wire n_818;
wire n_1685;
wire n_779;
wire n_594;
wire n_1877;
wire n_1397;
wire n_1052;
wire n_272;
wire n_1333;
wire n_1306;
wire n_1849;
wire n_833;
wire n_1426;
wire n_879;
wire n_1117;
wire n_422;
wire n_1269;
wire n_1303;
wire n_1547;
wire n_1438;
wire n_1541;
wire n_597;
wire n_1047;
wire n_1472;
wire n_1593;
wire n_1050;
wire n_566;
wire n_1201;
wire n_1288;
wire n_858;
wire n_1185;
wire n_335;
wire n_1035;
wire n_1143;
wire n_344;
wire n_426;
wire n_433;
wire n_398;
wire n_210;
wire n_1090;
wire n_1367;
wire n_253;
wire n_928;
wire n_1153;
wire n_271;
wire n_465;
wire n_825;
wire n_1103;
wire n_732;
wire n_1565;
wire n_1192;
wire n_224;
wire n_894;
wire n_1380;
wire n_1624;
wire n_1801;
wire n_420;
wire n_1291;
wire n_562;
wire n_748;
wire n_510;
wire n_1045;
wire n_256;
wire n_1160;
wire n_1882;
wire n_1023;
wire n_1881;
wire n_988;
wire n_330;
wire n_914;
wire n_400;
wire n_689;
wire n_1116;
wire n_282;
wire n_328;
wire n_368;
wire n_467;
wire n_1511;
wire n_1422;
wire n_644;
wire n_1197;
wire n_276;
wire n_497;
wire n_1165;
wire n_1641;
wire n_538;
wire n_1517;
wire n_576;
wire n_843;
wire n_511;
wire n_455;
wire n_429;
wire n_588;
wire n_638;
wire n_1307;
wire n_1128;
wire n_1671;
wire n_1417;
wire n_1048;
wire n_775;
wire n_667;
wire n_1049;
wire n_869;
wire n_846;
wire n_1398;
wire n_1356;
wire n_1341;
wire n_1504;
wire n_1773;
wire n_1440;
wire n_1370;
wire n_1603;
wire n_305;
wire n_312;
wire n_728;
wire n_413;
wire n_715;
wire n_889;
wire n_1066;
wire n_1549;
wire n_935;
wire n_685;
wire n_911;
wire n_361;
wire n_623;
wire n_1712;
wire n_1403;
wire n_1065;
wire n_453;
wire n_1534;
wire n_810;
wire n_1290;
wire n_617;
wire n_543;
wire n_1362;
wire n_1559;
wire n_236;
wire n_601;
wire n_683;
wire n_565;
wire n_628;
wire n_1300;
wire n_743;
wire n_1194;
wire n_1647;
wire n_1546;
wire n_1420;
wire n_907;
wire n_1454;
wire n_660;
wire n_464;
wire n_962;
wire n_941;
wire n_1210;
wire n_847;
wire n_747;
wire n_1622;
wire n_1135;
wire n_918;
wire n_1885;
wire n_639;
wire n_452;
wire n_673;
wire n_1038;
wire n_414;
wire n_571;
wire n_1521;
wire n_1694;
wire n_284;
wire n_593;
wire n_1695;
wire n_1164;
wire n_609;
wire n_1193;
wire n_1345;
wire n_613;
wire n_1022;
wire n_1336;
wire n_1033;
wire n_1774;
wire n_409;
wire n_519;
wire n_384;
wire n_1166;
wire n_1056;
wire n_526;
wire n_1767;
wire n_1040;
wire n_674;
wire n_1158;
wire n_316;
wire n_1444;
wire n_1803;
wire n_820;
wire n_1749;
wire n_872;
wire n_1653;
wire n_254;
wire n_1157;
wire n_1584;
wire n_234;
wire n_848;
wire n_1664;
wire n_280;
wire n_629;
wire n_1739;
wire n_1814;
wire n_532;
wire n_1789;
wire n_763;
wire n_540;
wire n_216;
wire n_692;
wire n_1857;
wire n_984;
wire n_1687;
wire n_223;
wire n_1552;
wire n_750;
wire n_834;
wire n_1612;
wire n_800;
wire n_1816;
wire n_1756;
wire n_1606;
wire n_395;
wire n_621;
wire n_1587;
wire n_213;
wire n_1772;
wire n_1014;
wire n_724;
wire n_1427;
wire n_1481;
wire n_493;
wire n_1311;
wire n_1589;
wire n_1100;
wire n_585;
wire n_875;
wire n_1617;
wire n_827;
wire n_697;
wire n_622;
wire n_1626;
wire n_1335;
wire n_1715;
wire n_296;
wire n_880;
wire n_793;
wire n_1175;
wire n_751;
wire n_1027;
wire n_1070;
wire n_1621;
wire n_739;
wire n_1485;
wire n_1028;
wire n_1221;
wire n_530;
wire n_1785;
wire n_792;
wire n_1262;
wire n_580;
wire n_1579;
wire n_494;
wire n_434;
wire n_975;
wire n_229;
wire n_394;
wire n_923;
wire n_1645;
wire n_1124;
wire n_1381;
wire n_1494;
wire n_932;
wire n_1893;
wire n_1183;
wire n_1326;
wire n_1805;
wire n_981;
wire n_1110;
wire n_1758;
wire n_243;
wire n_1407;
wire n_1204;
wire n_1554;
wire n_994;
wire n_1360;
wire n_973;
wire n_268;
wire n_972;
wire n_856;
wire n_1248;
wire n_1176;
wire n_1564;
wire n_1054;
wire n_508;
wire n_1679;
wire n_1858;
wire n_353;
wire n_1678;
wire n_1482;
wire n_1361;
wire n_1601;
wire n_1057;
wire n_191;
wire n_1834;
wire n_1011;
wire n_978;
wire n_1520;
wire n_1509;
wire n_828;
wire n_322;
wire n_1411;
wire n_1359;
wire n_558;
wire n_1721;
wire n_653;
wire n_1445;
wire n_1317;
wire n_783;
wire n_556;
wire n_1127;
wire n_1536;
wire n_1471;
wire n_1008;
wire n_332;
wire n_581;
wire n_294;
wire n_1024;
wire n_830;
wire n_987;
wire n_936;
wire n_1620;
wire n_1385;
wire n_1525;
wire n_541;
wire n_499;
wire n_1775;
wire n_788;
wire n_908;
wire n_1036;
wire n_341;
wire n_1270;
wire n_1167;
wire n_1272;
wire n_549;
wire n_591;
wire n_969;
wire n_919;
wire n_1663;
wire n_1625;
wire n_318;
wire n_1458;
wire n_244;
wire n_679;
wire n_1630;
wire n_220;
wire n_663;
wire n_1720;
wire n_443;
wire n_1412;
wire n_1738;
wire n_1550;
wire n_528;
wire n_1358;
wire n_1200;
wire n_387;
wire n_406;
wire n_826;
wire n_1735;
wire n_1788;
wire n_391;
wire n_940;
wire n_1537;
wire n_1077;
wire n_607;
wire n_956;
wire n_445;
wire n_765;
wire n_1809;
wire n_1843;
wire n_1268;
wire n_385;
wire n_917;
wire n_1271;
wire n_372;
wire n_1530;
wire n_631;
wire n_399;
wire n_1170;
wire n_1261;
wire n_702;
wire n_857;
wire n_898;
wire n_363;
wire n_968;
wire n_1067;
wire n_1235;
wire n_1323;
wire n_1462;
wire n_1064;
wire n_633;
wire n_900;
wire n_1446;
wire n_1282;
wire n_1701;
wire n_1093;
wire n_1551;
wire n_1755;
wire n_1285;
wire n_193;
wire n_733;
wire n_761;
wire n_731;
wire n_336;
wire n_1813;
wire n_315;
wire n_311;
wire n_1452;
wire n_1573;
wire n_668;
wire n_758;
wire n_1106;
wire n_648;
wire n_784;
wire n_269;
wire n_816;
wire n_1322;
wire n_1473;
wire n_835;
wire n_446;
wire n_1076;
wire n_1348;
wire n_753;
wire n_1770;
wire n_701;
wire n_1003;
wire n_1125;
wire n_1710;
wire n_1865;
wire n_309;
wire n_1344;
wire n_1390;
wire n_401;
wire n_485;
wire n_1792;
wire n_504;
wire n_483;
wire n_435;
wire n_1141;
wire n_1629;
wire n_291;
wire n_1640;
wire n_822;
wire n_1094;
wire n_840;
wire n_1459;
wire n_1510;
wire n_1099;
wire n_839;
wire n_1754;
wire n_759;
wire n_567;
wire n_369;
wire n_240;
wire n_1727;
wire n_1575;
wire n_1848;
wire n_1892;
wire n_1172;
wire n_614;
wire n_1212;
wire n_831;
wire n_778;
wire n_1619;
wire n_188;
wire n_323;
wire n_550;
wire n_1315;
wire n_1660;
wire n_997;
wire n_635;
wire n_694;
wire n_1643;
wire n_1320;
wire n_1113;
wire n_248;
wire n_1152;
wire n_1845;
wire n_921;
wire n_1615;
wire n_1236;
wire n_228;
wire n_1265;
wire n_1576;
wire n_1470;
wire n_671;
wire n_1533;
wire n_1806;
wire n_1409;
wire n_1148;
wire n_1684;
wire n_1588;
wire n_1673;
wire n_1334;
wire n_654;
wire n_1275;
wire n_488;
wire n_904;
wire n_505;
wire n_1696;
wire n_498;
wire n_1875;
wire n_1059;
wire n_684;
wire n_1039;
wire n_539;
wire n_1150;
wire n_977;
wire n_449;
wire n_392;
wire n_1628;
wire n_1289;
wire n_1831;
wire n_1497;
wire n_1866;
wire n_459;
wire n_1136;
wire n_1782;
wire n_458;
wire n_1190;
wire n_1600;
wire n_1144;
wire n_383;
wire n_838;
wire n_1558;
wire n_1316;
wire n_950;
wire n_1017;
wire n_711;
wire n_734;
wire n_723;
wire n_1393;
wire n_658;
wire n_630;
wire n_1369;
wire n_362;
wire n_310;
wire n_1781;
wire n_709;
wire n_809;
wire n_1686;
wire n_235;
wire n_881;
wire n_1019;
wire n_1477;
wire n_1777;
wire n_662;
wire n_641;
wire n_910;
wire n_290;
wire n_741;
wire n_939;
wire n_1410;
wire n_371;
wire n_199;
wire n_217;
wire n_1114;
wire n_1325;
wire n_1742;
wire n_708;
wire n_308;
wire n_1223;
wire n_201;
wire n_1768;
wire n_572;
wire n_1199;
wire n_865;
wire n_1273;
wire n_1041;
wire n_993;
wire n_1862;
wire n_948;
wire n_922;
wire n_1004;
wire n_1810;
wire n_448;
wire n_1347;
wire n_860;
wire n_1043;
wire n_255;
wire n_450;
wire n_1764;
wire n_896;
wire n_1737;
wire n_1479;
wire n_1613;
wire n_902;
wire n_1031;
wire n_1723;
wire n_1638;
wire n_853;
wire n_716;
wire n_1571;
wire n_1698;
wire n_196;
wire n_1337;
wire n_774;
wire n_933;
wire n_1779;
wire n_596;
wire n_954;
wire n_1168;
wire n_1821;
wire n_219;
wire n_1310;
wire n_231;
wire n_656;
wire n_492;
wire n_574;
wire n_664;
wire n_252;
wire n_1591;
wire n_1229;
wire n_1683;
wire n_1896;
wire n_1732;
wire n_415;
wire n_1280;
wire n_544;
wire n_1516;
wire n_1186;
wire n_1705;
wire n_599;
wire n_768;
wire n_1091;
wire n_537;
wire n_1063;
wire n_991;
wire n_389;
wire n_1724;
wire n_1670;
wire n_1707;
wire n_1799;
wire n_1126;
wire n_195;
wire n_1846;
wire n_938;
wire n_1891;
wire n_1328;
wire n_895;
wire n_304;
wire n_1639;
wire n_583;
wire n_1302;
wire n_1000;
wire n_313;
wire n_626;
wire n_378;
wire n_1581;
wire n_946;
wire n_757;
wire n_375;
wire n_1655;
wire n_1818;
wire n_1146;
wire n_1634;
wire n_1203;
wire n_998;
wire n_1699;
wire n_1598;
wire n_472;
wire n_937;
wire n_1474;
wire n_265;
wire n_1583;
wire n_1604;
wire n_208;
wire n_1631;
wire n_1702;
wire n_275;
wire n_1794;
wire n_1375;
wire n_204;
wire n_1232;
wire n_996;
wire n_1211;
wire n_1368;
wire n_963;
wire n_1264;
wire n_1082;
wire n_1725;
wire n_496;
wire n_1827;
wire n_866;
wire n_246;
wire n_925;
wire n_1752;
wire n_1313;
wire n_1001;
wire n_1722;
wire n_1115;
wire n_1339;
wire n_1002;
wire n_1644;
wire n_1051;
wire n_719;
wire n_263;
wire n_1102;
wire n_360;
wire n_1129;
wire n_1252;
wire n_250;
wire n_1464;
wire n_1296;
wire n_773;
wire n_1010;
wire n_882;
wire n_1249;
wire n_803;
wire n_1871;
wire n_329;
wire n_718;
wire n_1434;
wire n_340;
wire n_1569;
wire n_289;
wire n_548;
wire n_523;
wire n_1662;
wire n_457;
wire n_1299;
wire n_1870;
wire n_782;
wire n_364;
wire n_258;
wire n_431;
wire n_1861;
wire n_1228;
wire n_1244;
wire n_1796;
wire n_411;
wire n_484;
wire n_849;
wire n_1820;
wire n_357;
wire n_412;
wire n_1251;
wire n_447;
wire n_1421;
wire n_1762;
wire n_1233;
wire n_1808;
wire n_1574;
wire n_1672;
wire n_1635;
wire n_1704;
wire n_893;
wire n_1582;
wire n_841;
wire n_886;
wire n_1069;
wire n_359;
wire n_1308;
wire n_573;
wire n_796;
wire n_531;
wire n_1730;
wire n_1374;
wire n_1451;
wire n_1487;
wire n_675;

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_180),
.Y(n_186)
);

CKINVDCx5p33_ASAP7_75t_R g187 ( 
.A(n_105),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_58),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_2),
.Y(n_189)
);

CKINVDCx5p33_ASAP7_75t_R g190 ( 
.A(n_51),
.Y(n_190)
);

INVx2_ASAP7_75t_SL g191 ( 
.A(n_119),
.Y(n_191)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_57),
.Y(n_192)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_147),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_106),
.Y(n_194)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_74),
.Y(n_195)
);

BUFx10_ASAP7_75t_L g196 ( 
.A(n_37),
.Y(n_196)
);

INVx1_ASAP7_75t_SL g197 ( 
.A(n_120),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_176),
.Y(n_198)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_41),
.Y(n_199)
);

CKINVDCx5p33_ASAP7_75t_R g200 ( 
.A(n_85),
.Y(n_200)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_185),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_157),
.Y(n_202)
);

CKINVDCx5p33_ASAP7_75t_R g203 ( 
.A(n_3),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_117),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_66),
.Y(n_205)
);

CKINVDCx5p33_ASAP7_75t_R g206 ( 
.A(n_40),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_64),
.Y(n_207)
);

CKINVDCx5p33_ASAP7_75t_R g208 ( 
.A(n_171),
.Y(n_208)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_44),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_14),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_113),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_115),
.Y(n_213)
);

INVx2_ASAP7_75t_L g214 ( 
.A(n_70),
.Y(n_214)
);

HB1xp67_ASAP7_75t_L g215 ( 
.A(n_84),
.Y(n_215)
);

CKINVDCx5p33_ASAP7_75t_R g216 ( 
.A(n_23),
.Y(n_216)
);

INVx1_ASAP7_75t_SL g217 ( 
.A(n_132),
.Y(n_217)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_182),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_148),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_86),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_63),
.Y(n_221)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_135),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_97),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_152),
.Y(n_224)
);

CKINVDCx5p33_ASAP7_75t_R g225 ( 
.A(n_145),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_24),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_90),
.Y(n_227)
);

CKINVDCx5p33_ASAP7_75t_R g228 ( 
.A(n_100),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_183),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_17),
.Y(n_230)
);

CKINVDCx5p33_ASAP7_75t_R g231 ( 
.A(n_43),
.Y(n_231)
);

CKINVDCx5p33_ASAP7_75t_R g232 ( 
.A(n_17),
.Y(n_232)
);

CKINVDCx5p33_ASAP7_75t_R g233 ( 
.A(n_96),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_52),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_159),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_23),
.Y(n_236)
);

INVx1_ASAP7_75t_L g237 ( 
.A(n_137),
.Y(n_237)
);

CKINVDCx5p33_ASAP7_75t_R g238 ( 
.A(n_149),
.Y(n_238)
);

CKINVDCx5p33_ASAP7_75t_R g239 ( 
.A(n_140),
.Y(n_239)
);

INVx2_ASAP7_75t_L g240 ( 
.A(n_126),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g241 ( 
.A(n_67),
.Y(n_241)
);

CKINVDCx5p33_ASAP7_75t_R g242 ( 
.A(n_31),
.Y(n_242)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_168),
.Y(n_243)
);

CKINVDCx5p33_ASAP7_75t_R g244 ( 
.A(n_61),
.Y(n_244)
);

CKINVDCx5p33_ASAP7_75t_R g245 ( 
.A(n_61),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_55),
.Y(n_246)
);

CKINVDCx5p33_ASAP7_75t_R g247 ( 
.A(n_36),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_110),
.Y(n_248)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_101),
.Y(n_249)
);

BUFx8_ASAP7_75t_SL g250 ( 
.A(n_173),
.Y(n_250)
);

CKINVDCx5p33_ASAP7_75t_R g251 ( 
.A(n_43),
.Y(n_251)
);

CKINVDCx5p33_ASAP7_75t_R g252 ( 
.A(n_111),
.Y(n_252)
);

CKINVDCx5p33_ASAP7_75t_R g253 ( 
.A(n_5),
.Y(n_253)
);

CKINVDCx5p33_ASAP7_75t_R g254 ( 
.A(n_45),
.Y(n_254)
);

CKINVDCx5p33_ASAP7_75t_R g255 ( 
.A(n_62),
.Y(n_255)
);

CKINVDCx5p33_ASAP7_75t_R g256 ( 
.A(n_14),
.Y(n_256)
);

CKINVDCx5p33_ASAP7_75t_R g257 ( 
.A(n_146),
.Y(n_257)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_112),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_163),
.Y(n_259)
);

CKINVDCx5p33_ASAP7_75t_R g260 ( 
.A(n_35),
.Y(n_260)
);

BUFx2_ASAP7_75t_L g261 ( 
.A(n_22),
.Y(n_261)
);

CKINVDCx5p33_ASAP7_75t_R g262 ( 
.A(n_18),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_36),
.Y(n_263)
);

CKINVDCx5p33_ASAP7_75t_R g264 ( 
.A(n_127),
.Y(n_264)
);

CKINVDCx5p33_ASAP7_75t_R g265 ( 
.A(n_69),
.Y(n_265)
);

HB1xp67_ASAP7_75t_L g266 ( 
.A(n_172),
.Y(n_266)
);

CKINVDCx5p33_ASAP7_75t_R g267 ( 
.A(n_72),
.Y(n_267)
);

CKINVDCx5p33_ASAP7_75t_R g268 ( 
.A(n_1),
.Y(n_268)
);

BUFx5_ASAP7_75t_L g269 ( 
.A(n_133),
.Y(n_269)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_0),
.Y(n_270)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_76),
.Y(n_271)
);

CKINVDCx5p33_ASAP7_75t_R g272 ( 
.A(n_181),
.Y(n_272)
);

INVx2_ASAP7_75t_L g273 ( 
.A(n_12),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_54),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_107),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_19),
.Y(n_276)
);

CKINVDCx5p33_ASAP7_75t_R g277 ( 
.A(n_33),
.Y(n_277)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_114),
.Y(n_278)
);

CKINVDCx5p33_ASAP7_75t_R g279 ( 
.A(n_26),
.Y(n_279)
);

BUFx8_ASAP7_75t_SL g280 ( 
.A(n_0),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_91),
.Y(n_281)
);

CKINVDCx5p33_ASAP7_75t_R g282 ( 
.A(n_89),
.Y(n_282)
);

CKINVDCx5p33_ASAP7_75t_R g283 ( 
.A(n_49),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_34),
.Y(n_284)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_174),
.Y(n_285)
);

CKINVDCx14_ASAP7_75t_R g286 ( 
.A(n_37),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g287 ( 
.A(n_40),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_130),
.Y(n_288)
);

BUFx10_ASAP7_75t_L g289 ( 
.A(n_118),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_162),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_158),
.Y(n_291)
);

BUFx8_ASAP7_75t_SL g292 ( 
.A(n_103),
.Y(n_292)
);

CKINVDCx5p33_ASAP7_75t_R g293 ( 
.A(n_38),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_53),
.Y(n_294)
);

CKINVDCx5p33_ASAP7_75t_R g295 ( 
.A(n_136),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_33),
.Y(n_296)
);

CKINVDCx5p33_ASAP7_75t_R g297 ( 
.A(n_6),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_131),
.Y(n_298)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_121),
.Y(n_299)
);

INVx2_ASAP7_75t_SL g300 ( 
.A(n_57),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g301 ( 
.A(n_45),
.Y(n_301)
);

CKINVDCx5p33_ASAP7_75t_R g302 ( 
.A(n_34),
.Y(n_302)
);

CKINVDCx5p33_ASAP7_75t_R g303 ( 
.A(n_129),
.Y(n_303)
);

CKINVDCx16_ASAP7_75t_R g304 ( 
.A(n_164),
.Y(n_304)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_175),
.Y(n_305)
);

BUFx2_ASAP7_75t_L g306 ( 
.A(n_9),
.Y(n_306)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_48),
.Y(n_307)
);

CKINVDCx5p33_ASAP7_75t_R g308 ( 
.A(n_54),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_35),
.Y(n_309)
);

CKINVDCx5p33_ASAP7_75t_R g310 ( 
.A(n_39),
.Y(n_310)
);

INVx1_ASAP7_75t_SL g311 ( 
.A(n_53),
.Y(n_311)
);

CKINVDCx5p33_ASAP7_75t_R g312 ( 
.A(n_21),
.Y(n_312)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_160),
.Y(n_313)
);

CKINVDCx5p33_ASAP7_75t_R g314 ( 
.A(n_8),
.Y(n_314)
);

CKINVDCx5p33_ASAP7_75t_R g315 ( 
.A(n_108),
.Y(n_315)
);

CKINVDCx5p33_ASAP7_75t_R g316 ( 
.A(n_178),
.Y(n_316)
);

INVx1_ASAP7_75t_L g317 ( 
.A(n_92),
.Y(n_317)
);

INVx2_ASAP7_75t_L g318 ( 
.A(n_124),
.Y(n_318)
);

CKINVDCx16_ASAP7_75t_R g319 ( 
.A(n_30),
.Y(n_319)
);

CKINVDCx5p33_ASAP7_75t_R g320 ( 
.A(n_122),
.Y(n_320)
);

CKINVDCx5p33_ASAP7_75t_R g321 ( 
.A(n_4),
.Y(n_321)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_13),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_30),
.Y(n_323)
);

BUFx5_ASAP7_75t_L g324 ( 
.A(n_75),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_16),
.Y(n_325)
);

INVx1_ASAP7_75t_SL g326 ( 
.A(n_46),
.Y(n_326)
);

CKINVDCx5p33_ASAP7_75t_R g327 ( 
.A(n_109),
.Y(n_327)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_20),
.Y(n_328)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_93),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_9),
.Y(n_330)
);

CKINVDCx5p33_ASAP7_75t_R g331 ( 
.A(n_44),
.Y(n_331)
);

CKINVDCx20_ASAP7_75t_R g332 ( 
.A(n_80),
.Y(n_332)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_62),
.Y(n_333)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_83),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_139),
.Y(n_335)
);

CKINVDCx5p33_ASAP7_75t_R g336 ( 
.A(n_94),
.Y(n_336)
);

CKINVDCx5p33_ASAP7_75t_R g337 ( 
.A(n_42),
.Y(n_337)
);

CKINVDCx5p33_ASAP7_75t_R g338 ( 
.A(n_104),
.Y(n_338)
);

BUFx2_ASAP7_75t_L g339 ( 
.A(n_169),
.Y(n_339)
);

CKINVDCx5p33_ASAP7_75t_R g340 ( 
.A(n_21),
.Y(n_340)
);

CKINVDCx5p33_ASAP7_75t_R g341 ( 
.A(n_10),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g342 ( 
.A(n_24),
.Y(n_342)
);

CKINVDCx5p33_ASAP7_75t_R g343 ( 
.A(n_18),
.Y(n_343)
);

CKINVDCx5p33_ASAP7_75t_R g344 ( 
.A(n_177),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_165),
.Y(n_345)
);

CKINVDCx5p33_ASAP7_75t_R g346 ( 
.A(n_12),
.Y(n_346)
);

CKINVDCx5p33_ASAP7_75t_R g347 ( 
.A(n_125),
.Y(n_347)
);

CKINVDCx5p33_ASAP7_75t_R g348 ( 
.A(n_73),
.Y(n_348)
);

INVx2_ASAP7_75t_SL g349 ( 
.A(n_51),
.Y(n_349)
);

CKINVDCx5p33_ASAP7_75t_R g350 ( 
.A(n_55),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_95),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_8),
.Y(n_352)
);

INVx2_ASAP7_75t_SL g353 ( 
.A(n_81),
.Y(n_353)
);

INVx2_ASAP7_75t_SL g354 ( 
.A(n_65),
.Y(n_354)
);

CKINVDCx5p33_ASAP7_75t_R g355 ( 
.A(n_29),
.Y(n_355)
);

CKINVDCx5p33_ASAP7_75t_R g356 ( 
.A(n_166),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_52),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_26),
.Y(n_358)
);

CKINVDCx5p33_ASAP7_75t_R g359 ( 
.A(n_142),
.Y(n_359)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_184),
.Y(n_360)
);

CKINVDCx5p33_ASAP7_75t_R g361 ( 
.A(n_170),
.Y(n_361)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_151),
.Y(n_362)
);

BUFx2_ASAP7_75t_L g363 ( 
.A(n_150),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_167),
.Y(n_364)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_4),
.Y(n_365)
);

CKINVDCx5p33_ASAP7_75t_R g366 ( 
.A(n_56),
.Y(n_366)
);

CKINVDCx5p33_ASAP7_75t_R g367 ( 
.A(n_59),
.Y(n_367)
);

CKINVDCx5p33_ASAP7_75t_R g368 ( 
.A(n_99),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_41),
.Y(n_369)
);

CKINVDCx5p33_ASAP7_75t_R g370 ( 
.A(n_47),
.Y(n_370)
);

CKINVDCx5p33_ASAP7_75t_R g371 ( 
.A(n_280),
.Y(n_371)
);

NOR2xp33_ASAP7_75t_L g372 ( 
.A(n_339),
.B(n_1),
.Y(n_372)
);

CKINVDCx5p33_ASAP7_75t_R g373 ( 
.A(n_250),
.Y(n_373)
);

CKINVDCx5p33_ASAP7_75t_R g374 ( 
.A(n_292),
.Y(n_374)
);

INVxp67_ASAP7_75t_SL g375 ( 
.A(n_301),
.Y(n_375)
);

INVx1_ASAP7_75t_L g376 ( 
.A(n_358),
.Y(n_376)
);

INVx1_ASAP7_75t_L g377 ( 
.A(n_358),
.Y(n_377)
);

CKINVDCx20_ASAP7_75t_R g378 ( 
.A(n_286),
.Y(n_378)
);

CKINVDCx5p33_ASAP7_75t_R g379 ( 
.A(n_319),
.Y(n_379)
);

INVx1_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g381 ( 
.A(n_363),
.B(n_2),
.Y(n_381)
);

CKINVDCx20_ASAP7_75t_R g382 ( 
.A(n_193),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g383 ( 
.A(n_261),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_358),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_358),
.Y(n_385)
);

HB1xp67_ASAP7_75t_L g386 ( 
.A(n_306),
.Y(n_386)
);

CKINVDCx5p33_ASAP7_75t_R g387 ( 
.A(n_198),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g388 ( 
.A(n_304),
.Y(n_388)
);

CKINVDCx5p33_ASAP7_75t_R g389 ( 
.A(n_212),
.Y(n_389)
);

CKINVDCx20_ASAP7_75t_R g390 ( 
.A(n_224),
.Y(n_390)
);

CKINVDCx5p33_ASAP7_75t_R g391 ( 
.A(n_241),
.Y(n_391)
);

INVx1_ASAP7_75t_L g392 ( 
.A(n_246),
.Y(n_392)
);

INVxp67_ASAP7_75t_SL g393 ( 
.A(n_301),
.Y(n_393)
);

HB1xp67_ASAP7_75t_L g394 ( 
.A(n_188),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_246),
.Y(n_395)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_273),
.Y(n_396)
);

INVx1_ASAP7_75t_L g397 ( 
.A(n_273),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_357),
.Y(n_398)
);

INVxp67_ASAP7_75t_SL g399 ( 
.A(n_357),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_269),
.Y(n_400)
);

CKINVDCx20_ASAP7_75t_R g401 ( 
.A(n_288),
.Y(n_401)
);

BUFx2_ASAP7_75t_L g402 ( 
.A(n_188),
.Y(n_402)
);

INVxp67_ASAP7_75t_SL g403 ( 
.A(n_369),
.Y(n_403)
);

CKINVDCx5p33_ASAP7_75t_R g404 ( 
.A(n_329),
.Y(n_404)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_332),
.Y(n_405)
);

CKINVDCx20_ASAP7_75t_R g406 ( 
.A(n_345),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_369),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g408 ( 
.A(n_209),
.Y(n_408)
);

INVx1_ASAP7_75t_L g409 ( 
.A(n_195),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_195),
.Y(n_410)
);

CKINVDCx5p33_ASAP7_75t_R g411 ( 
.A(n_232),
.Y(n_411)
);

CKINVDCx5p33_ASAP7_75t_R g412 ( 
.A(n_236),
.Y(n_412)
);

INVxp67_ASAP7_75t_L g413 ( 
.A(n_300),
.Y(n_413)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_342),
.Y(n_414)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_214),
.Y(n_415)
);

INVx1_ASAP7_75t_L g416 ( 
.A(n_214),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_289),
.Y(n_417)
);

INVx1_ASAP7_75t_L g418 ( 
.A(n_222),
.Y(n_418)
);

INVxp33_ASAP7_75t_L g419 ( 
.A(n_192),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_222),
.Y(n_420)
);

CKINVDCx5p33_ASAP7_75t_R g421 ( 
.A(n_242),
.Y(n_421)
);

HB1xp67_ASAP7_75t_L g422 ( 
.A(n_189),
.Y(n_422)
);

INVxp33_ASAP7_75t_SL g423 ( 
.A(n_189),
.Y(n_423)
);

INVxp67_ASAP7_75t_L g424 ( 
.A(n_300),
.Y(n_424)
);

CKINVDCx20_ASAP7_75t_R g425 ( 
.A(n_289),
.Y(n_425)
);

INVx1_ASAP7_75t_L g426 ( 
.A(n_240),
.Y(n_426)
);

CKINVDCx20_ASAP7_75t_R g427 ( 
.A(n_289),
.Y(n_427)
);

CKINVDCx5p33_ASAP7_75t_R g428 ( 
.A(n_244),
.Y(n_428)
);

BUFx2_ASAP7_75t_L g429 ( 
.A(n_190),
.Y(n_429)
);

CKINVDCx5p33_ASAP7_75t_R g430 ( 
.A(n_245),
.Y(n_430)
);

CKINVDCx5p33_ASAP7_75t_R g431 ( 
.A(n_247),
.Y(n_431)
);

INVx1_ASAP7_75t_L g432 ( 
.A(n_240),
.Y(n_432)
);

CKINVDCx20_ASAP7_75t_R g433 ( 
.A(n_196),
.Y(n_433)
);

CKINVDCx5p33_ASAP7_75t_R g434 ( 
.A(n_251),
.Y(n_434)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_190),
.B(n_3),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_318),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_318),
.Y(n_437)
);

NOR2xp33_ASAP7_75t_L g438 ( 
.A(n_215),
.B(n_5),
.Y(n_438)
);

HB1xp67_ASAP7_75t_L g439 ( 
.A(n_203),
.Y(n_439)
);

CKINVDCx5p33_ASAP7_75t_R g440 ( 
.A(n_253),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_196),
.Y(n_441)
);

BUFx2_ASAP7_75t_SL g442 ( 
.A(n_191),
.Y(n_442)
);

INVx1_ASAP7_75t_L g443 ( 
.A(n_199),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_234),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_263),
.Y(n_445)
);

CKINVDCx5p33_ASAP7_75t_R g446 ( 
.A(n_254),
.Y(n_446)
);

CKINVDCx5p33_ASAP7_75t_R g447 ( 
.A(n_255),
.Y(n_447)
);

INVxp33_ASAP7_75t_SL g448 ( 
.A(n_203),
.Y(n_448)
);

HB1xp67_ASAP7_75t_L g449 ( 
.A(n_206),
.Y(n_449)
);

CKINVDCx5p33_ASAP7_75t_R g450 ( 
.A(n_256),
.Y(n_450)
);

CKINVDCx5p33_ASAP7_75t_R g451 ( 
.A(n_260),
.Y(n_451)
);

CKINVDCx5p33_ASAP7_75t_R g452 ( 
.A(n_262),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_196),
.Y(n_453)
);

CKINVDCx5p33_ASAP7_75t_R g454 ( 
.A(n_268),
.Y(n_454)
);

CKINVDCx20_ASAP7_75t_R g455 ( 
.A(n_206),
.Y(n_455)
);

CKINVDCx5p33_ASAP7_75t_R g456 ( 
.A(n_277),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_270),
.Y(n_457)
);

INVx2_ASAP7_75t_L g458 ( 
.A(n_269),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_274),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_276),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_269),
.Y(n_461)
);

CKINVDCx5p33_ASAP7_75t_R g462 ( 
.A(n_279),
.Y(n_462)
);

CKINVDCx20_ASAP7_75t_R g463 ( 
.A(n_211),
.Y(n_463)
);

CKINVDCx5p33_ASAP7_75t_R g464 ( 
.A(n_283),
.Y(n_464)
);

BUFx2_ASAP7_75t_L g465 ( 
.A(n_211),
.Y(n_465)
);

CKINVDCx5p33_ASAP7_75t_R g466 ( 
.A(n_387),
.Y(n_466)
);

BUFx6f_ASAP7_75t_L g467 ( 
.A(n_400),
.Y(n_467)
);

CKINVDCx5p33_ASAP7_75t_R g468 ( 
.A(n_389),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_400),
.Y(n_469)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_376),
.Y(n_470)
);

INVx2_ASAP7_75t_L g471 ( 
.A(n_400),
.Y(n_471)
);

CKINVDCx5p33_ASAP7_75t_R g472 ( 
.A(n_391),
.Y(n_472)
);

CKINVDCx5p33_ASAP7_75t_R g473 ( 
.A(n_404),
.Y(n_473)
);

BUFx2_ASAP7_75t_L g474 ( 
.A(n_455),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_377),
.Y(n_475)
);

CKINVDCx5p33_ASAP7_75t_R g476 ( 
.A(n_373),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_377),
.Y(n_477)
);

BUFx6f_ASAP7_75t_L g478 ( 
.A(n_458),
.Y(n_478)
);

INVx1_ASAP7_75t_L g479 ( 
.A(n_380),
.Y(n_479)
);

CKINVDCx5p33_ASAP7_75t_R g480 ( 
.A(n_374),
.Y(n_480)
);

HB1xp67_ASAP7_75t_L g481 ( 
.A(n_402),
.Y(n_481)
);

INVx3_ASAP7_75t_L g482 ( 
.A(n_458),
.Y(n_482)
);

NAND2xp5_ASAP7_75t_L g483 ( 
.A(n_409),
.B(n_266),
.Y(n_483)
);

OA21x2_ASAP7_75t_L g484 ( 
.A1(n_380),
.A2(n_202),
.B(n_201),
.Y(n_484)
);

HB1xp67_ASAP7_75t_L g485 ( 
.A(n_402),
.Y(n_485)
);

INVx1_ASAP7_75t_L g486 ( 
.A(n_384),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_384),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_385),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g489 ( 
.A(n_408),
.Y(n_489)
);

CKINVDCx5p33_ASAP7_75t_R g490 ( 
.A(n_382),
.Y(n_490)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_442),
.B(n_191),
.Y(n_491)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_385),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_442),
.B(n_353),
.Y(n_493)
);

INVx1_ASAP7_75t_L g494 ( 
.A(n_409),
.Y(n_494)
);

BUFx3_ASAP7_75t_L g495 ( 
.A(n_458),
.Y(n_495)
);

CKINVDCx5p33_ASAP7_75t_R g496 ( 
.A(n_390),
.Y(n_496)
);

CKINVDCx5p33_ASAP7_75t_R g497 ( 
.A(n_401),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_410),
.Y(n_498)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_381),
.B(n_353),
.Y(n_499)
);

INVx2_ASAP7_75t_L g500 ( 
.A(n_461),
.Y(n_500)
);

HB1xp67_ASAP7_75t_L g501 ( 
.A(n_429),
.Y(n_501)
);

INVx2_ASAP7_75t_L g502 ( 
.A(n_461),
.Y(n_502)
);

CKINVDCx5p33_ASAP7_75t_R g503 ( 
.A(n_405),
.Y(n_503)
);

CKINVDCx5p33_ASAP7_75t_R g504 ( 
.A(n_406),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_L g505 ( 
.A(n_410),
.B(n_205),
.Y(n_505)
);

CKINVDCx20_ASAP7_75t_R g506 ( 
.A(n_414),
.Y(n_506)
);

AND2x2_ASAP7_75t_SL g507 ( 
.A(n_381),
.B(n_207),
.Y(n_507)
);

CKINVDCx5p33_ASAP7_75t_R g508 ( 
.A(n_371),
.Y(n_508)
);

CKINVDCx20_ASAP7_75t_R g509 ( 
.A(n_378),
.Y(n_509)
);

INVx2_ASAP7_75t_L g510 ( 
.A(n_461),
.Y(n_510)
);

CKINVDCx5p33_ASAP7_75t_R g511 ( 
.A(n_411),
.Y(n_511)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_415),
.Y(n_512)
);

CKINVDCx5p33_ASAP7_75t_R g513 ( 
.A(n_412),
.Y(n_513)
);

INVx2_ASAP7_75t_L g514 ( 
.A(n_415),
.Y(n_514)
);

NOR2xp33_ASAP7_75t_L g515 ( 
.A(n_375),
.B(n_354),
.Y(n_515)
);

CKINVDCx5p33_ASAP7_75t_R g516 ( 
.A(n_421),
.Y(n_516)
);

CKINVDCx5p33_ASAP7_75t_R g517 ( 
.A(n_428),
.Y(n_517)
);

INVx2_ASAP7_75t_L g518 ( 
.A(n_416),
.Y(n_518)
);

CKINVDCx5p33_ASAP7_75t_R g519 ( 
.A(n_430),
.Y(n_519)
);

CKINVDCx5p33_ASAP7_75t_R g520 ( 
.A(n_431),
.Y(n_520)
);

AND3x2_ASAP7_75t_L g521 ( 
.A(n_386),
.B(n_296),
.C(n_294),
.Y(n_521)
);

CKINVDCx5p33_ASAP7_75t_R g522 ( 
.A(n_434),
.Y(n_522)
);

BUFx6f_ASAP7_75t_L g523 ( 
.A(n_416),
.Y(n_523)
);

INVx2_ASAP7_75t_L g524 ( 
.A(n_418),
.Y(n_524)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_418),
.Y(n_525)
);

INVx2_ASAP7_75t_L g526 ( 
.A(n_420),
.Y(n_526)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_420),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g528 ( 
.A(n_426),
.B(n_210),
.Y(n_528)
);

CKINVDCx5p33_ASAP7_75t_R g529 ( 
.A(n_440),
.Y(n_529)
);

BUFx3_ASAP7_75t_L g530 ( 
.A(n_426),
.Y(n_530)
);

BUFx2_ASAP7_75t_L g531 ( 
.A(n_463),
.Y(n_531)
);

NAND2xp5_ASAP7_75t_L g532 ( 
.A(n_432),
.B(n_436),
.Y(n_532)
);

INVx2_ASAP7_75t_L g533 ( 
.A(n_432),
.Y(n_533)
);

INVx2_ASAP7_75t_L g534 ( 
.A(n_436),
.Y(n_534)
);

INVx1_ASAP7_75t_L g535 ( 
.A(n_437),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_437),
.Y(n_536)
);

CKINVDCx5p33_ASAP7_75t_R g537 ( 
.A(n_446),
.Y(n_537)
);

BUFx6f_ASAP7_75t_L g538 ( 
.A(n_392),
.Y(n_538)
);

CKINVDCx5p33_ASAP7_75t_R g539 ( 
.A(n_447),
.Y(n_539)
);

CKINVDCx5p33_ASAP7_75t_R g540 ( 
.A(n_450),
.Y(n_540)
);

AND2x2_ASAP7_75t_L g541 ( 
.A(n_399),
.B(n_349),
.Y(n_541)
);

CKINVDCx5p33_ASAP7_75t_R g542 ( 
.A(n_451),
.Y(n_542)
);

INVx2_ASAP7_75t_L g543 ( 
.A(n_392),
.Y(n_543)
);

AND2x2_ASAP7_75t_L g544 ( 
.A(n_481),
.B(n_388),
.Y(n_544)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_530),
.Y(n_545)
);

INVx2_ASAP7_75t_L g546 ( 
.A(n_523),
.Y(n_546)
);

INVx2_ASAP7_75t_L g547 ( 
.A(n_471),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_L g548 ( 
.A(n_491),
.B(n_388),
.Y(n_548)
);

NAND2xp5_ASAP7_75t_SL g549 ( 
.A(n_507),
.B(n_452),
.Y(n_549)
);

NAND2xp33_ASAP7_75t_L g550 ( 
.A(n_511),
.B(n_454),
.Y(n_550)
);

AND2x6_ASAP7_75t_L g551 ( 
.A(n_491),
.B(n_218),
.Y(n_551)
);

AND2x2_ASAP7_75t_SL g552 ( 
.A(n_507),
.B(n_372),
.Y(n_552)
);

NAND2xp5_ASAP7_75t_SL g553 ( 
.A(n_507),
.B(n_456),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_530),
.Y(n_554)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_530),
.Y(n_555)
);

INVx2_ASAP7_75t_L g556 ( 
.A(n_523),
.Y(n_556)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_494),
.Y(n_557)
);

NAND2xp33_ASAP7_75t_L g558 ( 
.A(n_513),
.B(n_516),
.Y(n_558)
);

AOI22xp33_ASAP7_75t_L g559 ( 
.A1(n_494),
.A2(n_438),
.B1(n_419),
.B2(n_349),
.Y(n_559)
);

NOR2xp33_ASAP7_75t_L g560 ( 
.A(n_493),
.B(n_423),
.Y(n_560)
);

INVx4_ASAP7_75t_L g561 ( 
.A(n_517),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_493),
.B(n_462),
.Y(n_562)
);

INVxp67_ASAP7_75t_SL g563 ( 
.A(n_495),
.Y(n_563)
);

NOR2xp33_ASAP7_75t_L g564 ( 
.A(n_499),
.B(n_448),
.Y(n_564)
);

INVx2_ASAP7_75t_SL g565 ( 
.A(n_519),
.Y(n_565)
);

BUFx6f_ASAP7_75t_L g566 ( 
.A(n_467),
.Y(n_566)
);

INVx1_ASAP7_75t_L g567 ( 
.A(n_498),
.Y(n_567)
);

INVx2_ASAP7_75t_L g568 ( 
.A(n_471),
.Y(n_568)
);

INVx1_ASAP7_75t_L g569 ( 
.A(n_498),
.Y(n_569)
);

BUFx2_ASAP7_75t_L g570 ( 
.A(n_520),
.Y(n_570)
);

NOR2xp33_ASAP7_75t_L g571 ( 
.A(n_499),
.B(n_393),
.Y(n_571)
);

INVx1_ASAP7_75t_SL g572 ( 
.A(n_489),
.Y(n_572)
);

INVxp67_ASAP7_75t_SL g573 ( 
.A(n_495),
.Y(n_573)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_512),
.Y(n_574)
);

NOR2xp33_ASAP7_75t_L g575 ( 
.A(n_515),
.B(n_464),
.Y(n_575)
);

NAND2xp33_ASAP7_75t_L g576 ( 
.A(n_522),
.B(n_186),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_515),
.B(n_429),
.Y(n_577)
);

INVx3_ASAP7_75t_L g578 ( 
.A(n_523),
.Y(n_578)
);

INVxp67_ASAP7_75t_L g579 ( 
.A(n_481),
.Y(n_579)
);

NAND2xp33_ASAP7_75t_L g580 ( 
.A(n_529),
.B(n_186),
.Y(n_580)
);

OR2x2_ASAP7_75t_L g581 ( 
.A(n_485),
.B(n_465),
.Y(n_581)
);

BUFx6f_ASAP7_75t_L g582 ( 
.A(n_467),
.Y(n_582)
);

INVx2_ASAP7_75t_L g583 ( 
.A(n_471),
.Y(n_583)
);

INVx1_ASAP7_75t_L g584 ( 
.A(n_512),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_525),
.Y(n_585)
);

NAND2xp5_ASAP7_75t_SL g586 ( 
.A(n_467),
.B(n_223),
.Y(n_586)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_525),
.Y(n_587)
);

INVx1_ASAP7_75t_L g588 ( 
.A(n_527),
.Y(n_588)
);

INVx1_ASAP7_75t_SL g589 ( 
.A(n_506),
.Y(n_589)
);

BUFx3_ASAP7_75t_L g590 ( 
.A(n_495),
.Y(n_590)
);

AND2x4_ASAP7_75t_L g591 ( 
.A(n_541),
.B(n_403),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g592 ( 
.A(n_467),
.B(n_227),
.Y(n_592)
);

NOR2xp33_ASAP7_75t_L g593 ( 
.A(n_541),
.B(n_465),
.Y(n_593)
);

BUFx3_ASAP7_75t_L g594 ( 
.A(n_500),
.Y(n_594)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_541),
.B(n_413),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_SL g596 ( 
.A1(n_483),
.A2(n_383),
.B1(n_413),
.B2(n_424),
.Y(n_596)
);

OAI22x1_ASAP7_75t_L g597 ( 
.A1(n_474),
.A2(n_435),
.B1(n_379),
.B2(n_394),
.Y(n_597)
);

INVx2_ASAP7_75t_SL g598 ( 
.A(n_537),
.Y(n_598)
);

INVx1_ASAP7_75t_SL g599 ( 
.A(n_474),
.Y(n_599)
);

INVx2_ASAP7_75t_L g600 ( 
.A(n_500),
.Y(n_600)
);

NOR2xp33_ASAP7_75t_L g601 ( 
.A(n_483),
.B(n_422),
.Y(n_601)
);

NAND2xp5_ASAP7_75t_L g602 ( 
.A(n_469),
.B(n_482),
.Y(n_602)
);

NOR2xp33_ASAP7_75t_L g603 ( 
.A(n_527),
.B(n_439),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_535),
.Y(n_604)
);

BUFx10_ASAP7_75t_L g605 ( 
.A(n_508),
.Y(n_605)
);

INVx2_ASAP7_75t_L g606 ( 
.A(n_500),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_535),
.Y(n_607)
);

BUFx3_ASAP7_75t_L g608 ( 
.A(n_502),
.Y(n_608)
);

NAND2x1p5_ASAP7_75t_L g609 ( 
.A(n_523),
.B(n_443),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_476),
.Y(n_610)
);

OR2x6_ASAP7_75t_L g611 ( 
.A(n_531),
.B(n_485),
.Y(n_611)
);

INVx1_ASAP7_75t_L g612 ( 
.A(n_532),
.Y(n_612)
);

AND2x2_ASAP7_75t_L g613 ( 
.A(n_501),
.B(n_449),
.Y(n_613)
);

NAND2xp5_ASAP7_75t_L g614 ( 
.A(n_469),
.B(n_443),
.Y(n_614)
);

INVx2_ASAP7_75t_L g615 ( 
.A(n_502),
.Y(n_615)
);

NAND2xp5_ASAP7_75t_L g616 ( 
.A(n_469),
.B(n_444),
.Y(n_616)
);

OR2x2_ASAP7_75t_L g617 ( 
.A(n_501),
.B(n_435),
.Y(n_617)
);

NAND2xp5_ASAP7_75t_SL g618 ( 
.A(n_467),
.B(n_478),
.Y(n_618)
);

INVx1_ASAP7_75t_L g619 ( 
.A(n_532),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_470),
.Y(n_620)
);

NAND2xp5_ASAP7_75t_L g621 ( 
.A(n_469),
.B(n_444),
.Y(n_621)
);

AOI22xp33_ASAP7_75t_L g622 ( 
.A1(n_514),
.A2(n_323),
.B1(n_309),
.B2(n_322),
.Y(n_622)
);

OAI22xp33_ASAP7_75t_L g623 ( 
.A1(n_539),
.A2(n_326),
.B1(n_307),
.B2(n_311),
.Y(n_623)
);

INVx1_ASAP7_75t_L g624 ( 
.A(n_470),
.Y(n_624)
);

OR2x2_ASAP7_75t_L g625 ( 
.A(n_531),
.B(n_540),
.Y(n_625)
);

NAND2xp5_ASAP7_75t_L g626 ( 
.A(n_482),
.B(n_445),
.Y(n_626)
);

OR2x6_ASAP7_75t_L g627 ( 
.A(n_505),
.B(n_445),
.Y(n_627)
);

NOR2xp33_ASAP7_75t_L g628 ( 
.A(n_482),
.B(n_457),
.Y(n_628)
);

NAND2xp33_ASAP7_75t_R g629 ( 
.A(n_542),
.B(n_457),
.Y(n_629)
);

INVx2_ASAP7_75t_SL g630 ( 
.A(n_466),
.Y(n_630)
);

BUFx4f_ASAP7_75t_L g631 ( 
.A(n_538),
.Y(n_631)
);

INVx2_ASAP7_75t_L g632 ( 
.A(n_502),
.Y(n_632)
);

NAND2xp5_ASAP7_75t_SL g633 ( 
.A(n_467),
.B(n_235),
.Y(n_633)
);

NAND2xp5_ASAP7_75t_L g634 ( 
.A(n_482),
.B(n_459),
.Y(n_634)
);

OR2x2_ASAP7_75t_L g635 ( 
.A(n_468),
.B(n_472),
.Y(n_635)
);

INVx6_ASAP7_75t_L g636 ( 
.A(n_523),
.Y(n_636)
);

NAND2xp33_ASAP7_75t_L g637 ( 
.A(n_480),
.B(n_187),
.Y(n_637)
);

NOR2xp33_ASAP7_75t_L g638 ( 
.A(n_505),
.B(n_528),
.Y(n_638)
);

NAND2xp5_ASAP7_75t_SL g639 ( 
.A(n_467),
.B(n_237),
.Y(n_639)
);

AND2x2_ASAP7_75t_L g640 ( 
.A(n_473),
.B(n_417),
.Y(n_640)
);

BUFx3_ASAP7_75t_L g641 ( 
.A(n_510),
.Y(n_641)
);

INVx1_ASAP7_75t_L g642 ( 
.A(n_475),
.Y(n_642)
);

NOR2xp33_ASAP7_75t_SL g643 ( 
.A(n_490),
.B(n_425),
.Y(n_643)
);

INVx2_ASAP7_75t_L g644 ( 
.A(n_510),
.Y(n_644)
);

INVx5_ASAP7_75t_L g645 ( 
.A(n_478),
.Y(n_645)
);

INVx4_ASAP7_75t_L g646 ( 
.A(n_478),
.Y(n_646)
);

OR2x2_ASAP7_75t_L g647 ( 
.A(n_496),
.B(n_459),
.Y(n_647)
);

NAND2xp5_ASAP7_75t_SL g648 ( 
.A(n_478),
.B(n_243),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_477),
.Y(n_649)
);

INVx2_ASAP7_75t_L g650 ( 
.A(n_510),
.Y(n_650)
);

NAND2xp5_ASAP7_75t_L g651 ( 
.A(n_514),
.B(n_460),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_478),
.Y(n_652)
);

AND2x2_ASAP7_75t_L g653 ( 
.A(n_497),
.B(n_427),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_477),
.Y(n_654)
);

INVx1_ASAP7_75t_SL g655 ( 
.A(n_503),
.Y(n_655)
);

NAND2xp5_ASAP7_75t_SL g656 ( 
.A(n_478),
.B(n_248),
.Y(n_656)
);

INVx1_ASAP7_75t_SL g657 ( 
.A(n_504),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_478),
.Y(n_658)
);

INVx1_ASAP7_75t_L g659 ( 
.A(n_479),
.Y(n_659)
);

AOI22xp5_ASAP7_75t_L g660 ( 
.A1(n_528),
.A2(n_293),
.B1(n_370),
.B2(n_297),
.Y(n_660)
);

NOR3xp33_ASAP7_75t_L g661 ( 
.A(n_543),
.B(n_226),
.C(n_216),
.Y(n_661)
);

NAND2xp5_ASAP7_75t_L g662 ( 
.A(n_514),
.B(n_460),
.Y(n_662)
);

NAND3xp33_ASAP7_75t_SL g663 ( 
.A(n_509),
.B(n_226),
.C(n_216),
.Y(n_663)
);

NAND2xp5_ASAP7_75t_L g664 ( 
.A(n_518),
.B(n_197),
.Y(n_664)
);

INVx4_ASAP7_75t_L g665 ( 
.A(n_523),
.Y(n_665)
);

HB1xp67_ASAP7_75t_L g666 ( 
.A(n_509),
.Y(n_666)
);

CKINVDCx16_ASAP7_75t_R g667 ( 
.A(n_523),
.Y(n_667)
);

NOR2xp33_ASAP7_75t_L g668 ( 
.A(n_518),
.B(n_395),
.Y(n_668)
);

INVx1_ASAP7_75t_L g669 ( 
.A(n_479),
.Y(n_669)
);

NAND2xp33_ASAP7_75t_L g670 ( 
.A(n_538),
.B(n_187),
.Y(n_670)
);

OR2x6_ASAP7_75t_L g671 ( 
.A(n_543),
.B(n_395),
.Y(n_671)
);

OR2x2_ASAP7_75t_L g672 ( 
.A(n_543),
.B(n_230),
.Y(n_672)
);

NAND2xp5_ASAP7_75t_SL g673 ( 
.A(n_538),
.B(n_249),
.Y(n_673)
);

OAI22xp33_ASAP7_75t_L g674 ( 
.A1(n_518),
.A2(n_337),
.B1(n_340),
.B2(n_341),
.Y(n_674)
);

INVx4_ASAP7_75t_SL g675 ( 
.A(n_538),
.Y(n_675)
);

INVx1_ASAP7_75t_L g676 ( 
.A(n_486),
.Y(n_676)
);

INVx3_ASAP7_75t_L g677 ( 
.A(n_538),
.Y(n_677)
);

INVx4_ASAP7_75t_SL g678 ( 
.A(n_538),
.Y(n_678)
);

NAND2xp5_ASAP7_75t_L g679 ( 
.A(n_524),
.B(n_217),
.Y(n_679)
);

INVx2_ASAP7_75t_L g680 ( 
.A(n_538),
.Y(n_680)
);

AOI22xp33_ASAP7_75t_L g681 ( 
.A1(n_524),
.A2(n_325),
.B1(n_328),
.B2(n_330),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_526),
.B(n_194),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_L g683 ( 
.A(n_486),
.B(n_200),
.Y(n_683)
);

AND2x2_ASAP7_75t_L g684 ( 
.A(n_526),
.B(n_433),
.Y(n_684)
);

NAND2xp5_ASAP7_75t_SL g685 ( 
.A(n_536),
.B(n_258),
.Y(n_685)
);

INVx1_ASAP7_75t_SL g686 ( 
.A(n_521),
.Y(n_686)
);

INVxp67_ASAP7_75t_L g687 ( 
.A(n_526),
.Y(n_687)
);

NOR2xp33_ASAP7_75t_L g688 ( 
.A(n_533),
.B(n_396),
.Y(n_688)
);

NAND2xp5_ASAP7_75t_SL g689 ( 
.A(n_533),
.B(n_271),
.Y(n_689)
);

INVx2_ASAP7_75t_SL g690 ( 
.A(n_521),
.Y(n_690)
);

INVx2_ASAP7_75t_SL g691 ( 
.A(n_536),
.Y(n_691)
);

BUFx3_ASAP7_75t_L g692 ( 
.A(n_533),
.Y(n_692)
);

AOI22xp33_ASAP7_75t_L g693 ( 
.A1(n_552),
.A2(n_536),
.B1(n_534),
.B2(n_484),
.Y(n_693)
);

OAI22xp5_ASAP7_75t_L g694 ( 
.A1(n_552),
.A2(n_331),
.B1(n_231),
.B2(n_230),
.Y(n_694)
);

OAI22xp33_ASAP7_75t_L g695 ( 
.A1(n_627),
.A2(n_352),
.B1(n_365),
.B2(n_333),
.Y(n_695)
);

NAND2xp5_ASAP7_75t_L g696 ( 
.A(n_638),
.B(n_534),
.Y(n_696)
);

AOI21xp5_ASAP7_75t_L g697 ( 
.A1(n_638),
.A2(n_484),
.B(n_487),
.Y(n_697)
);

NAND2xp5_ASAP7_75t_L g698 ( 
.A(n_560),
.B(n_534),
.Y(n_698)
);

INVx2_ASAP7_75t_L g699 ( 
.A(n_594),
.Y(n_699)
);

NAND2xp5_ASAP7_75t_L g700 ( 
.A(n_560),
.B(n_487),
.Y(n_700)
);

AND2x4_ASAP7_75t_L g701 ( 
.A(n_561),
.B(n_441),
.Y(n_701)
);

NAND2xp5_ASAP7_75t_L g702 ( 
.A(n_575),
.B(n_488),
.Y(n_702)
);

NOR2xp33_ASAP7_75t_SL g703 ( 
.A(n_561),
.B(n_635),
.Y(n_703)
);

NOR2x1p5_ASAP7_75t_L g704 ( 
.A(n_625),
.B(n_581),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_SL g705 ( 
.A(n_667),
.B(n_200),
.Y(n_705)
);

OAI21xp33_ASAP7_75t_L g706 ( 
.A1(n_577),
.A2(n_321),
.B(n_231),
.Y(n_706)
);

AND2x2_ASAP7_75t_L g707 ( 
.A(n_613),
.B(n_593),
.Y(n_707)
);

NAND2xp5_ASAP7_75t_SL g708 ( 
.A(n_562),
.B(n_204),
.Y(n_708)
);

AND2x6_ASAP7_75t_SL g709 ( 
.A(n_611),
.B(n_396),
.Y(n_709)
);

NAND2xp5_ASAP7_75t_L g710 ( 
.A(n_575),
.B(n_488),
.Y(n_710)
);

OAI22xp5_ASAP7_75t_SL g711 ( 
.A1(n_617),
.A2(n_453),
.B1(n_331),
.B2(n_321),
.Y(n_711)
);

NOR3xp33_ASAP7_75t_L g712 ( 
.A(n_549),
.B(n_340),
.C(n_337),
.Y(n_712)
);

INVx2_ASAP7_75t_L g713 ( 
.A(n_608),
.Y(n_713)
);

INVx2_ASAP7_75t_L g714 ( 
.A(n_641),
.Y(n_714)
);

NAND2xp5_ASAP7_75t_L g715 ( 
.A(n_577),
.B(n_492),
.Y(n_715)
);

AND2x2_ASAP7_75t_L g716 ( 
.A(n_593),
.B(n_397),
.Y(n_716)
);

NAND2xp5_ASAP7_75t_L g717 ( 
.A(n_612),
.B(n_492),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_L g718 ( 
.A(n_619),
.B(n_204),
.Y(n_718)
);

NOR2xp67_ASAP7_75t_L g719 ( 
.A(n_565),
.B(n_397),
.Y(n_719)
);

NAND2xp5_ASAP7_75t_L g720 ( 
.A(n_601),
.B(n_551),
.Y(n_720)
);

NOR2xp33_ASAP7_75t_L g721 ( 
.A(n_548),
.B(n_284),
.Y(n_721)
);

NAND2xp5_ASAP7_75t_L g722 ( 
.A(n_601),
.B(n_208),
.Y(n_722)
);

INVx2_ASAP7_75t_SL g723 ( 
.A(n_647),
.Y(n_723)
);

AND2x2_ASAP7_75t_L g724 ( 
.A(n_544),
.B(n_398),
.Y(n_724)
);

NAND3xp33_ASAP7_75t_L g725 ( 
.A(n_629),
.B(n_350),
.C(n_346),
.Y(n_725)
);

NAND3xp33_ASAP7_75t_L g726 ( 
.A(n_629),
.B(n_550),
.C(n_576),
.Y(n_726)
);

NAND2xp5_ASAP7_75t_L g727 ( 
.A(n_551),
.B(n_208),
.Y(n_727)
);

INVx2_ASAP7_75t_L g728 ( 
.A(n_641),
.Y(n_728)
);

INVx2_ASAP7_75t_L g729 ( 
.A(n_692),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_651),
.Y(n_730)
);

INVx2_ASAP7_75t_L g731 ( 
.A(n_590),
.Y(n_731)
);

OAI22xp5_ASAP7_75t_L g732 ( 
.A1(n_549),
.A2(n_350),
.B1(n_346),
.B2(n_367),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_662),
.Y(n_733)
);

INVx2_ASAP7_75t_L g734 ( 
.A(n_590),
.Y(n_734)
);

NOR2xp33_ASAP7_75t_L g735 ( 
.A(n_553),
.B(n_287),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_620),
.Y(n_736)
);

OR2x2_ASAP7_75t_L g737 ( 
.A(n_599),
.B(n_341),
.Y(n_737)
);

NAND2xp33_ASAP7_75t_L g738 ( 
.A(n_551),
.B(n_213),
.Y(n_738)
);

NAND2xp5_ASAP7_75t_L g739 ( 
.A(n_551),
.B(n_213),
.Y(n_739)
);

BUFx5_ASAP7_75t_L g740 ( 
.A(n_551),
.Y(n_740)
);

NAND2xp5_ASAP7_75t_L g741 ( 
.A(n_595),
.B(n_219),
.Y(n_741)
);

A2O1A1Ixp33_ASAP7_75t_L g742 ( 
.A1(n_595),
.A2(n_334),
.B(n_275),
.C(n_285),
.Y(n_742)
);

INVx5_ASAP7_75t_L g743 ( 
.A(n_566),
.Y(n_743)
);

NAND2xp5_ASAP7_75t_L g744 ( 
.A(n_591),
.B(n_219),
.Y(n_744)
);

NAND2xp5_ASAP7_75t_L g745 ( 
.A(n_591),
.B(n_220),
.Y(n_745)
);

O2A1O1Ixp5_ASAP7_75t_L g746 ( 
.A1(n_553),
.A2(n_360),
.B(n_317),
.C(n_313),
.Y(n_746)
);

INVx2_ASAP7_75t_L g747 ( 
.A(n_547),
.Y(n_747)
);

NAND2xp5_ASAP7_75t_L g748 ( 
.A(n_627),
.B(n_220),
.Y(n_748)
);

NOR2xp33_ASAP7_75t_L g749 ( 
.A(n_564),
.B(n_302),
.Y(n_749)
);

INVx1_ASAP7_75t_L g750 ( 
.A(n_624),
.Y(n_750)
);

OAI22xp5_ASAP7_75t_L g751 ( 
.A1(n_564),
.A2(n_355),
.B1(n_343),
.B2(n_367),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_570),
.Y(n_752)
);

NAND2xp5_ASAP7_75t_L g753 ( 
.A(n_627),
.B(n_221),
.Y(n_753)
);

INVx2_ASAP7_75t_SL g754 ( 
.A(n_684),
.Y(n_754)
);

INVxp67_ASAP7_75t_L g755 ( 
.A(n_572),
.Y(n_755)
);

OAI22xp5_ASAP7_75t_L g756 ( 
.A1(n_579),
.A2(n_366),
.B1(n_343),
.B2(n_355),
.Y(n_756)
);

NAND2xp5_ASAP7_75t_L g757 ( 
.A(n_571),
.B(n_221),
.Y(n_757)
);

NOR2xp33_ASAP7_75t_L g758 ( 
.A(n_571),
.B(n_308),
.Y(n_758)
);

BUFx6f_ASAP7_75t_L g759 ( 
.A(n_566),
.Y(n_759)
);

NOR2xp33_ASAP7_75t_R g760 ( 
.A(n_558),
.B(n_605),
.Y(n_760)
);

BUFx6f_ASAP7_75t_L g761 ( 
.A(n_566),
.Y(n_761)
);

NAND2xp5_ASAP7_75t_L g762 ( 
.A(n_628),
.B(n_225),
.Y(n_762)
);

HB1xp67_ASAP7_75t_L g763 ( 
.A(n_611),
.Y(n_763)
);

NAND2xp5_ASAP7_75t_L g764 ( 
.A(n_628),
.B(n_225),
.Y(n_764)
);

AOI22xp33_ASAP7_75t_L g765 ( 
.A1(n_622),
.A2(n_484),
.B1(n_354),
.B2(n_398),
.Y(n_765)
);

HB1xp67_ASAP7_75t_L g766 ( 
.A(n_611),
.Y(n_766)
);

INVx2_ASAP7_75t_SL g767 ( 
.A(n_589),
.Y(n_767)
);

CKINVDCx5p33_ASAP7_75t_R g768 ( 
.A(n_605),
.Y(n_768)
);

AND2x4_ASAP7_75t_L g769 ( 
.A(n_690),
.B(n_407),
.Y(n_769)
);

NAND2xp5_ASAP7_75t_L g770 ( 
.A(n_603),
.B(n_228),
.Y(n_770)
);

BUFx5_ASAP7_75t_L g771 ( 
.A(n_545),
.Y(n_771)
);

NAND2xp5_ASAP7_75t_SL g772 ( 
.A(n_566),
.B(n_582),
.Y(n_772)
);

NAND2xp5_ASAP7_75t_SL g773 ( 
.A(n_582),
.B(n_598),
.Y(n_773)
);

NAND2xp5_ASAP7_75t_L g774 ( 
.A(n_603),
.B(n_228),
.Y(n_774)
);

BUFx5_ASAP7_75t_L g775 ( 
.A(n_554),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_642),
.Y(n_776)
);

HB1xp67_ASAP7_75t_L g777 ( 
.A(n_666),
.Y(n_777)
);

INVx1_ASAP7_75t_L g778 ( 
.A(n_649),
.Y(n_778)
);

INVx1_ASAP7_75t_SL g779 ( 
.A(n_655),
.Y(n_779)
);

INVxp67_ASAP7_75t_SL g780 ( 
.A(n_563),
.Y(n_780)
);

AND2x2_ASAP7_75t_L g781 ( 
.A(n_630),
.B(n_407),
.Y(n_781)
);

NAND2xp5_ASAP7_75t_L g782 ( 
.A(n_687),
.B(n_229),
.Y(n_782)
);

NAND2xp5_ASAP7_75t_L g783 ( 
.A(n_557),
.B(n_229),
.Y(n_783)
);

INVx2_ASAP7_75t_SL g784 ( 
.A(n_672),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_568),
.Y(n_785)
);

A2O1A1Ixp33_ASAP7_75t_L g786 ( 
.A1(n_668),
.A2(n_366),
.B(n_298),
.C(n_305),
.Y(n_786)
);

INVx1_ASAP7_75t_SL g787 ( 
.A(n_657),
.Y(n_787)
);

INVx2_ASAP7_75t_L g788 ( 
.A(n_568),
.Y(n_788)
);

OAI22xp5_ASAP7_75t_L g789 ( 
.A1(n_559),
.A2(n_310),
.B1(n_312),
.B2(n_314),
.Y(n_789)
);

NOR2xp33_ASAP7_75t_L g790 ( 
.A(n_567),
.B(n_316),
.Y(n_790)
);

AOI22xp5_ASAP7_75t_L g791 ( 
.A1(n_683),
.A2(n_580),
.B1(n_559),
.B2(n_661),
.Y(n_791)
);

NAND2xp5_ASAP7_75t_L g792 ( 
.A(n_569),
.B(n_574),
.Y(n_792)
);

NAND2xp5_ASAP7_75t_L g793 ( 
.A(n_584),
.B(n_316),
.Y(n_793)
);

AOI22xp5_ASAP7_75t_L g794 ( 
.A1(n_691),
.A2(n_347),
.B1(n_368),
.B2(n_320),
.Y(n_794)
);

INVx1_ASAP7_75t_L g795 ( 
.A(n_654),
.Y(n_795)
);

INVx2_ASAP7_75t_L g796 ( 
.A(n_583),
.Y(n_796)
);

OAI22xp5_ASAP7_75t_L g797 ( 
.A1(n_585),
.A2(n_347),
.B1(n_368),
.B2(n_320),
.Y(n_797)
);

NAND2xp5_ASAP7_75t_L g798 ( 
.A(n_587),
.B(n_327),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_SL g799 ( 
.A(n_582),
.B(n_327),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_588),
.B(n_336),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_604),
.B(n_336),
.Y(n_801)
);

NOR2xp33_ASAP7_75t_L g802 ( 
.A(n_607),
.B(n_338),
.Y(n_802)
);

BUFx6f_ASAP7_75t_L g803 ( 
.A(n_582),
.Y(n_803)
);

AND2x2_ASAP7_75t_SL g804 ( 
.A(n_622),
.B(n_484),
.Y(n_804)
);

A2O1A1Ixp33_ASAP7_75t_L g805 ( 
.A1(n_659),
.A2(n_278),
.B(n_364),
.C(n_362),
.Y(n_805)
);

INVx3_ASAP7_75t_L g806 ( 
.A(n_609),
.Y(n_806)
);

CKINVDCx14_ASAP7_75t_R g807 ( 
.A(n_610),
.Y(n_807)
);

AOI22xp33_ASAP7_75t_L g808 ( 
.A1(n_681),
.A2(n_484),
.B1(n_290),
.B2(n_299),
.Y(n_808)
);

AOI22xp33_ASAP7_75t_L g809 ( 
.A1(n_681),
.A2(n_335),
.B1(n_351),
.B2(n_269),
.Y(n_809)
);

NAND2xp5_ASAP7_75t_L g810 ( 
.A(n_664),
.B(n_338),
.Y(n_810)
);

NAND2xp5_ASAP7_75t_L g811 ( 
.A(n_679),
.B(n_344),
.Y(n_811)
);

NAND2xp5_ASAP7_75t_SL g812 ( 
.A(n_646),
.B(n_344),
.Y(n_812)
);

INVx2_ASAP7_75t_L g813 ( 
.A(n_583),
.Y(n_813)
);

NOR2xp33_ASAP7_75t_L g814 ( 
.A(n_555),
.B(n_348),
.Y(n_814)
);

NAND2xp33_ASAP7_75t_L g815 ( 
.A(n_602),
.B(n_348),
.Y(n_815)
);

INVx1_ASAP7_75t_L g816 ( 
.A(n_669),
.Y(n_816)
);

NAND2xp5_ASAP7_75t_L g817 ( 
.A(n_573),
.B(n_356),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_L g818 ( 
.A(n_671),
.B(n_356),
.Y(n_818)
);

INVxp67_ASAP7_75t_L g819 ( 
.A(n_643),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_676),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_671),
.Y(n_821)
);

NAND2xp5_ASAP7_75t_L g822 ( 
.A(n_671),
.B(n_614),
.Y(n_822)
);

NAND2xp5_ASAP7_75t_L g823 ( 
.A(n_616),
.B(n_359),
.Y(n_823)
);

BUFx6f_ASAP7_75t_L g824 ( 
.A(n_646),
.Y(n_824)
);

NAND2xp5_ASAP7_75t_SL g825 ( 
.A(n_631),
.B(n_359),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_631),
.B(n_361),
.Y(n_826)
);

NAND2xp5_ASAP7_75t_SL g827 ( 
.A(n_665),
.B(n_361),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_621),
.Y(n_828)
);

NAND2xp5_ASAP7_75t_L g829 ( 
.A(n_626),
.B(n_233),
.Y(n_829)
);

INVx2_ASAP7_75t_L g830 ( 
.A(n_600),
.Y(n_830)
);

NOR2xp67_ASAP7_75t_L g831 ( 
.A(n_663),
.B(n_640),
.Y(n_831)
);

INVx3_ASAP7_75t_L g832 ( 
.A(n_609),
.Y(n_832)
);

NAND2xp5_ASAP7_75t_L g833 ( 
.A(n_634),
.B(n_238),
.Y(n_833)
);

NOR2xp67_ASAP7_75t_L g834 ( 
.A(n_660),
.B(n_239),
.Y(n_834)
);

INVx2_ASAP7_75t_L g835 ( 
.A(n_600),
.Y(n_835)
);

INVxp67_ASAP7_75t_L g836 ( 
.A(n_653),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_668),
.Y(n_837)
);

AND2x2_ASAP7_75t_L g838 ( 
.A(n_610),
.B(n_6),
.Y(n_838)
);

NAND2xp5_ASAP7_75t_L g839 ( 
.A(n_682),
.B(n_252),
.Y(n_839)
);

NAND2xp5_ASAP7_75t_L g840 ( 
.A(n_606),
.B(n_257),
.Y(n_840)
);

INVx8_ASAP7_75t_L g841 ( 
.A(n_645),
.Y(n_841)
);

AND2x6_ASAP7_75t_SL g842 ( 
.A(n_688),
.B(n_7),
.Y(n_842)
);

INVx2_ASAP7_75t_SL g843 ( 
.A(n_686),
.Y(n_843)
);

BUFx6f_ASAP7_75t_L g844 ( 
.A(n_636),
.Y(n_844)
);

NAND2xp5_ASAP7_75t_L g845 ( 
.A(n_606),
.B(n_281),
.Y(n_845)
);

NAND2xp5_ASAP7_75t_L g846 ( 
.A(n_615),
.B(n_272),
.Y(n_846)
);

AOI22xp33_ASAP7_75t_L g847 ( 
.A1(n_623),
.A2(n_674),
.B1(n_688),
.B2(n_632),
.Y(n_847)
);

A2O1A1Ixp33_ASAP7_75t_L g848 ( 
.A1(n_615),
.A2(n_259),
.B(n_264),
.C(n_265),
.Y(n_848)
);

NOR2xp33_ASAP7_75t_L g849 ( 
.A(n_665),
.B(n_7),
.Y(n_849)
);

INVx2_ASAP7_75t_L g850 ( 
.A(n_632),
.Y(n_850)
);

INVx2_ASAP7_75t_SL g851 ( 
.A(n_685),
.Y(n_851)
);

INVx2_ASAP7_75t_SL g852 ( 
.A(n_685),
.Y(n_852)
);

INVx2_ASAP7_75t_L g853 ( 
.A(n_644),
.Y(n_853)
);

O2A1O1Ixp33_ASAP7_75t_L g854 ( 
.A1(n_674),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_854)
);

INVx1_ASAP7_75t_L g855 ( 
.A(n_644),
.Y(n_855)
);

AND2x2_ASAP7_75t_L g856 ( 
.A(n_637),
.B(n_11),
.Y(n_856)
);

NAND2xp5_ASAP7_75t_L g857 ( 
.A(n_749),
.B(n_650),
.Y(n_857)
);

AOI21xp5_ASAP7_75t_L g858 ( 
.A1(n_696),
.A2(n_618),
.B(n_652),
.Y(n_858)
);

AOI21xp5_ASAP7_75t_L g859 ( 
.A1(n_698),
.A2(n_618),
.B(n_652),
.Y(n_859)
);

AOI21xp5_ASAP7_75t_L g860 ( 
.A1(n_772),
.A2(n_658),
.B(n_578),
.Y(n_860)
);

AOI21xp5_ASAP7_75t_L g861 ( 
.A1(n_772),
.A2(n_658),
.B(n_578),
.Y(n_861)
);

AND2x2_ASAP7_75t_L g862 ( 
.A(n_707),
.B(n_597),
.Y(n_862)
);

OAI21x1_ASAP7_75t_L g863 ( 
.A1(n_697),
.A2(n_680),
.B(n_650),
.Y(n_863)
);

NAND2xp5_ASAP7_75t_L g864 ( 
.A(n_749),
.B(n_715),
.Y(n_864)
);

AND2x4_ASAP7_75t_L g865 ( 
.A(n_769),
.B(n_843),
.Y(n_865)
);

AOI21xp5_ASAP7_75t_L g866 ( 
.A1(n_702),
.A2(n_677),
.B(n_670),
.Y(n_866)
);

OAI22xp5_ASAP7_75t_L g867 ( 
.A1(n_720),
.A2(n_710),
.B1(n_837),
.B2(n_700),
.Y(n_867)
);

OR2x2_ASAP7_75t_L g868 ( 
.A(n_723),
.B(n_623),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_736),
.Y(n_869)
);

A2O1A1Ixp33_ASAP7_75t_L g870 ( 
.A1(n_758),
.A2(n_689),
.B(n_680),
.C(n_677),
.Y(n_870)
);

OAI21xp5_ASAP7_75t_L g871 ( 
.A1(n_693),
.A2(n_556),
.B(n_546),
.Y(n_871)
);

NAND2xp5_ASAP7_75t_L g872 ( 
.A(n_758),
.B(n_596),
.Y(n_872)
);

AOI21xp5_ASAP7_75t_L g873 ( 
.A1(n_717),
.A2(n_645),
.B(n_586),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_750),
.Y(n_874)
);

NAND2xp5_ASAP7_75t_L g875 ( 
.A(n_722),
.B(n_689),
.Y(n_875)
);

NAND2xp5_ASAP7_75t_L g876 ( 
.A(n_721),
.B(n_645),
.Y(n_876)
);

AOI21xp5_ASAP7_75t_L g877 ( 
.A1(n_780),
.A2(n_645),
.B(n_586),
.Y(n_877)
);

OAI21xp5_ASAP7_75t_L g878 ( 
.A1(n_693),
.A2(n_592),
.B(n_633),
.Y(n_878)
);

OAI21xp5_ASAP7_75t_L g879 ( 
.A1(n_828),
.A2(n_592),
.B(n_633),
.Y(n_879)
);

AOI21x1_ASAP7_75t_L g880 ( 
.A1(n_855),
.A2(n_656),
.B(n_648),
.Y(n_880)
);

NAND2xp5_ASAP7_75t_L g881 ( 
.A(n_721),
.B(n_636),
.Y(n_881)
);

NAND2xp5_ASAP7_75t_SL g882 ( 
.A(n_740),
.B(n_675),
.Y(n_882)
);

A2O1A1Ixp33_ASAP7_75t_L g883 ( 
.A1(n_735),
.A2(n_673),
.B(n_656),
.C(n_648),
.Y(n_883)
);

O2A1O1Ixp33_ASAP7_75t_L g884 ( 
.A1(n_694),
.A2(n_673),
.B(n_639),
.C(n_19),
.Y(n_884)
);

AOI21xp5_ASAP7_75t_L g885 ( 
.A1(n_780),
.A2(n_639),
.B(n_267),
.Y(n_885)
);

INVxp67_ASAP7_75t_L g886 ( 
.A(n_767),
.Y(n_886)
);

OAI22xp5_ASAP7_75t_L g887 ( 
.A1(n_791),
.A2(n_636),
.B1(n_291),
.B2(n_295),
.Y(n_887)
);

NAND2xp5_ASAP7_75t_L g888 ( 
.A(n_716),
.B(n_678),
.Y(n_888)
);

AOI21xp5_ASAP7_75t_L g889 ( 
.A1(n_792),
.A2(n_315),
.B(n_303),
.Y(n_889)
);

OAI22xp5_ASAP7_75t_L g890 ( 
.A1(n_770),
.A2(n_282),
.B1(n_16),
.B2(n_20),
.Y(n_890)
);

INVx3_ASAP7_75t_L g891 ( 
.A(n_841),
.Y(n_891)
);

OAI21xp33_ASAP7_75t_L g892 ( 
.A1(n_774),
.A2(n_15),
.B(n_22),
.Y(n_892)
);

INVxp67_ASAP7_75t_SL g893 ( 
.A(n_759),
.Y(n_893)
);

AO21x1_ASAP7_75t_L g894 ( 
.A1(n_735),
.A2(n_678),
.B(n_675),
.Y(n_894)
);

O2A1O1Ixp33_ASAP7_75t_L g895 ( 
.A1(n_706),
.A2(n_751),
.B(n_786),
.C(n_741),
.Y(n_895)
);

NAND2xp5_ASAP7_75t_SL g896 ( 
.A(n_740),
.B(n_678),
.Y(n_896)
);

NAND2xp5_ASAP7_75t_L g897 ( 
.A(n_769),
.B(n_675),
.Y(n_897)
);

O2A1O1Ixp33_ASAP7_75t_L g898 ( 
.A1(n_786),
.A2(n_15),
.B(n_25),
.C(n_27),
.Y(n_898)
);

AOI21xp33_ASAP7_75t_L g899 ( 
.A1(n_757),
.A2(n_25),
.B(n_27),
.Y(n_899)
);

NAND2x1p5_ASAP7_75t_L g900 ( 
.A(n_806),
.B(n_82),
.Y(n_900)
);

AOI21xp5_ASAP7_75t_L g901 ( 
.A1(n_839),
.A2(n_826),
.B(n_825),
.Y(n_901)
);

NOR2xp33_ASAP7_75t_L g902 ( 
.A(n_754),
.B(n_28),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_729),
.Y(n_903)
);

NAND2xp5_ASAP7_75t_SL g904 ( 
.A(n_740),
.B(n_324),
.Y(n_904)
);

NAND2xp5_ASAP7_75t_L g905 ( 
.A(n_730),
.B(n_28),
.Y(n_905)
);

NOR2xp33_ASAP7_75t_SL g906 ( 
.A(n_779),
.B(n_324),
.Y(n_906)
);

NAND2xp5_ASAP7_75t_L g907 ( 
.A(n_733),
.B(n_29),
.Y(n_907)
);

AND2x2_ASAP7_75t_L g908 ( 
.A(n_787),
.B(n_31),
.Y(n_908)
);

NAND2xp5_ASAP7_75t_L g909 ( 
.A(n_847),
.B(n_32),
.Y(n_909)
);

NAND2xp5_ASAP7_75t_L g910 ( 
.A(n_847),
.B(n_32),
.Y(n_910)
);

NAND2xp5_ASAP7_75t_SL g911 ( 
.A(n_740),
.B(n_324),
.Y(n_911)
);

AOI21xp5_ASAP7_75t_L g912 ( 
.A1(n_773),
.A2(n_324),
.B(n_269),
.Y(n_912)
);

NAND2xp5_ASAP7_75t_L g913 ( 
.A(n_724),
.B(n_38),
.Y(n_913)
);

NAND2xp5_ASAP7_75t_L g914 ( 
.A(n_718),
.B(n_39),
.Y(n_914)
);

AOI33xp33_ASAP7_75t_L g915 ( 
.A1(n_695),
.A2(n_42),
.A3(n_46),
.B1(n_47),
.B2(n_48),
.B3(n_49),
.Y(n_915)
);

AOI21xp5_ASAP7_75t_L g916 ( 
.A1(n_773),
.A2(n_324),
.B(n_123),
.Y(n_916)
);

NAND2xp5_ASAP7_75t_SL g917 ( 
.A(n_740),
.B(n_50),
.Y(n_917)
);

HB1xp67_ASAP7_75t_L g918 ( 
.A(n_763),
.Y(n_918)
);

INVx4_ASAP7_75t_L g919 ( 
.A(n_841),
.Y(n_919)
);

AOI21xp5_ASAP7_75t_L g920 ( 
.A1(n_812),
.A2(n_116),
.B(n_161),
.Y(n_920)
);

NAND2xp5_ASAP7_75t_L g921 ( 
.A(n_790),
.B(n_50),
.Y(n_921)
);

AOI21xp5_ASAP7_75t_L g922 ( 
.A1(n_812),
.A2(n_817),
.B(n_827),
.Y(n_922)
);

AOI21xp5_ASAP7_75t_L g923 ( 
.A1(n_827),
.A2(n_102),
.B(n_156),
.Y(n_923)
);

NOR2xp33_ASAP7_75t_L g924 ( 
.A(n_703),
.B(n_56),
.Y(n_924)
);

INVx3_ASAP7_75t_L g925 ( 
.A(n_841),
.Y(n_925)
);

OAI21x1_ASAP7_75t_L g926 ( 
.A1(n_747),
.A2(n_128),
.B(n_155),
.Y(n_926)
);

AOI22xp5_ASAP7_75t_L g927 ( 
.A1(n_726),
.A2(n_58),
.B1(n_59),
.B2(n_60),
.Y(n_927)
);

AND2x2_ASAP7_75t_L g928 ( 
.A(n_704),
.B(n_60),
.Y(n_928)
);

OAI21xp5_ASAP7_75t_L g929 ( 
.A1(n_822),
.A2(n_68),
.B(n_71),
.Y(n_929)
);

NAND3xp33_ASAP7_75t_SL g930 ( 
.A(n_752),
.B(n_77),
.C(n_78),
.Y(n_930)
);

AND2x4_ASAP7_75t_L g931 ( 
.A(n_763),
.B(n_87),
.Y(n_931)
);

INVx2_ASAP7_75t_L g932 ( 
.A(n_699),
.Y(n_932)
);

NAND2xp5_ASAP7_75t_L g933 ( 
.A(n_790),
.B(n_88),
.Y(n_933)
);

AOI21xp5_ASAP7_75t_L g934 ( 
.A1(n_829),
.A2(n_98),
.B(n_134),
.Y(n_934)
);

NAND2x1p5_ASAP7_75t_L g935 ( 
.A(n_806),
.B(n_138),
.Y(n_935)
);

O2A1O1Ixp33_ASAP7_75t_L g936 ( 
.A1(n_732),
.A2(n_141),
.B(n_143),
.C(n_144),
.Y(n_936)
);

AOI21xp5_ASAP7_75t_L g937 ( 
.A1(n_833),
.A2(n_153),
.B(n_154),
.Y(n_937)
);

O2A1O1Ixp33_ASAP7_75t_L g938 ( 
.A1(n_789),
.A2(n_179),
.B(n_712),
.C(n_742),
.Y(n_938)
);

NAND2xp5_ASAP7_75t_L g939 ( 
.A(n_802),
.B(n_784),
.Y(n_939)
);

AOI21xp5_ASAP7_75t_L g940 ( 
.A1(n_738),
.A2(n_708),
.B(n_764),
.Y(n_940)
);

AOI21xp5_ASAP7_75t_L g941 ( 
.A1(n_708),
.A2(n_762),
.B(n_799),
.Y(n_941)
);

NAND2xp5_ASAP7_75t_L g942 ( 
.A(n_802),
.B(n_781),
.Y(n_942)
);

INVx3_ASAP7_75t_L g943 ( 
.A(n_844),
.Y(n_943)
);

BUFx3_ASAP7_75t_L g944 ( 
.A(n_768),
.Y(n_944)
);

AOI21xp5_ASAP7_75t_L g945 ( 
.A1(n_799),
.A2(n_823),
.B(n_782),
.Y(n_945)
);

AOI21xp5_ASAP7_75t_L g946 ( 
.A1(n_824),
.A2(n_820),
.B(n_778),
.Y(n_946)
);

NAND2xp5_ASAP7_75t_L g947 ( 
.A(n_776),
.B(n_795),
.Y(n_947)
);

O2A1O1Ixp33_ASAP7_75t_L g948 ( 
.A1(n_712),
.A2(n_695),
.B(n_854),
.C(n_816),
.Y(n_948)
);

NOR2xp33_ASAP7_75t_L g949 ( 
.A(n_836),
.B(n_819),
.Y(n_949)
);

AOI21xp5_ASAP7_75t_L g950 ( 
.A1(n_824),
.A2(n_815),
.B(n_793),
.Y(n_950)
);

OAI21xp5_ASAP7_75t_L g951 ( 
.A1(n_727),
.A2(n_739),
.B(n_746),
.Y(n_951)
);

NAND2xp5_ASAP7_75t_L g952 ( 
.A(n_851),
.B(n_852),
.Y(n_952)
);

AOI21xp5_ASAP7_75t_L g953 ( 
.A1(n_824),
.A2(n_783),
.B(n_798),
.Y(n_953)
);

OAI321xp33_ASAP7_75t_L g954 ( 
.A1(n_809),
.A2(n_711),
.A3(n_856),
.B1(n_756),
.B2(n_725),
.C(n_836),
.Y(n_954)
);

AOI21xp5_ASAP7_75t_L g955 ( 
.A1(n_824),
.A2(n_801),
.B(n_800),
.Y(n_955)
);

CKINVDCx10_ASAP7_75t_R g956 ( 
.A(n_807),
.Y(n_956)
);

BUFx8_ASAP7_75t_L g957 ( 
.A(n_701),
.Y(n_957)
);

AOI21xp5_ASAP7_75t_L g958 ( 
.A1(n_840),
.A2(n_846),
.B(n_845),
.Y(n_958)
);

AND2x2_ASAP7_75t_L g959 ( 
.A(n_819),
.B(n_766),
.Y(n_959)
);

INVx2_ASAP7_75t_SL g960 ( 
.A(n_766),
.Y(n_960)
);

NAND2xp5_ASAP7_75t_L g961 ( 
.A(n_810),
.B(n_811),
.Y(n_961)
);

CKINVDCx10_ASAP7_75t_R g962 ( 
.A(n_842),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_821),
.Y(n_963)
);

NAND2xp5_ASAP7_75t_L g964 ( 
.A(n_744),
.B(n_745),
.Y(n_964)
);

INVx2_ASAP7_75t_L g965 ( 
.A(n_785),
.Y(n_965)
);

AOI21xp5_ASAP7_75t_L g966 ( 
.A1(n_759),
.A2(n_803),
.B(n_761),
.Y(n_966)
);

AOI21xp5_ASAP7_75t_L g967 ( 
.A1(n_759),
.A2(n_803),
.B(n_761),
.Y(n_967)
);

NAND2xp5_ASAP7_75t_SL g968 ( 
.A(n_740),
.B(n_771),
.Y(n_968)
);

O2A1O1Ixp33_ASAP7_75t_L g969 ( 
.A1(n_848),
.A2(n_797),
.B(n_753),
.C(n_748),
.Y(n_969)
);

NOR2x1p5_ASAP7_75t_L g970 ( 
.A(n_701),
.B(n_737),
.Y(n_970)
);

AOI21xp5_ASAP7_75t_L g971 ( 
.A1(n_759),
.A2(n_803),
.B(n_761),
.Y(n_971)
);

INVx2_ASAP7_75t_L g972 ( 
.A(n_713),
.Y(n_972)
);

AND2x2_ASAP7_75t_L g973 ( 
.A(n_755),
.B(n_777),
.Y(n_973)
);

HB1xp67_ASAP7_75t_L g974 ( 
.A(n_777),
.Y(n_974)
);

AO22x1_ASAP7_75t_L g975 ( 
.A1(n_755),
.A2(n_838),
.B1(n_818),
.B2(n_709),
.Y(n_975)
);

NAND2xp5_ASAP7_75t_SL g976 ( 
.A(n_771),
.B(n_775),
.Y(n_976)
);

AOI21xp5_ASAP7_75t_L g977 ( 
.A1(n_761),
.A2(n_803),
.B(n_796),
.Y(n_977)
);

NOR3xp33_ASAP7_75t_L g978 ( 
.A(n_831),
.B(n_719),
.C(n_805),
.Y(n_978)
);

BUFx3_ASAP7_75t_L g979 ( 
.A(n_844),
.Y(n_979)
);

A2O1A1Ixp33_ASAP7_75t_L g980 ( 
.A1(n_849),
.A2(n_814),
.B(n_809),
.C(n_834),
.Y(n_980)
);

INVx1_ASAP7_75t_SL g981 ( 
.A(n_760),
.Y(n_981)
);

O2A1O1Ixp33_ASAP7_75t_L g982 ( 
.A1(n_848),
.A2(n_705),
.B(n_814),
.C(n_849),
.Y(n_982)
);

AOI21xp5_ASAP7_75t_L g983 ( 
.A1(n_788),
.A2(n_853),
.B(n_830),
.Y(n_983)
);

NAND2xp33_ASAP7_75t_L g984 ( 
.A(n_760),
.B(n_775),
.Y(n_984)
);

AOI21xp5_ASAP7_75t_L g985 ( 
.A1(n_813),
.A2(n_850),
.B(n_835),
.Y(n_985)
);

INVxp67_ASAP7_75t_L g986 ( 
.A(n_705),
.Y(n_986)
);

AOI21xp5_ASAP7_75t_L g987 ( 
.A1(n_731),
.A2(n_734),
.B(n_728),
.Y(n_987)
);

OAI22xp5_ASAP7_75t_L g988 ( 
.A1(n_808),
.A2(n_832),
.B1(n_804),
.B2(n_765),
.Y(n_988)
);

NAND2xp5_ASAP7_75t_L g989 ( 
.A(n_714),
.B(n_765),
.Y(n_989)
);

AOI21xp5_ASAP7_75t_L g990 ( 
.A1(n_743),
.A2(n_832),
.B(n_844),
.Y(n_990)
);

INVx4_ASAP7_75t_L g991 ( 
.A(n_743),
.Y(n_991)
);

INVx1_ASAP7_75t_L g992 ( 
.A(n_844),
.Y(n_992)
);

OAI22xp5_ASAP7_75t_L g993 ( 
.A1(n_808),
.A2(n_804),
.B1(n_743),
.B2(n_794),
.Y(n_993)
);

AOI21xp5_ASAP7_75t_L g994 ( 
.A1(n_743),
.A2(n_771),
.B(n_775),
.Y(n_994)
);

NAND2xp5_ASAP7_75t_L g995 ( 
.A(n_771),
.B(n_775),
.Y(n_995)
);

NAND2xp5_ASAP7_75t_L g996 ( 
.A(n_771),
.B(n_775),
.Y(n_996)
);

INVx2_ASAP7_75t_L g997 ( 
.A(n_771),
.Y(n_997)
);

NAND3xp33_ASAP7_75t_L g998 ( 
.A(n_775),
.B(n_749),
.C(n_560),
.Y(n_998)
);

NOR2xp67_ASAP7_75t_L g999 ( 
.A(n_768),
.B(n_561),
.Y(n_999)
);

NAND2xp5_ASAP7_75t_SL g1000 ( 
.A(n_740),
.B(n_720),
.Y(n_1000)
);

AOI21xp5_ASAP7_75t_L g1001 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1001)
);

AOI21xp5_ASAP7_75t_L g1002 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1002)
);

INVxp67_ASAP7_75t_L g1003 ( 
.A(n_767),
.Y(n_1003)
);

AOI21xp5_ASAP7_75t_L g1004 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1004)
);

NAND2xp5_ASAP7_75t_L g1005 ( 
.A(n_749),
.B(n_638),
.Y(n_1005)
);

AOI21xp5_ASAP7_75t_L g1006 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1006)
);

NAND2x1p5_ASAP7_75t_L g1007 ( 
.A(n_806),
.B(n_832),
.Y(n_1007)
);

OAI22xp5_ASAP7_75t_L g1008 ( 
.A1(n_720),
.A2(n_552),
.B1(n_749),
.B2(n_710),
.Y(n_1008)
);

NAND2xp5_ASAP7_75t_L g1009 ( 
.A(n_749),
.B(n_638),
.Y(n_1009)
);

A2O1A1Ixp33_ASAP7_75t_L g1010 ( 
.A1(n_749),
.A2(n_720),
.B(n_758),
.C(n_638),
.Y(n_1010)
);

AND2x2_ASAP7_75t_L g1011 ( 
.A(n_707),
.B(n_544),
.Y(n_1011)
);

HB1xp67_ASAP7_75t_L g1012 ( 
.A(n_763),
.Y(n_1012)
);

AND2x4_ASAP7_75t_L g1013 ( 
.A(n_769),
.B(n_561),
.Y(n_1013)
);

OAI22x1_ASAP7_75t_L g1014 ( 
.A1(n_749),
.A2(n_704),
.B1(n_791),
.B2(n_766),
.Y(n_1014)
);

NAND2xp5_ASAP7_75t_L g1015 ( 
.A(n_749),
.B(n_638),
.Y(n_1015)
);

OR2x2_ASAP7_75t_L g1016 ( 
.A(n_723),
.B(n_572),
.Y(n_1016)
);

OAI22xp5_ASAP7_75t_L g1017 ( 
.A1(n_720),
.A2(n_552),
.B1(n_749),
.B2(n_710),
.Y(n_1017)
);

AOI21xp5_ASAP7_75t_L g1018 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1018)
);

OAI21xp5_ASAP7_75t_L g1019 ( 
.A1(n_697),
.A2(n_696),
.B(n_698),
.Y(n_1019)
);

OAI21x1_ASAP7_75t_L g1020 ( 
.A1(n_697),
.A2(n_693),
.B(n_658),
.Y(n_1020)
);

INVx2_ASAP7_75t_SL g1021 ( 
.A(n_767),
.Y(n_1021)
);

NAND2xp5_ASAP7_75t_L g1022 ( 
.A(n_749),
.B(n_638),
.Y(n_1022)
);

OAI21xp5_ASAP7_75t_L g1023 ( 
.A1(n_697),
.A2(n_696),
.B(n_698),
.Y(n_1023)
);

AOI21xp5_ASAP7_75t_L g1024 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1024)
);

NAND2xp5_ASAP7_75t_L g1025 ( 
.A(n_749),
.B(n_638),
.Y(n_1025)
);

NAND2xp5_ASAP7_75t_L g1026 ( 
.A(n_749),
.B(n_638),
.Y(n_1026)
);

AOI21xp5_ASAP7_75t_L g1027 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1027)
);

AOI21x1_ASAP7_75t_L g1028 ( 
.A1(n_772),
.A2(n_618),
.B(n_697),
.Y(n_1028)
);

BUFx8_ASAP7_75t_L g1029 ( 
.A(n_701),
.Y(n_1029)
);

AOI21xp5_ASAP7_75t_L g1030 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1030)
);

AOI21xp5_ASAP7_75t_L g1031 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1031)
);

NOR2xp33_ASAP7_75t_L g1032 ( 
.A(n_749),
.B(n_560),
.Y(n_1032)
);

AOI21xp5_ASAP7_75t_L g1033 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1033)
);

BUFx2_ASAP7_75t_L g1034 ( 
.A(n_755),
.Y(n_1034)
);

AOI21xp5_ASAP7_75t_L g1035 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1035)
);

AOI21xp5_ASAP7_75t_L g1036 ( 
.A1(n_696),
.A2(n_698),
.B(n_772),
.Y(n_1036)
);

NAND2xp5_ASAP7_75t_L g1037 ( 
.A(n_749),
.B(n_638),
.Y(n_1037)
);

NAND2xp5_ASAP7_75t_L g1038 ( 
.A(n_749),
.B(n_638),
.Y(n_1038)
);

OAI22xp5_ASAP7_75t_L g1039 ( 
.A1(n_720),
.A2(n_552),
.B1(n_749),
.B2(n_710),
.Y(n_1039)
);

INVx1_ASAP7_75t_L g1040 ( 
.A(n_869),
.Y(n_1040)
);

OAI21x1_ASAP7_75t_L g1041 ( 
.A1(n_1020),
.A2(n_863),
.B(n_1028),
.Y(n_1041)
);

INVx1_ASAP7_75t_L g1042 ( 
.A(n_874),
.Y(n_1042)
);

AOI21x1_ASAP7_75t_L g1043 ( 
.A1(n_941),
.A2(n_1000),
.B(n_940),
.Y(n_1043)
);

OAI21xp5_ASAP7_75t_L g1044 ( 
.A1(n_1032),
.A2(n_1010),
.B(n_1009),
.Y(n_1044)
);

OAI21x1_ASAP7_75t_L g1045 ( 
.A1(n_994),
.A2(n_968),
.B(n_976),
.Y(n_1045)
);

AOI21xp5_ASAP7_75t_L g1046 ( 
.A1(n_1005),
.A2(n_1022),
.B(n_1015),
.Y(n_1046)
);

OAI21x1_ASAP7_75t_L g1047 ( 
.A1(n_968),
.A2(n_976),
.B(n_858),
.Y(n_1047)
);

AO31x2_ASAP7_75t_L g1048 ( 
.A1(n_870),
.A2(n_1010),
.A3(n_883),
.B(n_1017),
.Y(n_1048)
);

CKINVDCx12_ASAP7_75t_R g1049 ( 
.A(n_1016),
.Y(n_1049)
);

INVxp67_ASAP7_75t_L g1050 ( 
.A(n_974),
.Y(n_1050)
);

NOR2xp33_ASAP7_75t_L g1051 ( 
.A(n_1032),
.B(n_1025),
.Y(n_1051)
);

NAND2xp5_ASAP7_75t_L g1052 ( 
.A(n_1026),
.B(n_1037),
.Y(n_1052)
);

BUFx3_ASAP7_75t_L g1053 ( 
.A(n_957),
.Y(n_1053)
);

AND2x2_ASAP7_75t_L g1054 ( 
.A(n_1011),
.B(n_973),
.Y(n_1054)
);

OAI21xp5_ASAP7_75t_L g1055 ( 
.A1(n_1038),
.A2(n_864),
.B(n_1008),
.Y(n_1055)
);

OAI21xp5_ASAP7_75t_L g1056 ( 
.A1(n_1039),
.A2(n_867),
.B(n_1001),
.Y(n_1056)
);

AND2x2_ASAP7_75t_L g1057 ( 
.A(n_974),
.B(n_970),
.Y(n_1057)
);

NAND2xp5_ASAP7_75t_L g1058 ( 
.A(n_942),
.B(n_949),
.Y(n_1058)
);

OAI21x1_ASAP7_75t_L g1059 ( 
.A1(n_995),
.A2(n_996),
.B(n_859),
.Y(n_1059)
);

AOI21xp5_ASAP7_75t_L g1060 ( 
.A1(n_1019),
.A2(n_1023),
.B(n_857),
.Y(n_1060)
);

NAND2xp5_ASAP7_75t_L g1061 ( 
.A(n_949),
.B(n_939),
.Y(n_1061)
);

NAND2xp5_ASAP7_75t_L g1062 ( 
.A(n_1013),
.B(n_872),
.Y(n_1062)
);

NAND2xp5_ASAP7_75t_L g1063 ( 
.A(n_1013),
.B(n_961),
.Y(n_1063)
);

AOI21x1_ASAP7_75t_L g1064 ( 
.A1(n_1000),
.A2(n_901),
.B(n_922),
.Y(n_1064)
);

AND2x2_ASAP7_75t_L g1065 ( 
.A(n_1034),
.B(n_868),
.Y(n_1065)
);

NAND2xp5_ASAP7_75t_L g1066 ( 
.A(n_865),
.B(n_964),
.Y(n_1066)
);

OAI21xp5_ASAP7_75t_L g1067 ( 
.A1(n_1002),
.A2(n_1006),
.B(n_1004),
.Y(n_1067)
);

NAND2xp5_ASAP7_75t_L g1068 ( 
.A(n_865),
.B(n_947),
.Y(n_1068)
);

OAI21x1_ASAP7_75t_L g1069 ( 
.A1(n_860),
.A2(n_861),
.B(n_966),
.Y(n_1069)
);

CKINVDCx20_ASAP7_75t_R g1070 ( 
.A(n_957),
.Y(n_1070)
);

OA22x2_ASAP7_75t_L g1071 ( 
.A1(n_862),
.A2(n_986),
.B1(n_1014),
.B2(n_918),
.Y(n_1071)
);

OAI21x1_ASAP7_75t_L g1072 ( 
.A1(n_967),
.A2(n_971),
.B(n_880),
.Y(n_1072)
);

AOI21xp5_ASAP7_75t_SL g1073 ( 
.A1(n_980),
.A2(n_993),
.B(n_988),
.Y(n_1073)
);

BUFx6f_ASAP7_75t_L g1074 ( 
.A(n_919),
.Y(n_1074)
);

BUFx2_ASAP7_75t_L g1075 ( 
.A(n_1029),
.Y(n_1075)
);

AOI21xp5_ASAP7_75t_L g1076 ( 
.A1(n_1018),
.A2(n_1033),
.B(n_1035),
.Y(n_1076)
);

INVxp67_ASAP7_75t_L g1077 ( 
.A(n_918),
.Y(n_1077)
);

AOI21xp5_ASAP7_75t_L g1078 ( 
.A1(n_1024),
.A2(n_1027),
.B(n_1030),
.Y(n_1078)
);

AND2x2_ASAP7_75t_L g1079 ( 
.A(n_959),
.B(n_1012),
.Y(n_1079)
);

OAI21x1_ASAP7_75t_L g1080 ( 
.A1(n_926),
.A2(n_977),
.B(n_871),
.Y(n_1080)
);

INVxp67_ASAP7_75t_L g1081 ( 
.A(n_1012),
.Y(n_1081)
);

AO21x1_ASAP7_75t_L g1082 ( 
.A1(n_982),
.A2(n_933),
.B(n_921),
.Y(n_1082)
);

AOI21xp5_ASAP7_75t_L g1083 ( 
.A1(n_1031),
.A2(n_1036),
.B(n_876),
.Y(n_1083)
);

INVx2_ASAP7_75t_SL g1084 ( 
.A(n_1029),
.Y(n_1084)
);

OAI21x1_ASAP7_75t_L g1085 ( 
.A1(n_904),
.A2(n_911),
.B(n_896),
.Y(n_1085)
);

AOI22xp33_ASAP7_75t_L g1086 ( 
.A1(n_909),
.A2(n_910),
.B1(n_924),
.B2(n_892),
.Y(n_1086)
);

OAI21x1_ASAP7_75t_L g1087 ( 
.A1(n_904),
.A2(n_911),
.B(n_882),
.Y(n_1087)
);

AND2x4_ASAP7_75t_L g1088 ( 
.A(n_931),
.B(n_960),
.Y(n_1088)
);

BUFx3_ASAP7_75t_L g1089 ( 
.A(n_944),
.Y(n_1089)
);

OAI21x1_ASAP7_75t_L g1090 ( 
.A1(n_882),
.A2(n_896),
.B(n_946),
.Y(n_1090)
);

AND2x4_ASAP7_75t_L g1091 ( 
.A(n_931),
.B(n_981),
.Y(n_1091)
);

NAND2xp5_ASAP7_75t_L g1092 ( 
.A(n_986),
.B(n_902),
.Y(n_1092)
);

INVx2_ASAP7_75t_SL g1093 ( 
.A(n_956),
.Y(n_1093)
);

AOI21xp5_ASAP7_75t_L g1094 ( 
.A1(n_998),
.A2(n_958),
.B(n_881),
.Y(n_1094)
);

AOI22xp5_ASAP7_75t_L g1095 ( 
.A1(n_924),
.A2(n_928),
.B1(n_978),
.B2(n_902),
.Y(n_1095)
);

NAND2xp5_ASAP7_75t_L g1096 ( 
.A(n_952),
.B(n_913),
.Y(n_1096)
);

OAI21x1_ASAP7_75t_L g1097 ( 
.A1(n_983),
.A2(n_985),
.B(n_912),
.Y(n_1097)
);

HB1xp67_ASAP7_75t_L g1098 ( 
.A(n_897),
.Y(n_1098)
);

OAI21xp5_ASAP7_75t_L g1099 ( 
.A1(n_870),
.A2(n_875),
.B(n_866),
.Y(n_1099)
);

OAI21x1_ASAP7_75t_L g1100 ( 
.A1(n_997),
.A2(n_916),
.B(n_955),
.Y(n_1100)
);

AND2x2_ASAP7_75t_L g1101 ( 
.A(n_908),
.B(n_886),
.Y(n_1101)
);

NAND2xp5_ASAP7_75t_L g1102 ( 
.A(n_948),
.B(n_886),
.Y(n_1102)
);

AOI21xp5_ASAP7_75t_L g1103 ( 
.A1(n_953),
.A2(n_945),
.B(n_984),
.Y(n_1103)
);

OAI21x1_ASAP7_75t_SL g1104 ( 
.A1(n_938),
.A2(n_969),
.B(n_895),
.Y(n_1104)
);

OAI21xp5_ASAP7_75t_L g1105 ( 
.A1(n_905),
.A2(n_907),
.B(n_951),
.Y(n_1105)
);

INVx3_ASAP7_75t_SL g1106 ( 
.A(n_944),
.Y(n_1106)
);

OAI21xp5_ASAP7_75t_SL g1107 ( 
.A1(n_927),
.A2(n_890),
.B(n_898),
.Y(n_1107)
);

AOI21xp5_ASAP7_75t_L g1108 ( 
.A1(n_950),
.A2(n_980),
.B(n_888),
.Y(n_1108)
);

NAND2xp5_ASAP7_75t_L g1109 ( 
.A(n_1003),
.B(n_963),
.Y(n_1109)
);

AOI21xp33_ASAP7_75t_L g1110 ( 
.A1(n_954),
.A2(n_884),
.B(n_914),
.Y(n_1110)
);

A2O1A1Ixp33_ASAP7_75t_L g1111 ( 
.A1(n_915),
.A2(n_899),
.B(n_883),
.C(n_936),
.Y(n_1111)
);

NAND2xp5_ASAP7_75t_L g1112 ( 
.A(n_1003),
.B(n_1021),
.Y(n_1112)
);

BUFx12f_ASAP7_75t_L g1113 ( 
.A(n_919),
.Y(n_1113)
);

NAND2xp5_ASAP7_75t_SL g1114 ( 
.A(n_917),
.B(n_879),
.Y(n_1114)
);

NOR2xp33_ASAP7_75t_SL g1115 ( 
.A(n_999),
.B(n_906),
.Y(n_1115)
);

AOI21xp5_ASAP7_75t_L g1116 ( 
.A1(n_873),
.A2(n_893),
.B(n_877),
.Y(n_1116)
);

OAI21xp5_ASAP7_75t_L g1117 ( 
.A1(n_987),
.A2(n_878),
.B(n_885),
.Y(n_1117)
);

AOI21xp5_ASAP7_75t_L g1118 ( 
.A1(n_893),
.A2(n_917),
.B(n_929),
.Y(n_1118)
);

AND3x4_ASAP7_75t_L g1119 ( 
.A(n_978),
.B(n_962),
.C(n_979),
.Y(n_1119)
);

OAI21x1_ASAP7_75t_L g1120 ( 
.A1(n_894),
.A2(n_990),
.B(n_937),
.Y(n_1120)
);

INVx2_ASAP7_75t_SL g1121 ( 
.A(n_979),
.Y(n_1121)
);

AOI21xp5_ASAP7_75t_L g1122 ( 
.A1(n_889),
.A2(n_934),
.B(n_887),
.Y(n_1122)
);

AOI21x1_ASAP7_75t_L g1123 ( 
.A1(n_920),
.A2(n_923),
.B(n_989),
.Y(n_1123)
);

OAI21x1_ASAP7_75t_L g1124 ( 
.A1(n_900),
.A2(n_935),
.B(n_965),
.Y(n_1124)
);

AND2x2_ASAP7_75t_L g1125 ( 
.A(n_975),
.B(n_915),
.Y(n_1125)
);

CKINVDCx20_ASAP7_75t_R g1126 ( 
.A(n_992),
.Y(n_1126)
);

OA22x2_ASAP7_75t_L g1127 ( 
.A1(n_903),
.A2(n_972),
.B1(n_932),
.B2(n_943),
.Y(n_1127)
);

AOI21xp5_ASAP7_75t_L g1128 ( 
.A1(n_943),
.A2(n_991),
.B(n_930),
.Y(n_1128)
);

OAI21x1_ASAP7_75t_L g1129 ( 
.A1(n_900),
.A2(n_935),
.B(n_1007),
.Y(n_1129)
);

OR2x6_ASAP7_75t_L g1130 ( 
.A(n_1007),
.B(n_991),
.Y(n_1130)
);

BUFx2_ASAP7_75t_L g1131 ( 
.A(n_891),
.Y(n_1131)
);

NAND2xp5_ASAP7_75t_L g1132 ( 
.A(n_891),
.B(n_925),
.Y(n_1132)
);

AO21x2_ASAP7_75t_L g1133 ( 
.A1(n_925),
.A2(n_870),
.B(n_1019),
.Y(n_1133)
);

INVx3_ASAP7_75t_L g1134 ( 
.A(n_919),
.Y(n_1134)
);

NAND2xp5_ASAP7_75t_L g1135 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1135)
);

OAI21x1_ASAP7_75t_L g1136 ( 
.A1(n_1020),
.A2(n_863),
.B(n_1028),
.Y(n_1136)
);

NAND2xp5_ASAP7_75t_SL g1137 ( 
.A(n_1010),
.B(n_1008),
.Y(n_1137)
);

A2O1A1Ixp33_ASAP7_75t_L g1138 ( 
.A1(n_1032),
.A2(n_1009),
.B(n_1015),
.C(n_1005),
.Y(n_1138)
);

AO31x2_ASAP7_75t_L g1139 ( 
.A1(n_870),
.A2(n_1010),
.A3(n_883),
.B(n_1008),
.Y(n_1139)
);

AOI21xp5_ASAP7_75t_L g1140 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1140)
);

AOI21xp5_ASAP7_75t_L g1141 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1141)
);

AND2x2_ASAP7_75t_SL g1142 ( 
.A(n_924),
.B(n_1032),
.Y(n_1142)
);

A2O1A1Ixp33_ASAP7_75t_L g1143 ( 
.A1(n_1032),
.A2(n_1009),
.B(n_1015),
.C(n_1005),
.Y(n_1143)
);

AOI21xp5_ASAP7_75t_L g1144 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1144)
);

NAND2xp5_ASAP7_75t_L g1145 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1145)
);

AOI21xp33_ASAP7_75t_L g1146 ( 
.A1(n_1032),
.A2(n_749),
.B(n_720),
.Y(n_1146)
);

O2A1O1Ixp5_ASAP7_75t_L g1147 ( 
.A1(n_1032),
.A2(n_1010),
.B(n_1017),
.C(n_1008),
.Y(n_1147)
);

AOI21xp5_ASAP7_75t_SL g1148 ( 
.A1(n_1010),
.A2(n_867),
.B(n_980),
.Y(n_1148)
);

INVx1_ASAP7_75t_L g1149 ( 
.A(n_869),
.Y(n_1149)
);

OAI21xp33_ASAP7_75t_SL g1150 ( 
.A1(n_1032),
.A2(n_1009),
.B(n_1005),
.Y(n_1150)
);

OAI22xp5_ASAP7_75t_L g1151 ( 
.A1(n_1032),
.A2(n_1009),
.B1(n_1022),
.B2(n_1005),
.Y(n_1151)
);

BUFx2_ASAP7_75t_L g1152 ( 
.A(n_1034),
.Y(n_1152)
);

NAND3xp33_ASAP7_75t_SL g1153 ( 
.A(n_1032),
.B(n_1009),
.C(n_1005),
.Y(n_1153)
);

OAI22xp5_ASAP7_75t_L g1154 ( 
.A1(n_1032),
.A2(n_1009),
.B1(n_1022),
.B2(n_1005),
.Y(n_1154)
);

INVx4_ASAP7_75t_L g1155 ( 
.A(n_919),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_869),
.Y(n_1156)
);

NAND3xp33_ASAP7_75t_L g1157 ( 
.A(n_1032),
.B(n_1009),
.C(n_1005),
.Y(n_1157)
);

INVx1_ASAP7_75t_L g1158 ( 
.A(n_869),
.Y(n_1158)
);

OAI21xp5_ASAP7_75t_L g1159 ( 
.A1(n_1032),
.A2(n_1010),
.B(n_1009),
.Y(n_1159)
);

AOI21xp5_ASAP7_75t_L g1160 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1160)
);

AOI21xp5_ASAP7_75t_L g1161 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1161)
);

INVx1_ASAP7_75t_L g1162 ( 
.A(n_869),
.Y(n_1162)
);

AOI21xp33_ASAP7_75t_L g1163 ( 
.A1(n_1032),
.A2(n_749),
.B(n_720),
.Y(n_1163)
);

NAND2xp5_ASAP7_75t_L g1164 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1164)
);

NAND2xp5_ASAP7_75t_L g1165 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1165)
);

INVx1_ASAP7_75t_SL g1166 ( 
.A(n_1034),
.Y(n_1166)
);

OAI21xp5_ASAP7_75t_L g1167 ( 
.A1(n_1032),
.A2(n_1010),
.B(n_1009),
.Y(n_1167)
);

OAI21xp33_ASAP7_75t_SL g1168 ( 
.A1(n_1032),
.A2(n_1009),
.B(n_1005),
.Y(n_1168)
);

CKINVDCx11_ASAP7_75t_R g1169 ( 
.A(n_944),
.Y(n_1169)
);

AOI21xp5_ASAP7_75t_L g1170 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1170)
);

OAI21x1_ASAP7_75t_L g1171 ( 
.A1(n_1020),
.A2(n_863),
.B(n_1028),
.Y(n_1171)
);

AND2x2_ASAP7_75t_SL g1172 ( 
.A(n_924),
.B(n_1032),
.Y(n_1172)
);

HB1xp67_ASAP7_75t_L g1173 ( 
.A(n_974),
.Y(n_1173)
);

NAND2xp5_ASAP7_75t_L g1174 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1174)
);

AOI21xp5_ASAP7_75t_L g1175 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1175)
);

OAI21x1_ASAP7_75t_SL g1176 ( 
.A1(n_994),
.A2(n_946),
.B(n_938),
.Y(n_1176)
);

AOI222xp33_ASAP7_75t_L g1177 ( 
.A1(n_1032),
.A2(n_711),
.B1(n_623),
.B2(n_435),
.C1(n_707),
.C2(n_749),
.Y(n_1177)
);

AOI21xp5_ASAP7_75t_L g1178 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1178)
);

AOI21xp5_ASAP7_75t_L g1179 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1179)
);

AOI21xp5_ASAP7_75t_L g1180 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1180)
);

INVx1_ASAP7_75t_L g1181 ( 
.A(n_869),
.Y(n_1181)
);

AND2x4_ASAP7_75t_L g1182 ( 
.A(n_1013),
.B(n_919),
.Y(n_1182)
);

AOI21x1_ASAP7_75t_SL g1183 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1183)
);

INVx1_ASAP7_75t_L g1184 ( 
.A(n_869),
.Y(n_1184)
);

AO31x2_ASAP7_75t_L g1185 ( 
.A1(n_870),
.A2(n_1010),
.A3(n_883),
.B(n_1008),
.Y(n_1185)
);

AO21x1_ASAP7_75t_L g1186 ( 
.A1(n_1008),
.A2(n_1039),
.B(n_1017),
.Y(n_1186)
);

AOI21xp5_ASAP7_75t_L g1187 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1187)
);

NOR2xp33_ASAP7_75t_L g1188 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1188)
);

AOI21xp5_ASAP7_75t_L g1189 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1189)
);

NOR2xp33_ASAP7_75t_L g1190 ( 
.A(n_1032),
.B(n_1005),
.Y(n_1190)
);

INVx4_ASAP7_75t_L g1191 ( 
.A(n_919),
.Y(n_1191)
);

CKINVDCx5p33_ASAP7_75t_R g1192 ( 
.A(n_956),
.Y(n_1192)
);

AOI21xp5_ASAP7_75t_L g1193 ( 
.A1(n_1005),
.A2(n_1015),
.B(n_1009),
.Y(n_1193)
);

A2O1A1Ixp33_ASAP7_75t_L g1194 ( 
.A1(n_1032),
.A2(n_1009),
.B(n_1015),
.C(n_1005),
.Y(n_1194)
);

NAND2xp5_ASAP7_75t_L g1195 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_1192),
.Y(n_1196)
);

NOR2xp33_ASAP7_75t_L g1197 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1197)
);

BUFx6f_ASAP7_75t_L g1198 ( 
.A(n_1182),
.Y(n_1198)
);

BUFx6f_ASAP7_75t_L g1199 ( 
.A(n_1182),
.Y(n_1199)
);

NAND2xp5_ASAP7_75t_SL g1200 ( 
.A(n_1142),
.B(n_1172),
.Y(n_1200)
);

AND2x2_ASAP7_75t_L g1201 ( 
.A(n_1054),
.B(n_1142),
.Y(n_1201)
);

INVx3_ASAP7_75t_L g1202 ( 
.A(n_1130),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_1192),
.Y(n_1203)
);

AND2x2_ASAP7_75t_L g1204 ( 
.A(n_1172),
.B(n_1065),
.Y(n_1204)
);

CKINVDCx6p67_ASAP7_75t_R g1205 ( 
.A(n_1053),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_1040),
.Y(n_1206)
);

INVxp67_ASAP7_75t_L g1207 ( 
.A(n_1152),
.Y(n_1207)
);

OAI22xp33_ASAP7_75t_L g1208 ( 
.A1(n_1095),
.A2(n_1135),
.B1(n_1145),
.B2(n_1164),
.Y(n_1208)
);

AOI22xp33_ASAP7_75t_SL g1209 ( 
.A1(n_1190),
.A2(n_1125),
.B1(n_1177),
.B2(n_1071),
.Y(n_1209)
);

OAI22xp5_ASAP7_75t_L g1210 ( 
.A1(n_1190),
.A2(n_1174),
.B1(n_1165),
.B2(n_1154),
.Y(n_1210)
);

AOI22xp33_ASAP7_75t_SL g1211 ( 
.A1(n_1071),
.A2(n_1151),
.B1(n_1157),
.B2(n_1126),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_1042),
.Y(n_1212)
);

AND2x2_ASAP7_75t_L g1213 ( 
.A(n_1079),
.B(n_1173),
.Y(n_1213)
);

INVxp67_ASAP7_75t_SL g1214 ( 
.A(n_1050),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_L g1215 ( 
.A(n_1138),
.B(n_1143),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1138),
.B(n_1143),
.Y(n_1216)
);

AOI21xp5_ASAP7_75t_L g1217 ( 
.A1(n_1148),
.A2(n_1159),
.B(n_1044),
.Y(n_1217)
);

CKINVDCx20_ASAP7_75t_R g1218 ( 
.A(n_1070),
.Y(n_1218)
);

NAND2x1p5_ASAP7_75t_L g1219 ( 
.A(n_1182),
.B(n_1089),
.Y(n_1219)
);

NAND2xp5_ASAP7_75t_L g1220 ( 
.A(n_1052),
.B(n_1058),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_L g1221 ( 
.A(n_1113),
.Y(n_1221)
);

NOR2xp33_ASAP7_75t_L g1222 ( 
.A(n_1153),
.B(n_1061),
.Y(n_1222)
);

HB1xp67_ASAP7_75t_L g1223 ( 
.A(n_1173),
.Y(n_1223)
);

INVx3_ASAP7_75t_SL g1224 ( 
.A(n_1070),
.Y(n_1224)
);

INVx1_ASAP7_75t_SL g1225 ( 
.A(n_1057),
.Y(n_1225)
);

INVxp67_ASAP7_75t_SL g1226 ( 
.A(n_1050),
.Y(n_1226)
);

HB1xp67_ASAP7_75t_L g1227 ( 
.A(n_1077),
.Y(n_1227)
);

INVx2_ASAP7_75t_SL g1228 ( 
.A(n_1053),
.Y(n_1228)
);

AOI21xp5_ASAP7_75t_L g1229 ( 
.A1(n_1167),
.A2(n_1056),
.B(n_1055),
.Y(n_1229)
);

OAI21x1_ASAP7_75t_L g1230 ( 
.A1(n_1041),
.A2(n_1171),
.B(n_1136),
.Y(n_1230)
);

NAND2xp5_ASAP7_75t_L g1231 ( 
.A(n_1194),
.B(n_1046),
.Y(n_1231)
);

A2O1A1Ixp33_ASAP7_75t_L g1232 ( 
.A1(n_1146),
.A2(n_1163),
.B(n_1150),
.C(n_1168),
.Y(n_1232)
);

BUFx6f_ASAP7_75t_L g1233 ( 
.A(n_1113),
.Y(n_1233)
);

BUFx12f_ASAP7_75t_L g1234 ( 
.A(n_1169),
.Y(n_1234)
);

NAND2xp5_ASAP7_75t_L g1235 ( 
.A(n_1194),
.B(n_1153),
.Y(n_1235)
);

INVx2_ASAP7_75t_SL g1236 ( 
.A(n_1106),
.Y(n_1236)
);

NAND2xp5_ASAP7_75t_L g1237 ( 
.A(n_1063),
.B(n_1140),
.Y(n_1237)
);

INVxp67_ASAP7_75t_L g1238 ( 
.A(n_1101),
.Y(n_1238)
);

AND2x4_ASAP7_75t_L g1239 ( 
.A(n_1089),
.B(n_1091),
.Y(n_1239)
);

AND2x2_ASAP7_75t_L g1240 ( 
.A(n_1077),
.B(n_1081),
.Y(n_1240)
);

AOI21xp5_ASAP7_75t_L g1241 ( 
.A1(n_1141),
.A2(n_1193),
.B(n_1189),
.Y(n_1241)
);

CKINVDCx20_ASAP7_75t_R g1242 ( 
.A(n_1169),
.Y(n_1242)
);

BUFx6f_ASAP7_75t_L g1243 ( 
.A(n_1074),
.Y(n_1243)
);

INVx5_ASAP7_75t_L g1244 ( 
.A(n_1130),
.Y(n_1244)
);

OA21x2_ASAP7_75t_L g1245 ( 
.A1(n_1067),
.A2(n_1083),
.B(n_1076),
.Y(n_1245)
);

NAND2xp5_ASAP7_75t_L g1246 ( 
.A(n_1144),
.B(n_1160),
.Y(n_1246)
);

OAI22xp5_ASAP7_75t_SL g1247 ( 
.A1(n_1119),
.A2(n_1126),
.B1(n_1102),
.B2(n_1106),
.Y(n_1247)
);

NAND2xp5_ASAP7_75t_SL g1248 ( 
.A(n_1161),
.B(n_1170),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_1093),
.Y(n_1249)
);

NOR4xp25_ASAP7_75t_SL g1250 ( 
.A(n_1107),
.B(n_1137),
.C(n_1111),
.D(n_1110),
.Y(n_1250)
);

NAND2xp5_ASAP7_75t_L g1251 ( 
.A(n_1175),
.B(n_1178),
.Y(n_1251)
);

OAI21x1_ASAP7_75t_L g1252 ( 
.A1(n_1080),
.A2(n_1072),
.B(n_1120),
.Y(n_1252)
);

BUFx6f_ASAP7_75t_L g1253 ( 
.A(n_1074),
.Y(n_1253)
);

OR2x6_ASAP7_75t_L g1254 ( 
.A(n_1073),
.B(n_1091),
.Y(n_1254)
);

NAND2xp5_ASAP7_75t_L g1255 ( 
.A(n_1179),
.B(n_1180),
.Y(n_1255)
);

AND2x4_ASAP7_75t_L g1256 ( 
.A(n_1088),
.B(n_1155),
.Y(n_1256)
);

AND2x2_ASAP7_75t_L g1257 ( 
.A(n_1081),
.B(n_1088),
.Y(n_1257)
);

NOR2xp33_ASAP7_75t_L g1258 ( 
.A(n_1062),
.B(n_1092),
.Y(n_1258)
);

NAND2xp5_ASAP7_75t_L g1259 ( 
.A(n_1187),
.B(n_1086),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1149),
.Y(n_1260)
);

AOI22xp33_ASAP7_75t_L g1261 ( 
.A1(n_1086),
.A2(n_1186),
.B1(n_1066),
.B2(n_1068),
.Y(n_1261)
);

AOI21xp5_ASAP7_75t_L g1262 ( 
.A1(n_1060),
.A2(n_1147),
.B(n_1137),
.Y(n_1262)
);

BUFx6f_ASAP7_75t_L g1263 ( 
.A(n_1074),
.Y(n_1263)
);

OAI22xp5_ASAP7_75t_L g1264 ( 
.A1(n_1111),
.A2(n_1096),
.B1(n_1156),
.B2(n_1184),
.Y(n_1264)
);

OR2x6_ASAP7_75t_SL g1265 ( 
.A(n_1112),
.B(n_1109),
.Y(n_1265)
);

INVx2_ASAP7_75t_SL g1266 ( 
.A(n_1075),
.Y(n_1266)
);

AOI21xp5_ASAP7_75t_SL g1267 ( 
.A1(n_1105),
.A2(n_1118),
.B(n_1114),
.Y(n_1267)
);

INVx1_ASAP7_75t_L g1268 ( 
.A(n_1158),
.Y(n_1268)
);

INVx1_ASAP7_75t_L g1269 ( 
.A(n_1162),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_1181),
.B(n_1084),
.Y(n_1270)
);

AOI21xp5_ASAP7_75t_SL g1271 ( 
.A1(n_1114),
.A2(n_1117),
.B(n_1128),
.Y(n_1271)
);

AND2x4_ASAP7_75t_L g1272 ( 
.A(n_1155),
.B(n_1191),
.Y(n_1272)
);

OAI22xp5_ASAP7_75t_L g1273 ( 
.A1(n_1119),
.A2(n_1147),
.B1(n_1099),
.B2(n_1131),
.Y(n_1273)
);

AOI21xp5_ASAP7_75t_L g1274 ( 
.A1(n_1094),
.A2(n_1082),
.B(n_1103),
.Y(n_1274)
);

INVx3_ASAP7_75t_SL g1275 ( 
.A(n_1191),
.Y(n_1275)
);

OR2x2_ASAP7_75t_L g1276 ( 
.A(n_1121),
.B(n_1098),
.Y(n_1276)
);

A2O1A1Ixp33_ASAP7_75t_L g1277 ( 
.A1(n_1122),
.A2(n_1108),
.B(n_1129),
.C(n_1115),
.Y(n_1277)
);

NAND2xp5_ASAP7_75t_L g1278 ( 
.A(n_1098),
.B(n_1134),
.Y(n_1278)
);

OAI221xp5_ASAP7_75t_L g1279 ( 
.A1(n_1123),
.A2(n_1116),
.B1(n_1132),
.B2(n_1104),
.C(n_1134),
.Y(n_1279)
);

A2O1A1Ixp33_ASAP7_75t_SL g1280 ( 
.A1(n_1078),
.A2(n_1183),
.B(n_1064),
.C(n_1043),
.Y(n_1280)
);

AND2x4_ASAP7_75t_L g1281 ( 
.A(n_1124),
.B(n_1133),
.Y(n_1281)
);

OR2x2_ASAP7_75t_L g1282 ( 
.A(n_1049),
.B(n_1185),
.Y(n_1282)
);

INVx2_ASAP7_75t_SL g1283 ( 
.A(n_1127),
.Y(n_1283)
);

AND2x4_ASAP7_75t_L g1284 ( 
.A(n_1133),
.B(n_1090),
.Y(n_1284)
);

INVx2_ASAP7_75t_L g1285 ( 
.A(n_1127),
.Y(n_1285)
);

BUFx2_ASAP7_75t_L g1286 ( 
.A(n_1048),
.Y(n_1286)
);

AND2x2_ASAP7_75t_L g1287 ( 
.A(n_1048),
.B(n_1139),
.Y(n_1287)
);

INVx2_ASAP7_75t_SL g1288 ( 
.A(n_1085),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_L g1289 ( 
.A(n_1183),
.B(n_1176),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1097),
.Y(n_1290)
);

BUFx6f_ASAP7_75t_L g1291 ( 
.A(n_1047),
.Y(n_1291)
);

NOR2x1_ASAP7_75t_SL g1292 ( 
.A(n_1087),
.B(n_1045),
.Y(n_1292)
);

AOI21xp33_ASAP7_75t_SL g1293 ( 
.A1(n_1100),
.A2(n_1059),
.B(n_1069),
.Y(n_1293)
);

INVx3_ASAP7_75t_L g1294 ( 
.A(n_1048),
.Y(n_1294)
);

BUFx12f_ASAP7_75t_L g1295 ( 
.A(n_1048),
.Y(n_1295)
);

OAI22xp5_ASAP7_75t_L g1296 ( 
.A1(n_1139),
.A2(n_1142),
.B1(n_1172),
.B2(n_1051),
.Y(n_1296)
);

NAND2xp5_ASAP7_75t_L g1297 ( 
.A(n_1185),
.B(n_1051),
.Y(n_1297)
);

NAND2xp5_ASAP7_75t_L g1298 ( 
.A(n_1185),
.B(n_1051),
.Y(n_1298)
);

AND2x2_ASAP7_75t_L g1299 ( 
.A(n_1185),
.B(n_1054),
.Y(n_1299)
);

INVx1_ASAP7_75t_L g1300 ( 
.A(n_1040),
.Y(n_1300)
);

OAI22xp5_ASAP7_75t_L g1301 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1188),
.B2(n_1051),
.Y(n_1301)
);

AOI21xp5_ASAP7_75t_L g1302 ( 
.A1(n_1148),
.A2(n_1010),
.B(n_1044),
.Y(n_1302)
);

AND2x2_ASAP7_75t_L g1303 ( 
.A(n_1054),
.B(n_1011),
.Y(n_1303)
);

OAI21xp5_ASAP7_75t_L g1304 ( 
.A1(n_1147),
.A2(n_1032),
.B(n_1010),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_L g1305 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1305)
);

NAND2xp5_ASAP7_75t_L g1306 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1306)
);

AND2x2_ASAP7_75t_L g1307 ( 
.A(n_1054),
.B(n_1011),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_1040),
.Y(n_1308)
);

AND2x4_ASAP7_75t_L g1309 ( 
.A(n_1182),
.B(n_1089),
.Y(n_1309)
);

INVx4_ASAP7_75t_L g1310 ( 
.A(n_1106),
.Y(n_1310)
);

INVx5_ASAP7_75t_L g1311 ( 
.A(n_1130),
.Y(n_1311)
);

AOI21xp5_ASAP7_75t_L g1312 ( 
.A1(n_1148),
.A2(n_1010),
.B(n_1044),
.Y(n_1312)
);

BUFx12f_ASAP7_75t_L g1313 ( 
.A(n_1192),
.Y(n_1313)
);

AND2x4_ASAP7_75t_L g1314 ( 
.A(n_1182),
.B(n_1089),
.Y(n_1314)
);

NAND2xp5_ASAP7_75t_L g1315 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1315)
);

OR2x2_ASAP7_75t_L g1316 ( 
.A(n_1054),
.B(n_1166),
.Y(n_1316)
);

INVx2_ASAP7_75t_SL g1317 ( 
.A(n_1053),
.Y(n_1317)
);

OAI21xp33_ASAP7_75t_L g1318 ( 
.A1(n_1051),
.A2(n_1032),
.B(n_1188),
.Y(n_1318)
);

AOI22xp5_ASAP7_75t_L g1319 ( 
.A1(n_1142),
.A2(n_1032),
.B1(n_1172),
.B2(n_1177),
.Y(n_1319)
);

OAI22xp5_ASAP7_75t_L g1320 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1188),
.B2(n_1051),
.Y(n_1320)
);

BUFx10_ASAP7_75t_L g1321 ( 
.A(n_1192),
.Y(n_1321)
);

CKINVDCx6p67_ASAP7_75t_R g1322 ( 
.A(n_1053),
.Y(n_1322)
);

AND2x4_ASAP7_75t_L g1323 ( 
.A(n_1182),
.B(n_1089),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_L g1324 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1324)
);

NAND2xp5_ASAP7_75t_SL g1325 ( 
.A(n_1142),
.B(n_1172),
.Y(n_1325)
);

OAI22xp5_ASAP7_75t_L g1326 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1188),
.B2(n_1051),
.Y(n_1326)
);

INVx1_ASAP7_75t_L g1327 ( 
.A(n_1040),
.Y(n_1327)
);

INVx1_ASAP7_75t_L g1328 ( 
.A(n_1040),
.Y(n_1328)
);

CKINVDCx5p33_ASAP7_75t_R g1329 ( 
.A(n_1192),
.Y(n_1329)
);

OAI21xp5_ASAP7_75t_L g1330 ( 
.A1(n_1147),
.A2(n_1032),
.B(n_1010),
.Y(n_1330)
);

OAI22xp5_ASAP7_75t_L g1331 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1188),
.B2(n_1051),
.Y(n_1331)
);

NAND2xp5_ASAP7_75t_L g1332 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1332)
);

O2A1O1Ixp33_ASAP7_75t_L g1333 ( 
.A1(n_1051),
.A2(n_1032),
.B(n_1009),
.C(n_1015),
.Y(n_1333)
);

AOI22xp5_ASAP7_75t_L g1334 ( 
.A1(n_1142),
.A2(n_1032),
.B1(n_1172),
.B2(n_1177),
.Y(n_1334)
);

BUFx3_ASAP7_75t_L g1335 ( 
.A(n_1106),
.Y(n_1335)
);

NAND2xp5_ASAP7_75t_L g1336 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1336)
);

AOI22xp5_ASAP7_75t_L g1337 ( 
.A1(n_1142),
.A2(n_1032),
.B1(n_1172),
.B2(n_1177),
.Y(n_1337)
);

OAI22xp5_ASAP7_75t_L g1338 ( 
.A1(n_1142),
.A2(n_1172),
.B1(n_1188),
.B2(n_1051),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1040),
.Y(n_1339)
);

INVx5_ASAP7_75t_L g1340 ( 
.A(n_1130),
.Y(n_1340)
);

NAND2xp5_ASAP7_75t_L g1341 ( 
.A(n_1051),
.B(n_1188),
.Y(n_1341)
);

OAI21xp5_ASAP7_75t_L g1342 ( 
.A1(n_1147),
.A2(n_1032),
.B(n_1010),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_SL g1343 ( 
.A(n_1142),
.B(n_1172),
.Y(n_1343)
);

INVx2_ASAP7_75t_SL g1344 ( 
.A(n_1053),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1206),
.Y(n_1345)
);

INVx1_ASAP7_75t_SL g1346 ( 
.A(n_1316),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_1254),
.Y(n_1347)
);

BUFx3_ASAP7_75t_L g1348 ( 
.A(n_1335),
.Y(n_1348)
);

CKINVDCx5p33_ASAP7_75t_R g1349 ( 
.A(n_1218),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1212),
.Y(n_1350)
);

OAI21x1_ASAP7_75t_L g1351 ( 
.A1(n_1252),
.A2(n_1274),
.B(n_1230),
.Y(n_1351)
);

OAI22xp5_ASAP7_75t_L g1352 ( 
.A1(n_1319),
.A2(n_1337),
.B1(n_1334),
.B2(n_1197),
.Y(n_1352)
);

AOI22xp5_ASAP7_75t_L g1353 ( 
.A1(n_1209),
.A2(n_1320),
.B1(n_1326),
.B2(n_1301),
.Y(n_1353)
);

OAI21x1_ASAP7_75t_L g1354 ( 
.A1(n_1241),
.A2(n_1262),
.B(n_1290),
.Y(n_1354)
);

INVx5_ASAP7_75t_L g1355 ( 
.A(n_1254),
.Y(n_1355)
);

BUFx6f_ASAP7_75t_SL g1356 ( 
.A(n_1321),
.Y(n_1356)
);

AOI22xp33_ASAP7_75t_L g1357 ( 
.A1(n_1211),
.A2(n_1296),
.B1(n_1331),
.B2(n_1301),
.Y(n_1357)
);

CKINVDCx8_ASAP7_75t_R g1358 ( 
.A(n_1309),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1260),
.Y(n_1359)
);

BUFx3_ASAP7_75t_L g1360 ( 
.A(n_1309),
.Y(n_1360)
);

AOI22xp33_ASAP7_75t_L g1361 ( 
.A1(n_1296),
.A2(n_1326),
.B1(n_1331),
.B2(n_1320),
.Y(n_1361)
);

INVx1_ASAP7_75t_L g1362 ( 
.A(n_1268),
.Y(n_1362)
);

HB1xp67_ASAP7_75t_L g1363 ( 
.A(n_1213),
.Y(n_1363)
);

AOI22xp33_ASAP7_75t_L g1364 ( 
.A1(n_1338),
.A2(n_1318),
.B1(n_1295),
.B2(n_1208),
.Y(n_1364)
);

AND2x2_ASAP7_75t_L g1365 ( 
.A(n_1299),
.B(n_1297),
.Y(n_1365)
);

INVx1_ASAP7_75t_L g1366 ( 
.A(n_1269),
.Y(n_1366)
);

AOI22xp33_ASAP7_75t_SL g1367 ( 
.A1(n_1338),
.A2(n_1273),
.B1(n_1247),
.B2(n_1210),
.Y(n_1367)
);

BUFx3_ASAP7_75t_L g1368 ( 
.A(n_1314),
.Y(n_1368)
);

AOI22xp33_ASAP7_75t_SL g1369 ( 
.A1(n_1273),
.A2(n_1210),
.B1(n_1222),
.B2(n_1342),
.Y(n_1369)
);

HB1xp67_ASAP7_75t_L g1370 ( 
.A(n_1223),
.Y(n_1370)
);

INVx1_ASAP7_75t_L g1371 ( 
.A(n_1300),
.Y(n_1371)
);

BUFx2_ASAP7_75t_L g1372 ( 
.A(n_1284),
.Y(n_1372)
);

OAI21x1_ASAP7_75t_L g1373 ( 
.A1(n_1248),
.A2(n_1246),
.B(n_1251),
.Y(n_1373)
);

INVx1_ASAP7_75t_L g1374 ( 
.A(n_1308),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_1327),
.Y(n_1375)
);

AOI22xp33_ASAP7_75t_SL g1376 ( 
.A1(n_1304),
.A2(n_1342),
.B1(n_1330),
.B2(n_1217),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_1328),
.Y(n_1377)
);

AOI22xp5_ASAP7_75t_L g1378 ( 
.A1(n_1258),
.A2(n_1343),
.B1(n_1200),
.B2(n_1325),
.Y(n_1378)
);

HB1xp67_ASAP7_75t_L g1379 ( 
.A(n_1240),
.Y(n_1379)
);

CKINVDCx5p33_ASAP7_75t_R g1380 ( 
.A(n_1196),
.Y(n_1380)
);

INVx3_ASAP7_75t_SL g1381 ( 
.A(n_1203),
.Y(n_1381)
);

OA21x2_ASAP7_75t_L g1382 ( 
.A1(n_1229),
.A2(n_1302),
.B(n_1312),
.Y(n_1382)
);

AND2x6_ASAP7_75t_L g1383 ( 
.A(n_1285),
.B(n_1202),
.Y(n_1383)
);

AND2x2_ASAP7_75t_L g1384 ( 
.A(n_1297),
.B(n_1298),
.Y(n_1384)
);

AOI22xp33_ASAP7_75t_L g1385 ( 
.A1(n_1282),
.A2(n_1204),
.B1(n_1283),
.B2(n_1201),
.Y(n_1385)
);

INVx1_ASAP7_75t_L g1386 ( 
.A(n_1339),
.Y(n_1386)
);

AND2x2_ASAP7_75t_L g1387 ( 
.A(n_1298),
.B(n_1287),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1214),
.Y(n_1388)
);

INVx1_ASAP7_75t_L g1389 ( 
.A(n_1226),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1286),
.B(n_1235),
.Y(n_1390)
);

INVx1_ASAP7_75t_L g1391 ( 
.A(n_1227),
.Y(n_1391)
);

INVx3_ASAP7_75t_L g1392 ( 
.A(n_1284),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1276),
.Y(n_1393)
);

BUFx2_ASAP7_75t_L g1394 ( 
.A(n_1294),
.Y(n_1394)
);

AND2x4_ASAP7_75t_L g1395 ( 
.A(n_1244),
.B(n_1311),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_1278),
.Y(n_1396)
);

AOI22xp33_ASAP7_75t_L g1397 ( 
.A1(n_1303),
.A2(n_1307),
.B1(n_1261),
.B2(n_1315),
.Y(n_1397)
);

INVx1_ASAP7_75t_L g1398 ( 
.A(n_1264),
.Y(n_1398)
);

INVx5_ASAP7_75t_L g1399 ( 
.A(n_1311),
.Y(n_1399)
);

BUFx6f_ASAP7_75t_L g1400 ( 
.A(n_1198),
.Y(n_1400)
);

AOI22xp5_ASAP7_75t_L g1401 ( 
.A1(n_1305),
.A2(n_1306),
.B1(n_1341),
.B2(n_1332),
.Y(n_1401)
);

BUFx2_ASAP7_75t_R g1402 ( 
.A(n_1329),
.Y(n_1402)
);

INVx1_ASAP7_75t_L g1403 ( 
.A(n_1264),
.Y(n_1403)
);

INVx1_ASAP7_75t_L g1404 ( 
.A(n_1257),
.Y(n_1404)
);

OAI21x1_ASAP7_75t_L g1405 ( 
.A1(n_1246),
.A2(n_1255),
.B(n_1251),
.Y(n_1405)
);

BUFx8_ASAP7_75t_SL g1406 ( 
.A(n_1313),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1237),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_1238),
.Y(n_1408)
);

OAI21xp5_ASAP7_75t_L g1409 ( 
.A1(n_1333),
.A2(n_1304),
.B(n_1330),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1259),
.Y(n_1410)
);

NAND2xp5_ASAP7_75t_L g1411 ( 
.A(n_1195),
.B(n_1315),
.Y(n_1411)
);

INVx2_ASAP7_75t_L g1412 ( 
.A(n_1281),
.Y(n_1412)
);

CKINVDCx20_ASAP7_75t_R g1413 ( 
.A(n_1242),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1270),
.Y(n_1414)
);

INVx1_ASAP7_75t_L g1415 ( 
.A(n_1255),
.Y(n_1415)
);

AO21x2_ASAP7_75t_L g1416 ( 
.A1(n_1293),
.A2(n_1232),
.B(n_1277),
.Y(n_1416)
);

AOI22xp33_ASAP7_75t_L g1417 ( 
.A1(n_1195),
.A2(n_1336),
.B1(n_1324),
.B2(n_1225),
.Y(n_1417)
);

INVx1_ASAP7_75t_L g1418 ( 
.A(n_1231),
.Y(n_1418)
);

BUFx2_ASAP7_75t_L g1419 ( 
.A(n_1291),
.Y(n_1419)
);

INVx2_ASAP7_75t_L g1420 ( 
.A(n_1245),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_1231),
.Y(n_1421)
);

OAI22xp5_ASAP7_75t_L g1422 ( 
.A1(n_1324),
.A2(n_1336),
.B1(n_1250),
.B2(n_1216),
.Y(n_1422)
);

AO21x1_ASAP7_75t_L g1423 ( 
.A1(n_1215),
.A2(n_1216),
.B(n_1289),
.Y(n_1423)
);

AO21x2_ASAP7_75t_L g1424 ( 
.A1(n_1280),
.A2(n_1271),
.B(n_1267),
.Y(n_1424)
);

INVx3_ASAP7_75t_L g1425 ( 
.A(n_1291),
.Y(n_1425)
);

NAND2xp5_ASAP7_75t_L g1426 ( 
.A(n_1220),
.B(n_1207),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1225),
.Y(n_1427)
);

INVx2_ASAP7_75t_SL g1428 ( 
.A(n_1340),
.Y(n_1428)
);

OAI22xp33_ASAP7_75t_L g1429 ( 
.A1(n_1265),
.A2(n_1215),
.B1(n_1224),
.B2(n_1266),
.Y(n_1429)
);

INVx1_ASAP7_75t_L g1430 ( 
.A(n_1239),
.Y(n_1430)
);

INVx2_ASAP7_75t_L g1431 ( 
.A(n_1288),
.Y(n_1431)
);

HB1xp67_ASAP7_75t_L g1432 ( 
.A(n_1314),
.Y(n_1432)
);

INVx1_ASAP7_75t_L g1433 ( 
.A(n_1239),
.Y(n_1433)
);

INVx1_ASAP7_75t_L g1434 ( 
.A(n_1219),
.Y(n_1434)
);

INVx1_ASAP7_75t_L g1435 ( 
.A(n_1219),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1323),
.Y(n_1436)
);

BUFx6f_ASAP7_75t_L g1437 ( 
.A(n_1198),
.Y(n_1437)
);

INVx1_ASAP7_75t_L g1438 ( 
.A(n_1323),
.Y(n_1438)
);

CKINVDCx11_ASAP7_75t_R g1439 ( 
.A(n_1321),
.Y(n_1439)
);

AOI22xp33_ASAP7_75t_L g1440 ( 
.A1(n_1340),
.A2(n_1344),
.B1(n_1317),
.B2(n_1228),
.Y(n_1440)
);

AND2x2_ASAP7_75t_L g1441 ( 
.A(n_1250),
.B(n_1199),
.Y(n_1441)
);

BUFx2_ASAP7_75t_SL g1442 ( 
.A(n_1310),
.Y(n_1442)
);

CKINVDCx11_ASAP7_75t_R g1443 ( 
.A(n_1234),
.Y(n_1443)
);

BUFx4f_ASAP7_75t_SL g1444 ( 
.A(n_1205),
.Y(n_1444)
);

OAI21x1_ASAP7_75t_L g1445 ( 
.A1(n_1292),
.A2(n_1279),
.B(n_1291),
.Y(n_1445)
);

INVx2_ASAP7_75t_SL g1446 ( 
.A(n_1243),
.Y(n_1446)
);

HB1xp67_ASAP7_75t_L g1447 ( 
.A(n_1243),
.Y(n_1447)
);

AOI22xp33_ASAP7_75t_SL g1448 ( 
.A1(n_1199),
.A2(n_1256),
.B1(n_1233),
.B2(n_1221),
.Y(n_1448)
);

INVx3_ASAP7_75t_L g1449 ( 
.A(n_1253),
.Y(n_1449)
);

INVx1_ASAP7_75t_L g1450 ( 
.A(n_1253),
.Y(n_1450)
);

OR2x6_ASAP7_75t_L g1451 ( 
.A(n_1221),
.B(n_1233),
.Y(n_1451)
);

AOI22xp33_ASAP7_75t_L g1452 ( 
.A1(n_1256),
.A2(n_1322),
.B1(n_1233),
.B2(n_1221),
.Y(n_1452)
);

INVx4_ASAP7_75t_L g1453 ( 
.A(n_1253),
.Y(n_1453)
);

INVx2_ASAP7_75t_L g1454 ( 
.A(n_1263),
.Y(n_1454)
);

INVx1_ASAP7_75t_L g1455 ( 
.A(n_1236),
.Y(n_1455)
);

INVx2_ASAP7_75t_L g1456 ( 
.A(n_1272),
.Y(n_1456)
);

BUFx2_ASAP7_75t_L g1457 ( 
.A(n_1310),
.Y(n_1457)
);

BUFx3_ASAP7_75t_L g1458 ( 
.A(n_1275),
.Y(n_1458)
);

OR2x6_ASAP7_75t_L g1459 ( 
.A(n_1249),
.B(n_1073),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1206),
.Y(n_1460)
);

BUFx2_ASAP7_75t_L g1461 ( 
.A(n_1284),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1206),
.Y(n_1462)
);

AOI22xp33_ASAP7_75t_L g1463 ( 
.A1(n_1319),
.A2(n_1177),
.B1(n_1172),
.B2(n_1142),
.Y(n_1463)
);

AOI222xp33_ASAP7_75t_L g1464 ( 
.A1(n_1197),
.A2(n_1142),
.B1(n_1172),
.B2(n_623),
.C1(n_711),
.C2(n_1032),
.Y(n_1464)
);

AOI21x1_ASAP7_75t_L g1465 ( 
.A1(n_1274),
.A2(n_1083),
.B(n_1078),
.Y(n_1465)
);

INVx1_ASAP7_75t_L g1466 ( 
.A(n_1206),
.Y(n_1466)
);

AOI21x1_ASAP7_75t_L g1467 ( 
.A1(n_1274),
.A2(n_1083),
.B(n_1078),
.Y(n_1467)
);

INVx3_ASAP7_75t_L g1468 ( 
.A(n_1425),
.Y(n_1468)
);

BUFx6f_ASAP7_75t_L g1469 ( 
.A(n_1347),
.Y(n_1469)
);

INVx3_ASAP7_75t_L g1470 ( 
.A(n_1425),
.Y(n_1470)
);

AND2x2_ASAP7_75t_L g1471 ( 
.A(n_1365),
.B(n_1387),
.Y(n_1471)
);

OAI21x1_ASAP7_75t_L g1472 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1351),
.Y(n_1472)
);

NOR2xp33_ASAP7_75t_L g1473 ( 
.A(n_1401),
.B(n_1349),
.Y(n_1473)
);

BUFx2_ASAP7_75t_SL g1474 ( 
.A(n_1358),
.Y(n_1474)
);

OAI21x1_ASAP7_75t_L g1475 ( 
.A1(n_1465),
.A2(n_1467),
.B(n_1354),
.Y(n_1475)
);

AND2x2_ASAP7_75t_L g1476 ( 
.A(n_1365),
.B(n_1387),
.Y(n_1476)
);

BUFx2_ASAP7_75t_SL g1477 ( 
.A(n_1358),
.Y(n_1477)
);

INVx1_ASAP7_75t_L g1478 ( 
.A(n_1415),
.Y(n_1478)
);

INVx2_ASAP7_75t_L g1479 ( 
.A(n_1420),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1410),
.Y(n_1480)
);

OA21x2_ASAP7_75t_L g1481 ( 
.A1(n_1405),
.A2(n_1373),
.B(n_1423),
.Y(n_1481)
);

INVx3_ASAP7_75t_L g1482 ( 
.A(n_1445),
.Y(n_1482)
);

BUFx2_ASAP7_75t_L g1483 ( 
.A(n_1419),
.Y(n_1483)
);

INVx1_ASAP7_75t_L g1484 ( 
.A(n_1384),
.Y(n_1484)
);

INVx2_ASAP7_75t_L g1485 ( 
.A(n_1382),
.Y(n_1485)
);

NOR2xp33_ASAP7_75t_L g1486 ( 
.A(n_1349),
.B(n_1411),
.Y(n_1486)
);

INVx2_ASAP7_75t_L g1487 ( 
.A(n_1382),
.Y(n_1487)
);

HB1xp67_ASAP7_75t_L g1488 ( 
.A(n_1370),
.Y(n_1488)
);

INVx1_ASAP7_75t_L g1489 ( 
.A(n_1407),
.Y(n_1489)
);

AO21x2_ASAP7_75t_L g1490 ( 
.A1(n_1353),
.A2(n_1409),
.B(n_1431),
.Y(n_1490)
);

INVx1_ASAP7_75t_L g1491 ( 
.A(n_1418),
.Y(n_1491)
);

AO21x2_ASAP7_75t_L g1492 ( 
.A1(n_1431),
.A2(n_1416),
.B(n_1421),
.Y(n_1492)
);

AND2x4_ASAP7_75t_L g1493 ( 
.A(n_1355),
.B(n_1392),
.Y(n_1493)
);

NAND4xp25_ASAP7_75t_L g1494 ( 
.A(n_1464),
.B(n_1369),
.C(n_1367),
.D(n_1463),
.Y(n_1494)
);

OR2x2_ASAP7_75t_L g1495 ( 
.A(n_1390),
.B(n_1363),
.Y(n_1495)
);

INVx1_ASAP7_75t_L g1496 ( 
.A(n_1398),
.Y(n_1496)
);

HB1xp67_ASAP7_75t_L g1497 ( 
.A(n_1379),
.Y(n_1497)
);

INVx1_ASAP7_75t_L g1498 ( 
.A(n_1403),
.Y(n_1498)
);

BUFx3_ASAP7_75t_L g1499 ( 
.A(n_1372),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_1394),
.Y(n_1500)
);

AOI22xp33_ASAP7_75t_L g1501 ( 
.A1(n_1352),
.A2(n_1357),
.B1(n_1397),
.B2(n_1364),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1394),
.Y(n_1502)
);

INVx1_ASAP7_75t_L g1503 ( 
.A(n_1345),
.Y(n_1503)
);

INVx1_ASAP7_75t_L g1504 ( 
.A(n_1350),
.Y(n_1504)
);

BUFx2_ASAP7_75t_L g1505 ( 
.A(n_1419),
.Y(n_1505)
);

AND2x2_ASAP7_75t_L g1506 ( 
.A(n_1390),
.B(n_1372),
.Y(n_1506)
);

HB1xp67_ASAP7_75t_L g1507 ( 
.A(n_1388),
.Y(n_1507)
);

INVx4_ASAP7_75t_L g1508 ( 
.A(n_1355),
.Y(n_1508)
);

AND2x2_ASAP7_75t_L g1509 ( 
.A(n_1461),
.B(n_1361),
.Y(n_1509)
);

BUFx3_ASAP7_75t_L g1510 ( 
.A(n_1461),
.Y(n_1510)
);

AOI21x1_ASAP7_75t_L g1511 ( 
.A1(n_1445),
.A2(n_1423),
.B(n_1422),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_1359),
.Y(n_1512)
);

OR2x2_ASAP7_75t_L g1513 ( 
.A(n_1389),
.B(n_1396),
.Y(n_1513)
);

INVx1_ASAP7_75t_L g1514 ( 
.A(n_1362),
.Y(n_1514)
);

AND2x2_ASAP7_75t_L g1515 ( 
.A(n_1376),
.B(n_1366),
.Y(n_1515)
);

INVx1_ASAP7_75t_L g1516 ( 
.A(n_1371),
.Y(n_1516)
);

INVx1_ASAP7_75t_L g1517 ( 
.A(n_1374),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_1391),
.Y(n_1518)
);

AND2x2_ASAP7_75t_L g1519 ( 
.A(n_1375),
.B(n_1377),
.Y(n_1519)
);

AND2x2_ASAP7_75t_L g1520 ( 
.A(n_1386),
.B(n_1460),
.Y(n_1520)
);

AND2x2_ASAP7_75t_L g1521 ( 
.A(n_1462),
.B(n_1466),
.Y(n_1521)
);

AND2x2_ASAP7_75t_L g1522 ( 
.A(n_1404),
.B(n_1412),
.Y(n_1522)
);

HB1xp67_ASAP7_75t_L g1523 ( 
.A(n_1393),
.Y(n_1523)
);

OR2x2_ASAP7_75t_L g1524 ( 
.A(n_1427),
.B(n_1346),
.Y(n_1524)
);

HB1xp67_ASAP7_75t_L g1525 ( 
.A(n_1408),
.Y(n_1525)
);

HB1xp67_ASAP7_75t_SL g1526 ( 
.A(n_1348),
.Y(n_1526)
);

AND2x2_ASAP7_75t_L g1527 ( 
.A(n_1414),
.B(n_1441),
.Y(n_1527)
);

INVx2_ASAP7_75t_SL g1528 ( 
.A(n_1424),
.Y(n_1528)
);

INVx1_ASAP7_75t_L g1529 ( 
.A(n_1383),
.Y(n_1529)
);

AND2x4_ASAP7_75t_L g1530 ( 
.A(n_1459),
.B(n_1399),
.Y(n_1530)
);

AOI21x1_ASAP7_75t_L g1531 ( 
.A1(n_1457),
.A2(n_1459),
.B(n_1447),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1459),
.Y(n_1532)
);

AND2x2_ASAP7_75t_L g1533 ( 
.A(n_1417),
.B(n_1459),
.Y(n_1533)
);

AOI21xp5_ASAP7_75t_SL g1534 ( 
.A1(n_1395),
.A2(n_1360),
.B(n_1368),
.Y(n_1534)
);

OA21x2_ASAP7_75t_L g1535 ( 
.A1(n_1385),
.A2(n_1378),
.B(n_1454),
.Y(n_1535)
);

INVx2_ASAP7_75t_L g1536 ( 
.A(n_1434),
.Y(n_1536)
);

INVxp67_ASAP7_75t_L g1537 ( 
.A(n_1488),
.Y(n_1537)
);

AOI22xp5_ASAP7_75t_L g1538 ( 
.A1(n_1494),
.A2(n_1429),
.B1(n_1426),
.B2(n_1432),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1497),
.B(n_1457),
.Y(n_1539)
);

INVx2_ASAP7_75t_L g1540 ( 
.A(n_1479),
.Y(n_1540)
);

AOI22xp5_ASAP7_75t_L g1541 ( 
.A1(n_1494),
.A2(n_1436),
.B1(n_1438),
.B2(n_1448),
.Y(n_1541)
);

AND2x2_ASAP7_75t_L g1542 ( 
.A(n_1471),
.B(n_1456),
.Y(n_1542)
);

AND2x2_ASAP7_75t_L g1543 ( 
.A(n_1471),
.B(n_1456),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_1503),
.Y(n_1544)
);

INVx1_ASAP7_75t_L g1545 ( 
.A(n_1503),
.Y(n_1545)
);

HB1xp67_ASAP7_75t_L g1546 ( 
.A(n_1518),
.Y(n_1546)
);

AND2x2_ASAP7_75t_L g1547 ( 
.A(n_1476),
.B(n_1455),
.Y(n_1547)
);

OAI22xp5_ASAP7_75t_L g1548 ( 
.A1(n_1501),
.A2(n_1413),
.B1(n_1440),
.B2(n_1348),
.Y(n_1548)
);

AND2x2_ASAP7_75t_L g1549 ( 
.A(n_1476),
.B(n_1450),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_1504),
.Y(n_1550)
);

INVx2_ASAP7_75t_SL g1551 ( 
.A(n_1499),
.Y(n_1551)
);

INVx1_ASAP7_75t_L g1552 ( 
.A(n_1504),
.Y(n_1552)
);

BUFx6f_ASAP7_75t_L g1553 ( 
.A(n_1530),
.Y(n_1553)
);

AND2x2_ASAP7_75t_L g1554 ( 
.A(n_1506),
.B(n_1449),
.Y(n_1554)
);

BUFx2_ASAP7_75t_L g1555 ( 
.A(n_1499),
.Y(n_1555)
);

AOI22xp33_ASAP7_75t_L g1556 ( 
.A1(n_1533),
.A2(n_1430),
.B1(n_1433),
.B2(n_1435),
.Y(n_1556)
);

AND2x2_ASAP7_75t_L g1557 ( 
.A(n_1506),
.B(n_1449),
.Y(n_1557)
);

AND2x2_ASAP7_75t_L g1558 ( 
.A(n_1484),
.B(n_1449),
.Y(n_1558)
);

INVxp67_ASAP7_75t_L g1559 ( 
.A(n_1473),
.Y(n_1559)
);

AND2x4_ASAP7_75t_SL g1560 ( 
.A(n_1530),
.B(n_1508),
.Y(n_1560)
);

OAI211xp5_ASAP7_75t_SL g1561 ( 
.A1(n_1486),
.A2(n_1439),
.B(n_1443),
.C(n_1452),
.Y(n_1561)
);

AOI221xp5_ASAP7_75t_L g1562 ( 
.A1(n_1515),
.A2(n_1356),
.B1(n_1458),
.B2(n_1446),
.C(n_1442),
.Y(n_1562)
);

OR2x2_ASAP7_75t_L g1563 ( 
.A(n_1495),
.B(n_1507),
.Y(n_1563)
);

AND2x2_ASAP7_75t_L g1564 ( 
.A(n_1495),
.B(n_1509),
.Y(n_1564)
);

OAI22xp5_ASAP7_75t_L g1565 ( 
.A1(n_1526),
.A2(n_1413),
.B1(n_1458),
.B2(n_1356),
.Y(n_1565)
);

AND2x2_ASAP7_75t_L g1566 ( 
.A(n_1509),
.B(n_1453),
.Y(n_1566)
);

OAI21xp33_ASAP7_75t_SL g1567 ( 
.A1(n_1534),
.A2(n_1453),
.B(n_1428),
.Y(n_1567)
);

AND2x2_ASAP7_75t_L g1568 ( 
.A(n_1519),
.B(n_1453),
.Y(n_1568)
);

OAI22xp5_ASAP7_75t_L g1569 ( 
.A1(n_1526),
.A2(n_1356),
.B1(n_1451),
.B2(n_1444),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_L g1570 ( 
.A(n_1523),
.B(n_1368),
.Y(n_1570)
);

OR2x2_ASAP7_75t_L g1571 ( 
.A(n_1510),
.B(n_1513),
.Y(n_1571)
);

AND2x2_ASAP7_75t_L g1572 ( 
.A(n_1519),
.B(n_1400),
.Y(n_1572)
);

INVx1_ASAP7_75t_SL g1573 ( 
.A(n_1483),
.Y(n_1573)
);

HB1xp67_ASAP7_75t_L g1574 ( 
.A(n_1525),
.Y(n_1574)
);

HB1xp67_ASAP7_75t_L g1575 ( 
.A(n_1500),
.Y(n_1575)
);

NAND2xp5_ASAP7_75t_L g1576 ( 
.A(n_1520),
.B(n_1451),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1520),
.B(n_1400),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1500),
.Y(n_1578)
);

HB1xp67_ASAP7_75t_L g1579 ( 
.A(n_1502),
.Y(n_1579)
);

AND2x2_ASAP7_75t_L g1580 ( 
.A(n_1521),
.B(n_1400),
.Y(n_1580)
);

BUFx2_ASAP7_75t_L g1581 ( 
.A(n_1483),
.Y(n_1581)
);

OR2x2_ASAP7_75t_L g1582 ( 
.A(n_1513),
.B(n_1437),
.Y(n_1582)
);

INVx3_ASAP7_75t_L g1583 ( 
.A(n_1482),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1489),
.B(n_1437),
.Y(n_1584)
);

AND2x4_ASAP7_75t_L g1585 ( 
.A(n_1532),
.B(n_1493),
.Y(n_1585)
);

AOI22xp33_ASAP7_75t_L g1586 ( 
.A1(n_1548),
.A2(n_1533),
.B1(n_1490),
.B2(n_1535),
.Y(n_1586)
);

NAND2xp5_ASAP7_75t_L g1587 ( 
.A(n_1546),
.B(n_1490),
.Y(n_1587)
);

AOI22xp33_ASAP7_75t_L g1588 ( 
.A1(n_1548),
.A2(n_1490),
.B1(n_1535),
.B2(n_1527),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1574),
.B(n_1490),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1564),
.B(n_1480),
.Y(n_1590)
);

NAND2xp5_ASAP7_75t_L g1591 ( 
.A(n_1564),
.B(n_1480),
.Y(n_1591)
);

NAND2xp5_ASAP7_75t_L g1592 ( 
.A(n_1537),
.B(n_1563),
.Y(n_1592)
);

AOI22xp33_ASAP7_75t_SL g1593 ( 
.A1(n_1559),
.A2(n_1535),
.B1(n_1474),
.B2(n_1477),
.Y(n_1593)
);

NAND2xp5_ASAP7_75t_L g1594 ( 
.A(n_1563),
.B(n_1478),
.Y(n_1594)
);

INVx2_ASAP7_75t_SL g1595 ( 
.A(n_1581),
.Y(n_1595)
);

NAND3xp33_ASAP7_75t_L g1596 ( 
.A(n_1538),
.B(n_1489),
.C(n_1478),
.Y(n_1596)
);

AOI22xp33_ASAP7_75t_L g1597 ( 
.A1(n_1556),
.A2(n_1535),
.B1(n_1527),
.B2(n_1522),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1565),
.B(n_1439),
.Y(n_1598)
);

INVx1_ASAP7_75t_L g1599 ( 
.A(n_1544),
.Y(n_1599)
);

AND2x2_ASAP7_75t_L g1600 ( 
.A(n_1554),
.B(n_1557),
.Y(n_1600)
);

INVx2_ASAP7_75t_L g1601 ( 
.A(n_1540),
.Y(n_1601)
);

AND2x2_ASAP7_75t_L g1602 ( 
.A(n_1554),
.B(n_1505),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_L g1603 ( 
.A(n_1547),
.B(n_1496),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1547),
.B(n_1496),
.Y(n_1604)
);

NAND2xp5_ASAP7_75t_L g1605 ( 
.A(n_1542),
.B(n_1498),
.Y(n_1605)
);

AOI22xp33_ASAP7_75t_L g1606 ( 
.A1(n_1541),
.A2(n_1535),
.B1(n_1522),
.B2(n_1536),
.Y(n_1606)
);

NAND2xp5_ASAP7_75t_L g1607 ( 
.A(n_1542),
.B(n_1543),
.Y(n_1607)
);

OAI21xp5_ASAP7_75t_SL g1608 ( 
.A1(n_1562),
.A2(n_1538),
.B(n_1561),
.Y(n_1608)
);

NAND2xp5_ASAP7_75t_L g1609 ( 
.A(n_1543),
.B(n_1498),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1573),
.B(n_1491),
.Y(n_1610)
);

NAND2xp5_ASAP7_75t_L g1611 ( 
.A(n_1573),
.B(n_1491),
.Y(n_1611)
);

NAND2xp5_ASAP7_75t_L g1612 ( 
.A(n_1539),
.B(n_1512),
.Y(n_1612)
);

AND2x2_ASAP7_75t_L g1613 ( 
.A(n_1557),
.B(n_1549),
.Y(n_1613)
);

OAI21xp5_ASAP7_75t_SL g1614 ( 
.A1(n_1569),
.A2(n_1511),
.B(n_1531),
.Y(n_1614)
);

NAND3xp33_ASAP7_75t_L g1615 ( 
.A(n_1584),
.B(n_1516),
.C(n_1514),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1549),
.B(n_1571),
.Y(n_1616)
);

AOI21xp5_ASAP7_75t_L g1617 ( 
.A1(n_1567),
.A2(n_1534),
.B(n_1528),
.Y(n_1617)
);

AND2x2_ASAP7_75t_L g1618 ( 
.A(n_1572),
.B(n_1505),
.Y(n_1618)
);

AND2x4_ASAP7_75t_L g1619 ( 
.A(n_1585),
.B(n_1531),
.Y(n_1619)
);

NAND2xp5_ASAP7_75t_L g1620 ( 
.A(n_1571),
.B(n_1512),
.Y(n_1620)
);

AND2x2_ASAP7_75t_L g1621 ( 
.A(n_1577),
.B(n_1481),
.Y(n_1621)
);

NAND4xp25_ASAP7_75t_L g1622 ( 
.A(n_1541),
.B(n_1517),
.C(n_1516),
.D(n_1524),
.Y(n_1622)
);

OAI22xp5_ASAP7_75t_L g1623 ( 
.A1(n_1570),
.A2(n_1511),
.B1(n_1517),
.B2(n_1468),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1568),
.B(n_1524),
.Y(n_1624)
);

NAND2xp5_ASAP7_75t_L g1625 ( 
.A(n_1568),
.B(n_1492),
.Y(n_1625)
);

OA21x2_ASAP7_75t_L g1626 ( 
.A1(n_1540),
.A2(n_1472),
.B(n_1475),
.Y(n_1626)
);

NAND2xp5_ASAP7_75t_L g1627 ( 
.A(n_1577),
.B(n_1492),
.Y(n_1627)
);

AND2x2_ASAP7_75t_SL g1628 ( 
.A(n_1560),
.B(n_1508),
.Y(n_1628)
);

NAND2xp5_ASAP7_75t_L g1629 ( 
.A(n_1580),
.B(n_1492),
.Y(n_1629)
);

NAND3xp33_ASAP7_75t_L g1630 ( 
.A(n_1575),
.B(n_1485),
.C(n_1487),
.Y(n_1630)
);

NOR2xp67_ASAP7_75t_L g1631 ( 
.A(n_1583),
.B(n_1528),
.Y(n_1631)
);

NAND2xp5_ASAP7_75t_L g1632 ( 
.A(n_1558),
.B(n_1578),
.Y(n_1632)
);

NOR2xp33_ASAP7_75t_L g1633 ( 
.A(n_1576),
.B(n_1381),
.Y(n_1633)
);

AND2x2_ASAP7_75t_L g1634 ( 
.A(n_1566),
.B(n_1481),
.Y(n_1634)
);

NAND2xp5_ASAP7_75t_SL g1635 ( 
.A(n_1567),
.B(n_1469),
.Y(n_1635)
);

OAI21xp5_ASAP7_75t_SL g1636 ( 
.A1(n_1560),
.A2(n_1482),
.B(n_1529),
.Y(n_1636)
);

OAI211xp5_ASAP7_75t_SL g1637 ( 
.A1(n_1583),
.A2(n_1443),
.B(n_1468),
.C(n_1470),
.Y(n_1637)
);

NAND2xp5_ASAP7_75t_L g1638 ( 
.A(n_1558),
.B(n_1492),
.Y(n_1638)
);

AND2x4_ASAP7_75t_L g1639 ( 
.A(n_1619),
.B(n_1583),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1587),
.B(n_1579),
.Y(n_1640)
);

INVx1_ASAP7_75t_L g1641 ( 
.A(n_1599),
.Y(n_1641)
);

INVx2_ASAP7_75t_L g1642 ( 
.A(n_1626),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1599),
.Y(n_1643)
);

INVx2_ASAP7_75t_L g1644 ( 
.A(n_1626),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1634),
.B(n_1555),
.Y(n_1645)
);

NAND2xp5_ASAP7_75t_L g1646 ( 
.A(n_1589),
.B(n_1544),
.Y(n_1646)
);

INVxp67_ASAP7_75t_L g1647 ( 
.A(n_1623),
.Y(n_1647)
);

NAND2xp5_ASAP7_75t_L g1648 ( 
.A(n_1621),
.B(n_1545),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1626),
.Y(n_1649)
);

INVx2_ASAP7_75t_SL g1650 ( 
.A(n_1628),
.Y(n_1650)
);

OR2x2_ASAP7_75t_L g1651 ( 
.A(n_1638),
.B(n_1625),
.Y(n_1651)
);

INVx2_ASAP7_75t_L g1652 ( 
.A(n_1626),
.Y(n_1652)
);

INVx1_ASAP7_75t_L g1653 ( 
.A(n_1620),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1615),
.Y(n_1654)
);

OR2x2_ASAP7_75t_L g1655 ( 
.A(n_1627),
.B(n_1629),
.Y(n_1655)
);

OR2x2_ASAP7_75t_L g1656 ( 
.A(n_1594),
.B(n_1590),
.Y(n_1656)
);

AND2x2_ASAP7_75t_L g1657 ( 
.A(n_1613),
.B(n_1600),
.Y(n_1657)
);

INVx2_ASAP7_75t_L g1658 ( 
.A(n_1601),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1615),
.Y(n_1659)
);

NAND2xp5_ASAP7_75t_L g1660 ( 
.A(n_1610),
.B(n_1545),
.Y(n_1660)
);

INVx1_ASAP7_75t_SL g1661 ( 
.A(n_1595),
.Y(n_1661)
);

AND2x4_ASAP7_75t_L g1662 ( 
.A(n_1619),
.B(n_1583),
.Y(n_1662)
);

NOR2x1_ASAP7_75t_SL g1663 ( 
.A(n_1635),
.B(n_1553),
.Y(n_1663)
);

OR2x2_ASAP7_75t_L g1664 ( 
.A(n_1591),
.B(n_1592),
.Y(n_1664)
);

NAND2xp5_ASAP7_75t_SL g1665 ( 
.A(n_1628),
.B(n_1551),
.Y(n_1665)
);

HB1xp67_ASAP7_75t_L g1666 ( 
.A(n_1630),
.Y(n_1666)
);

BUFx2_ASAP7_75t_L g1667 ( 
.A(n_1628),
.Y(n_1667)
);

HB1xp67_ASAP7_75t_L g1668 ( 
.A(n_1630),
.Y(n_1668)
);

OR2x2_ASAP7_75t_L g1669 ( 
.A(n_1595),
.B(n_1582),
.Y(n_1669)
);

OR2x2_ASAP7_75t_L g1670 ( 
.A(n_1612),
.B(n_1550),
.Y(n_1670)
);

NAND2xp5_ASAP7_75t_L g1671 ( 
.A(n_1611),
.B(n_1550),
.Y(n_1671)
);

INVx2_ASAP7_75t_L g1672 ( 
.A(n_1619),
.Y(n_1672)
);

HB1xp67_ASAP7_75t_L g1673 ( 
.A(n_1632),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1605),
.Y(n_1674)
);

NAND2x1p5_ASAP7_75t_L g1675 ( 
.A(n_1617),
.B(n_1508),
.Y(n_1675)
);

HB1xp67_ASAP7_75t_L g1676 ( 
.A(n_1602),
.Y(n_1676)
);

NOR2x1p5_ASAP7_75t_SL g1677 ( 
.A(n_1642),
.B(n_1644),
.Y(n_1677)
);

INVx1_ASAP7_75t_L g1678 ( 
.A(n_1641),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1654),
.B(n_1659),
.Y(n_1679)
);

INVx1_ASAP7_75t_L g1680 ( 
.A(n_1641),
.Y(n_1680)
);

NAND2xp5_ASAP7_75t_L g1681 ( 
.A(n_1654),
.B(n_1603),
.Y(n_1681)
);

INVx1_ASAP7_75t_L g1682 ( 
.A(n_1643),
.Y(n_1682)
);

INVx3_ASAP7_75t_L g1683 ( 
.A(n_1639),
.Y(n_1683)
);

NOR3x1_ASAP7_75t_L g1684 ( 
.A(n_1667),
.B(n_1608),
.C(n_1636),
.Y(n_1684)
);

OR2x6_ASAP7_75t_L g1685 ( 
.A(n_1675),
.B(n_1596),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1643),
.Y(n_1686)
);

INVx1_ASAP7_75t_SL g1687 ( 
.A(n_1661),
.Y(n_1687)
);

INVx1_ASAP7_75t_L g1688 ( 
.A(n_1670),
.Y(n_1688)
);

INVx2_ASAP7_75t_SL g1689 ( 
.A(n_1669),
.Y(n_1689)
);

INVx2_ASAP7_75t_L g1690 ( 
.A(n_1658),
.Y(n_1690)
);

AND2x2_ASAP7_75t_L g1691 ( 
.A(n_1657),
.B(n_1618),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_L g1692 ( 
.A(n_1659),
.B(n_1604),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1653),
.B(n_1609),
.Y(n_1693)
);

AOI22xp5_ASAP7_75t_L g1694 ( 
.A1(n_1647),
.A2(n_1622),
.B1(n_1596),
.B2(n_1593),
.Y(n_1694)
);

OR2x2_ASAP7_75t_L g1695 ( 
.A(n_1648),
.B(n_1664),
.Y(n_1695)
);

INVxp33_ASAP7_75t_L g1696 ( 
.A(n_1663),
.Y(n_1696)
);

INVx1_ASAP7_75t_L g1697 ( 
.A(n_1670),
.Y(n_1697)
);

INVx2_ASAP7_75t_L g1698 ( 
.A(n_1658),
.Y(n_1698)
);

INVx1_ASAP7_75t_L g1699 ( 
.A(n_1670),
.Y(n_1699)
);

AOI211xp5_ASAP7_75t_L g1700 ( 
.A1(n_1647),
.A2(n_1622),
.B(n_1614),
.C(n_1636),
.Y(n_1700)
);

NAND2xp5_ASAP7_75t_L g1701 ( 
.A(n_1653),
.B(n_1624),
.Y(n_1701)
);

INVx1_ASAP7_75t_L g1702 ( 
.A(n_1660),
.Y(n_1702)
);

AND2x2_ASAP7_75t_L g1703 ( 
.A(n_1657),
.B(n_1602),
.Y(n_1703)
);

AND2x2_ASAP7_75t_L g1704 ( 
.A(n_1657),
.B(n_1633),
.Y(n_1704)
);

OR2x2_ASAP7_75t_L g1705 ( 
.A(n_1648),
.B(n_1616),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1660),
.Y(n_1706)
);

INVx1_ASAP7_75t_L g1707 ( 
.A(n_1671),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1671),
.Y(n_1708)
);

OAI21xp33_ASAP7_75t_L g1709 ( 
.A1(n_1666),
.A2(n_1668),
.B(n_1640),
.Y(n_1709)
);

INVx1_ASAP7_75t_L g1710 ( 
.A(n_1674),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1658),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1674),
.Y(n_1712)
);

NAND2xp5_ASAP7_75t_L g1713 ( 
.A(n_1673),
.B(n_1552),
.Y(n_1713)
);

AOI211xp5_ASAP7_75t_L g1714 ( 
.A1(n_1666),
.A2(n_1598),
.B(n_1637),
.C(n_1631),
.Y(n_1714)
);

OR2x2_ASAP7_75t_L g1715 ( 
.A(n_1664),
.B(n_1607),
.Y(n_1715)
);

AND2x2_ASAP7_75t_L g1716 ( 
.A(n_1667),
.B(n_1551),
.Y(n_1716)
);

NAND2xp5_ASAP7_75t_L g1717 ( 
.A(n_1679),
.B(n_1668),
.Y(n_1717)
);

AND2x4_ASAP7_75t_L g1718 ( 
.A(n_1685),
.B(n_1663),
.Y(n_1718)
);

HB1xp67_ASAP7_75t_L g1719 ( 
.A(n_1710),
.Y(n_1719)
);

AND2x2_ASAP7_75t_L g1720 ( 
.A(n_1684),
.B(n_1672),
.Y(n_1720)
);

INVx1_ASAP7_75t_L g1721 ( 
.A(n_1678),
.Y(n_1721)
);

INVx1_ASAP7_75t_L g1722 ( 
.A(n_1678),
.Y(n_1722)
);

AND2x2_ASAP7_75t_L g1723 ( 
.A(n_1691),
.B(n_1667),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_L g1724 ( 
.A(n_1712),
.B(n_1646),
.Y(n_1724)
);

INVx2_ASAP7_75t_L g1725 ( 
.A(n_1690),
.Y(n_1725)
);

AND2x2_ASAP7_75t_L g1726 ( 
.A(n_1691),
.B(n_1672),
.Y(n_1726)
);

INVxp67_ASAP7_75t_SL g1727 ( 
.A(n_1694),
.Y(n_1727)
);

INVx1_ASAP7_75t_L g1728 ( 
.A(n_1686),
.Y(n_1728)
);

INVx2_ASAP7_75t_L g1729 ( 
.A(n_1690),
.Y(n_1729)
);

BUFx2_ASAP7_75t_L g1730 ( 
.A(n_1685),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1686),
.Y(n_1731)
);

INVx1_ASAP7_75t_L g1732 ( 
.A(n_1680),
.Y(n_1732)
);

OR2x2_ASAP7_75t_L g1733 ( 
.A(n_1695),
.B(n_1640),
.Y(n_1733)
);

HB1xp67_ASAP7_75t_L g1734 ( 
.A(n_1688),
.Y(n_1734)
);

AND2x2_ASAP7_75t_L g1735 ( 
.A(n_1700),
.B(n_1672),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1709),
.A2(n_1586),
.B1(n_1588),
.B2(n_1606),
.Y(n_1736)
);

AND2x2_ASAP7_75t_L g1737 ( 
.A(n_1703),
.B(n_1672),
.Y(n_1737)
);

INVx1_ASAP7_75t_L g1738 ( 
.A(n_1682),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1703),
.B(n_1696),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1702),
.B(n_1646),
.Y(n_1740)
);

AND2x2_ASAP7_75t_L g1741 ( 
.A(n_1696),
.B(n_1639),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1697),
.Y(n_1742)
);

NOR2xp33_ASAP7_75t_L g1743 ( 
.A(n_1704),
.B(n_1406),
.Y(n_1743)
);

AND2x4_ASAP7_75t_L g1744 ( 
.A(n_1685),
.B(n_1650),
.Y(n_1744)
);

AND2x2_ASAP7_75t_L g1745 ( 
.A(n_1685),
.B(n_1639),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1746)
);

AND2x2_ASAP7_75t_L g1747 ( 
.A(n_1683),
.B(n_1639),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1697),
.Y(n_1748)
);

AND2x2_ASAP7_75t_L g1749 ( 
.A(n_1704),
.B(n_1676),
.Y(n_1749)
);

AND2x2_ASAP7_75t_L g1750 ( 
.A(n_1683),
.B(n_1689),
.Y(n_1750)
);

INVx1_ASAP7_75t_SL g1751 ( 
.A(n_1687),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1713),
.Y(n_1752)
);

NAND2xp5_ASAP7_75t_L g1753 ( 
.A(n_1706),
.B(n_1656),
.Y(n_1753)
);

NAND2xp5_ASAP7_75t_L g1754 ( 
.A(n_1707),
.B(n_1656),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1699),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1693),
.Y(n_1756)
);

INVx1_ASAP7_75t_L g1757 ( 
.A(n_1708),
.Y(n_1757)
);

AND2x2_ASAP7_75t_L g1758 ( 
.A(n_1689),
.B(n_1662),
.Y(n_1758)
);

OR2x2_ASAP7_75t_L g1759 ( 
.A(n_1695),
.B(n_1664),
.Y(n_1759)
);

AND2x4_ASAP7_75t_L g1760 ( 
.A(n_1677),
.B(n_1650),
.Y(n_1760)
);

INVxp33_ASAP7_75t_SL g1761 ( 
.A(n_1743),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1727),
.B(n_1681),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1750),
.Y(n_1763)
);

INVxp67_ASAP7_75t_SL g1764 ( 
.A(n_1727),
.Y(n_1764)
);

AO21x2_ASAP7_75t_L g1765 ( 
.A1(n_1717),
.A2(n_1644),
.B(n_1642),
.Y(n_1765)
);

INVx3_ASAP7_75t_L g1766 ( 
.A(n_1718),
.Y(n_1766)
);

BUFx3_ASAP7_75t_L g1767 ( 
.A(n_1751),
.Y(n_1767)
);

OR2x2_ASAP7_75t_L g1768 ( 
.A(n_1759),
.B(n_1692),
.Y(n_1768)
);

CKINVDCx16_ASAP7_75t_R g1769 ( 
.A(n_1751),
.Y(n_1769)
);

INVx1_ASAP7_75t_SL g1770 ( 
.A(n_1730),
.Y(n_1770)
);

NOR2xp33_ASAP7_75t_L g1771 ( 
.A(n_1759),
.B(n_1406),
.Y(n_1771)
);

HB1xp67_ASAP7_75t_L g1772 ( 
.A(n_1719),
.Y(n_1772)
);

INVx1_ASAP7_75t_L g1773 ( 
.A(n_1721),
.Y(n_1773)
);

AND2x2_ASAP7_75t_L g1774 ( 
.A(n_1749),
.B(n_1716),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1721),
.Y(n_1775)
);

NAND2xp5_ASAP7_75t_L g1776 ( 
.A(n_1756),
.B(n_1715),
.Y(n_1776)
);

NOR2x1p5_ASAP7_75t_L g1777 ( 
.A(n_1718),
.B(n_1720),
.Y(n_1777)
);

AND2x2_ASAP7_75t_L g1778 ( 
.A(n_1749),
.B(n_1716),
.Y(n_1778)
);

INVx3_ASAP7_75t_L g1779 ( 
.A(n_1718),
.Y(n_1779)
);

AND2x4_ASAP7_75t_L g1780 ( 
.A(n_1718),
.B(n_1744),
.Y(n_1780)
);

BUFx2_ASAP7_75t_L g1781 ( 
.A(n_1735),
.Y(n_1781)
);

AOI22xp33_ASAP7_75t_L g1782 ( 
.A1(n_1736),
.A2(n_1597),
.B1(n_1655),
.B2(n_1651),
.Y(n_1782)
);

NAND2xp5_ASAP7_75t_L g1783 ( 
.A(n_1756),
.B(n_1715),
.Y(n_1783)
);

AOI22xp33_ASAP7_75t_L g1784 ( 
.A1(n_1735),
.A2(n_1655),
.B1(n_1651),
.B2(n_1649),
.Y(n_1784)
);

INVx2_ASAP7_75t_SL g1785 ( 
.A(n_1718),
.Y(n_1785)
);

NAND2xp5_ASAP7_75t_SL g1786 ( 
.A(n_1744),
.B(n_1714),
.Y(n_1786)
);

AND2x2_ASAP7_75t_L g1787 ( 
.A(n_1739),
.B(n_1662),
.Y(n_1787)
);

INVx1_ASAP7_75t_L g1788 ( 
.A(n_1722),
.Y(n_1788)
);

INVx3_ASAP7_75t_L g1789 ( 
.A(n_1744),
.Y(n_1789)
);

CKINVDCx16_ASAP7_75t_R g1790 ( 
.A(n_1735),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_L g1791 ( 
.A(n_1752),
.B(n_1757),
.Y(n_1791)
);

AOI22x1_ASAP7_75t_L g1792 ( 
.A1(n_1730),
.A2(n_1381),
.B1(n_1380),
.B2(n_1650),
.Y(n_1792)
);

AND2x2_ASAP7_75t_L g1793 ( 
.A(n_1739),
.B(n_1662),
.Y(n_1793)
);

OR2x6_ASAP7_75t_L g1794 ( 
.A(n_1760),
.B(n_1677),
.Y(n_1794)
);

HB1xp67_ASAP7_75t_L g1795 ( 
.A(n_1734),
.Y(n_1795)
);

OR2x2_ASAP7_75t_L g1796 ( 
.A(n_1717),
.B(n_1705),
.Y(n_1796)
);

INVx2_ASAP7_75t_L g1797 ( 
.A(n_1767),
.Y(n_1797)
);

AOI22xp5_ASAP7_75t_L g1798 ( 
.A1(n_1790),
.A2(n_1720),
.B1(n_1760),
.B2(n_1739),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1769),
.B(n_1752),
.Y(n_1799)
);

AOI21xp5_ASAP7_75t_L g1800 ( 
.A1(n_1764),
.A2(n_1720),
.B(n_1744),
.Y(n_1800)
);

NAND2xp5_ASAP7_75t_L g1801 ( 
.A(n_1769),
.B(n_1755),
.Y(n_1801)
);

OAI31xp33_ASAP7_75t_L g1802 ( 
.A1(n_1764),
.A2(n_1760),
.A3(n_1744),
.B(n_1745),
.Y(n_1802)
);

OR2x2_ASAP7_75t_L g1803 ( 
.A(n_1781),
.B(n_1733),
.Y(n_1803)
);

INVx1_ASAP7_75t_L g1804 ( 
.A(n_1773),
.Y(n_1804)
);

INVx2_ASAP7_75t_L g1805 ( 
.A(n_1767),
.Y(n_1805)
);

INVx1_ASAP7_75t_L g1806 ( 
.A(n_1773),
.Y(n_1806)
);

OAI22xp5_ASAP7_75t_L g1807 ( 
.A1(n_1790),
.A2(n_1745),
.B1(n_1723),
.B2(n_1760),
.Y(n_1807)
);

AOI221xp5_ASAP7_75t_L g1808 ( 
.A1(n_1781),
.A2(n_1760),
.B1(n_1642),
.B2(n_1652),
.C(n_1649),
.Y(n_1808)
);

AOI22xp5_ASAP7_75t_L g1809 ( 
.A1(n_1782),
.A2(n_1725),
.B1(n_1729),
.B2(n_1755),
.Y(n_1809)
);

INVxp67_ASAP7_75t_L g1810 ( 
.A(n_1767),
.Y(n_1810)
);

INVx1_ASAP7_75t_L g1811 ( 
.A(n_1775),
.Y(n_1811)
);

OAI22xp33_ASAP7_75t_L g1812 ( 
.A1(n_1762),
.A2(n_1733),
.B1(n_1757),
.B2(n_1675),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1775),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1788),
.Y(n_1814)
);

INVx1_ASAP7_75t_L g1815 ( 
.A(n_1788),
.Y(n_1815)
);

INVx2_ASAP7_75t_SL g1816 ( 
.A(n_1777),
.Y(n_1816)
);

OAI21xp5_ASAP7_75t_L g1817 ( 
.A1(n_1786),
.A2(n_1750),
.B(n_1745),
.Y(n_1817)
);

INVx1_ASAP7_75t_L g1818 ( 
.A(n_1795),
.Y(n_1818)
);

INVx1_ASAP7_75t_SL g1819 ( 
.A(n_1761),
.Y(n_1819)
);

NAND2xp33_ASAP7_75t_SL g1820 ( 
.A(n_1777),
.B(n_1750),
.Y(n_1820)
);

OAI22xp33_ASAP7_75t_SL g1821 ( 
.A1(n_1794),
.A2(n_1762),
.B1(n_1785),
.B2(n_1770),
.Y(n_1821)
);

OAI221xp5_ASAP7_75t_L g1822 ( 
.A1(n_1784),
.A2(n_1742),
.B1(n_1748),
.B2(n_1652),
.C(n_1644),
.Y(n_1822)
);

NOR2xp33_ASAP7_75t_L g1823 ( 
.A(n_1819),
.B(n_1771),
.Y(n_1823)
);

NAND2xp5_ASAP7_75t_L g1824 ( 
.A(n_1810),
.B(n_1770),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1810),
.Y(n_1825)
);

OR2x2_ASAP7_75t_L g1826 ( 
.A(n_1803),
.B(n_1768),
.Y(n_1826)
);

NAND2xp5_ASAP7_75t_L g1827 ( 
.A(n_1797),
.B(n_1772),
.Y(n_1827)
);

AO21x1_ASAP7_75t_L g1828 ( 
.A1(n_1821),
.A2(n_1780),
.B(n_1791),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_L g1829 ( 
.A(n_1805),
.B(n_1763),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1800),
.B(n_1763),
.Y(n_1830)
);

NOR2xp67_ASAP7_75t_SL g1831 ( 
.A(n_1801),
.B(n_1380),
.Y(n_1831)
);

AND2x2_ASAP7_75t_L g1832 ( 
.A(n_1817),
.B(n_1774),
.Y(n_1832)
);

INVx1_ASAP7_75t_SL g1833 ( 
.A(n_1820),
.Y(n_1833)
);

NAND2xp5_ASAP7_75t_L g1834 ( 
.A(n_1800),
.B(n_1774),
.Y(n_1834)
);

NAND2xp5_ASAP7_75t_L g1835 ( 
.A(n_1818),
.B(n_1799),
.Y(n_1835)
);

OAI21xp5_ASAP7_75t_SL g1836 ( 
.A1(n_1798),
.A2(n_1780),
.B(n_1789),
.Y(n_1836)
);

INVx1_ASAP7_75t_L g1837 ( 
.A(n_1804),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1806),
.Y(n_1838)
);

NAND2xp33_ASAP7_75t_SL g1839 ( 
.A(n_1816),
.B(n_1785),
.Y(n_1839)
);

NAND2xp5_ASAP7_75t_L g1840 ( 
.A(n_1809),
.B(n_1778),
.Y(n_1840)
);

AND2x2_ASAP7_75t_L g1841 ( 
.A(n_1807),
.B(n_1778),
.Y(n_1841)
);

INVx1_ASAP7_75t_L g1842 ( 
.A(n_1811),
.Y(n_1842)
);

INVx1_ASAP7_75t_L g1843 ( 
.A(n_1824),
.Y(n_1843)
);

AOI211xp5_ASAP7_75t_L g1844 ( 
.A1(n_1828),
.A2(n_1802),
.B(n_1812),
.C(n_1820),
.Y(n_1844)
);

O2A1O1Ixp5_ASAP7_75t_L g1845 ( 
.A1(n_1834),
.A2(n_1839),
.B(n_1830),
.C(n_1840),
.Y(n_1845)
);

AOI221xp5_ASAP7_75t_L g1846 ( 
.A1(n_1833),
.A2(n_1822),
.B1(n_1808),
.B2(n_1835),
.C(n_1812),
.Y(n_1846)
);

NAND4xp25_ASAP7_75t_L g1847 ( 
.A(n_1823),
.B(n_1814),
.C(n_1815),
.D(n_1813),
.Y(n_1847)
);

OAI221xp5_ASAP7_75t_L g1848 ( 
.A1(n_1836),
.A2(n_1794),
.B1(n_1785),
.B2(n_1779),
.C(n_1766),
.Y(n_1848)
);

NOR4xp75_ASAP7_75t_L g1849 ( 
.A(n_1827),
.B(n_1829),
.C(n_1841),
.D(n_1832),
.Y(n_1849)
);

AOI221xp5_ASAP7_75t_L g1850 ( 
.A1(n_1837),
.A2(n_1765),
.B1(n_1791),
.B2(n_1789),
.C(n_1776),
.Y(n_1850)
);

AOI22xp5_ASAP7_75t_L g1851 ( 
.A1(n_1823),
.A2(n_1794),
.B1(n_1765),
.B2(n_1780),
.Y(n_1851)
);

AOI211xp5_ASAP7_75t_L g1852 ( 
.A1(n_1839),
.A2(n_1780),
.B(n_1766),
.C(n_1779),
.Y(n_1852)
);

NOR3xp33_ASAP7_75t_L g1853 ( 
.A(n_1825),
.B(n_1789),
.C(n_1779),
.Y(n_1853)
);

OAI22xp5_ASAP7_75t_L g1854 ( 
.A1(n_1826),
.A2(n_1794),
.B1(n_1792),
.B2(n_1789),
.Y(n_1854)
);

AND4x1_ASAP7_75t_L g1855 ( 
.A(n_1845),
.B(n_1831),
.C(n_1841),
.D(n_1838),
.Y(n_1855)
);

NAND4xp25_ASAP7_75t_SL g1856 ( 
.A(n_1844),
.B(n_1842),
.C(n_1787),
.D(n_1793),
.Y(n_1856)
);

AOI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1846),
.A2(n_1794),
.B(n_1783),
.Y(n_1857)
);

NAND4xp75_ASAP7_75t_L g1858 ( 
.A(n_1843),
.B(n_1783),
.C(n_1776),
.D(n_1787),
.Y(n_1858)
);

NOR3xp33_ASAP7_75t_L g1859 ( 
.A(n_1848),
.B(n_1779),
.C(n_1766),
.Y(n_1859)
);

NAND5xp2_ASAP7_75t_L g1860 ( 
.A(n_1852),
.B(n_1793),
.C(n_1741),
.D(n_1723),
.E(n_1758),
.Y(n_1860)
);

NAND4xp25_ASAP7_75t_L g1861 ( 
.A(n_1853),
.B(n_1850),
.C(n_1847),
.D(n_1851),
.Y(n_1861)
);

INVx1_ASAP7_75t_SL g1862 ( 
.A(n_1849),
.Y(n_1862)
);

AOI211xp5_ASAP7_75t_L g1863 ( 
.A1(n_1854),
.A2(n_1766),
.B(n_1796),
.C(n_1768),
.Y(n_1863)
);

AND2x2_ASAP7_75t_L g1864 ( 
.A(n_1843),
.B(n_1758),
.Y(n_1864)
);

NOR3xp33_ASAP7_75t_L g1865 ( 
.A(n_1845),
.B(n_1796),
.C(n_1729),
.Y(n_1865)
);

AOI22xp33_ASAP7_75t_L g1866 ( 
.A1(n_1856),
.A2(n_1865),
.B1(n_1862),
.B2(n_1857),
.Y(n_1866)
);

NAND3xp33_ASAP7_75t_SL g1867 ( 
.A(n_1855),
.B(n_1741),
.C(n_1758),
.Y(n_1867)
);

NOR2xp67_ASAP7_75t_SL g1868 ( 
.A(n_1858),
.B(n_1402),
.Y(n_1868)
);

AOI211xp5_ASAP7_75t_L g1869 ( 
.A1(n_1861),
.A2(n_1741),
.B(n_1742),
.C(n_1748),
.Y(n_1869)
);

AOI32xp33_ASAP7_75t_L g1870 ( 
.A1(n_1863),
.A2(n_1737),
.A3(n_1726),
.B1(n_1765),
.B2(n_1747),
.Y(n_1870)
);

NOR3xp33_ASAP7_75t_SL g1871 ( 
.A(n_1860),
.B(n_1665),
.C(n_1753),
.Y(n_1871)
);

NOR2xp33_ASAP7_75t_L g1872 ( 
.A(n_1864),
.B(n_1732),
.Y(n_1872)
);

NOR2xp33_ASAP7_75t_R g1873 ( 
.A(n_1859),
.B(n_1732),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_SL g1874 ( 
.A1(n_1873),
.A2(n_1765),
.B1(n_1792),
.B2(n_1729),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1872),
.Y(n_1875)
);

NOR2xp67_ASAP7_75t_L g1876 ( 
.A(n_1867),
.B(n_1722),
.Y(n_1876)
);

INVx1_ASAP7_75t_L g1877 ( 
.A(n_1869),
.Y(n_1877)
);

NAND2xp5_ASAP7_75t_L g1878 ( 
.A(n_1866),
.B(n_1753),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1868),
.A2(n_1725),
.B1(n_1731),
.B2(n_1728),
.Y(n_1879)
);

INVx1_ASAP7_75t_L g1880 ( 
.A(n_1871),
.Y(n_1880)
);

NOR4xp75_ASAP7_75t_L g1881 ( 
.A(n_1878),
.B(n_1870),
.C(n_1754),
.D(n_1747),
.Y(n_1881)
);

CKINVDCx5p33_ASAP7_75t_R g1882 ( 
.A(n_1875),
.Y(n_1882)
);

NAND3xp33_ASAP7_75t_SL g1883 ( 
.A(n_1880),
.B(n_1725),
.C(n_1754),
.Y(n_1883)
);

OAI22xp5_ASAP7_75t_L g1884 ( 
.A1(n_1879),
.A2(n_1731),
.B1(n_1728),
.B2(n_1738),
.Y(n_1884)
);

AND2x4_ASAP7_75t_L g1885 ( 
.A(n_1877),
.B(n_1746),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1876),
.Y(n_1886)
);

XNOR2xp5_ASAP7_75t_L g1887 ( 
.A(n_1881),
.B(n_1874),
.Y(n_1887)
);

AND2x2_ASAP7_75t_L g1888 ( 
.A(n_1885),
.B(n_1726),
.Y(n_1888)
);

AND2x2_ASAP7_75t_L g1889 ( 
.A(n_1882),
.B(n_1746),
.Y(n_1889)
);

OR3x1_ASAP7_75t_L g1890 ( 
.A(n_1887),
.B(n_1886),
.C(n_1883),
.Y(n_1890)
);

OAI221xp5_ASAP7_75t_L g1891 ( 
.A1(n_1890),
.A2(n_1884),
.B1(n_1889),
.B2(n_1888),
.C(n_1724),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1891),
.B(n_1888),
.Y(n_1892)
);

AOI21xp5_ASAP7_75t_L g1893 ( 
.A1(n_1891),
.A2(n_1724),
.B(n_1738),
.Y(n_1893)
);

AOI22xp5_ASAP7_75t_L g1894 ( 
.A1(n_1892),
.A2(n_1893),
.B1(n_1737),
.B2(n_1726),
.Y(n_1894)
);

AOI21xp33_ASAP7_75t_L g1895 ( 
.A1(n_1892),
.A2(n_1711),
.B(n_1698),
.Y(n_1895)
);

AOI21x1_ASAP7_75t_L g1896 ( 
.A1(n_1894),
.A2(n_1747),
.B(n_1746),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1895),
.A2(n_1740),
.B(n_1737),
.Y(n_1897)
);

AOI21xp5_ASAP7_75t_L g1898 ( 
.A1(n_1897),
.A2(n_1740),
.B(n_1644),
.Y(n_1898)
);

AOI322xp5_ASAP7_75t_L g1899 ( 
.A1(n_1898),
.A2(n_1896),
.A3(n_1642),
.B1(n_1652),
.B2(n_1649),
.C1(n_1698),
.C2(n_1711),
.Y(n_1899)
);

AOI221xp5_ASAP7_75t_L g1900 ( 
.A1(n_1899),
.A2(n_1649),
.B1(n_1652),
.B2(n_1661),
.C(n_1701),
.Y(n_1900)
);

AOI211xp5_ASAP7_75t_L g1901 ( 
.A1(n_1900),
.A2(n_1665),
.B(n_1705),
.C(n_1645),
.Y(n_1901)
);


endmodule