module real_jpeg_2222_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_384;
wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_366;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_353;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_348;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_393;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_378;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_387;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_372;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_383;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_402;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_386;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_395;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_357;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_380;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_397;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_391;
wire n_401;
wire n_148;
wire n_373;
wire n_396;
wire n_392;
wire n_196;
wire n_375;
wire n_330;
wire n_298;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_385;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_343;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_400;
wire n_174;
wire n_388;
wire n_255;
wire n_243;
wire n_299;
wire n_352;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_379;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_351;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_51;
wire n_205;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_389;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;
wire n_364;

INVx2_ASAP7_75t_L g110 ( 
.A(n_0),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_1),
.B(n_24),
.Y(n_55)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_1),
.B(n_36),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_1),
.B(n_29),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_1),
.B(n_46),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_1),
.B(n_108),
.Y(n_169)
);

INVx1_ASAP7_75t_L g176 ( 
.A(n_1),
.Y(n_176)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_2),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g181 ( 
.A(n_2),
.B(n_58),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_2),
.B(n_108),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_2),
.B(n_77),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_2),
.B(n_132),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g345 ( 
.A(n_2),
.B(n_24),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_3),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_4),
.B(n_29),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g180 ( 
.A(n_4),
.B(n_46),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_4),
.B(n_58),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_4),
.B(n_36),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_4),
.B(n_77),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_4),
.B(n_108),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_4),
.B(n_132),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_4),
.B(n_24),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_5),
.B(n_36),
.Y(n_149)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_5),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_5),
.B(n_29),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_5),
.B(n_46),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_5),
.B(n_58),
.Y(n_261)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

BUFx10_ASAP7_75t_L g77 ( 
.A(n_8),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_9),
.B(n_24),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_29),
.Y(n_67)
);

AND2x2_ASAP7_75t_L g71 ( 
.A(n_9),
.B(n_46),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_9),
.B(n_58),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g119 ( 
.A(n_9),
.B(n_77),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_9),
.B(n_108),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_9),
.B(n_132),
.Y(n_219)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_11),
.B(n_24),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_11),
.B(n_36),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_11),
.B(n_29),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_11),
.B(n_46),
.Y(n_102)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_11),
.B(n_58),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_11),
.B(n_132),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_11),
.B(n_108),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_11),
.B(n_77),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_12),
.B(n_29),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_12),
.B(n_36),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_12),
.B(n_46),
.Y(n_190)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_12),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_12),
.B(n_58),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_12),
.B(n_77),
.Y(n_262)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_14),
.B(n_29),
.Y(n_28)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_14),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_14),
.B(n_46),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_14),
.B(n_58),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_14),
.B(n_77),
.Y(n_76)
);

AND2x2_ASAP7_75t_SL g107 ( 
.A(n_14),
.B(n_108),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_14),
.B(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_14),
.B(n_24),
.Y(n_133)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_15),
.Y(n_59)
);

XOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_86),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_85),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_60),
.Y(n_18)
);

OR2x2_ASAP7_75t_L g85 ( 
.A(n_19),
.B(n_60),
.Y(n_85)
);

XOR2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_47),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_SL g20 ( 
.A1(n_21),
.A2(n_22),
.B1(n_39),
.B2(n_40),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_L g22 ( 
.A1(n_23),
.A2(n_26),
.B1(n_27),
.B2(n_38),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_23),
.Y(n_38)
);

MAJIxp5_ASAP7_75t_L g70 ( 
.A(n_23),
.B(n_71),
.C(n_72),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_23),
.A2(n_38),
.B1(n_125),
.B2(n_127),
.Y(n_124)
);

INVx4_ASAP7_75t_L g157 ( 
.A(n_24),
.Y(n_157)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

BUFx24_ASAP7_75t_SL g406 ( 
.A(n_27),
.Y(n_406)
);

HAxp5_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_32),
.CON(n_27),
.SN(n_27)
);

MAJIxp5_ASAP7_75t_L g40 ( 
.A(n_28),
.B(n_41),
.C(n_44),
.Y(n_40)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_28),
.A2(n_44),
.B1(n_45),
.B2(n_51),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_28),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_28),
.A2(n_51),
.B1(n_328),
.B2(n_329),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g341 ( 
.A(n_28),
.B(n_329),
.C(n_330),
.Y(n_341)
);

INVx4_ASAP7_75t_L g202 ( 
.A(n_29),
.Y(n_202)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_32),
.A2(n_33),
.B1(n_352),
.B2(n_353),
.Y(n_351)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_33),
.B(n_107),
.C(n_131),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_34),
.B(n_35),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_35),
.B(n_43),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_35),
.B(n_165),
.Y(n_313)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_36),
.Y(n_35)
);

BUFx12f_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

OAI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_41),
.A2(n_42),
.B1(n_49),
.B2(n_50),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_41),
.A2(n_42),
.B1(n_122),
.B2(n_123),
.Y(n_121)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_42),
.B(n_99),
.C(n_101),
.Y(n_98)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_44),
.A2(n_45),
.B1(n_56),
.B2(n_57),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g208 ( 
.A1(n_44),
.A2(n_45),
.B1(n_209),
.B2(n_210),
.Y(n_208)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g53 ( 
.A(n_45),
.B(n_54),
.C(n_56),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_45),
.B(n_100),
.C(n_209),
.Y(n_314)
);

INVx3_ASAP7_75t_SL g164 ( 
.A(n_46),
.Y(n_164)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_48),
.B(n_52),
.C(n_53),
.Y(n_47)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_48),
.B(n_84),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_52),
.B(n_53),
.Y(n_84)
);

OAI22xp5_ASAP7_75t_SL g79 ( 
.A1(n_54),
.A2(n_55),
.B1(n_80),
.B2(n_81),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_55),
.Y(n_54)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_56),
.A2(n_57),
.B1(n_75),
.B2(n_76),
.Y(n_97)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_56),
.A2(n_57),
.B1(n_119),
.B2(n_159),
.Y(n_158)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

MAJIxp5_ASAP7_75t_L g74 ( 
.A(n_57),
.B(n_75),
.C(n_78),
.Y(n_74)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_57),
.B(n_119),
.C(n_155),
.Y(n_199)
);

INVx4_ASAP7_75t_L g310 ( 
.A(n_58),
.Y(n_310)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_82),
.C(n_83),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_61),
.A2(n_62),
.B1(n_135),
.B2(n_136),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g61 ( 
.A(n_62),
.Y(n_61)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_63),
.B(n_74),
.C(n_79),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_63),
.A2(n_64),
.B1(n_92),
.B2(n_93),
.Y(n_91)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_64),
.Y(n_63)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_65),
.B(n_70),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_66),
.A2(n_67),
.B1(n_68),
.B2(n_69),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_66),
.B(n_69),
.C(n_70),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g344 ( 
.A1(n_66),
.A2(n_67),
.B1(n_345),
.B2(n_346),
.Y(n_344)
);

OAI22xp5_ASAP7_75t_SL g370 ( 
.A1(n_66),
.A2(n_67),
.B1(n_133),
.B2(n_371),
.Y(n_370)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g128 ( 
.A(n_67),
.B(n_129),
.C(n_133),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_67),
.B(n_343),
.C(n_346),
.Y(n_367)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_69),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_71),
.A2(n_72),
.B1(n_73),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_71),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g311 ( 
.A1(n_71),
.A2(n_126),
.B1(n_312),
.B2(n_313),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g343 ( 
.A(n_71),
.B(n_309),
.C(n_313),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_73),
.Y(n_72)
);

XNOR2xp5_ASAP7_75t_SL g92 ( 
.A(n_74),
.B(n_79),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g103 ( 
.A(n_75),
.B(n_104),
.C(n_106),
.Y(n_103)
);

OAI22xp5_ASAP7_75t_L g116 ( 
.A1(n_75),
.A2(n_76),
.B1(n_106),
.B2(n_107),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_75),
.A2(n_76),
.B1(n_180),
.B2(n_186),
.Y(n_185)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

MAJIxp5_ASAP7_75t_L g179 ( 
.A(n_76),
.B(n_180),
.C(n_181),
.Y(n_179)
);

INVx13_ASAP7_75t_L g204 ( 
.A(n_77),
.Y(n_204)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_78),
.B(n_97),
.Y(n_96)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_81),
.Y(n_80)
);

XNOR2xp5_ASAP7_75t_SL g135 ( 
.A(n_82),
.B(n_83),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_137),
.B(n_401),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_89),
.B(n_134),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g402 ( 
.A(n_89),
.B(n_134),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_94),
.C(n_111),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g386 ( 
.A1(n_90),
.A2(n_91),
.B1(n_94),
.B2(n_387),
.Y(n_386)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_92),
.Y(n_93)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_94),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_95),
.B(n_98),
.C(n_103),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g391 ( 
.A1(n_95),
.A2(n_96),
.B1(n_392),
.B2(n_393),
.Y(n_391)
);

CKINVDCx16_ASAP7_75t_R g95 ( 
.A(n_96),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_SL g392 ( 
.A(n_98),
.B(n_103),
.Y(n_392)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_99),
.A2(n_100),
.B1(n_101),
.B2(n_102),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_99),
.A2(n_100),
.B1(n_207),
.B2(n_208),
.Y(n_206)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_104),
.A2(n_105),
.B1(n_115),
.B2(n_116),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_105),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_106),
.A2(n_107),
.B1(n_219),
.B2(n_222),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_106),
.A2(n_107),
.B1(n_131),
.B2(n_243),
.Y(n_352)
);

CKINVDCx20_ASAP7_75t_R g106 ( 
.A(n_107),
.Y(n_106)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_109),
.B(n_224),
.Y(n_265)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g385 ( 
.A(n_111),
.B(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_124),
.C(n_128),
.Y(n_111)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_112),
.B(n_390),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g112 ( 
.A(n_113),
.B(n_117),
.C(n_121),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g362 ( 
.A1(n_113),
.A2(n_114),
.B1(n_363),
.B2(n_364),
.Y(n_362)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_SL g363 ( 
.A(n_117),
.B(n_121),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_119),
.C(n_120),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g357 ( 
.A(n_118),
.B(n_120),
.Y(n_357)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_119),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_119),
.A2(n_159),
.B1(n_357),
.B2(n_358),
.Y(n_356)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_123),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g390 ( 
.A(n_124),
.B(n_128),
.Y(n_390)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_125),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g368 ( 
.A1(n_129),
.A2(n_130),
.B1(n_369),
.B2(n_370),
.Y(n_368)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_130),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_131),
.B(n_147),
.Y(n_146)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_131),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_131),
.A2(n_241),
.B1(n_242),
.B2(n_243),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g316 ( 
.A1(n_131),
.A2(n_147),
.B1(n_177),
.B2(n_243),
.Y(n_316)
);

INVx2_ASAP7_75t_L g175 ( 
.A(n_132),
.Y(n_175)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_133),
.Y(n_371)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_135),
.Y(n_136)
);

AOI21xp5_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_383),
.B(n_398),
.Y(n_137)
);

OAI31xp33_ASAP7_75t_L g138 ( 
.A1(n_139),
.A2(n_333),
.A3(n_372),
.B(n_377),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g139 ( 
.A(n_140),
.B(n_301),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_225),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_193),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g379 ( 
.A(n_142),
.B(n_193),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_160),
.C(n_183),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_143),
.B(n_298),
.Y(n_297)
);

BUFx24_ASAP7_75t_SL g403 ( 
.A(n_143),
.Y(n_403)
);

FAx1_ASAP7_75t_SL g143 ( 
.A(n_144),
.B(n_150),
.CI(n_154),
.CON(n_143),
.SN(n_143)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_144),
.B(n_150),
.C(n_154),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g144 ( 
.A(n_145),
.B(n_148),
.C(n_149),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_145),
.A2(n_146),
.B1(n_293),
.B2(n_294),
.Y(n_292)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

O2A1O1Ixp33_ASAP7_75t_L g355 ( 
.A1(n_146),
.A2(n_177),
.B(n_243),
.C(n_317),
.Y(n_355)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_147),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_L g191 ( 
.A1(n_147),
.A2(n_174),
.B1(n_177),
.B2(n_192),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_SL g294 ( 
.A(n_148),
.B(n_149),
.Y(n_294)
);

OAI21xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B(n_153),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_L g153 ( 
.A(n_151),
.B(n_152),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_153),
.A2(n_214),
.B1(n_215),
.B2(n_216),
.Y(n_213)
);

CKINVDCx20_ASAP7_75t_R g215 ( 
.A(n_153),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_155),
.B(n_158),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_157),
.Y(n_155)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_156),
.B(n_175),
.Y(n_270)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_156),
.B(n_204),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_157),
.B(n_224),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_160),
.B(n_183),
.Y(n_298)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_161),
.A2(n_162),
.B1(n_171),
.B2(n_182),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g195 ( 
.A(n_161),
.B(n_172),
.C(n_179),
.Y(n_195)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

XOR2xp5_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_166),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g214 ( 
.A(n_163),
.B(n_168),
.C(n_170),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_165),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_L g201 ( 
.A(n_165),
.B(n_202),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_167),
.A2(n_168),
.B1(n_169),
.B2(n_170),
.Y(n_166)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_167),
.Y(n_170)
);

CKINVDCx16_ASAP7_75t_R g168 ( 
.A(n_169),
.Y(n_168)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_171),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_173),
.B1(n_178),
.B2(n_179),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g173 ( 
.A(n_174),
.B(n_177),
.Y(n_173)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_174),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_176),
.B(n_204),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_176),
.B(n_310),
.Y(n_309)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_179),
.Y(n_178)
);

CKINVDCx14_ASAP7_75t_R g186 ( 
.A(n_180),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_181),
.B(n_185),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_184),
.B(n_187),
.C(n_191),
.Y(n_183)
);

FAx1_ASAP7_75t_SL g288 ( 
.A(n_184),
.B(n_187),
.CI(n_191),
.CON(n_288),
.SN(n_288)
);

MAJIxp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_189),
.C(n_190),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g236 ( 
.A(n_188),
.B(n_190),
.Y(n_236)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_189),
.B(n_236),
.Y(n_235)
);

BUFx24_ASAP7_75t_SL g405 ( 
.A(n_193),
.Y(n_405)
);

FAx1_ASAP7_75t_SL g193 ( 
.A(n_194),
.B(n_211),
.CI(n_212),
.CON(n_193),
.SN(n_193)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_194),
.B(n_211),
.C(n_212),
.Y(n_332)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_196),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_195),
.B(n_198),
.C(n_205),
.Y(n_304)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_197),
.A2(n_198),
.B1(n_205),
.B2(n_206),
.Y(n_196)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_199),
.B(n_200),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_199),
.B(n_201),
.C(n_203),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_203),
.Y(n_200)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_208),
.Y(n_207)
);

CKINVDCx16_ASAP7_75t_R g210 ( 
.A(n_209),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g212 ( 
.A(n_213),
.B(n_217),
.Y(n_212)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_214),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_214),
.B(n_215),
.C(n_217),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_219),
.A2(n_220),
.B1(n_221),
.B2(n_222),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g222 ( 
.A(n_219),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g331 ( 
.A(n_219),
.B(n_221),
.C(n_223),
.Y(n_331)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_221),
.Y(n_220)
);

AOI21xp5_ASAP7_75t_SL g225 ( 
.A1(n_226),
.A2(n_296),
.B(n_300),
.Y(n_225)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_227),
.A2(n_284),
.B(n_295),
.Y(n_226)
);

AOI21xp5_ASAP7_75t_L g227 ( 
.A1(n_228),
.A2(n_256),
.B(n_283),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_247),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_229),
.B(n_247),
.Y(n_283)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_230),
.B(n_239),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_235),
.B1(n_237),
.B2(n_238),
.Y(n_230)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_231),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_233),
.C(n_234),
.Y(n_231)
);

FAx1_ASAP7_75t_SL g248 ( 
.A(n_232),
.B(n_233),
.CI(n_234),
.CON(n_248),
.SN(n_248)
);

CKINVDCx16_ASAP7_75t_R g238 ( 
.A(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g285 ( 
.A(n_235),
.B(n_237),
.C(n_239),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_SL g239 ( 
.A(n_240),
.B(n_244),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_240),
.B(n_245),
.C(n_246),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g240 ( 
.A(n_241),
.B(n_243),
.Y(n_240)
);

CKINVDCx16_ASAP7_75t_R g241 ( 
.A(n_242),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_248),
.B(n_249),
.C(n_255),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g279 ( 
.A(n_248),
.B(n_280),
.Y(n_279)
);

BUFx24_ASAP7_75t_SL g410 ( 
.A(n_248),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_L g280 ( 
.A1(n_249),
.A2(n_250),
.B1(n_255),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_250),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g250 ( 
.A(n_251),
.B(n_253),
.Y(n_250)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_251),
.A2(n_252),
.B1(n_253),
.B2(n_254),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_252),
.Y(n_251)
);

CKINVDCx16_ASAP7_75t_R g253 ( 
.A(n_254),
.Y(n_253)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_255),
.Y(n_281)
);

OAI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_277),
.B(n_282),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_258),
.A2(n_268),
.B(n_276),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g258 ( 
.A(n_259),
.B(n_264),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_259),
.B(n_264),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_260),
.B(n_263),
.Y(n_259)
);

XNOR2xp5_ASAP7_75t_L g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_262),
.C(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_L g269 ( 
.A(n_265),
.B(n_270),
.Y(n_269)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_266),
.B1(n_267),
.B2(n_274),
.Y(n_273)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_265),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

OAI21xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_271),
.B(n_275),
.Y(n_268)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_273),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_272),
.B(n_273),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_278),
.B(n_279),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_278),
.B(n_279),
.Y(n_282)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_285),
.B(n_286),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_SL g295 ( 
.A(n_285),
.B(n_286),
.Y(n_295)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_287),
.A2(n_288),
.B1(n_289),
.B2(n_290),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_287),
.B(n_291),
.C(n_292),
.Y(n_299)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

BUFx24_ASAP7_75t_SL g411 ( 
.A(n_288),
.Y(n_411)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_290),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

CKINVDCx16_ASAP7_75t_R g293 ( 
.A(n_294),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_SL g296 ( 
.A(n_297),
.B(n_299),
.Y(n_296)
);

NOR2xp33_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_299),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_302),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g378 ( 
.A1(n_302),
.A2(n_379),
.B(n_380),
.Y(n_378)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_303),
.B(n_332),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_303),
.B(n_332),
.Y(n_380)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_304),
.B(n_305),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_304),
.B(n_306),
.C(n_319),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_318),
.B2(n_319),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_307),
.Y(n_306)
);

BUFx24_ASAP7_75t_SL g404 ( 
.A(n_307),
.Y(n_404)
);

FAx1_ASAP7_75t_SL g307 ( 
.A(n_308),
.B(n_314),
.CI(n_315),
.CON(n_307),
.SN(n_307)
);

MAJIxp5_ASAP7_75t_L g339 ( 
.A(n_308),
.B(n_314),
.C(n_315),
.Y(n_339)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_311),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

OAI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_320),
.B(n_324),
.C(n_325),
.Y(n_348)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

XNOR2xp5_ASAP7_75t_SL g323 ( 
.A(n_324),
.B(n_325),
.Y(n_323)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_326),
.A2(n_327),
.B1(n_330),
.B2(n_331),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_327),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_329),
.Y(n_328)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_331),
.Y(n_330)
);

INVxp33_ASAP7_75t_L g333 ( 
.A(n_334),
.Y(n_333)
);

A2O1A1O1Ixp25_ASAP7_75t_SL g377 ( 
.A1(n_334),
.A2(n_373),
.B(n_378),
.C(n_381),
.D(n_382),
.Y(n_377)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_335),
.B(n_359),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_335),
.B(n_359),
.Y(n_382)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_336),
.B(n_348),
.C(n_349),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g375 ( 
.A1(n_336),
.A2(n_337),
.B1(n_349),
.B2(n_350),
.Y(n_375)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_338),
.A2(n_339),
.B1(n_340),
.B2(n_347),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_338),
.B(n_341),
.C(n_342),
.Y(n_360)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_339),
.Y(n_338)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_340),
.Y(n_347)
);

XNOR2xp5_ASAP7_75t_SL g340 ( 
.A(n_341),
.B(n_342),
.Y(n_340)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_343),
.B(n_344),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g346 ( 
.A(n_345),
.Y(n_346)
);

XOR2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_375),
.Y(n_374)
);

CKINVDCx14_ASAP7_75t_R g349 ( 
.A(n_350),
.Y(n_349)
);

XNOR2xp5_ASAP7_75t_SL g350 ( 
.A(n_351),
.B(n_354),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g366 ( 
.A(n_351),
.B(n_355),
.C(n_356),
.Y(n_366)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_352),
.Y(n_353)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_355),
.B(n_356),
.Y(n_354)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_357),
.Y(n_358)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_360),
.B(n_361),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_360),
.B(n_362),
.C(n_365),
.Y(n_397)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_362),
.B(n_365),
.Y(n_361)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_363),
.Y(n_364)
);

BUFx24_ASAP7_75t_SL g408 ( 
.A(n_365),
.Y(n_408)
);

FAx1_ASAP7_75t_SL g365 ( 
.A(n_366),
.B(n_367),
.CI(n_368),
.CON(n_365),
.SN(n_365)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_366),
.B(n_367),
.C(n_368),
.Y(n_394)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_370),
.Y(n_369)
);

INVx1_ASAP7_75t_L g372 ( 
.A(n_373),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_SL g373 ( 
.A(n_374),
.B(n_376),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_374),
.B(n_376),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_L g383 ( 
.A(n_384),
.B(n_395),
.Y(n_383)
);

OAI21xp5_ASAP7_75t_L g398 ( 
.A1(n_384),
.A2(n_399),
.B(n_400),
.Y(n_398)
);

NOR2xp33_ASAP7_75t_SL g384 ( 
.A(n_385),
.B(n_388),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_385),
.B(n_388),
.Y(n_400)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_389),
.B(n_391),
.C(n_394),
.Y(n_388)
);

FAx1_ASAP7_75t_SL g396 ( 
.A(n_389),
.B(n_391),
.CI(n_394),
.CON(n_396),
.SN(n_396)
);

INVx1_ASAP7_75t_L g393 ( 
.A(n_392),
.Y(n_393)
);

NOR2xp33_ASAP7_75t_SL g395 ( 
.A(n_396),
.B(n_397),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_396),
.B(n_397),
.Y(n_399)
);

BUFx24_ASAP7_75t_SL g409 ( 
.A(n_396),
.Y(n_409)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);


endmodule