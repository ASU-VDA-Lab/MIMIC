module fake_jpeg_953_n_583 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_583);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_583;

wire n_529;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_547;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_570;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_384;
wire n_296;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_358;
wire n_312;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_568;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_17),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_7),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_17),
.Y(n_21)
);

CKINVDCx16_ASAP7_75t_R g22 ( 
.A(n_16),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_16),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_9),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_2),
.Y(n_28)
);

CKINVDCx14_ASAP7_75t_R g29 ( 
.A(n_11),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_14),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_11),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

INVx4_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_5),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_2),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_0),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_4),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx8_ASAP7_75t_L g45 ( 
.A(n_0),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_10),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g47 ( 
.A(n_7),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_4),
.B(n_3),
.Y(n_48)
);

INVx11_ASAP7_75t_SL g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_14),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_8),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_17),
.Y(n_52)
);

INVx8_ASAP7_75t_L g53 ( 
.A(n_8),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_12),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_0),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_3),
.Y(n_56)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_57),
.Y(n_129)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_26),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_58),
.Y(n_136)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_49),
.Y(n_59)
);

BUFx10_ASAP7_75t_L g176 ( 
.A(n_59),
.Y(n_176)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx4_ASAP7_75t_SL g174 ( 
.A(n_60),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_18),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_61),
.B(n_80),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_9),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_62),
.B(n_65),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g141 ( 
.A(n_63),
.Y(n_141)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_37),
.Y(n_64)
);

INVx3_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_23),
.B(n_9),
.Y(n_65)
);

INVx3_ASAP7_75t_L g66 ( 
.A(n_33),
.Y(n_66)
);

INVx3_ASAP7_75t_L g165 ( 
.A(n_66),
.Y(n_165)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_26),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g150 ( 
.A(n_67),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_23),
.B(n_9),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_68),
.B(n_71),
.Y(n_149)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_33),
.Y(n_69)
);

INVx5_ASAP7_75t_L g171 ( 
.A(n_69),
.Y(n_171)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_33),
.Y(n_70)
);

INVx6_ASAP7_75t_L g175 ( 
.A(n_70),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_19),
.B(n_10),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_38),
.Y(n_72)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_72),
.Y(n_128)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_38),
.Y(n_73)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_73),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_19),
.B(n_10),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_75),
.B(n_84),
.Y(n_189)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_33),
.Y(n_76)
);

INVx3_ASAP7_75t_L g168 ( 
.A(n_76),
.Y(n_168)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_30),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_77),
.Y(n_173)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_53),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g167 ( 
.A(n_78),
.Y(n_167)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_35),
.Y(n_79)
);

INVx3_ASAP7_75t_L g210 ( 
.A(n_79),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_38),
.B(n_10),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_30),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g185 ( 
.A(n_81),
.Y(n_185)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_35),
.Y(n_82)
);

INVx3_ASAP7_75t_L g216 ( 
.A(n_82),
.Y(n_216)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_49),
.Y(n_83)
);

INVx4_ASAP7_75t_L g151 ( 
.A(n_83),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_20),
.B(n_7),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_33),
.Y(n_85)
);

INVx2_ASAP7_75t_L g131 ( 
.A(n_85),
.Y(n_131)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_33),
.Y(n_86)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_86),
.Y(n_155)
);

INVx11_ASAP7_75t_L g87 ( 
.A(n_35),
.Y(n_87)
);

INVx11_ASAP7_75t_L g162 ( 
.A(n_87),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_20),
.B(n_7),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_SL g193 ( 
.A(n_88),
.B(n_98),
.Y(n_193)
);

INVx8_ASAP7_75t_L g89 ( 
.A(n_41),
.Y(n_89)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_89),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_30),
.Y(n_90)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_90),
.Y(n_187)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_30),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g201 ( 
.A(n_91),
.Y(n_201)
);

INVx2_ASAP7_75t_SL g92 ( 
.A(n_21),
.Y(n_92)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_92),
.Y(n_161)
);

INVx8_ASAP7_75t_L g93 ( 
.A(n_41),
.Y(n_93)
);

INVx6_ASAP7_75t_L g200 ( 
.A(n_93),
.Y(n_200)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_41),
.Y(n_94)
);

INVx2_ASAP7_75t_L g132 ( 
.A(n_94),
.Y(n_132)
);

INVx6_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g209 ( 
.A(n_95),
.Y(n_209)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_53),
.Y(n_96)
);

BUFx3_ASAP7_75t_L g181 ( 
.A(n_96),
.Y(n_181)
);

BUFx3_ASAP7_75t_L g97 ( 
.A(n_53),
.Y(n_97)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_97),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_25),
.B(n_12),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_22),
.Y(n_99)
);

INVxp67_ASAP7_75t_L g134 ( 
.A(n_99),
.Y(n_134)
);

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_45),
.Y(n_100)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_100),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_40),
.Y(n_101)
);

INVx6_ASAP7_75t_L g203 ( 
.A(n_101),
.Y(n_203)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_41),
.Y(n_102)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_102),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_40),
.Y(n_103)
);

INVx6_ASAP7_75t_L g207 ( 
.A(n_103),
.Y(n_207)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_104),
.Y(n_139)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_45),
.Y(n_105)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_105),
.Y(n_140)
);

BUFx6f_ASAP7_75t_L g106 ( 
.A(n_40),
.Y(n_106)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_106),
.Y(n_170)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_47),
.Y(n_107)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g108 ( 
.A(n_47),
.Y(n_108)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_108),
.Y(n_145)
);

INVx11_ASAP7_75t_L g109 ( 
.A(n_22),
.Y(n_109)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_109),
.Y(n_156)
);

BUFx12f_ASAP7_75t_L g110 ( 
.A(n_45),
.Y(n_110)
);

BUFx12_ASAP7_75t_L g183 ( 
.A(n_110),
.Y(n_183)
);

INVx8_ASAP7_75t_L g111 ( 
.A(n_42),
.Y(n_111)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_111),
.Y(n_157)
);

INVx4_ASAP7_75t_L g112 ( 
.A(n_42),
.Y(n_112)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_112),
.Y(n_160)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_47),
.Y(n_113)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_113),
.Y(n_163)
);

INVx11_ASAP7_75t_L g114 ( 
.A(n_29),
.Y(n_114)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_114),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx2_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_47),
.Y(n_116)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_116),
.Y(n_166)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_54),
.Y(n_117)
);

INVx2_ASAP7_75t_L g169 ( 
.A(n_117),
.Y(n_169)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_42),
.Y(n_118)
);

INVx2_ASAP7_75t_L g179 ( 
.A(n_118),
.Y(n_179)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_54),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

BUFx4f_ASAP7_75t_SL g120 ( 
.A(n_54),
.Y(n_120)
);

INVx6_ASAP7_75t_SL g184 ( 
.A(n_120),
.Y(n_184)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_54),
.Y(n_121)
);

INVx2_ASAP7_75t_L g188 ( 
.A(n_121),
.Y(n_188)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_21),
.Y(n_122)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_122),
.Y(n_192)
);

INVx8_ASAP7_75t_L g123 ( 
.A(n_55),
.Y(n_123)
);

INVx2_ASAP7_75t_L g195 ( 
.A(n_123),
.Y(n_195)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_21),
.Y(n_124)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_124),
.Y(n_202)
);

INVx3_ASAP7_75t_L g125 ( 
.A(n_24),
.Y(n_125)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_125),
.Y(n_206)
);

BUFx6f_ASAP7_75t_L g126 ( 
.A(n_24),
.Y(n_126)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_126),
.Y(n_212)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_63),
.A2(n_55),
.B1(n_56),
.B2(n_28),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_127),
.A2(n_133),
.B1(n_135),
.B2(n_146),
.Y(n_226)
);

AOI22xp33_ASAP7_75t_SL g133 ( 
.A1(n_59),
.A2(n_56),
.B1(n_51),
.B2(n_44),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_67),
.A2(n_25),
.B1(n_52),
.B2(n_50),
.Y(n_135)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_59),
.A2(n_27),
.B1(n_51),
.B2(n_44),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g147 ( 
.A1(n_58),
.A2(n_52),
.B1(n_50),
.B2(n_46),
.Y(n_147)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_147),
.A2(n_172),
.B1(n_182),
.B2(n_194),
.Y(n_242)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_92),
.Y(n_153)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_153),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_57),
.B(n_46),
.C(n_43),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_158),
.B(n_148),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_95),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_159),
.A2(n_177),
.B1(n_208),
.B2(n_116),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g172 ( 
.A1(n_117),
.A2(n_34),
.B1(n_31),
.B2(n_32),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_74),
.A2(n_39),
.B1(n_36),
.B2(n_43),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_78),
.A2(n_36),
.B1(n_39),
.B2(n_44),
.Y(n_178)
);

OR2x2_ASAP7_75t_L g269 ( 
.A(n_178),
.B(n_191),
.Y(n_269)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_124),
.Y(n_180)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_180),
.Y(n_268)
);

AOI22xp33_ASAP7_75t_SL g182 ( 
.A1(n_87),
.A2(n_56),
.B1(n_51),
.B2(n_28),
.Y(n_182)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_126),
.Y(n_190)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_190),
.Y(n_274)
);

AOI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_97),
.A2(n_28),
.B1(n_27),
.B2(n_24),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_SL g194 ( 
.A1(n_99),
.A2(n_109),
.B1(n_83),
.B2(n_110),
.Y(n_194)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_123),
.Y(n_196)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_196),
.Y(n_276)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_112),
.Y(n_198)
);

INVx1_ASAP7_75t_SL g250 ( 
.A(n_198),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_100),
.B(n_27),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_199),
.B(n_205),
.Y(n_218)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_89),
.Y(n_204)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_204),
.B(n_214),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_100),
.B(n_6),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_77),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_208)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_110),
.A2(n_6),
.B1(n_1),
.B2(n_2),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_211),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_245)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_93),
.Y(n_214)
);

INVx2_ASAP7_75t_L g215 ( 
.A(n_81),
.Y(n_215)
);

INVx2_ASAP7_75t_L g238 ( 
.A(n_215),
.Y(n_238)
);

AND2x2_ASAP7_75t_L g217 ( 
.A(n_69),
.B(n_13),
.Y(n_217)
);

NOR2xp33_ASAP7_75t_SL g227 ( 
.A(n_217),
.B(n_0),
.Y(n_227)
);

INVx4_ASAP7_75t_L g219 ( 
.A(n_175),
.Y(n_219)
);

INVx4_ASAP7_75t_L g302 ( 
.A(n_219),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_120),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_220),
.B(n_227),
.Y(n_333)
);

AND2x2_ASAP7_75t_L g300 ( 
.A(n_221),
.B(n_270),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_202),
.A2(n_103),
.B1(n_108),
.B2(n_107),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_222),
.A2(n_225),
.B1(n_236),
.B2(n_272),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_164),
.Y(n_224)
);

BUFx3_ASAP7_75t_L g306 ( 
.A(n_224),
.Y(n_306)
);

AOI22xp33_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_106),
.B1(n_101),
.B2(n_91),
.Y(n_225)
);

CKINVDCx16_ASAP7_75t_R g228 ( 
.A(n_184),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g307 ( 
.A(n_228),
.B(n_232),
.Y(n_307)
);

INVx5_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

INVx4_ASAP7_75t_L g323 ( 
.A(n_229),
.Y(n_323)
);

BUFx2_ASAP7_75t_L g230 ( 
.A(n_152),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g296 ( 
.A(n_230),
.Y(n_296)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_199),
.A2(n_111),
.B1(n_70),
.B2(n_90),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g310 ( 
.A(n_231),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_197),
.Y(n_232)
);

INVx3_ASAP7_75t_L g233 ( 
.A(n_151),
.Y(n_233)
);

INVx4_ASAP7_75t_L g340 ( 
.A(n_233),
.Y(n_340)
);

AOI22xp33_ASAP7_75t_SL g234 ( 
.A1(n_161),
.A2(n_1),
.B1(n_3),
.B2(n_4),
.Y(n_234)
);

INVxp67_ASAP7_75t_L g321 ( 
.A(n_234),
.Y(n_321)
);

AOI22xp33_ASAP7_75t_SL g235 ( 
.A1(n_149),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g330 ( 
.A(n_235),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_142),
.A2(n_5),
.B1(n_13),
.B2(n_14),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_143),
.B(n_5),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_237),
.B(n_278),
.Y(n_295)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_141),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g312 ( 
.A(n_239),
.Y(n_312)
);

BUFx2_ASAP7_75t_L g240 ( 
.A(n_167),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_240),
.Y(n_341)
);

INVx4_ASAP7_75t_L g241 ( 
.A(n_175),
.Y(n_241)
);

INVx3_ASAP7_75t_L g299 ( 
.A(n_241),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_140),
.Y(n_243)
);

INVxp67_ASAP7_75t_L g336 ( 
.A(n_243),
.Y(n_336)
);

INVx3_ASAP7_75t_L g244 ( 
.A(n_171),
.Y(n_244)
);

INVx3_ASAP7_75t_L g329 ( 
.A(n_244),
.Y(n_329)
);

AOI22xp33_ASAP7_75t_SL g331 ( 
.A1(n_245),
.A2(n_247),
.B1(n_279),
.B2(n_284),
.Y(n_331)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_169),
.Y(n_246)
);

INVx2_ASAP7_75t_L g316 ( 
.A(n_246),
.Y(n_316)
);

INVx11_ASAP7_75t_L g247 ( 
.A(n_162),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_L g248 ( 
.A1(n_142),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g328 ( 
.A1(n_248),
.A2(n_259),
.B1(n_263),
.B2(n_264),
.Y(n_328)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_213),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g322 ( 
.A(n_249),
.Y(n_322)
);

INVx6_ASAP7_75t_L g251 ( 
.A(n_141),
.Y(n_251)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_251),
.Y(n_325)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_197),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_252),
.B(n_261),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g253 ( 
.A(n_205),
.B(n_15),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g315 ( 
.A(n_253),
.B(n_236),
.C(n_270),
.Y(n_315)
);

INVx4_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx2_ASAP7_75t_L g326 ( 
.A(n_254),
.Y(n_326)
);

A2O1A1Ixp33_ASAP7_75t_L g255 ( 
.A1(n_189),
.A2(n_18),
.B(n_149),
.C(n_193),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_255),
.B(n_218),
.Y(n_345)
);

INVx5_ASAP7_75t_L g256 ( 
.A(n_170),
.Y(n_256)
);

INVx2_ASAP7_75t_L g346 ( 
.A(n_256),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g257 ( 
.A(n_137),
.Y(n_257)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_257),
.Y(n_337)
);

INVx2_ASAP7_75t_L g258 ( 
.A(n_132),
.Y(n_258)
);

INVx1_ASAP7_75t_L g344 ( 
.A(n_258),
.Y(n_344)
);

OAI22xp33_ASAP7_75t_L g259 ( 
.A1(n_182),
.A2(n_18),
.B1(n_146),
.B2(n_133),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g260 ( 
.A(n_181),
.Y(n_260)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_260),
.Y(n_298)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_200),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g263 ( 
.A1(n_127),
.A2(n_211),
.B1(n_128),
.B2(n_166),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_195),
.A2(n_217),
.B1(n_194),
.B2(n_207),
.Y(n_264)
);

INVx2_ASAP7_75t_L g265 ( 
.A(n_138),
.Y(n_265)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_265),
.Y(n_309)
);

INVx2_ASAP7_75t_L g266 ( 
.A(n_139),
.Y(n_266)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_266),
.Y(n_311)
);

INVx3_ASAP7_75t_L g267 ( 
.A(n_157),
.Y(n_267)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_267),
.Y(n_339)
);

CKINVDCx20_ASAP7_75t_R g271 ( 
.A(n_136),
.Y(n_271)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_271),
.B(n_280),
.Y(n_317)
);

AOI22xp33_ASAP7_75t_L g272 ( 
.A1(n_130),
.A2(n_192),
.B1(n_206),
.B2(n_163),
.Y(n_272)
);

OAI22xp5_ASAP7_75t_L g273 ( 
.A1(n_203),
.A2(n_207),
.B1(n_145),
.B2(n_144),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_273),
.A2(n_294),
.B1(n_287),
.B2(n_293),
.Y(n_350)
);

INVx2_ASAP7_75t_L g275 ( 
.A(n_179),
.Y(n_275)
);

INVx1_ASAP7_75t_L g347 ( 
.A(n_275),
.Y(n_347)
);

INVx2_ASAP7_75t_L g277 ( 
.A(n_188),
.Y(n_277)
);

INVx1_ASAP7_75t_L g349 ( 
.A(n_277),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_131),
.B(n_156),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_SL g279 ( 
.A1(n_174),
.A2(n_216),
.B1(n_210),
.B2(n_129),
.Y(n_279)
);

CKINVDCx20_ASAP7_75t_R g280 ( 
.A(n_136),
.Y(n_280)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_155),
.Y(n_281)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_281),
.B(n_282),
.Y(n_304)
);

INVx2_ASAP7_75t_L g282 ( 
.A(n_160),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_134),
.B(n_174),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_283),
.B(n_285),
.Y(n_319)
);

INVx8_ASAP7_75t_L g284 ( 
.A(n_150),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_186),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g286 ( 
.A1(n_209),
.A2(n_173),
.B1(n_150),
.B2(n_154),
.Y(n_286)
);

OAI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_286),
.A2(n_222),
.B1(n_289),
.B2(n_221),
.Y(n_318)
);

BUFx2_ASAP7_75t_L g287 ( 
.A(n_170),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g314 ( 
.A(n_287),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_165),
.B(n_168),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_288),
.B(n_253),
.Y(n_305)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_134),
.A2(n_209),
.B1(n_173),
.B2(n_154),
.Y(n_289)
);

MAJx2_ASAP7_75t_L g303 ( 
.A(n_289),
.B(n_263),
.C(n_286),
.Y(n_303)
);

INVx4_ASAP7_75t_L g290 ( 
.A(n_203),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g324 ( 
.A(n_290),
.B(n_291),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g291 ( 
.A(n_185),
.B(n_187),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g292 ( 
.A(n_176),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_292),
.B(n_293),
.Y(n_332)
);

INVx2_ASAP7_75t_L g293 ( 
.A(n_185),
.Y(n_293)
);

OAI22xp5_ASAP7_75t_L g294 ( 
.A1(n_187),
.A2(n_201),
.B1(n_183),
.B2(n_176),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_226),
.A2(n_201),
.B1(n_183),
.B2(n_176),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g392 ( 
.A(n_301),
.Y(n_392)
);

CKINVDCx14_ASAP7_75t_R g359 ( 
.A(n_303),
.Y(n_359)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_305),
.B(n_315),
.Y(n_385)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_237),
.B(n_253),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g352 ( 
.A(n_313),
.B(n_320),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_297),
.B1(n_328),
.B2(n_300),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_270),
.B(n_278),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_288),
.B(n_255),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g365 ( 
.A(n_327),
.B(n_348),
.Y(n_365)
);

AOI22xp33_ASAP7_75t_L g334 ( 
.A1(n_242),
.A2(n_269),
.B1(n_268),
.B2(n_274),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g384 ( 
.A1(n_334),
.A2(n_339),
.B1(n_304),
.B2(n_347),
.Y(n_384)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_276),
.B(n_262),
.Y(n_335)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_335),
.B(n_343),
.Y(n_354)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_259),
.A2(n_269),
.B(n_224),
.Y(n_338)
);

AOI22xp33_ASAP7_75t_SL g382 ( 
.A1(n_338),
.A2(n_342),
.B1(n_298),
.B2(n_341),
.Y(n_382)
);

AOI22xp33_ASAP7_75t_SL g342 ( 
.A1(n_254),
.A2(n_260),
.B1(n_244),
.B2(n_241),
.Y(n_342)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_223),
.Y(n_343)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_345),
.B(n_313),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g348 ( 
.A(n_258),
.B(n_275),
.Y(n_348)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_350),
.Y(n_355)
);

OAI22xp5_ASAP7_75t_SL g351 ( 
.A1(n_300),
.A2(n_328),
.B1(n_338),
.B2(n_327),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_351),
.A2(n_363),
.B1(n_366),
.B2(n_373),
.Y(n_402)
);

OAI22xp5_ASAP7_75t_L g412 ( 
.A1(n_353),
.A2(n_368),
.B1(n_374),
.B2(n_377),
.Y(n_412)
);

AOI22xp5_ASAP7_75t_SL g356 ( 
.A1(n_330),
.A2(n_240),
.B1(n_256),
.B2(n_219),
.Y(n_356)
);

OAI21xp5_ASAP7_75t_L g397 ( 
.A1(n_356),
.A2(n_362),
.B(n_364),
.Y(n_397)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_348),
.Y(n_357)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_357),
.Y(n_394)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_324),
.Y(n_358)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_358),
.Y(n_395)
);

CKINVDCx20_ASAP7_75t_R g360 ( 
.A(n_308),
.Y(n_360)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_360),
.B(n_367),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_SL g410 ( 
.A(n_361),
.B(n_371),
.Y(n_410)
);

AOI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_330),
.A2(n_229),
.B1(n_230),
.B2(n_267),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_300),
.A2(n_290),
.B1(n_251),
.B2(n_246),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_SL g364 ( 
.A1(n_310),
.A2(n_249),
.B1(n_281),
.B2(n_250),
.Y(n_364)
);

OAI22xp5_ASAP7_75t_SL g366 ( 
.A1(n_320),
.A2(n_238),
.B1(n_239),
.B2(n_265),
.Y(n_366)
);

CKINVDCx20_ASAP7_75t_R g367 ( 
.A(n_317),
.Y(n_367)
);

AOI22xp5_ASAP7_75t_L g368 ( 
.A1(n_318),
.A2(n_238),
.B1(n_266),
.B2(n_277),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_SL g369 ( 
.A1(n_310),
.A2(n_321),
.B1(n_319),
.B2(n_297),
.Y(n_369)
);

OR2x2_ASAP7_75t_L g424 ( 
.A(n_369),
.B(n_384),
.Y(n_424)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_309),
.Y(n_370)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_370),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_307),
.B(n_250),
.Y(n_371)
);

NAND2xp5_ASAP7_75t_L g372 ( 
.A(n_295),
.B(n_285),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_372),
.B(n_376),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_301),
.A2(n_284),
.B1(n_282),
.B2(n_233),
.Y(n_373)
);

AOI22xp5_ASAP7_75t_L g374 ( 
.A1(n_295),
.A2(n_247),
.B1(n_315),
.B2(n_305),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_309),
.Y(n_375)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_375),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g376 ( 
.A(n_304),
.Y(n_376)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_303),
.A2(n_350),
.B1(n_345),
.B2(n_321),
.Y(n_377)
);

BUFx2_ASAP7_75t_SL g378 ( 
.A(n_298),
.Y(n_378)
);

AOI22xp33_ASAP7_75t_SL g406 ( 
.A1(n_378),
.A2(n_382),
.B1(n_340),
.B2(n_302),
.Y(n_406)
);

INVx2_ASAP7_75t_L g379 ( 
.A(n_325),
.Y(n_379)
);

INVx1_ASAP7_75t_L g401 ( 
.A(n_379),
.Y(n_401)
);

OAI22xp5_ASAP7_75t_SL g380 ( 
.A1(n_331),
.A2(n_333),
.B1(n_332),
.B2(n_314),
.Y(n_380)
);

AOI22xp5_ASAP7_75t_L g405 ( 
.A1(n_380),
.A2(n_388),
.B1(n_336),
.B2(n_299),
.Y(n_405)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_311),
.Y(n_381)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_381),
.Y(n_407)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_349),
.B(n_347),
.C(n_311),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g404 ( 
.A(n_383),
.B(n_336),
.C(n_326),
.Y(n_404)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_349),
.Y(n_386)
);

INVx1_ASAP7_75t_L g415 ( 
.A(n_386),
.Y(n_415)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_304),
.Y(n_387)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_387),
.Y(n_419)
);

OAI22xp5_ASAP7_75t_SL g388 ( 
.A1(n_325),
.A2(n_329),
.B1(n_344),
.B2(n_346),
.Y(n_388)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_316),
.Y(n_389)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_389),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g390 ( 
.A1(n_346),
.A2(n_339),
.B1(n_326),
.B2(n_299),
.Y(n_390)
);

OAI22xp5_ASAP7_75t_SL g411 ( 
.A1(n_390),
.A2(n_355),
.B1(n_368),
.B2(n_375),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_337),
.B(n_316),
.Y(n_391)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_391),
.B(n_393),
.Y(n_416)
);

CKINVDCx20_ASAP7_75t_R g393 ( 
.A(n_296),
.Y(n_393)
);

CKINVDCx20_ASAP7_75t_R g399 ( 
.A(n_391),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g441 ( 
.A(n_399),
.B(n_421),
.Y(n_441)
);

FAx1_ASAP7_75t_L g400 ( 
.A(n_359),
.B(n_329),
.CI(n_323),
.CON(n_400),
.SN(n_400)
);

OAI21xp5_ASAP7_75t_SL g432 ( 
.A1(n_400),
.A2(n_403),
.B(n_406),
.Y(n_432)
);

AOI21xp5_ASAP7_75t_L g403 ( 
.A1(n_382),
.A2(n_323),
.B(n_340),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g447 ( 
.A(n_404),
.B(n_389),
.C(n_379),
.Y(n_447)
);

AOI22xp5_ASAP7_75t_L g437 ( 
.A1(n_405),
.A2(n_418),
.B1(n_425),
.B2(n_366),
.Y(n_437)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_385),
.B(n_322),
.Y(n_408)
);

XNOR2xp5_ASAP7_75t_SL g445 ( 
.A(n_408),
.B(n_386),
.Y(n_445)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_411),
.Y(n_436)
);

AOI21xp5_ASAP7_75t_L g413 ( 
.A1(n_359),
.A2(n_302),
.B(n_322),
.Y(n_413)
);

OAI21xp5_ASAP7_75t_SL g443 ( 
.A1(n_413),
.A2(n_414),
.B(n_428),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g414 ( 
.A1(n_392),
.A2(n_306),
.B(n_312),
.Y(n_414)
);

AOI32xp33_ASAP7_75t_L g417 ( 
.A1(n_351),
.A2(n_306),
.A3(n_312),
.B1(n_365),
.B2(n_358),
.Y(n_417)
);

INVxp67_ASAP7_75t_L g460 ( 
.A(n_417),
.Y(n_460)
);

OAI22xp5_ASAP7_75t_SL g418 ( 
.A1(n_353),
.A2(n_365),
.B1(n_369),
.B2(n_377),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_357),
.B(n_372),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_L g440 ( 
.A(n_420),
.B(n_367),
.Y(n_440)
);

CKINVDCx20_ASAP7_75t_R g421 ( 
.A(n_354),
.Y(n_421)
);

INVx1_ASAP7_75t_L g423 ( 
.A(n_370),
.Y(n_423)
);

INVx1_ASAP7_75t_L g451 ( 
.A(n_423),
.Y(n_451)
);

OAI22xp5_ASAP7_75t_SL g425 ( 
.A1(n_369),
.A2(n_355),
.B1(n_374),
.B2(n_352),
.Y(n_425)
);

AO21x2_ASAP7_75t_L g427 ( 
.A1(n_373),
.A2(n_384),
.B(n_363),
.Y(n_427)
);

INVx1_ASAP7_75t_SL g444 ( 
.A(n_427),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_SL g428 ( 
.A1(n_385),
.A2(n_361),
.B(n_352),
.Y(n_428)
);

OAI22xp5_ASAP7_75t_SL g429 ( 
.A1(n_424),
.A2(n_376),
.B1(n_380),
.B2(n_360),
.Y(n_429)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_429),
.A2(n_431),
.B1(n_433),
.B2(n_438),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g430 ( 
.A(n_428),
.B(n_371),
.Y(n_430)
);

XOR2xp5_ASAP7_75t_L g477 ( 
.A(n_430),
.B(n_445),
.Y(n_477)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_424),
.A2(n_356),
.B1(n_362),
.B2(n_387),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g433 ( 
.A1(n_427),
.A2(n_402),
.B1(n_400),
.B2(n_420),
.Y(n_433)
);

CKINVDCx16_ASAP7_75t_R g434 ( 
.A(n_416),
.Y(n_434)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_434),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_L g435 ( 
.A(n_408),
.B(n_383),
.Y(n_435)
);

MAJIxp5_ASAP7_75t_L g467 ( 
.A(n_435),
.B(n_439),
.C(n_447),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_437),
.A2(n_442),
.B1(n_449),
.B2(n_454),
.Y(n_463)
);

OAI22xp5_ASAP7_75t_SL g438 ( 
.A1(n_427),
.A2(n_402),
.B1(n_400),
.B2(n_394),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g439 ( 
.A(n_425),
.B(n_383),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g474 ( 
.A(n_440),
.B(n_456),
.Y(n_474)
);

AOI22xp5_ASAP7_75t_L g442 ( 
.A1(n_412),
.A2(n_393),
.B1(n_378),
.B2(n_381),
.Y(n_442)
);

XNOR2xp5_ASAP7_75t_SL g489 ( 
.A(n_445),
.B(n_429),
.Y(n_489)
);

OAI22xp5_ASAP7_75t_SL g446 ( 
.A1(n_427),
.A2(n_356),
.B1(n_362),
.B2(n_364),
.Y(n_446)
);

AOI22xp5_ASAP7_75t_SL g479 ( 
.A1(n_446),
.A2(n_450),
.B1(n_431),
.B2(n_444),
.Y(n_479)
);

NAND2xp5_ASAP7_75t_L g448 ( 
.A(n_399),
.B(n_354),
.Y(n_448)
);

INVx1_ASAP7_75t_L g472 ( 
.A(n_448),
.Y(n_472)
);

AOI22xp5_ASAP7_75t_L g449 ( 
.A1(n_418),
.A2(n_388),
.B1(n_390),
.B2(n_394),
.Y(n_449)
);

OAI22xp5_ASAP7_75t_SL g450 ( 
.A1(n_427),
.A2(n_409),
.B1(n_405),
.B2(n_413),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_L g452 ( 
.A1(n_409),
.A2(n_403),
.B(n_416),
.Y(n_452)
);

OAI21xp5_ASAP7_75t_SL g470 ( 
.A1(n_452),
.A2(n_415),
.B(n_423),
.Y(n_470)
);

INVx1_ASAP7_75t_L g453 ( 
.A(n_396),
.Y(n_453)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_453),
.Y(n_476)
);

AOI22xp5_ASAP7_75t_L g454 ( 
.A1(n_411),
.A2(n_397),
.B1(n_419),
.B2(n_417),
.Y(n_454)
);

MAJIxp5_ASAP7_75t_L g455 ( 
.A(n_404),
.B(n_395),
.C(n_419),
.Y(n_455)
);

MAJIxp5_ASAP7_75t_L g468 ( 
.A(n_455),
.B(n_398),
.C(n_407),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g456 ( 
.A(n_426),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_L g457 ( 
.A(n_421),
.B(n_395),
.Y(n_457)
);

INVx1_ASAP7_75t_L g483 ( 
.A(n_457),
.Y(n_483)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_396),
.Y(n_458)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_458),
.Y(n_484)
);

CKINVDCx20_ASAP7_75t_R g459 ( 
.A(n_422),
.Y(n_459)
);

NAND2xp5_ASAP7_75t_L g487 ( 
.A(n_459),
.B(n_458),
.Y(n_487)
);

CKINVDCx20_ASAP7_75t_R g461 ( 
.A(n_457),
.Y(n_461)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_461),
.B(n_464),
.Y(n_492)
);

OAI22xp5_ASAP7_75t_L g462 ( 
.A1(n_444),
.A2(n_397),
.B1(n_414),
.B2(n_410),
.Y(n_462)
);

OAI22xp5_ASAP7_75t_L g498 ( 
.A1(n_462),
.A2(n_471),
.B1(n_453),
.B2(n_451),
.Y(n_498)
);

OAI21xp5_ASAP7_75t_L g464 ( 
.A1(n_443),
.A2(n_410),
.B(n_407),
.Y(n_464)
);

CKINVDCx16_ASAP7_75t_R g466 ( 
.A(n_441),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g513 ( 
.A(n_466),
.B(n_478),
.Y(n_513)
);

MAJIxp5_ASAP7_75t_L g497 ( 
.A(n_468),
.B(n_475),
.C(n_486),
.Y(n_497)
);

XOR2xp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_398),
.Y(n_469)
);

XOR2xp5_ASAP7_75t_L g509 ( 
.A(n_469),
.B(n_467),
.Y(n_509)
);

AOI21xp5_ASAP7_75t_L g490 ( 
.A1(n_470),
.A2(n_473),
.B(n_482),
.Y(n_490)
);

OAI22xp5_ASAP7_75t_L g471 ( 
.A1(n_444),
.A2(n_415),
.B1(n_422),
.B2(n_401),
.Y(n_471)
);

NAND2xp33_ASAP7_75t_SL g473 ( 
.A(n_443),
.B(n_401),
.Y(n_473)
);

MAJIxp5_ASAP7_75t_L g475 ( 
.A(n_435),
.B(n_455),
.C(n_447),
.Y(n_475)
);

XNOR2x1_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_469),
.Y(n_505)
);

INVxp67_ASAP7_75t_L g478 ( 
.A(n_452),
.Y(n_478)
);

OAI22xp5_ASAP7_75t_SL g495 ( 
.A1(n_479),
.A2(n_442),
.B1(n_432),
.B2(n_450),
.Y(n_495)
);

CKINVDCx20_ASAP7_75t_R g480 ( 
.A(n_441),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_480),
.B(n_485),
.Y(n_504)
);

OAI21xp5_ASAP7_75t_SL g482 ( 
.A1(n_432),
.A2(n_460),
.B(n_454),
.Y(n_482)
);

OAI22xp5_ASAP7_75t_SL g485 ( 
.A1(n_436),
.A2(n_437),
.B1(n_449),
.B2(n_434),
.Y(n_485)
);

MAJIxp5_ASAP7_75t_L g486 ( 
.A(n_430),
.B(n_440),
.C(n_448),
.Y(n_486)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_487),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_436),
.B(n_459),
.Y(n_488)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_488),
.Y(n_508)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_489),
.B(n_477),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_466),
.B(n_480),
.Y(n_491)
);

INVx1_ASAP7_75t_L g530 ( 
.A(n_491),
.Y(n_530)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_468),
.B(n_456),
.Y(n_493)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_493),
.Y(n_516)
);

OA21x2_ASAP7_75t_L g494 ( 
.A1(n_473),
.A2(n_433),
.B(n_438),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g523 ( 
.A1(n_494),
.A2(n_495),
.B1(n_498),
.B2(n_463),
.Y(n_523)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_486),
.B(n_451),
.Y(n_496)
);

INVx1_ASAP7_75t_L g520 ( 
.A(n_496),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g499 ( 
.A(n_467),
.B(n_446),
.C(n_475),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g514 ( 
.A(n_499),
.B(n_477),
.C(n_489),
.Y(n_514)
);

OAI22xp5_ASAP7_75t_L g500 ( 
.A1(n_481),
.A2(n_461),
.B1(n_483),
.B2(n_479),
.Y(n_500)
);

OAI22xp5_ASAP7_75t_L g515 ( 
.A1(n_500),
.A2(n_503),
.B1(n_507),
.B2(n_481),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g501 ( 
.A(n_474),
.B(n_470),
.Y(n_501)
);

INVx1_ASAP7_75t_L g521 ( 
.A(n_501),
.Y(n_521)
);

CKINVDCx20_ASAP7_75t_R g503 ( 
.A(n_487),
.Y(n_503)
);

XNOR2xp5_ASAP7_75t_SL g517 ( 
.A(n_505),
.B(n_506),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_SL g507 ( 
.A1(n_462),
.A2(n_463),
.B1(n_465),
.B2(n_472),
.Y(n_507)
);

XOR2xp5_ASAP7_75t_L g519 ( 
.A(n_509),
.B(n_489),
.Y(n_519)
);

NOR2xp67_ASAP7_75t_R g510 ( 
.A(n_474),
.B(n_472),
.Y(n_510)
);

XNOR2x1_ASAP7_75t_L g522 ( 
.A(n_510),
.B(n_465),
.Y(n_522)
);

INVx1_ASAP7_75t_L g511 ( 
.A(n_483),
.Y(n_511)
);

INVx1_ASAP7_75t_L g525 ( 
.A(n_511),
.Y(n_525)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_476),
.Y(n_512)
);

INVx1_ASAP7_75t_L g526 ( 
.A(n_512),
.Y(n_526)
);

XNOR2xp5_ASAP7_75t_L g532 ( 
.A(n_514),
.B(n_518),
.Y(n_532)
);

AOI22xp5_ASAP7_75t_L g534 ( 
.A1(n_515),
.A2(n_523),
.B1(n_495),
.B2(n_494),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g518 ( 
.A(n_497),
.B(n_464),
.Y(n_518)
);

XOR2xp5_ASAP7_75t_L g536 ( 
.A(n_519),
.B(n_524),
.Y(n_536)
);

INVx1_ASAP7_75t_L g537 ( 
.A(n_522),
.Y(n_537)
);

XOR2xp5_ASAP7_75t_L g524 ( 
.A(n_509),
.B(n_482),
.Y(n_524)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_497),
.B(n_485),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_L g539 ( 
.A(n_527),
.B(n_528),
.Y(n_539)
);

MAJIxp5_ASAP7_75t_L g528 ( 
.A(n_499),
.B(n_488),
.C(n_471),
.Y(n_528)
);

HB1xp67_ASAP7_75t_L g529 ( 
.A(n_500),
.Y(n_529)
);

INVx1_ASAP7_75t_L g545 ( 
.A(n_529),
.Y(n_545)
);

MAJIxp5_ASAP7_75t_L g531 ( 
.A(n_528),
.B(n_505),
.C(n_506),
.Y(n_531)
);

MAJIxp5_ASAP7_75t_L g557 ( 
.A(n_531),
.B(n_533),
.C(n_541),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g533 ( 
.A(n_527),
.B(n_513),
.C(n_498),
.Y(n_533)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_534),
.A2(n_503),
.B1(n_508),
.B2(n_502),
.Y(n_552)
);

NOR2xp33_ASAP7_75t_L g535 ( 
.A(n_516),
.B(n_513),
.Y(n_535)
);

NOR2xp33_ASAP7_75t_SL g546 ( 
.A(n_535),
.B(n_540),
.Y(n_546)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_526),
.Y(n_538)
);

INVx1_ASAP7_75t_L g550 ( 
.A(n_538),
.Y(n_550)
);

BUFx24_ASAP7_75t_SL g540 ( 
.A(n_520),
.Y(n_540)
);

MAJIxp5_ASAP7_75t_L g541 ( 
.A(n_518),
.B(n_504),
.C(n_490),
.Y(n_541)
);

AOI22xp5_ASAP7_75t_L g542 ( 
.A1(n_521),
.A2(n_492),
.B1(n_501),
.B2(n_508),
.Y(n_542)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_542),
.Y(n_555)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_523),
.A2(n_492),
.B(n_490),
.Y(n_543)
);

OR2x2_ASAP7_75t_L g551 ( 
.A(n_543),
.B(n_494),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g544 ( 
.A(n_514),
.B(n_524),
.C(n_519),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g554 ( 
.A(n_544),
.B(n_517),
.Y(n_554)
);

XNOR2xp5_ASAP7_75t_L g547 ( 
.A(n_532),
.B(n_530),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_547),
.B(n_549),
.Y(n_560)
);

XOR2xp5_ASAP7_75t_L g548 ( 
.A(n_536),
.B(n_517),
.Y(n_548)
);

XNOR2xp5_ASAP7_75t_L g559 ( 
.A(n_548),
.B(n_553),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g549 ( 
.A(n_532),
.B(n_504),
.Y(n_549)
);

INVxp67_ASAP7_75t_L g563 ( 
.A(n_551),
.Y(n_563)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_552),
.B(n_491),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g553 ( 
.A(n_541),
.B(n_522),
.Y(n_553)
);

NOR2xp33_ASAP7_75t_SL g558 ( 
.A(n_554),
.B(n_556),
.Y(n_558)
);

INVx1_ASAP7_75t_L g556 ( 
.A(n_545),
.Y(n_556)
);

AOI21x1_ASAP7_75t_L g561 ( 
.A1(n_555),
.A2(n_537),
.B(n_543),
.Y(n_561)
);

OAI21xp5_ASAP7_75t_SL g567 ( 
.A1(n_561),
.A2(n_562),
.B(n_566),
.Y(n_567)
);

AOI21xp5_ASAP7_75t_L g562 ( 
.A1(n_547),
.A2(n_539),
.B(n_533),
.Y(n_562)
);

NOR2xp67_ASAP7_75t_SL g564 ( 
.A(n_557),
.B(n_553),
.Y(n_564)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_564),
.Y(n_572)
);

NAND2xp5_ASAP7_75t_L g568 ( 
.A(n_565),
.B(n_563),
.Y(n_568)
);

OAI21xp5_ASAP7_75t_SL g566 ( 
.A1(n_551),
.A2(n_502),
.B(n_544),
.Y(n_566)
);

NAND2xp5_ASAP7_75t_L g575 ( 
.A(n_568),
.B(n_570),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_SL g569 ( 
.A(n_558),
.B(n_546),
.Y(n_569)
);

OR2x2_ASAP7_75t_L g576 ( 
.A(n_569),
.B(n_571),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g570 ( 
.A(n_560),
.B(n_550),
.Y(n_570)
);

NAND2xp5_ASAP7_75t_L g571 ( 
.A(n_563),
.B(n_552),
.Y(n_571)
);

XNOR2xp5_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_557),
.Y(n_573)
);

MAJIxp5_ASAP7_75t_L g577 ( 
.A(n_573),
.B(n_574),
.C(n_572),
.Y(n_577)
);

AOI321xp33_ASAP7_75t_SL g574 ( 
.A1(n_572),
.A2(n_510),
.A3(n_565),
.B1(n_549),
.B2(n_511),
.C(n_559),
.Y(n_574)
);

NAND4xp25_ASAP7_75t_L g579 ( 
.A(n_577),
.B(n_578),
.C(n_575),
.D(n_525),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g578 ( 
.A(n_576),
.B(n_559),
.C(n_531),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_579),
.B(n_512),
.C(n_484),
.Y(n_580)
);

AOI21xp5_ASAP7_75t_L g581 ( 
.A1(n_580),
.A2(n_476),
.B(n_484),
.Y(n_581)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_581),
.B(n_494),
.Y(n_582)
);

AOI21xp5_ASAP7_75t_L g583 ( 
.A1(n_582),
.A2(n_548),
.B(n_536),
.Y(n_583)
);


endmodule