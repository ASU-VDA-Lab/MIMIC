module fake_jpeg_6840_n_275 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_275);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_275;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_272;
wire n_171;
wire n_263;
wire n_119;
wire n_23;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_145;
wire n_20;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx4f_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_12),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

INVxp33_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_12),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

INVx13_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx3_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx16_ASAP7_75t_R g25 ( 
.A(n_6),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_7),
.Y(n_26)
);

BUFx3_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_13),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_28),
.B(n_30),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_21),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g31 ( 
.A(n_15),
.B(n_0),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_31),
.B(n_24),
.Y(n_44)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_21),
.Y(n_32)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_13),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_16),
.B(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_34),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_13),
.Y(n_35)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_35),
.Y(n_47)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_21),
.Y(n_36)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_36),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_13),
.Y(n_37)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_30),
.Y(n_40)
);

INVx5_ASAP7_75t_L g59 ( 
.A(n_40),
.Y(n_59)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_44),
.B(n_17),
.Y(n_66)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_45),
.Y(n_60)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_51),
.Y(n_55)
);

OAI22xp33_ASAP7_75t_L g48 ( 
.A1(n_31),
.A2(n_13),
.B1(n_18),
.B2(n_22),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_48),
.A2(n_14),
.B1(n_22),
.B2(n_33),
.Y(n_58)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_34),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_53),
.B(n_24),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_49),
.Y(n_54)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_54),
.Y(n_84)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_56),
.B(n_61),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_44),
.B(n_26),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_65),
.Y(n_86)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_58),
.A2(n_28),
.B1(n_52),
.B2(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_62),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_43),
.B(n_24),
.Y(n_63)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

A2O1A1Ixp33_ASAP7_75t_L g65 ( 
.A1(n_48),
.A2(n_14),
.B(n_22),
.C(n_17),
.Y(n_65)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_41),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_67),
.A2(n_71),
.B1(n_70),
.B2(n_68),
.Y(n_75)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_47),
.Y(n_68)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_68),
.Y(n_93)
);

AND2x2_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_28),
.Y(n_69)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_69),
.B(n_17),
.Y(n_76)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_47),
.Y(n_70)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_40),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_SL g72 ( 
.A(n_53),
.B(n_15),
.Y(n_72)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_72),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_45),
.Y(n_73)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_46),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_74),
.B(n_72),
.Y(n_96)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_63),
.Y(n_98)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_54),
.A2(n_52),
.B1(n_14),
.B2(n_50),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g110 ( 
.A1(n_80),
.A2(n_94),
.B1(n_26),
.B2(n_19),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g97 ( 
.A1(n_81),
.A2(n_89),
.B1(n_62),
.B2(n_70),
.Y(n_97)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_57),
.B(n_69),
.Y(n_85)
);

OAI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_85),
.A2(n_87),
.B(n_19),
.Y(n_106)
);

AND2x2_ASAP7_75t_L g87 ( 
.A(n_69),
.B(n_28),
.Y(n_87)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_65),
.A2(n_51),
.B1(n_50),
.B2(n_15),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_73),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_90),
.B(n_92),
.Y(n_101)
);

OA21x2_ASAP7_75t_L g91 ( 
.A1(n_65),
.A2(n_25),
.B(n_37),
.Y(n_91)
);

AOI21xp5_ASAP7_75t_L g100 ( 
.A1(n_91),
.A2(n_55),
.B(n_67),
.Y(n_100)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_73),
.Y(n_92)
);

INVxp67_ASAP7_75t_L g94 ( 
.A(n_55),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g95 ( 
.A1(n_86),
.A2(n_58),
.B1(n_66),
.B2(n_69),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_95),
.A2(n_105),
.B1(n_113),
.B2(n_87),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_L g119 ( 
.A(n_96),
.B(n_106),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_SL g117 ( 
.A1(n_97),
.A2(n_102),
.B1(n_107),
.B2(n_115),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_104),
.Y(n_120)
);

OR2x2_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_71),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g125 ( 
.A1(n_99),
.A2(n_100),
.B(n_106),
.Y(n_125)
);

AOI22xp5_ASAP7_75t_L g102 ( 
.A1(n_86),
.A2(n_61),
.B1(n_60),
.B2(n_59),
.Y(n_102)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_83),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_90),
.A2(n_60),
.B1(n_64),
.B2(n_59),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_89),
.A2(n_64),
.B1(n_59),
.B2(n_68),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_92),
.B(n_64),
.C(n_29),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_108),
.B(n_93),
.C(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_85),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_109),
.B(n_112),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g129 ( 
.A(n_110),
.Y(n_129)
);

BUFx2_ASAP7_75t_L g111 ( 
.A(n_77),
.Y(n_111)
);

BUFx2_ASAP7_75t_L g131 ( 
.A(n_111),
.Y(n_131)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_85),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g113 ( 
.A(n_74),
.B(n_29),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g114 ( 
.A1(n_79),
.A2(n_26),
.B1(n_19),
.B2(n_38),
.Y(n_114)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_87),
.A2(n_81),
.B1(n_91),
.B2(n_76),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_118),
.B(n_136),
.C(n_35),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_134),
.Y(n_151)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_105),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_121),
.B(n_132),
.Y(n_146)
);

INVx3_ASAP7_75t_L g122 ( 
.A(n_111),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_122),
.B(n_124),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_111),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_101),
.B(n_82),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_126),
.B(n_128),
.Y(n_139)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_127),
.A2(n_100),
.B(n_115),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_82),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_96),
.B(n_88),
.Y(n_130)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_130),
.Y(n_138)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_102),
.Y(n_132)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_107),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g158 ( 
.A(n_133),
.B(n_135),
.Y(n_158)
);

AOI322xp5_ASAP7_75t_L g134 ( 
.A1(n_113),
.A2(n_76),
.A3(n_88),
.B1(n_78),
.B2(n_91),
.C1(n_79),
.C2(n_94),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_108),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_109),
.B(n_78),
.C(n_93),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_113),
.B(n_112),
.Y(n_137)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_137),
.Y(n_141)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_103),
.B1(n_95),
.B2(n_97),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_140),
.A2(n_161),
.B1(n_123),
.B2(n_141),
.Y(n_178)
);

CKINVDCx16_ASAP7_75t_R g142 ( 
.A(n_120),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_142),
.B(n_154),
.Y(n_169)
);

XOR2xp5_ASAP7_75t_L g171 ( 
.A(n_143),
.B(n_149),
.Y(n_171)
);

XNOR2x1_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_98),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g166 ( 
.A(n_144),
.B(n_147),
.Y(n_166)
);

AO21x1_ASAP7_75t_SL g145 ( 
.A1(n_125),
.A2(n_103),
.B(n_99),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_145),
.B(n_20),
.Y(n_180)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_99),
.Y(n_147)
);

XNOR2x1_ASAP7_75t_L g148 ( 
.A(n_119),
.B(n_98),
.Y(n_148)
);

XNOR2xp5_ASAP7_75t_SL g174 ( 
.A(n_148),
.B(n_157),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_SL g149 ( 
.A1(n_116),
.A2(n_104),
.B(n_77),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g150 ( 
.A(n_118),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_150),
.B(n_160),
.Y(n_170)
);

XNOR2xp5_ASAP7_75t_L g153 ( 
.A(n_127),
.B(n_37),
.Y(n_153)
);

XOR2xp5_ASAP7_75t_L g179 ( 
.A(n_153),
.B(n_18),
.Y(n_179)
);

OAI22xp5_ASAP7_75t_SL g154 ( 
.A1(n_132),
.A2(n_38),
.B1(n_37),
.B2(n_35),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_155),
.B(n_133),
.C(n_129),
.Y(n_176)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_126),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_156),
.B(n_159),
.Y(n_168)
);

A2O1A1O1Ixp25_ASAP7_75t_L g157 ( 
.A1(n_137),
.A2(n_35),
.B(n_20),
.C(n_27),
.D(n_23),
.Y(n_157)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_128),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_130),
.B(n_56),
.Y(n_160)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_117),
.A2(n_18),
.B1(n_23),
.B2(n_21),
.Y(n_161)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_162),
.B(n_163),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g163 ( 
.A(n_149),
.Y(n_163)
);

INVx1_ASAP7_75t_L g164 ( 
.A(n_139),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_164),
.B(n_165),
.Y(n_196)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_139),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_151),
.B(n_136),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_173),
.Y(n_197)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_147),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_172),
.B(n_177),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_151),
.B(n_135),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_138),
.B(n_121),
.Y(n_175)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_175),
.Y(n_198)
);

MAJIxp5_ASAP7_75t_L g190 ( 
.A(n_176),
.B(n_179),
.C(n_183),
.Y(n_190)
);

NAND3xp33_ASAP7_75t_L g177 ( 
.A(n_148),
.B(n_123),
.C(n_27),
.Y(n_177)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_178),
.A2(n_181),
.B1(n_182),
.B2(n_154),
.Y(n_188)
);

INVx2_ASAP7_75t_L g200 ( 
.A(n_180),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_140),
.A2(n_122),
.B1(n_131),
.B2(n_124),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_147),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_155),
.B(n_124),
.C(n_131),
.Y(n_183)
);

XNOR2xp5_ASAP7_75t_L g184 ( 
.A(n_144),
.B(n_56),
.Y(n_184)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_184),
.B(n_20),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_176),
.A2(n_145),
.B1(n_161),
.B2(n_146),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_186),
.A2(n_192),
.B1(n_174),
.B2(n_23),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_SL g187 ( 
.A(n_166),
.B(n_150),
.Y(n_187)
);

MAJx2_ASAP7_75t_L g215 ( 
.A(n_187),
.B(n_199),
.C(n_0),
.Y(n_215)
);

OAI21xp5_ASAP7_75t_L g214 ( 
.A1(n_188),
.A2(n_23),
.B(n_20),
.Y(n_214)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_173),
.B(n_153),
.Y(n_189)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_189),
.B(n_201),
.C(n_203),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_170),
.A2(n_158),
.B1(n_181),
.B2(n_180),
.Y(n_192)
);

INVxp67_ASAP7_75t_L g193 ( 
.A(n_183),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_193),
.B(n_179),
.Y(n_206)
);

BUFx2_ASAP7_75t_L g194 ( 
.A(n_169),
.Y(n_194)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g195 ( 
.A1(n_178),
.A2(n_143),
.B1(n_157),
.B2(n_131),
.Y(n_195)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_195),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_167),
.B(n_171),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_171),
.A2(n_18),
.B1(n_1),
.B2(n_2),
.Y(n_202)
);

CKINVDCx16_ASAP7_75t_R g220 ( 
.A(n_202),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_184),
.B(n_27),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_200),
.A2(n_198),
.B1(n_193),
.B2(n_185),
.Y(n_204)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_204),
.A2(n_214),
.B1(n_216),
.B2(n_218),
.Y(n_225)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_206),
.B(n_215),
.C(n_203),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_196),
.B(n_168),
.Y(n_207)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_207),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g208 ( 
.A(n_191),
.B(n_11),
.Y(n_208)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_208),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_194),
.B(n_166),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g233 ( 
.A(n_209),
.Y(n_233)
);

AOI21xp5_ASAP7_75t_L g210 ( 
.A1(n_190),
.A2(n_174),
.B(n_27),
.Y(n_210)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_210),
.Y(n_229)
);

OAI22xp5_ASAP7_75t_SL g228 ( 
.A1(n_211),
.A2(n_219),
.B1(n_3),
.B2(n_4),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_199),
.B(n_0),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_212),
.B(n_3),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_187),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_216)
);

XNOR2x1_ASAP7_75t_L g218 ( 
.A(n_201),
.B(n_1),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g219 ( 
.A1(n_190),
.A2(n_1),
.B(n_2),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_204),
.B(n_207),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_230),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_223),
.B(n_231),
.C(n_213),
.Y(n_235)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_189),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_SL g240 ( 
.A(n_226),
.B(n_232),
.Y(n_240)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_209),
.B(n_197),
.Y(n_227)
);

AOI22x1_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_218),
.B1(n_215),
.B2(n_211),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_228),
.A2(n_214),
.B(n_5),
.Y(n_245)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_206),
.Y(n_230)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_213),
.B(n_197),
.C(n_210),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_205),
.B(n_3),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_234),
.B(n_220),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_235),
.B(n_241),
.C(n_4),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g253 ( 
.A1(n_237),
.A2(n_244),
.B(n_246),
.Y(n_253)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_238),
.Y(n_247)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_217),
.B1(n_220),
.B2(n_219),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_239),
.B(n_242),
.Y(n_248)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_231),
.B(n_216),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_223),
.B(n_212),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g243 ( 
.A(n_233),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_243),
.B(n_227),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g244 ( 
.A(n_224),
.B(n_217),
.Y(n_244)
);

OR2x2_ASAP7_75t_L g250 ( 
.A(n_245),
.B(n_228),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_222),
.B(n_4),
.Y(n_246)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_249),
.Y(n_261)
);

AND2x2_ASAP7_75t_L g258 ( 
.A(n_250),
.B(n_254),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_240),
.B(n_227),
.Y(n_251)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_251),
.Y(n_263)
);

AND2x2_ASAP7_75t_L g252 ( 
.A(n_241),
.B(n_229),
.Y(n_252)
);

AOI21xp5_ASAP7_75t_L g262 ( 
.A1(n_252),
.A2(n_255),
.B(n_8),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_237),
.A2(n_225),
.B1(n_229),
.B2(n_236),
.Y(n_254)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_243),
.A2(n_4),
.B(n_5),
.Y(n_255)
);

OAI21xp5_ASAP7_75t_L g260 ( 
.A1(n_256),
.A2(n_7),
.B(n_8),
.Y(n_260)
);

BUFx4f_ASAP7_75t_SL g257 ( 
.A(n_252),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_257),
.B(n_248),
.C(n_249),
.Y(n_264)
);

AOI22xp33_ASAP7_75t_L g259 ( 
.A1(n_253),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g266 ( 
.A1(n_259),
.A2(n_247),
.B1(n_9),
.B2(n_10),
.Y(n_266)
);

NOR3xp33_ASAP7_75t_SL g267 ( 
.A(n_260),
.B(n_9),
.C(n_10),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_262),
.B(n_9),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g269 ( 
.A1(n_264),
.A2(n_265),
.B(n_266),
.Y(n_269)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_258),
.B(n_250),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_SL g270 ( 
.A1(n_267),
.A2(n_268),
.B(n_261),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g272 ( 
.A(n_270),
.Y(n_272)
);

OAI21xp5_ASAP7_75t_L g271 ( 
.A1(n_269),
.A2(n_263),
.B(n_265),
.Y(n_271)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_271),
.A2(n_10),
.B(n_272),
.Y(n_273)
);

HB1xp67_ASAP7_75t_L g274 ( 
.A(n_273),
.Y(n_274)
);

FAx1_ASAP7_75t_SL g275 ( 
.A(n_274),
.B(n_10),
.CI(n_249),
.CON(n_275),
.SN(n_275)
);


endmodule