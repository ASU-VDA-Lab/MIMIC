module fake_jpeg_19387_n_263 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_263);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_263;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_223;
wire n_187;
wire n_21;
wire n_57;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_170;
wire n_162;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_217;
wire n_216;
wire n_184;
wire n_53;
wire n_33;
wire n_93;
wire n_54;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_258;
wire n_96;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_14),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

INVx6_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

BUFx8_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

CKINVDCx14_ASAP7_75t_R g24 ( 
.A(n_4),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_4),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_0),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_12),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_14),
.Y(n_30)
);

INVx11_ASAP7_75t_SL g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_3),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g33 ( 
.A(n_11),
.Y(n_33)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_15),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_20),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_35),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_20),
.Y(n_36)
);

INVx6_ASAP7_75t_L g48 ( 
.A(n_36),
.Y(n_48)
);

INVx6_ASAP7_75t_SL g37 ( 
.A(n_20),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_37),
.B(n_45),
.Y(n_51)
);

INVx3_ASAP7_75t_L g38 ( 
.A(n_20),
.Y(n_38)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_0),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_17),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_20),
.Y(n_40)
);

INVx6_ASAP7_75t_L g54 ( 
.A(n_40),
.Y(n_54)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_41),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_24),
.B(n_1),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_42),
.B(n_18),
.Y(n_55)
);

BUFx5_ASAP7_75t_L g43 ( 
.A(n_31),
.Y(n_43)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_43),
.Y(n_50)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_34),
.Y(n_44)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_44),
.Y(n_53)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_34),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g46 ( 
.A1(n_39),
.A2(n_19),
.B1(n_22),
.B2(n_28),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_46),
.A2(n_47),
.B1(n_49),
.B2(n_68),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g47 ( 
.A1(n_44),
.A2(n_19),
.B1(n_22),
.B2(n_28),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g49 ( 
.A1(n_45),
.A2(n_22),
.B1(n_28),
.B2(n_21),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g52 ( 
.A(n_41),
.B(n_17),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_SL g73 ( 
.A1(n_52),
.A2(n_67),
.B(n_58),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_SL g83 ( 
.A(n_55),
.B(n_62),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_56),
.B(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_42),
.B(n_27),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_63),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_35),
.B(n_34),
.Y(n_58)
);

INVx3_ASAP7_75t_L g60 ( 
.A(n_37),
.Y(n_60)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_60),
.Y(n_91)
);

MAJIxp5_ASAP7_75t_L g62 ( 
.A(n_38),
.B(n_35),
.C(n_40),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_37),
.B(n_27),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_38),
.B(n_26),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_17),
.Y(n_82)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_36),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_66),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_34),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_67),
.B(n_17),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_40),
.A2(n_22),
.B1(n_21),
.B2(n_25),
.Y(n_68)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_53),
.Y(n_70)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_53),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_71),
.B(n_76),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_73),
.B(n_16),
.Y(n_124)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_65),
.Y(n_74)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_74),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_56),
.A2(n_21),
.B1(n_30),
.B2(n_29),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g127 ( 
.A1(n_75),
.A2(n_72),
.B1(n_97),
.B2(n_101),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_50),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_60),
.A2(n_31),
.B1(n_18),
.B2(n_29),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g113 ( 
.A(n_77),
.Y(n_113)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_65),
.Y(n_79)
);

INVx4_ASAP7_75t_L g134 ( 
.A(n_79),
.Y(n_134)
);

NAND2xp33_ASAP7_75t_SL g80 ( 
.A(n_52),
.B(n_61),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g131 ( 
.A1(n_80),
.A2(n_105),
.B(n_5),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_82),
.B(n_100),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_48),
.A2(n_18),
.B1(n_32),
.B2(n_30),
.Y(n_84)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_84),
.A2(n_85),
.B1(n_87),
.B2(n_96),
.Y(n_111)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_61),
.Y(n_86)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_86),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_48),
.A2(n_25),
.B1(n_32),
.B2(n_26),
.Y(n_87)
);

OAI21xp33_ASAP7_75t_L g88 ( 
.A1(n_55),
.A2(n_1),
.B(n_2),
.Y(n_88)
);

A2O1A1Ixp33_ASAP7_75t_L g118 ( 
.A1(n_88),
.A2(n_1),
.B(n_2),
.C(n_5),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_89),
.B(n_93),
.Y(n_117)
);

OA22x2_ASAP7_75t_L g90 ( 
.A1(n_48),
.A2(n_54),
.B1(n_52),
.B2(n_46),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_90),
.A2(n_104),
.B1(n_43),
.B2(n_23),
.Y(n_107)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_59),
.Y(n_92)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_92),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_51),
.B(n_24),
.Y(n_93)
);

INVx1_ASAP7_75t_SL g94 ( 
.A(n_50),
.Y(n_94)
);

INVx1_ASAP7_75t_SL g123 ( 
.A(n_94),
.Y(n_123)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_49),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_95),
.B(n_102),
.Y(n_132)
);

INVx3_ASAP7_75t_SL g96 ( 
.A(n_59),
.Y(n_96)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_68),
.Y(n_97)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_97),
.Y(n_120)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

AOI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_54),
.A2(n_23),
.B1(n_17),
.B2(n_34),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g136 ( 
.A1(n_99),
.A2(n_14),
.B1(n_7),
.B2(n_8),
.Y(n_136)
);

CKINVDCx16_ASAP7_75t_R g100 ( 
.A(n_62),
.Y(n_100)
);

AND2x2_ASAP7_75t_SL g101 ( 
.A(n_47),
.B(n_43),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_101),
.B(n_16),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_54),
.B(n_33),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_55),
.B(n_33),
.Y(n_103)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_103),
.Y(n_121)
);

OA22x2_ASAP7_75t_L g104 ( 
.A1(n_53),
.A2(n_23),
.B1(n_17),
.B2(n_33),
.Y(n_104)
);

AOI21xp33_ASAP7_75t_L g105 ( 
.A1(n_55),
.A2(n_23),
.B(n_15),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_55),
.B(n_33),
.Y(n_106)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_106),
.Y(n_122)
);

AO22x1_ASAP7_75t_L g150 ( 
.A1(n_107),
.A2(n_112),
.B1(n_104),
.B2(n_80),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_95),
.A2(n_16),
.B1(n_23),
.B2(n_33),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_110),
.A2(n_127),
.B1(n_129),
.B2(n_133),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_118),
.Y(n_154)
);

XNOR2xp5_ASAP7_75t_SL g162 ( 
.A(n_124),
.B(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_78),
.B(n_16),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_137),
.Y(n_139)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_86),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_SL g148 ( 
.A(n_128),
.B(n_130),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_78),
.A2(n_90),
.B1(n_89),
.B2(n_101),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_79),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_90),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_133)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

INVx4_ASAP7_75t_L g144 ( 
.A(n_135),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_SL g141 ( 
.A1(n_136),
.A2(n_96),
.B1(n_85),
.B2(n_94),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g137 ( 
.A1(n_90),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_73),
.A2(n_6),
.B1(n_8),
.B2(n_9),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_138),
.B(n_75),
.Y(n_149)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_140),
.Y(n_170)
);

INVxp67_ASAP7_75t_L g168 ( 
.A(n_141),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_109),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_142),
.B(n_143),
.Y(n_189)
);

CKINVDCx20_ASAP7_75t_R g143 ( 
.A(n_108),
.Y(n_143)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_116),
.Y(n_145)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_145),
.Y(n_171)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_120),
.Y(n_146)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_146),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_121),
.B(n_83),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_147),
.B(n_156),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_149),
.B(n_150),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_125),
.B(n_83),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_152),
.B(n_157),
.Y(n_182)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_134),
.Y(n_153)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_153),
.Y(n_178)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_134),
.Y(n_155)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_155),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_122),
.B(n_76),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_129),
.B(n_124),
.Y(n_157)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_158),
.B(n_161),
.Y(n_184)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_127),
.Y(n_159)
);

CKINVDCx20_ASAP7_75t_R g180 ( 
.A(n_159),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g160 ( 
.A(n_119),
.B(n_70),
.C(n_71),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_160),
.B(n_165),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_112),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_110),
.Y(n_163)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_163),
.Y(n_185)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_115),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_164),
.A2(n_166),
.B(n_104),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_131),
.B(n_81),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_133),
.B(n_104),
.Y(n_166)
);

OAI21xp5_ASAP7_75t_L g167 ( 
.A1(n_154),
.A2(n_113),
.B(n_107),
.Y(n_167)
);

OAI21xp5_ASAP7_75t_L g206 ( 
.A1(n_167),
.A2(n_172),
.B(n_177),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_SL g169 ( 
.A1(n_140),
.A2(n_118),
.B(n_137),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_169),
.A2(n_172),
.B(n_175),
.Y(n_193)
);

AOI21xp5_ASAP7_75t_SL g172 ( 
.A1(n_159),
.A2(n_113),
.B(n_138),
.Y(n_172)
);

AOI21xp5_ASAP7_75t_L g175 ( 
.A1(n_157),
.A2(n_123),
.B(n_111),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_151),
.A2(n_123),
.B1(n_96),
.B2(n_92),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_176),
.A2(n_186),
.B1(n_187),
.B2(n_143),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g207 ( 
.A1(n_177),
.A2(n_150),
.B(n_155),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_166),
.A2(n_139),
.B1(n_163),
.B2(n_149),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_181),
.B(n_150),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g186 ( 
.A1(n_151),
.A2(n_126),
.B1(n_135),
.B2(n_115),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_139),
.A2(n_126),
.B1(n_98),
.B2(n_91),
.Y(n_187)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_168),
.A2(n_158),
.B(n_146),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_202),
.Y(n_219)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_191),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_192),
.A2(n_171),
.B1(n_178),
.B2(n_179),
.Y(n_215)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_171),
.Y(n_194)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_194),
.Y(n_222)
);

OAI21xp33_ASAP7_75t_L g195 ( 
.A1(n_170),
.A2(n_165),
.B(n_161),
.Y(n_195)
);

NOR2xp33_ASAP7_75t_SL g221 ( 
.A(n_195),
.B(n_208),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g196 ( 
.A(n_174),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_196),
.B(n_198),
.Y(n_220)
);

AND2x2_ASAP7_75t_L g197 ( 
.A(n_176),
.B(n_186),
.Y(n_197)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_197),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g198 ( 
.A(n_173),
.B(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_162),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_SL g216 ( 
.A(n_199),
.B(n_200),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_162),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_201),
.B(n_203),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g202 ( 
.A(n_182),
.B(n_152),
.Y(n_202)
);

XNOR2xp5_ASAP7_75t_L g203 ( 
.A(n_188),
.B(n_160),
.Y(n_203)
);

INVxp67_ASAP7_75t_L g204 ( 
.A(n_175),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_204),
.B(n_207),
.Y(n_213)
);

CKINVDCx16_ASAP7_75t_R g205 ( 
.A(n_174),
.Y(n_205)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_205),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g209 ( 
.A1(n_206),
.A2(n_167),
.B1(n_180),
.B2(n_185),
.Y(n_209)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_188),
.B(n_148),
.Y(n_208)
);

INVxp67_ASAP7_75t_L g233 ( 
.A(n_209),
.Y(n_233)
);

INVx8_ASAP7_75t_L g210 ( 
.A(n_190),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_210),
.B(n_193),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_201),
.A2(n_168),
.B1(n_187),
.B2(n_181),
.Y(n_214)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_214),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_SL g236 ( 
.A1(n_215),
.A2(n_217),
.B1(n_144),
.B2(n_164),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_197),
.A2(n_169),
.B1(n_179),
.B2(n_178),
.Y(n_217)
);

CKINVDCx16_ASAP7_75t_R g224 ( 
.A(n_220),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_224),
.B(n_225),
.Y(n_243)
);

XOR2xp5_ASAP7_75t_L g225 ( 
.A(n_216),
.B(n_199),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g226 ( 
.A1(n_221),
.A2(n_206),
.B1(n_204),
.B2(n_193),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_228),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g229 ( 
.A(n_211),
.B(n_203),
.Y(n_229)
);

AND2x2_ASAP7_75t_L g239 ( 
.A(n_229),
.B(n_235),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g230 ( 
.A1(n_213),
.A2(n_207),
.B(n_197),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g242 ( 
.A1(n_230),
.A2(n_212),
.B(n_216),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_217),
.A2(n_192),
.B1(n_202),
.B2(n_200),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g241 ( 
.A1(n_231),
.A2(n_232),
.B1(n_221),
.B2(n_211),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_212),
.B(n_145),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g234 ( 
.A1(n_223),
.A2(n_153),
.B1(n_144),
.B2(n_91),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_234),
.A2(n_215),
.B1(n_222),
.B2(n_218),
.Y(n_240)
);

BUFx10_ASAP7_75t_L g235 ( 
.A(n_218),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g238 ( 
.A1(n_236),
.A2(n_210),
.B1(n_219),
.B2(n_222),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_233),
.A2(n_213),
.B(n_223),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_237),
.B(n_238),
.Y(n_248)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_240),
.A2(n_241),
.B1(n_245),
.B2(n_236),
.Y(n_246)
);

OAI21xp5_ASAP7_75t_SL g249 ( 
.A1(n_242),
.A2(n_227),
.B(n_234),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_233),
.A2(n_69),
.B1(n_11),
.B2(n_12),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_246),
.A2(n_238),
.B1(n_237),
.B2(n_239),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_244),
.B(n_229),
.C(n_225),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_L g254 ( 
.A(n_247),
.B(n_249),
.Y(n_254)
);

NOR2xp67_ASAP7_75t_SL g250 ( 
.A(n_240),
.B(n_235),
.Y(n_250)
);

INVxp67_ASAP7_75t_L g252 ( 
.A(n_250),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g251 ( 
.A(n_243),
.B(n_235),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_251),
.B(n_239),
.Y(n_253)
);

INVxp67_ASAP7_75t_L g256 ( 
.A(n_253),
.Y(n_256)
);

AOI21xp5_ASAP7_75t_L g257 ( 
.A1(n_255),
.A2(n_248),
.B(n_239),
.Y(n_257)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_257),
.B(n_252),
.Y(n_260)
);

OAI21xp5_ASAP7_75t_SL g258 ( 
.A1(n_254),
.A2(n_248),
.B(n_235),
.Y(n_258)
);

MAJx2_ASAP7_75t_L g259 ( 
.A(n_258),
.B(n_252),
.C(n_13),
.Y(n_259)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_259),
.Y(n_261)
);

OAI21x1_ASAP7_75t_L g262 ( 
.A1(n_261),
.A2(n_256),
.B(n_260),
.Y(n_262)
);

XNOR2xp5_ASAP7_75t_L g263 ( 
.A(n_262),
.B(n_69),
.Y(n_263)
);


endmodule