module fake_aes_247_n_16 (n_3, n_1, n_2, n_0, n_16);
input n_3;
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
NAND2xp5_ASAP7_75t_SL g4 ( .A(n_0), .B(n_2), .Y(n_4) );
NAND3xp33_ASAP7_75t_L g5 ( .A(n_1), .B(n_0), .C(n_2), .Y(n_5) );
AND2x2_ASAP7_75t_SL g6 ( .A(n_2), .B(n_1), .Y(n_6) );
AND2x2_ASAP7_75t_L g7 ( .A(n_0), .B(n_3), .Y(n_7) );
INVx1_ASAP7_75t_L g8 ( .A(n_7), .Y(n_8) );
OR2x2_ASAP7_75t_L g9 ( .A(n_4), .B(n_5), .Y(n_9) );
INVx1_ASAP7_75t_L g10 ( .A(n_6), .Y(n_10) );
INVx1_ASAP7_75t_L g11 ( .A(n_8), .Y(n_11) );
AOI33xp33_ASAP7_75t_L g12 ( .A1(n_10), .A2(n_1), .A3(n_3), .B1(n_5), .B2(n_8), .B3(n_7), .Y(n_12) );
AND2x2_ASAP7_75t_L g13 ( .A(n_11), .B(n_9), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_11), .B(n_9), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_13), .Y(n_15) );
AOI22xp5_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_14), .B1(n_12), .B2(n_3), .Y(n_16) );
endmodule