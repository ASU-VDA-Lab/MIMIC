module fake_jpeg_21605_n_164 (n_13, n_21, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_14, n_40, n_19, n_18, n_20, n_35, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_12, n_32, n_8, n_15, n_7, n_164);

input n_13;
input n_21;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_164;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_51;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_155;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_106;
wire n_111;
wire n_143;
wire n_75;
wire n_122;
wire n_102;
wire n_99;
wire n_130;
wire n_121;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_78;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_107;
wire n_72;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_162;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_91;
wire n_93;
wire n_54;
wire n_161;
wire n_138;
wire n_101;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_153;
wire n_135;
wire n_62;
wire n_120;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_10),
.Y(n_48)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_1),
.Y(n_50)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_38),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_31),
.Y(n_52)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_41),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

INVx5_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

BUFx6f_ASAP7_75t_SL g56 ( 
.A(n_5),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_17),
.Y(n_58)
);

INVx8_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

CKINVDCx5p33_ASAP7_75t_R g60 ( 
.A(n_2),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g61 ( 
.A(n_25),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_11),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_46),
.Y(n_63)
);

INVx6_ASAP7_75t_SL g64 ( 
.A(n_47),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_8),
.Y(n_65)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_45),
.Y(n_67)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g69 ( 
.A(n_18),
.Y(n_69)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_39),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_0),
.B(n_5),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_10),
.Y(n_72)
);

BUFx12f_ASAP7_75t_L g73 ( 
.A(n_6),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_21),
.Y(n_75)
);

INVx13_ASAP7_75t_L g76 ( 
.A(n_35),
.Y(n_76)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_57),
.Y(n_77)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

INVx11_ASAP7_75t_L g78 ( 
.A(n_57),
.Y(n_78)
);

INVx6_ASAP7_75t_L g86 ( 
.A(n_78),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g79 ( 
.A(n_49),
.B(n_73),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_79),
.B(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_71),
.B(n_1),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_80),
.B(n_81),
.Y(n_84)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_60),
.Y(n_81)
);

INVx8_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx6_ASAP7_75t_L g94 ( 
.A(n_82),
.Y(n_94)
);

INVx4_ASAP7_75t_L g83 ( 
.A(n_58),
.Y(n_83)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_83),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_83),
.A2(n_55),
.B1(n_70),
.B2(n_59),
.Y(n_85)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_85),
.A2(n_82),
.B1(n_78),
.B2(n_94),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g87 ( 
.A(n_79),
.B(n_73),
.C(n_63),
.Y(n_87)
);

AND2x2_ASAP7_75t_L g97 ( 
.A(n_87),
.B(n_82),
.Y(n_97)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_83),
.Y(n_89)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_89),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_80),
.B(n_71),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_92),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_77),
.B(n_65),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g107 ( 
.A(n_93),
.B(n_50),
.Y(n_107)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_91),
.Y(n_95)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_95),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g121 ( 
.A1(n_96),
.A2(n_101),
.B1(n_103),
.B2(n_106),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_97),
.B(n_107),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_88),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_98),
.B(n_102),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_78),
.B1(n_75),
.B2(n_74),
.Y(n_101)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_88),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_91),
.A2(n_94),
.B1(n_89),
.B2(n_86),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_86),
.Y(n_104)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_104),
.Y(n_114)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_87),
.Y(n_105)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_105),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_84),
.A2(n_56),
.B1(n_51),
.B2(n_69),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g108 ( 
.A1(n_105),
.A2(n_54),
.B1(n_63),
.B2(n_67),
.Y(n_108)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_108),
.A2(n_117),
.B1(n_123),
.B2(n_7),
.Y(n_136)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_97),
.A2(n_54),
.B1(n_67),
.B2(n_52),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g135 ( 
.A1(n_109),
.A2(n_4),
.B1(n_6),
.B2(n_7),
.Y(n_135)
);

FAx1_ASAP7_75t_SL g111 ( 
.A(n_106),
.B(n_76),
.CI(n_68),
.CON(n_111),
.SN(n_111)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_111),
.B(n_112),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_103),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_62),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_113),
.B(n_116),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_100),
.B(n_48),
.Y(n_116)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_26),
.B1(n_32),
.B2(n_30),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_104),
.B(n_66),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_118),
.B(n_124),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_105),
.B(n_76),
.C(n_72),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_122),
.B(n_3),
.C(n_4),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_105),
.A2(n_64),
.B1(n_53),
.B2(n_61),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_99),
.B(n_2),
.Y(n_124)
);

XOR2xp5_ASAP7_75t_L g126 ( 
.A(n_110),
.B(n_19),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g145 ( 
.A(n_126),
.B(n_129),
.C(n_109),
.Y(n_145)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_120),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g146 ( 
.A(n_128),
.B(n_130),
.Y(n_146)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_115),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_119),
.A2(n_20),
.B1(n_42),
.B2(n_40),
.Y(n_131)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_131),
.A2(n_117),
.B1(n_111),
.B2(n_108),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_119),
.B(n_3),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_133),
.B(n_137),
.Y(n_139)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_114),
.Y(n_134)
);

INVx4_ASAP7_75t_L g141 ( 
.A(n_134),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g140 ( 
.A(n_135),
.B(n_136),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_122),
.B(n_8),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_SL g138 ( 
.A1(n_111),
.A2(n_9),
.B1(n_12),
.B2(n_13),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g144 ( 
.A(n_138),
.B(n_121),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g142 ( 
.A(n_127),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_144),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_143),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g150 ( 
.A(n_145),
.B(n_147),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_126),
.B(n_27),
.C(n_14),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g151 ( 
.A(n_146),
.B(n_132),
.Y(n_151)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_151),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_149),
.B(n_139),
.Y(n_152)
);

XNOR2xp5_ASAP7_75t_L g154 ( 
.A(n_152),
.B(n_129),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_154),
.B(n_150),
.C(n_153),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_155),
.B(n_131),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_156),
.B(n_135),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_157),
.Y(n_158)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_158),
.B(n_125),
.Y(n_159)
);

NOR3xp33_ASAP7_75t_L g160 ( 
.A(n_159),
.B(n_148),
.C(n_138),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_L g161 ( 
.A(n_160),
.B(n_144),
.C(n_140),
.Y(n_161)
);

AOI322xp5_ASAP7_75t_L g162 ( 
.A1(n_161),
.A2(n_143),
.A3(n_140),
.B1(n_16),
.B2(n_22),
.C1(n_23),
.C2(n_28),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_162),
.A2(n_141),
.B1(n_15),
.B2(n_29),
.Y(n_163)
);

XNOR2x2_ASAP7_75t_SL g164 ( 
.A(n_163),
.B(n_33),
.Y(n_164)
);


endmodule