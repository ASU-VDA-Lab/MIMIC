module fake_aes_6039_n_415 (n_53, n_45, n_20, n_2, n_38, n_44, n_54, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_3, n_18, n_32, n_0, n_41, n_1, n_35, n_55, n_12, n_9, n_17, n_14, n_10, n_15, n_56, n_42, n_24, n_19, n_21, n_6, n_4, n_51, n_29, n_43, n_7, n_40, n_27, n_39, n_415);
input n_53;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_54;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_3;
input n_18;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_12;
input n_9;
input n_17;
input n_14;
input n_10;
input n_15;
input n_56;
input n_42;
input n_24;
input n_19;
input n_21;
input n_6;
input n_4;
input n_51;
input n_29;
input n_43;
input n_7;
input n_40;
input n_27;
input n_39;
output n_415;
wire n_117;
wire n_361;
wire n_185;
wire n_57;
wire n_407;
wire n_284;
wire n_278;
wire n_60;
wire n_114;
wire n_94;
wire n_125;
wire n_161;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_229;
wire n_336;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_206;
wire n_288;
wire n_383;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_142;
wire n_232;
wire n_316;
wire n_211;
wire n_334;
wire n_389;
wire n_275;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_105;
wire n_227;
wire n_384;
wire n_231;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_228;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_150;
wire n_373;
wire n_301;
wire n_66;
wire n_222;
wire n_234;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_73;
wire n_119;
wire n_141;
wire n_97;
wire n_167;
wire n_171;
wire n_65;
wire n_196;
wire n_192;
wire n_312;
wire n_137;
wire n_277;
wire n_367;
wire n_250;
wire n_85;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_62;
wire n_255;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_241;
wire n_95;
wire n_238;
wire n_318;
wire n_293;
wire n_135;
wire n_393;
wire n_247;
wire n_381;
wire n_304;
wire n_399;
wire n_294;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_235;
wire n_243;
wire n_394;
wire n_331;
wire n_352;
wire n_268;
wire n_174;
wire n_248;
wire n_72;
wire n_299;
wire n_89;
wire n_338;
wire n_256;
wire n_67;
wire n_77;
wire n_404;
wire n_369;
wire n_172;
wire n_329;
wire n_251;
wire n_59;
wire n_218;
wire n_271;
wire n_302;
wire n_270;
wire n_362;
wire n_153;
wire n_61;
wire n_259;
wire n_308;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_224;
wire n_96;
wire n_219;
wire n_133;
wire n_149;
wire n_81;
wire n_69;
wire n_214;
wire n_204;
wire n_88;
wire n_107;
wire n_403;
wire n_254;
wire n_262;
wire n_239;
wire n_87;
wire n_379;
wire n_98;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_342;
wire n_370;
wire n_217;
wire n_139;
wire n_388;
wire n_193;
wire n_273;
wire n_390;
wire n_120;
wire n_70;
wire n_245;
wire n_90;
wire n_357;
wire n_260;
wire n_78;
wire n_201;
wire n_197;
wire n_317;
wire n_374;
wire n_111;
wire n_64;
wire n_265;
wire n_264;
wire n_200;
wire n_208;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_186;
wire n_364;
wire n_75;
wire n_376;
wire n_344;
wire n_136;
wire n_283;
wire n_76;
wire n_216;
wire n_147;
wire n_148;
wire n_212;
wire n_92;
wire n_396;
wire n_168;
wire n_398;
wire n_134;
wire n_233;
wire n_82;
wire n_106;
wire n_173;
wire n_327;
wire n_325;
wire n_349;
wire n_225;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_203;
wire n_102;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_121;
wire n_339;
wire n_240;
wire n_378;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_104;
wire n_74;
wire n_335;
wire n_272;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_156;
wire n_124;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_63;
wire n_71;
wire n_188;
wire n_377;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_58;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_371;
wire n_323;
wire n_347;
wire n_258;
wire n_253;
wire n_84;
wire n_266;
wire n_213;
wire n_182;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_176;
wire n_68;
wire n_123;
wire n_223;
wire n_372;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_332;
wire n_414;
wire n_350;
wire n_164;
wire n_175;
wire n_145;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx2_ASAP7_75t_L g57 ( .A(n_7), .Y(n_57) );
INVxp67_ASAP7_75t_SL g58 ( .A(n_1), .Y(n_58) );
CKINVDCx20_ASAP7_75t_R g59 ( .A(n_22), .Y(n_59) );
INVx1_ASAP7_75t_L g60 ( .A(n_50), .Y(n_60) );
INVx1_ASAP7_75t_L g61 ( .A(n_42), .Y(n_61) );
INVx1_ASAP7_75t_L g62 ( .A(n_20), .Y(n_62) );
INVxp33_ASAP7_75t_SL g63 ( .A(n_14), .Y(n_63) );
INVx1_ASAP7_75t_L g64 ( .A(n_33), .Y(n_64) );
INVx1_ASAP7_75t_L g65 ( .A(n_35), .Y(n_65) );
INVxp33_ASAP7_75t_SL g66 ( .A(n_15), .Y(n_66) );
INVx2_ASAP7_75t_L g67 ( .A(n_44), .Y(n_67) );
CKINVDCx14_ASAP7_75t_R g68 ( .A(n_37), .Y(n_68) );
INVxp67_ASAP7_75t_L g69 ( .A(n_6), .Y(n_69) );
CKINVDCx5p33_ASAP7_75t_R g70 ( .A(n_41), .Y(n_70) );
INVx1_ASAP7_75t_L g71 ( .A(n_29), .Y(n_71) );
INVx1_ASAP7_75t_L g72 ( .A(n_24), .Y(n_72) );
INVx2_ASAP7_75t_L g73 ( .A(n_30), .Y(n_73) );
HB1xp67_ASAP7_75t_L g74 ( .A(n_43), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_28), .Y(n_75) );
INVx2_ASAP7_75t_L g76 ( .A(n_19), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_49), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_5), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_55), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_10), .Y(n_80) );
CKINVDCx20_ASAP7_75t_R g81 ( .A(n_21), .Y(n_81) );
INVx2_ASAP7_75t_L g82 ( .A(n_14), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_23), .Y(n_83) );
INVx2_ASAP7_75t_L g84 ( .A(n_5), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_8), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_27), .Y(n_86) );
BUFx2_ASAP7_75t_L g87 ( .A(n_11), .Y(n_87) );
BUFx6f_ASAP7_75t_L g88 ( .A(n_13), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_26), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_11), .Y(n_90) );
INVxp33_ASAP7_75t_SL g91 ( .A(n_40), .Y(n_91) );
INVxp67_ASAP7_75t_SL g92 ( .A(n_1), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_52), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_9), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_57), .Y(n_95) );
INVx1_ASAP7_75t_L g96 ( .A(n_57), .Y(n_96) );
NOR2xp33_ASAP7_75t_R g97 ( .A(n_68), .B(n_34), .Y(n_97) );
BUFx2_ASAP7_75t_L g98 ( .A(n_87), .Y(n_98) );
NAND2xp5_ASAP7_75t_L g99 ( .A(n_87), .B(n_0), .Y(n_99) );
CKINVDCx5p33_ASAP7_75t_R g100 ( .A(n_59), .Y(n_100) );
CKINVDCx5p33_ASAP7_75t_R g101 ( .A(n_81), .Y(n_101) );
BUFx3_ASAP7_75t_L g102 ( .A(n_67), .Y(n_102) );
HB1xp67_ASAP7_75t_L g103 ( .A(n_57), .Y(n_103) );
BUFx6f_ASAP7_75t_L g104 ( .A(n_67), .Y(n_104) );
CKINVDCx5p33_ASAP7_75t_R g105 ( .A(n_80), .Y(n_105) );
NAND2xp33_ASAP7_75t_R g106 ( .A(n_91), .B(n_0), .Y(n_106) );
INVx2_ASAP7_75t_L g107 ( .A(n_67), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_90), .Y(n_108) );
AND2x4_ASAP7_75t_L g109 ( .A(n_76), .B(n_2), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_76), .Y(n_110) );
CKINVDCx5p33_ASAP7_75t_R g111 ( .A(n_63), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_76), .Y(n_112) );
BUFx6f_ASAP7_75t_L g113 ( .A(n_73), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_73), .Y(n_114) );
INVx1_ASAP7_75t_L g115 ( .A(n_82), .Y(n_115) );
CKINVDCx20_ASAP7_75t_R g116 ( .A(n_74), .Y(n_116) );
AND2x4_ASAP7_75t_L g117 ( .A(n_109), .B(n_82), .Y(n_117) );
CKINVDCx5p33_ASAP7_75t_R g118 ( .A(n_100), .Y(n_118) );
NAND2xp5_ASAP7_75t_L g119 ( .A(n_103), .B(n_60), .Y(n_119) );
BUFx6f_ASAP7_75t_L g120 ( .A(n_104), .Y(n_120) );
AO22x2_ASAP7_75t_L g121 ( .A1(n_109), .A2(n_75), .B1(n_93), .B2(n_60), .Y(n_121) );
BUFx3_ASAP7_75t_L g122 ( .A(n_109), .Y(n_122) );
INVx4_ASAP7_75t_L g123 ( .A(n_109), .Y(n_123) );
NAND2x1p5_ASAP7_75t_L g124 ( .A(n_102), .B(n_61), .Y(n_124) );
INVx4_ASAP7_75t_L g125 ( .A(n_102), .Y(n_125) );
AND2x6_ASAP7_75t_L g126 ( .A(n_102), .B(n_61), .Y(n_126) );
AND2x2_ASAP7_75t_L g127 ( .A(n_98), .B(n_82), .Y(n_127) );
INVx4_ASAP7_75t_L g128 ( .A(n_104), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_107), .Y(n_129) );
BUFx6f_ASAP7_75t_L g130 ( .A(n_104), .Y(n_130) );
AND2x2_ASAP7_75t_L g131 ( .A(n_98), .B(n_84), .Y(n_131) );
INVx1_ASAP7_75t_L g132 ( .A(n_107), .Y(n_132) );
NOR2xp33_ASAP7_75t_L g133 ( .A(n_103), .B(n_62), .Y(n_133) );
BUFx3_ASAP7_75t_L g134 ( .A(n_107), .Y(n_134) );
BUFx3_ASAP7_75t_L g135 ( .A(n_114), .Y(n_135) );
INVx3_ASAP7_75t_L g136 ( .A(n_114), .Y(n_136) );
AND2x6_ASAP7_75t_L g137 ( .A(n_99), .B(n_62), .Y(n_137) );
AND2x6_ASAP7_75t_L g138 ( .A(n_99), .B(n_64), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_114), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_104), .Y(n_140) );
INVxp67_ASAP7_75t_SL g141 ( .A(n_95), .Y(n_141) );
INVx1_ASAP7_75t_L g142 ( .A(n_123), .Y(n_142) );
BUFx6f_ASAP7_75t_L g143 ( .A(n_134), .Y(n_143) );
INVx2_ASAP7_75t_L g144 ( .A(n_134), .Y(n_144) );
OR2x6_ASAP7_75t_L g145 ( .A(n_121), .B(n_78), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g146 ( .A(n_119), .B(n_105), .Y(n_146) );
NAND2x1p5_ASAP7_75t_L g147 ( .A(n_123), .B(n_64), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_134), .Y(n_148) );
INVxp67_ASAP7_75t_L g149 ( .A(n_127), .Y(n_149) );
AO22x1_ASAP7_75t_L g150 ( .A1(n_137), .A2(n_66), .B1(n_92), .B2(n_58), .Y(n_150) );
BUFx2_ASAP7_75t_L g151 ( .A(n_121), .Y(n_151) );
NAND2xp5_ASAP7_75t_L g152 ( .A(n_119), .B(n_108), .Y(n_152) );
BUFx2_ASAP7_75t_L g153 ( .A(n_121), .Y(n_153) );
CKINVDCx5p33_ASAP7_75t_R g154 ( .A(n_118), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_135), .Y(n_155) );
INVx2_ASAP7_75t_SL g156 ( .A(n_121), .Y(n_156) );
AOI22xp33_ASAP7_75t_L g157 ( .A1(n_121), .A2(n_85), .B1(n_94), .B2(n_78), .Y(n_157) );
INVx1_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
INVx1_ASAP7_75t_L g159 ( .A(n_141), .Y(n_159) );
NOR3xp33_ASAP7_75t_SL g160 ( .A(n_133), .B(n_101), .C(n_111), .Y(n_160) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_133), .B(n_97), .Y(n_161) );
BUFx6f_ASAP7_75t_L g162 ( .A(n_135), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_117), .Y(n_163) );
INVxp67_ASAP7_75t_L g164 ( .A(n_127), .Y(n_164) );
INVx1_ASAP7_75t_L g165 ( .A(n_117), .Y(n_165) );
INVx1_ASAP7_75t_L g166 ( .A(n_117), .Y(n_166) );
BUFx6f_ASAP7_75t_L g167 ( .A(n_135), .Y(n_167) );
OR2x2_ASAP7_75t_L g168 ( .A(n_127), .B(n_69), .Y(n_168) );
NAND2xp5_ASAP7_75t_L g169 ( .A(n_123), .B(n_131), .Y(n_169) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_121), .A2(n_116), .B1(n_106), .B2(n_85), .Y(n_170) );
INVx1_ASAP7_75t_SL g171 ( .A(n_131), .Y(n_171) );
NAND2xp5_ASAP7_75t_L g172 ( .A(n_123), .B(n_97), .Y(n_172) );
NAND2xp5_ASAP7_75t_L g173 ( .A(n_123), .B(n_70), .Y(n_173) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_120), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_146), .B(n_137), .Y(n_175) );
BUFx2_ASAP7_75t_L g176 ( .A(n_145), .Y(n_176) );
AOI22xp5_ASAP7_75t_L g177 ( .A1(n_145), .A2(n_138), .B1(n_137), .B2(n_131), .Y(n_177) );
OAI21xp33_ASAP7_75t_L g178 ( .A1(n_152), .A2(n_122), .B(n_124), .Y(n_178) );
CKINVDCx5p33_ASAP7_75t_R g179 ( .A(n_154), .Y(n_179) );
OR2x6_ASAP7_75t_L g180 ( .A(n_145), .B(n_151), .Y(n_180) );
INVx4_ASAP7_75t_L g181 ( .A(n_145), .Y(n_181) );
NAND2xp5_ASAP7_75t_L g182 ( .A(n_169), .B(n_137), .Y(n_182) );
BUFx2_ASAP7_75t_L g183 ( .A(n_151), .Y(n_183) );
INVx1_ASAP7_75t_L g184 ( .A(n_158), .Y(n_184) );
INVx1_ASAP7_75t_L g185 ( .A(n_159), .Y(n_185) );
O2A1O1Ixp33_ASAP7_75t_L g186 ( .A1(n_149), .A2(n_122), .B(n_124), .C(n_117), .Y(n_186) );
NAND2x1p5_ASAP7_75t_L g187 ( .A(n_153), .B(n_125), .Y(n_187) );
INVx1_ASAP7_75t_L g188 ( .A(n_142), .Y(n_188) );
BUFx2_ASAP7_75t_L g189 ( .A(n_153), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_171), .B(n_124), .Y(n_190) );
CKINVDCx20_ASAP7_75t_R g191 ( .A(n_154), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g192 ( .A1(n_172), .A2(n_122), .B(n_117), .Y(n_192) );
OR2x2_ASAP7_75t_SL g193 ( .A(n_168), .B(n_106), .Y(n_193) );
OR2x6_ASAP7_75t_L g194 ( .A(n_156), .B(n_124), .Y(n_194) );
INVx1_ASAP7_75t_L g195 ( .A(n_142), .Y(n_195) );
AOI22xp33_ASAP7_75t_L g196 ( .A1(n_156), .A2(n_137), .B1(n_138), .B2(n_126), .Y(n_196) );
INVx3_ASAP7_75t_L g197 ( .A(n_143), .Y(n_197) );
OR2x2_ASAP7_75t_L g198 ( .A(n_168), .B(n_129), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_164), .B(n_137), .Y(n_199) );
INVx1_ASAP7_75t_SL g200 ( .A(n_147), .Y(n_200) );
BUFx2_ASAP7_75t_L g201 ( .A(n_147), .Y(n_201) );
NAND2xp5_ASAP7_75t_L g202 ( .A(n_161), .B(n_137), .Y(n_202) );
BUFx6f_ASAP7_75t_L g203 ( .A(n_143), .Y(n_203) );
AND2x4_ASAP7_75t_L g204 ( .A(n_163), .B(n_137), .Y(n_204) );
AOI22xp5_ASAP7_75t_L g205 ( .A1(n_170), .A2(n_138), .B1(n_137), .B2(n_125), .Y(n_205) );
AOI22xp5_ASAP7_75t_L g206 ( .A1(n_157), .A2(n_138), .B1(n_125), .B2(n_126), .Y(n_206) );
AOI22xp33_ASAP7_75t_SL g207 ( .A1(n_180), .A2(n_181), .B1(n_176), .B2(n_183), .Y(n_207) );
OAI21x1_ASAP7_75t_L g208 ( .A1(n_192), .A2(n_147), .B(n_73), .Y(n_208) );
AND2x2_ASAP7_75t_L g209 ( .A(n_180), .B(n_165), .Y(n_209) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_184), .B(n_166), .Y(n_210) );
INVx2_ASAP7_75t_L g211 ( .A(n_203), .Y(n_211) );
INVx4_ASAP7_75t_L g212 ( .A(n_180), .Y(n_212) );
AOI22xp33_ASAP7_75t_L g213 ( .A1(n_190), .A2(n_138), .B1(n_126), .B2(n_125), .Y(n_213) );
INVx2_ASAP7_75t_L g214 ( .A(n_203), .Y(n_214) );
AOI21xp5_ASAP7_75t_L g215 ( .A1(n_202), .A2(n_173), .B(n_144), .Y(n_215) );
BUFx2_ASAP7_75t_L g216 ( .A(n_181), .Y(n_216) );
OAI221xp5_ASAP7_75t_L g217 ( .A1(n_198), .A2(n_160), .B1(n_94), .B2(n_139), .C(n_132), .Y(n_217) );
AND2x2_ASAP7_75t_L g218 ( .A(n_190), .B(n_144), .Y(n_218) );
BUFx6f_ASAP7_75t_L g219 ( .A(n_203), .Y(n_219) );
BUFx2_ASAP7_75t_L g220 ( .A(n_181), .Y(n_220) );
NAND2xp5_ASAP7_75t_L g221 ( .A(n_185), .B(n_138), .Y(n_221) );
INVx2_ASAP7_75t_L g222 ( .A(n_203), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_201), .B(n_143), .Y(n_223) );
NAND2xp5_ASAP7_75t_L g224 ( .A(n_188), .B(n_138), .Y(n_224) );
AOI22xp33_ASAP7_75t_L g225 ( .A1(n_175), .A2(n_138), .B1(n_126), .B2(n_125), .Y(n_225) );
INVx1_ASAP7_75t_L g226 ( .A(n_195), .Y(n_226) );
NAND2xp33_ASAP7_75t_SL g227 ( .A(n_189), .B(n_143), .Y(n_227) );
AND2x2_ASAP7_75t_L g228 ( .A(n_194), .B(n_148), .Y(n_228) );
INVx1_ASAP7_75t_L g229 ( .A(n_182), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g230 ( .A(n_177), .B(n_138), .Y(n_230) );
AND2x2_ASAP7_75t_L g231 ( .A(n_194), .B(n_148), .Y(n_231) );
AND2x2_ASAP7_75t_L g232 ( .A(n_194), .B(n_155), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_199), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_212), .B(n_193), .Y(n_234) );
OAI22xp33_ASAP7_75t_L g235 ( .A1(n_217), .A2(n_191), .B1(n_179), .B2(n_200), .Y(n_235) );
BUFx6f_ASAP7_75t_L g236 ( .A(n_219), .Y(n_236) );
OAI22xp5_ASAP7_75t_L g237 ( .A1(n_212), .A2(n_205), .B1(n_187), .B2(n_186), .Y(n_237) );
INVx1_ASAP7_75t_L g238 ( .A(n_226), .Y(n_238) );
AND2x2_ASAP7_75t_L g239 ( .A(n_218), .B(n_187), .Y(n_239) );
BUFx4f_ASAP7_75t_SL g240 ( .A(n_212), .Y(n_240) );
OAI22xp5_ASAP7_75t_L g241 ( .A1(n_212), .A2(n_196), .B1(n_178), .B2(n_206), .Y(n_241) );
AOI22xp33_ASAP7_75t_L g242 ( .A1(n_217), .A2(n_209), .B1(n_212), .B2(n_229), .Y(n_242) );
INVx2_ASAP7_75t_L g243 ( .A(n_219), .Y(n_243) );
OR2x2_ASAP7_75t_L g244 ( .A(n_226), .B(n_218), .Y(n_244) );
A2O1A1Ixp33_ASAP7_75t_L g245 ( .A1(n_229), .A2(n_196), .B(n_204), .C(n_132), .Y(n_245) );
AND2x2_ASAP7_75t_L g246 ( .A(n_218), .B(n_204), .Y(n_246) );
OAI33xp33_ASAP7_75t_L g247 ( .A1(n_221), .A2(n_115), .A3(n_112), .B1(n_110), .B2(n_96), .B3(n_95), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_233), .B(n_204), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_210), .Y(n_249) );
INVx2_ASAP7_75t_SL g250 ( .A(n_216), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_210), .Y(n_251) );
OAI221xp5_ASAP7_75t_L g252 ( .A1(n_207), .A2(n_96), .B1(n_110), .B2(n_115), .C(n_112), .Y(n_252) );
AOI22xp33_ASAP7_75t_L g253 ( .A1(n_209), .A2(n_191), .B1(n_179), .B2(n_126), .Y(n_253) );
AO21x2_ASAP7_75t_L g254 ( .A1(n_215), .A2(n_65), .B(n_71), .Y(n_254) );
INVx2_ASAP7_75t_L g255 ( .A(n_219), .Y(n_255) );
HB1xp67_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
AOI221xp5_ASAP7_75t_L g257 ( .A1(n_235), .A2(n_150), .B1(n_84), .B2(n_233), .C(n_88), .Y(n_257) );
AND2x2_ASAP7_75t_L g258 ( .A(n_249), .B(n_223), .Y(n_258) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_242), .A2(n_209), .B1(n_230), .B2(n_207), .Y(n_259) );
OAI21xp5_ASAP7_75t_L g260 ( .A1(n_249), .A2(n_215), .B(n_208), .Y(n_260) );
AND2x2_ASAP7_75t_L g261 ( .A(n_251), .B(n_223), .Y(n_261) );
NOR2x1_ASAP7_75t_SL g262 ( .A(n_237), .B(n_219), .Y(n_262) );
AND2x4_ASAP7_75t_L g263 ( .A(n_243), .B(n_211), .Y(n_263) );
AO21x2_ASAP7_75t_L g264 ( .A1(n_254), .A2(n_208), .B(n_230), .Y(n_264) );
CKINVDCx5p33_ASAP7_75t_R g265 ( .A(n_240), .Y(n_265) );
INVxp67_ASAP7_75t_L g266 ( .A(n_244), .Y(n_266) );
OR2x6_ASAP7_75t_L g267 ( .A(n_237), .B(n_216), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g268 ( .A(n_238), .B(n_228), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g269 ( .A(n_239), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_243), .Y(n_270) );
AND2x2_ASAP7_75t_L g271 ( .A(n_244), .B(n_223), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_243), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_254), .Y(n_273) );
INVxp67_ASAP7_75t_L g274 ( .A(n_239), .Y(n_274) );
AOI22xp33_ASAP7_75t_L g275 ( .A1(n_252), .A2(n_221), .B1(n_220), .B2(n_227), .Y(n_275) );
OAI221xp5_ASAP7_75t_SL g276 ( .A1(n_252), .A2(n_213), .B1(n_225), .B2(n_224), .C(n_65), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_271), .B(n_254), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_273), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_273), .Y(n_279) );
AOI22xp33_ASAP7_75t_SL g280 ( .A1(n_269), .A2(n_234), .B1(n_250), .B2(n_241), .Y(n_280) );
AND2x2_ASAP7_75t_L g281 ( .A(n_271), .B(n_256), .Y(n_281) );
OAI21xp5_ASAP7_75t_SL g282 ( .A1(n_257), .A2(n_253), .B(n_241), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_266), .B(n_250), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_270), .Y(n_284) );
OAI33xp33_ASAP7_75t_L g285 ( .A1(n_266), .A2(n_71), .A3(n_72), .B1(n_75), .B2(n_77), .B3(n_79), .Y(n_285) );
BUFx2_ASAP7_75t_L g286 ( .A(n_267), .Y(n_286) );
INVx2_ASAP7_75t_L g287 ( .A(n_270), .Y(n_287) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_268), .B(n_255), .Y(n_288) );
OAI221xp5_ASAP7_75t_SL g289 ( .A1(n_257), .A2(n_248), .B1(n_246), .B2(n_213), .C(n_245), .Y(n_289) );
OAI33xp33_ASAP7_75t_L g290 ( .A1(n_268), .A2(n_72), .A3(n_77), .B1(n_79), .B2(n_83), .B3(n_86), .Y(n_290) );
AOI221xp5_ASAP7_75t_L g291 ( .A1(n_259), .A2(n_247), .B1(n_88), .B2(n_248), .C(n_246), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_258), .B(n_261), .Y(n_292) );
INVx2_ASAP7_75t_SL g293 ( .A(n_267), .Y(n_293) );
OA21x2_ASAP7_75t_L g294 ( .A1(n_260), .A2(n_255), .B(n_208), .Y(n_294) );
INVx2_ASAP7_75t_SL g295 ( .A(n_267), .Y(n_295) );
AND2x2_ASAP7_75t_L g296 ( .A(n_258), .B(n_236), .Y(n_296) );
AND2x2_ASAP7_75t_L g297 ( .A(n_261), .B(n_236), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_261), .B(n_236), .Y(n_298) );
AND2x2_ASAP7_75t_L g299 ( .A(n_270), .B(n_236), .Y(n_299) );
AND2x2_ASAP7_75t_L g300 ( .A(n_272), .B(n_236), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_272), .Y(n_301) );
AND2x2_ASAP7_75t_L g302 ( .A(n_281), .B(n_274), .Y(n_302) );
HB1xp67_ASAP7_75t_L g303 ( .A(n_284), .Y(n_303) );
OR2x2_ASAP7_75t_L g304 ( .A(n_292), .B(n_267), .Y(n_304) );
NAND4xp25_ASAP7_75t_L g305 ( .A(n_280), .B(n_275), .C(n_83), .D(n_86), .Y(n_305) );
AND2x2_ASAP7_75t_L g306 ( .A(n_281), .B(n_263), .Y(n_306) );
NAND5xp2_ASAP7_75t_SL g307 ( .A(n_282), .B(n_265), .C(n_275), .D(n_4), .E(n_6), .Y(n_307) );
AOI22xp33_ASAP7_75t_L g308 ( .A1(n_291), .A2(n_247), .B1(n_264), .B2(n_260), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g309 ( .A(n_277), .B(n_264), .Y(n_309) );
INVx1_ASAP7_75t_L g310 ( .A(n_283), .Y(n_310) );
AND2x2_ASAP7_75t_L g311 ( .A(n_277), .B(n_263), .Y(n_311) );
NOR2xp67_ASAP7_75t_SL g312 ( .A(n_286), .B(n_236), .Y(n_312) );
AND2x4_ASAP7_75t_L g313 ( .A(n_293), .B(n_262), .Y(n_313) );
NAND2xp5_ASAP7_75t_L g314 ( .A(n_283), .B(n_263), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_288), .B(n_278), .Y(n_315) );
NAND2x1p5_ASAP7_75t_L g316 ( .A(n_293), .B(n_219), .Y(n_316) );
INVx1_ASAP7_75t_SL g317 ( .A(n_296), .Y(n_317) );
OR2x2_ASAP7_75t_L g318 ( .A(n_298), .B(n_276), .Y(n_318) );
AOI22xp33_ASAP7_75t_SL g319 ( .A1(n_293), .A2(n_262), .B1(n_276), .B2(n_223), .Y(n_319) );
NOR3xp33_ASAP7_75t_L g320 ( .A(n_285), .B(n_89), .C(n_93), .Y(n_320) );
OR2x2_ASAP7_75t_L g321 ( .A(n_298), .B(n_301), .Y(n_321) );
AND2x2_ASAP7_75t_L g322 ( .A(n_296), .B(n_297), .Y(n_322) );
NOR2xp33_ASAP7_75t_L g323 ( .A(n_285), .B(n_2), .Y(n_323) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_279), .B(n_3), .Y(n_324) );
INVx2_ASAP7_75t_L g325 ( .A(n_287), .Y(n_325) );
AND2x4_ASAP7_75t_L g326 ( .A(n_295), .B(n_104), .Y(n_326) );
NOR2xp33_ASAP7_75t_L g327 ( .A(n_310), .B(n_290), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_315), .Y(n_328) );
INVx1_ASAP7_75t_SL g329 ( .A(n_317), .Y(n_329) );
O2A1O1Ixp33_ASAP7_75t_L g330 ( .A1(n_307), .A2(n_289), .B(n_290), .C(n_291), .Y(n_330) );
AND2x2_ASAP7_75t_L g331 ( .A(n_322), .B(n_295), .Y(n_331) );
AND2x2_ASAP7_75t_L g332 ( .A(n_311), .B(n_299), .Y(n_332) );
NAND2xp5_ASAP7_75t_SL g333 ( .A(n_319), .B(n_300), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_321), .Y(n_334) );
NOR2xp33_ASAP7_75t_L g335 ( .A(n_305), .B(n_3), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_306), .B(n_300), .Y(n_336) );
INVx1_ASAP7_75t_L g337 ( .A(n_314), .Y(n_337) );
INVx3_ASAP7_75t_L g338 ( .A(n_326), .Y(n_338) );
INVx1_ASAP7_75t_L g339 ( .A(n_324), .Y(n_339) );
OAI21xp33_ASAP7_75t_SL g340 ( .A1(n_304), .A2(n_232), .B(n_231), .Y(n_340) );
INVx1_ASAP7_75t_SL g341 ( .A(n_302), .Y(n_341) );
OAI22xp5_ASAP7_75t_L g342 ( .A1(n_319), .A2(n_294), .B1(n_222), .B2(n_214), .Y(n_342) );
NOR2xp67_ASAP7_75t_L g343 ( .A(n_303), .B(n_4), .Y(n_343) );
AOI22xp33_ASAP7_75t_L g344 ( .A1(n_323), .A2(n_294), .B1(n_232), .B2(n_231), .Y(n_344) );
NAND2xp5_ASAP7_75t_L g345 ( .A(n_309), .B(n_294), .Y(n_345) );
NOR2x1_ASAP7_75t_SL g346 ( .A(n_318), .B(n_219), .Y(n_346) );
AOI211xp5_ASAP7_75t_L g347 ( .A1(n_320), .A2(n_113), .B(n_140), .C(n_136), .Y(n_347) );
AOI32xp33_ASAP7_75t_L g348 ( .A1(n_320), .A2(n_12), .A3(n_13), .B1(n_15), .B2(n_16), .Y(n_348) );
INVx1_ASAP7_75t_L g349 ( .A(n_325), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_325), .Y(n_350) );
OAI32xp33_ASAP7_75t_L g351 ( .A1(n_316), .A2(n_17), .A3(n_18), .B1(n_19), .B2(n_136), .Y(n_351) );
NAND2xp5_ASAP7_75t_L g352 ( .A(n_308), .B(n_17), .Y(n_352) );
NAND2xp5_ASAP7_75t_SL g353 ( .A(n_313), .B(n_219), .Y(n_353) );
INVxp67_ASAP7_75t_L g354 ( .A(n_312), .Y(n_354) );
INVxp67_ASAP7_75t_L g355 ( .A(n_329), .Y(n_355) );
INVx1_ASAP7_75t_L g356 ( .A(n_334), .Y(n_356) );
XNOR2xp5_ASAP7_75t_L g357 ( .A(n_341), .B(n_18), .Y(n_357) );
INVxp67_ASAP7_75t_L g358 ( .A(n_328), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_332), .B(n_113), .Y(n_359) );
NAND2xp33_ASAP7_75t_SL g360 ( .A(n_333), .B(n_222), .Y(n_360) );
INVxp67_ASAP7_75t_L g361 ( .A(n_343), .Y(n_361) );
XNOR2xp5_ASAP7_75t_L g362 ( .A(n_331), .B(n_25), .Y(n_362) );
INVxp67_ASAP7_75t_L g363 ( .A(n_339), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_337), .Y(n_364) );
NOR2xp33_ASAP7_75t_L g365 ( .A(n_327), .B(n_31), .Y(n_365) );
AND2x2_ASAP7_75t_L g366 ( .A(n_336), .B(n_32), .Y(n_366) );
NAND2xp33_ASAP7_75t_SL g367 ( .A(n_338), .B(n_197), .Y(n_367) );
NAND3xp33_ASAP7_75t_L g368 ( .A(n_327), .B(n_120), .C(n_130), .Y(n_368) );
INVx3_ASAP7_75t_L g369 ( .A(n_338), .Y(n_369) );
A2O1A1Ixp33_ASAP7_75t_L g370 ( .A1(n_340), .A2(n_197), .B(n_38), .C(n_39), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_353), .B(n_36), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_349), .Y(n_372) );
INVx1_ASAP7_75t_L g373 ( .A(n_350), .Y(n_373) );
AND2x2_ASAP7_75t_L g374 ( .A(n_345), .B(n_130), .Y(n_374) );
OAI211xp5_ASAP7_75t_L g375 ( .A1(n_361), .A2(n_348), .B(n_330), .C(n_344), .Y(n_375) );
XNOR2xp5_ASAP7_75t_L g376 ( .A(n_357), .B(n_362), .Y(n_376) );
XNOR2x1_ASAP7_75t_L g377 ( .A(n_366), .B(n_342), .Y(n_377) );
OAI211xp5_ASAP7_75t_SL g378 ( .A1(n_363), .A2(n_344), .B(n_352), .C(n_335), .Y(n_378) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_358), .B(n_359), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_360), .A2(n_347), .B(n_354), .C(n_351), .Y(n_380) );
INVxp67_ASAP7_75t_L g381 ( .A(n_355), .Y(n_381) );
INVx1_ASAP7_75t_L g382 ( .A(n_364), .Y(n_382) );
NAND2xp5_ASAP7_75t_L g383 ( .A(n_372), .B(n_346), .Y(n_383) );
OAI21xp5_ASAP7_75t_L g384 ( .A1(n_370), .A2(n_128), .B(n_155), .Y(n_384) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_373), .B(n_130), .Y(n_385) );
AOI21xp5_ASAP7_75t_SL g386 ( .A1(n_370), .A2(n_45), .B(n_46), .Y(n_386) );
OAI22xp33_ASAP7_75t_SL g387 ( .A1(n_369), .A2(n_128), .B1(n_48), .B2(n_51), .Y(n_387) );
OAI322xp33_ASAP7_75t_L g388 ( .A1(n_356), .A2(n_120), .A3(n_128), .B1(n_167), .B2(n_162), .C1(n_143), .C2(n_56), .Y(n_388) );
NAND4xp75_ASAP7_75t_L g389 ( .A(n_365), .B(n_47), .C(n_53), .D(n_54), .Y(n_389) );
INVx2_ASAP7_75t_SL g390 ( .A(n_369), .Y(n_390) );
NOR2xp33_ASAP7_75t_R g391 ( .A(n_376), .B(n_367), .Y(n_391) );
NOR2x1_ASAP7_75t_L g392 ( .A(n_386), .B(n_368), .Y(n_392) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_382), .B(n_374), .Y(n_393) );
BUFx2_ASAP7_75t_L g394 ( .A(n_390), .Y(n_394) );
NOR2xp33_ASAP7_75t_R g395 ( .A(n_381), .B(n_371), .Y(n_395) );
BUFx2_ASAP7_75t_L g396 ( .A(n_383), .Y(n_396) );
NOR2x1_ASAP7_75t_L g397 ( .A(n_380), .B(n_374), .Y(n_397) );
OAI22xp33_ASAP7_75t_L g398 ( .A1(n_383), .A2(n_174), .B1(n_384), .B2(n_377), .Y(n_398) );
AOI221xp5_ASAP7_75t_L g399 ( .A1(n_388), .A2(n_375), .B1(n_378), .B2(n_358), .C(n_363), .Y(n_399) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_389), .A2(n_377), .B1(n_381), .B2(n_355), .Y(n_400) );
HB1xp67_ASAP7_75t_L g401 ( .A(n_385), .Y(n_401) );
AOI221xp5_ASAP7_75t_SL g402 ( .A1(n_387), .A2(n_381), .B1(n_361), .B2(n_355), .C(n_357), .Y(n_402) );
INVx1_ASAP7_75t_SL g403 ( .A(n_379), .Y(n_403) );
AOI22xp33_ASAP7_75t_R g404 ( .A1(n_391), .A2(n_395), .B1(n_401), .B2(n_402), .Y(n_404) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_399), .B(n_397), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_393), .Y(n_406) );
INVx1_ASAP7_75t_SL g407 ( .A(n_396), .Y(n_407) );
OAI222xp33_ASAP7_75t_L g408 ( .A1(n_404), .A2(n_400), .B1(n_398), .B2(n_394), .C1(n_403), .C2(n_392), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_406), .Y(n_409) );
INVx1_ASAP7_75t_L g410 ( .A(n_407), .Y(n_410) );
BUFx2_ASAP7_75t_L g411 ( .A(n_410), .Y(n_411) );
INVx1_ASAP7_75t_L g412 ( .A(n_409), .Y(n_412) );
INVx1_ASAP7_75t_L g413 ( .A(n_411), .Y(n_413) );
AOI22xp5_ASAP7_75t_L g414 ( .A1(n_413), .A2(n_405), .B1(n_411), .B2(n_409), .Y(n_414) );
AOI21xp5_ASAP7_75t_L g415 ( .A1(n_414), .A2(n_408), .B(n_412), .Y(n_415) );
endmodule