module fake_jpeg_21958_n_106 (n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_106);

input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_106;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_14;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_2),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_4),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_6),
.Y(n_18)
);

INVx4_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

BUFx10_ASAP7_75t_L g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_2),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_7),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx5_ASAP7_75t_SL g39 ( 
.A(n_23),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_12),
.B(n_0),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_24),
.B(n_29),
.Y(n_36)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_15),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_25),
.B(n_26),
.Y(n_32)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_17),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_17),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_27),
.Y(n_33)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_28),
.B(n_30),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g29 ( 
.A(n_12),
.B(n_0),
.Y(n_29)
);

INVx6_ASAP7_75t_L g30 ( 
.A(n_15),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g31 ( 
.A1(n_25),
.A2(n_19),
.B1(n_21),
.B2(n_16),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_31),
.B(n_30),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_29),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_35),
.B(n_38),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_27),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g48 ( 
.A(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_28),
.B(n_22),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_SL g40 ( 
.A(n_35),
.B(n_16),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_40),
.B(n_43),
.Y(n_63)
);

INVx11_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_41),
.B(n_47),
.Y(n_53)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_36),
.B(n_21),
.C(n_26),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_36),
.B(n_22),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_44),
.B(n_45),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_38),
.B(n_18),
.Y(n_45)
);

A2O1A1Ixp33_ASAP7_75t_L g46 ( 
.A1(n_32),
.A2(n_20),
.B(n_13),
.C(n_27),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g54 ( 
.A1(n_46),
.A2(n_49),
.B(n_34),
.Y(n_54)
);

INVx13_ASAP7_75t_L g47 ( 
.A(n_39),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_50),
.Y(n_62)
);

AND2x6_ASAP7_75t_L g51 ( 
.A(n_39),
.B(n_1),
.Y(n_51)
);

BUFx2_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_39),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g57 ( 
.A(n_52),
.B(n_34),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g68 ( 
.A1(n_54),
.A2(n_42),
.B(n_46),
.Y(n_68)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_43),
.A2(n_25),
.B1(n_30),
.B2(n_32),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_56),
.B(n_61),
.Y(n_71)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_50),
.Y(n_58)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_58),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_47),
.B(n_23),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g69 ( 
.A(n_59),
.B(n_60),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_47),
.B(n_52),
.Y(n_60)
);

AOI22xp5_ASAP7_75t_L g61 ( 
.A1(n_44),
.A2(n_26),
.B1(n_23),
.B2(n_21),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_55),
.B(n_40),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_65),
.B(n_67),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_55),
.B(n_42),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g77 ( 
.A1(n_68),
.A2(n_56),
.B1(n_61),
.B2(n_54),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_63),
.B(n_45),
.Y(n_70)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_70),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_58),
.B(n_41),
.Y(n_72)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_72),
.Y(n_78)
);

AND2x2_ASAP7_75t_L g73 ( 
.A(n_63),
.B(n_51),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_73),
.B(n_64),
.C(n_53),
.Y(n_80)
);

INVxp67_ASAP7_75t_SL g75 ( 
.A(n_69),
.Y(n_75)
);

INVxp33_ASAP7_75t_SL g88 ( 
.A(n_75),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_77),
.A2(n_71),
.B1(n_68),
.B2(n_73),
.Y(n_84)
);

XNOR2xp5_ASAP7_75t_L g85 ( 
.A(n_80),
.B(n_64),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_66),
.B(n_62),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_81),
.B(n_82),
.Y(n_86)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_70),
.Y(n_82)
);

AO221x1_ASAP7_75t_L g83 ( 
.A1(n_74),
.A2(n_62),
.B1(n_50),
.B2(n_48),
.C(n_33),
.Y(n_83)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_83),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g92 ( 
.A1(n_84),
.A2(n_89),
.B(n_48),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_85),
.B(n_20),
.C(n_11),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_80),
.A2(n_14),
.B1(n_13),
.B2(n_33),
.Y(n_89)
);

AOI322xp5_ASAP7_75t_L g90 ( 
.A1(n_85),
.A2(n_82),
.A3(n_79),
.B1(n_76),
.B2(n_78),
.C1(n_27),
.C2(n_14),
.Y(n_90)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_90),
.B(n_92),
.Y(n_95)
);

OAI321xp33_ASAP7_75t_L g91 ( 
.A1(n_88),
.A2(n_79),
.A3(n_76),
.B1(n_11),
.B2(n_20),
.C(n_33),
.Y(n_91)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_91),
.Y(n_98)
);

INVx1_ASAP7_75t_SL g93 ( 
.A(n_88),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_93),
.B(n_94),
.Y(n_97)
);

A2O1A1Ixp33_ASAP7_75t_L g96 ( 
.A1(n_92),
.A2(n_86),
.B(n_87),
.C(n_20),
.Y(n_96)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_96),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_97),
.B(n_98),
.C(n_95),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g102 ( 
.A(n_100),
.B(n_10),
.Y(n_102)
);

AOI211xp5_ASAP7_75t_L g101 ( 
.A1(n_96),
.A2(n_6),
.B(n_8),
.C(n_9),
.Y(n_101)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_101),
.A2(n_1),
.A3(n_3),
.B1(n_5),
.B2(n_8),
.C1(n_10),
.C2(n_99),
.Y(n_103)
);

MAJx2_ASAP7_75t_L g104 ( 
.A(n_102),
.B(n_103),
.C(n_1),
.Y(n_104)
);

OAI21xp5_ASAP7_75t_L g105 ( 
.A1(n_104),
.A2(n_100),
.B(n_3),
.Y(n_105)
);

XNOR2xp5_ASAP7_75t_L g106 ( 
.A(n_105),
.B(n_5),
.Y(n_106)
);


endmodule