module fake_jpeg_15377_n_144 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_144);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_144;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_141;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_142;
wire n_85;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_9),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_3),
.Y(n_16)
);

BUFx10_ASAP7_75t_L g17 ( 
.A(n_10),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_5),
.Y(n_18)
);

INVx11_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_2),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_12),
.B(n_7),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

BUFx5_ASAP7_75t_L g25 ( 
.A(n_3),
.Y(n_25)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_1),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_0),
.Y(n_28)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_29),
.B(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_21),
.B(n_0),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_30),
.B(n_35),
.Y(n_44)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_14),
.Y(n_31)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_31),
.Y(n_41)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_19),
.Y(n_32)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_32),
.Y(n_43)
);

INVx8_ASAP7_75t_L g33 ( 
.A(n_19),
.Y(n_33)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_33),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

OR2x2_ASAP7_75t_L g48 ( 
.A(n_34),
.B(n_37),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_21),
.B(n_1),
.Y(n_35)
);

INVx11_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_36),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_16),
.Y(n_37)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_39),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g40 ( 
.A1(n_36),
.A2(n_23),
.B1(n_27),
.B2(n_28),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_40),
.A2(n_13),
.B1(n_18),
.B2(n_24),
.Y(n_67)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

INVx3_ASAP7_75t_L g57 ( 
.A(n_42),
.Y(n_57)
);

INVx6_ASAP7_75t_SL g46 ( 
.A(n_31),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_47),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_34),
.B(n_23),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_51),
.B(n_20),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g50 ( 
.A(n_29),
.B(n_17),
.C(n_25),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g61 ( 
.A(n_50),
.B(n_35),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_L g51 ( 
.A1(n_34),
.A2(n_28),
.B(n_27),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_48),
.B(n_49),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_53),
.B(n_54),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_48),
.B(n_49),
.Y(n_54)
);

OAI22xp5_ASAP7_75t_SL g56 ( 
.A1(n_51),
.A2(n_36),
.B1(n_33),
.B2(n_32),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g78 ( 
.A1(n_56),
.A2(n_59),
.B1(n_43),
.B2(n_22),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_31),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_58),
.B(n_60),
.Y(n_82)
);

OAI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_45),
.A2(n_33),
.B1(n_20),
.B2(n_15),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_44),
.B(n_31),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_64),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g62 ( 
.A(n_44),
.B(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_62),
.B(n_63),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_13),
.Y(n_63)
);

A2O1A1Ixp33_ASAP7_75t_L g73 ( 
.A1(n_64),
.A2(n_22),
.B(n_18),
.C(n_24),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_15),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g72 ( 
.A(n_65),
.B(n_66),
.Y(n_72)
);

INVx1_ASAP7_75t_SL g66 ( 
.A(n_43),
.Y(n_66)
);

AOI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_67),
.A2(n_38),
.B1(n_41),
.B2(n_14),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_68),
.Y(n_77)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_68),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_70),
.B(n_71),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_52),
.Y(n_71)
);

OAI21xp5_ASAP7_75t_L g87 ( 
.A1(n_73),
.A2(n_53),
.B(n_54),
.Y(n_87)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_57),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_74),
.Y(n_97)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

HB1xp67_ASAP7_75t_L g86 ( 
.A(n_75),
.Y(n_86)
);

MAJIxp5_ASAP7_75t_L g98 ( 
.A(n_76),
.B(n_26),
.C(n_2),
.Y(n_98)
);

CKINVDCx14_ASAP7_75t_R g85 ( 
.A(n_78),
.Y(n_85)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_60),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_79),
.B(n_80),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g80 ( 
.A(n_55),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_56),
.A2(n_38),
.B1(n_50),
.B2(n_42),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_81),
.A2(n_29),
.B1(n_14),
.B2(n_17),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_84),
.A2(n_17),
.B1(n_25),
.B2(n_26),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_73),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_79),
.B(n_58),
.Y(n_88)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_88),
.B(n_89),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_SL g89 ( 
.A(n_83),
.B(n_61),
.Y(n_89)
);

INVxp67_ASAP7_75t_L g92 ( 
.A(n_72),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_92),
.B(n_74),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_69),
.B(n_66),
.Y(n_93)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_93),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_94),
.A2(n_95),
.B1(n_77),
.B2(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g96 ( 
.A(n_83),
.B(n_8),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_96),
.B(n_9),
.Y(n_100)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_98),
.B(n_81),
.C(n_82),
.Y(n_104)
);

XOR2xp5_ASAP7_75t_L g99 ( 
.A(n_88),
.B(n_76),
.Y(n_99)
);

XNOR2xp5_ASAP7_75t_L g113 ( 
.A(n_99),
.B(n_104),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_100),
.B(n_101),
.Y(n_120)
);

BUFx2_ASAP7_75t_L g101 ( 
.A(n_86),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_92),
.B(n_78),
.Y(n_102)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_102),
.Y(n_112)
);

AOI221xp5_ASAP7_75t_L g119 ( 
.A1(n_103),
.A2(n_109),
.B1(n_4),
.B2(n_6),
.C(n_11),
.Y(n_119)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_107),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_90),
.B(n_70),
.Y(n_108)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_108),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_89),
.B(n_77),
.C(n_4),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_110),
.A2(n_98),
.B1(n_87),
.B2(n_85),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_111),
.B(n_118),
.C(n_104),
.Y(n_122)
);

AOI21x1_ASAP7_75t_L g114 ( 
.A1(n_99),
.A2(n_94),
.B(n_97),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_114),
.B(n_119),
.Y(n_124)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_101),
.Y(n_117)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_117),
.Y(n_125)
);

OAI21xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_91),
.B(n_97),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_117),
.B(n_116),
.Y(n_121)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_121),
.Y(n_130)
);

MAJIxp5_ASAP7_75t_L g131 ( 
.A(n_122),
.B(n_127),
.C(n_113),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_120),
.Y(n_123)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_123),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_116),
.B(n_105),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g129 ( 
.A(n_126),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_115),
.B(n_110),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_125),
.A2(n_112),
.B1(n_114),
.B2(n_124),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_L g133 ( 
.A1(n_128),
.A2(n_131),
.B(n_121),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g137 ( 
.A(n_133),
.B(n_135),
.Y(n_137)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_130),
.Y(n_134)
);

OAI22xp5_ASAP7_75t_L g139 ( 
.A1(n_134),
.A2(n_136),
.B1(n_11),
.B2(n_12),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_129),
.B(n_111),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_SL g136 ( 
.A(n_132),
.B(n_113),
.Y(n_136)
);

XOR2xp5_ASAP7_75t_L g138 ( 
.A(n_133),
.B(n_129),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_1),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_139),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_140),
.B(n_137),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_142),
.B(n_138),
.Y(n_143)
);

XNOR2xp5_ASAP7_75t_L g144 ( 
.A(n_143),
.B(n_141),
.Y(n_144)
);


endmodule