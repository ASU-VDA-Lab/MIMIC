module fake_ibex_518_n_4419 (n_151, n_85, n_599, n_778, n_507, n_743, n_540, n_754, n_395, n_84, n_64, n_171, n_756, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_766, n_688, n_130, n_177, n_707, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_790, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_773, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_733, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_727, n_58, n_43, n_216, n_33, n_652, n_781, n_421, n_738, n_475, n_802, n_166, n_163, n_753, n_645, n_500, n_747, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_761, n_556, n_748, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_708, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_723, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_739, n_755, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_770, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_711, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_714, n_703, n_426, n_323, n_469, n_598, n_143, n_740, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_736, n_169, n_10, n_673, n_21, n_732, n_798, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_785, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_787, n_614, n_370, n_431, n_719, n_574, n_0, n_289, n_716, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_750, n_746, n_22, n_136, n_261, n_742, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_789, n_654, n_656, n_724, n_437, n_731, n_602, n_355, n_767, n_474, n_758, n_594, n_636, n_710, n_720, n_407, n_102, n_490, n_568, n_813, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_715, n_791, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_769, n_222, n_660, n_186, n_524, n_349, n_765, n_454, n_777, n_295, n_730, n_331, n_576, n_230, n_96, n_759, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_793, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_771, n_205, n_618, n_488, n_139, n_514, n_705, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_783, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_704, n_643, n_137, n_679, n_772, n_810, n_768, n_338, n_173, n_696, n_796, n_797, n_477, n_640, n_363, n_402, n_725, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_718, n_801, n_44, n_672, n_722, n_401, n_553, n_554, n_66, n_735, n_305, n_713, n_307, n_192, n_804, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_721, n_4, n_814, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_763, n_745, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_788, n_795, n_592, n_495, n_762, n_410, n_308, n_675, n_800, n_463, n_624, n_706, n_411, n_135, n_520, n_784, n_684, n_775, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_803, n_692, n_36, n_627, n_18, n_709, n_322, n_53, n_227, n_499, n_115, n_757, n_11, n_248, n_92, n_702, n_451, n_712, n_101, n_190, n_138, n_650, n_776, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_799, n_517, n_211, n_744, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_734, n_468, n_223, n_381, n_525, n_780, n_535, n_382, n_502, n_681, n_633, n_532, n_726, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_729, n_741, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_782, n_217, n_324, n_391, n_537, n_728, n_78, n_805, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_786, n_639, n_303, n_362, n_717, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_809, n_752, n_668, n_779, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_811, n_808, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_792, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_774, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_737, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_794, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_807, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_760, n_751, n_806, n_160, n_657, n_764, n_184, n_56, n_492, n_649, n_812, n_232, n_380, n_749, n_281, n_559, n_425, n_4419);

input n_151;
input n_85;
input n_599;
input n_778;
input n_507;
input n_743;
input n_540;
input n_754;
input n_395;
input n_84;
input n_64;
input n_171;
input n_756;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_766;
input n_688;
input n_130;
input n_177;
input n_707;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_790;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_773;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_733;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_727;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_781;
input n_421;
input n_738;
input n_475;
input n_802;
input n_166;
input n_163;
input n_753;
input n_645;
input n_500;
input n_747;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_761;
input n_556;
input n_748;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_708;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_723;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_739;
input n_755;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_770;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_711;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_714;
input n_703;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_740;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_736;
input n_169;
input n_10;
input n_673;
input n_21;
input n_732;
input n_798;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_785;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_787;
input n_614;
input n_370;
input n_431;
input n_719;
input n_574;
input n_0;
input n_289;
input n_716;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_750;
input n_746;
input n_22;
input n_136;
input n_261;
input n_742;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_789;
input n_654;
input n_656;
input n_724;
input n_437;
input n_731;
input n_602;
input n_355;
input n_767;
input n_474;
input n_758;
input n_594;
input n_636;
input n_710;
input n_720;
input n_407;
input n_102;
input n_490;
input n_568;
input n_813;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_715;
input n_791;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_769;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_765;
input n_454;
input n_777;
input n_295;
input n_730;
input n_331;
input n_576;
input n_230;
input n_96;
input n_759;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_793;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_771;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_705;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_783;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_704;
input n_643;
input n_137;
input n_679;
input n_772;
input n_810;
input n_768;
input n_338;
input n_173;
input n_696;
input n_796;
input n_797;
input n_477;
input n_640;
input n_363;
input n_402;
input n_725;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_718;
input n_801;
input n_44;
input n_672;
input n_722;
input n_401;
input n_553;
input n_554;
input n_66;
input n_735;
input n_305;
input n_713;
input n_307;
input n_192;
input n_804;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_721;
input n_4;
input n_814;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_763;
input n_745;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_788;
input n_795;
input n_592;
input n_495;
input n_762;
input n_410;
input n_308;
input n_675;
input n_800;
input n_463;
input n_624;
input n_706;
input n_411;
input n_135;
input n_520;
input n_784;
input n_684;
input n_775;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_803;
input n_692;
input n_36;
input n_627;
input n_18;
input n_709;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_757;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_712;
input n_101;
input n_190;
input n_138;
input n_650;
input n_776;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_799;
input n_517;
input n_211;
input n_744;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_734;
input n_468;
input n_223;
input n_381;
input n_525;
input n_780;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_726;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_729;
input n_741;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_782;
input n_217;
input n_324;
input n_391;
input n_537;
input n_728;
input n_78;
input n_805;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_786;
input n_639;
input n_303;
input n_362;
input n_717;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_809;
input n_752;
input n_668;
input n_779;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_811;
input n_808;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_792;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_774;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_737;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_794;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_807;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_760;
input n_751;
input n_806;
input n_160;
input n_657;
input n_764;
input n_184;
input n_56;
input n_492;
input n_649;
input n_812;
input n_232;
input n_380;
input n_749;
input n_281;
input n_559;
input n_425;

output n_4419;

wire n_1084;
wire n_4368;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_3853;
wire n_2512;
wire n_3590;
wire n_4056;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3610;
wire n_3911;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_4234;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_4146;
wire n_2835;
wire n_3915;
wire n_1100;
wire n_4158;
wire n_3559;
wire n_845;
wire n_4095;
wire n_2177;
wire n_1930;
wire n_2123;
wire n_4204;
wire n_4364;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2235;
wire n_1802;
wire n_2498;
wire n_3817;
wire n_3755;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_3812;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_909;
wire n_862;
wire n_2290;
wire n_3750;
wire n_3838;
wire n_957;
wire n_3255;
wire n_3272;
wire n_3674;
wire n_4249;
wire n_1652;
wire n_969;
wire n_1859;
wire n_1954;
wire n_2183;
wire n_4346;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_4159;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2682;
wire n_2640;
wire n_3605;
wire n_930;
wire n_4372;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_4004;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_3569;
wire n_4343;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_3819;
wire n_2598;
wire n_4353;
wire n_1722;
wire n_4371;
wire n_3931;
wire n_911;
wire n_2023;
wire n_2720;
wire n_3870;
wire n_4179;
wire n_3340;
wire n_2335;
wire n_1233;
wire n_2322;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3653;
wire n_3519;
wire n_4360;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_3843;
wire n_2139;
wire n_2847;
wire n_3693;
wire n_3033;
wire n_4399;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_1096;
wire n_2391;
wire n_2151;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3440;
wire n_3135;
wire n_3904;
wire n_4378;
wire n_850;
wire n_4169;
wire n_3175;
wire n_3729;
wire n_4239;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_3570;
wire n_879;
wire n_2179;
wire n_1957;
wire n_4197;
wire n_2188;
wire n_1144;
wire n_2359;
wire n_2360;
wire n_2506;
wire n_3984;
wire n_4233;
wire n_4369;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_3830;
wire n_3598;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_3721;
wire n_4418;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_3726;
wire n_4172;
wire n_1730;
wire n_4277;
wire n_1307;
wire n_875;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_1840;
wire n_3479;
wire n_2837;
wire n_3751;
wire n_989;
wire n_3262;
wire n_3407;
wire n_3804;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_3982;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_4201;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_4285;
wire n_1681;
wire n_2921;
wire n_4031;
wire n_3724;
wire n_939;
wire n_1636;
wire n_1687;
wire n_4120;
wire n_3192;
wire n_3533;
wire n_3896;
wire n_3753;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3566;
wire n_4065;
wire n_3469;
wire n_3170;
wire n_4155;
wire n_1922;
wire n_3890;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_2311;
wire n_1937;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_3839;
wire n_1654;
wire n_3577;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_3976;
wire n_824;
wire n_4304;
wire n_4348;
wire n_1945;
wire n_2638;
wire n_3939;
wire n_4160;
wire n_4382;
wire n_2860;
wire n_2448;
wire n_3631;
wire n_4002;
wire n_2015;
wire n_3807;
wire n_2537;
wire n_1130;
wire n_4246;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_3987;
wire n_3845;
wire n_3641;
wire n_2163;
wire n_3969;
wire n_1081;
wire n_2354;
wire n_3639;
wire n_3856;
wire n_1155;
wire n_1292;
wire n_3996;
wire n_4311;
wire n_2432;
wire n_2873;
wire n_3043;
wire n_1576;
wire n_1664;
wire n_4144;
wire n_2273;
wire n_3298;
wire n_1427;
wire n_852;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_4015;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_4211;
wire n_3264;
wire n_3204;
wire n_4119;
wire n_2003;
wire n_1970;
wire n_3671;
wire n_3946;
wire n_3727;
wire n_2621;
wire n_3620;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3881;
wire n_3949;
wire n_3507;
wire n_3884;
wire n_3103;
wire n_2839;
wire n_3926;
wire n_1030;
wire n_1698;
wire n_3688;
wire n_1094;
wire n_2462;
wire n_3770;
wire n_1496;
wire n_1910;
wire n_2333;
wire n_1663;
wire n_2436;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_1595;
wire n_2164;
wire n_3711;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_4349;
wire n_1886;
wire n_2269;
wire n_3748;
wire n_857;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_4389;
wire n_2685;
wire n_3197;
wire n_2846;
wire n_3668;
wire n_1955;
wire n_3699;
wire n_4312;
wire n_917;
wire n_2413;
wire n_2249;
wire n_2362;
wire n_968;
wire n_3148;
wire n_3022;
wire n_2822;
wire n_3766;
wire n_4014;
wire n_1253;
wire n_3707;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_4217;
wire n_4214;
wire n_1313;
wire n_3973;
wire n_4223;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3977;
wire n_3722;
wire n_3125;
wire n_2812;
wire n_3802;
wire n_3681;
wire n_2753;
wire n_3603;
wire n_1638;
wire n_4221;
wire n_2215;
wire n_1449;
wire n_1071;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_3882;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_3979;
wire n_3714;
wire n_3592;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_3565;
wire n_3883;
wire n_2906;
wire n_3097;
wire n_3030;
wire n_3943;
wire n_3809;
wire n_979;
wire n_1309;
wire n_1999;
wire n_3810;
wire n_3718;
wire n_1316;
wire n_1562;
wire n_3917;
wire n_1215;
wire n_3679;
wire n_3579;
wire n_2777;
wire n_2480;
wire n_3769;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_3910;
wire n_2813;
wire n_2147;
wire n_4295;
wire n_1716;
wire n_4238;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_3667;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_3822;
wire n_4171;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_3858;
wire n_4182;
wire n_1401;
wire n_4173;
wire n_3764;
wire n_3795;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_3765;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_4166;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_4259;
wire n_1561;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_3967;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_3842;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_3799;
wire n_2767;
wire n_3676;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_4060;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_1388;
wire n_2859;
wire n_2564;
wire n_3780;
wire n_3023;
wire n_1653;
wire n_4067;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_3762;
wire n_3965;
wire n_1969;
wire n_3798;
wire n_1296;
wire n_3060;
wire n_4124;
wire n_1326;
wire n_971;
wire n_1350;
wire n_3627;
wire n_906;
wire n_2957;
wire n_2586;
wire n_3958;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_4393;
wire n_978;
wire n_3777;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3916;
wire n_3381;
wire n_3630;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_3961;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_3618;
wire n_4078;
wire n_4283;
wire n_1794;
wire n_1423;
wire n_3836;
wire n_4174;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3732;
wire n_3779;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_3923;
wire n_4392;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3808;
wire n_4054;
wire n_3093;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_3716;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_4129;
wire n_4012;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_3567;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_4352;
wire n_3530;
wire n_1613;
wire n_820;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_3874;
wire n_4258;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_4290;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_3909;
wire n_3971;
wire n_1332;
wire n_2660;
wire n_4252;
wire n_2661;
wire n_4079;
wire n_4219;
wire n_2292;
wire n_3573;
wire n_3563;
wire n_3510;
wire n_3560;
wire n_4248;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_4240;
wire n_3652;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_3847;
wire n_4398;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_4055;
wire n_2693;
wire n_3194;
wire n_3607;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_3572;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_3887;
wire n_3963;
wire n_3800;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3951;
wire n_3355;
wire n_2529;
wire n_4126;
wire n_3583;
wire n_2019;
wire n_4103;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3832;
wire n_3508;
wire n_1003;
wire n_889;
wire n_3827;
wire n_2708;
wire n_3156;
wire n_4303;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_3698;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_4400;
wire n_2499;
wire n_3370;
wire n_4359;
wire n_1504;
wire n_3814;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_3888;
wire n_2069;
wire n_4331;
wire n_2602;
wire n_4090;
wire n_1441;
wire n_4105;
wire n_4206;
wire n_2028;
wire n_3309;
wire n_3678;
wire n_4136;
wire n_1924;
wire n_4216;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_4358;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_3968;
wire n_819;
wire n_3950;
wire n_4177;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_3471;
wire n_4098;
wire n_3117;
wire n_3320;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_3900;
wire n_1319;
wire n_4376;
wire n_4050;
wire n_1553;
wire n_3478;
wire n_3701;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_3756;
wire n_2828;
wire n_3754;
wire n_4156;
wire n_1964;
wire n_4411;
wire n_4408;
wire n_1090;
wire n_3720;
wire n_3374;
wire n_1196;
wire n_3704;
wire n_1182;
wire n_1271;
wire n_3811;
wire n_4074;
wire n_2416;
wire n_3633;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_4355;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_3694;
wire n_2052;
wire n_3690;
wire n_981;
wire n_3628;
wire n_3983;
wire n_2425;
wire n_2800;
wire n_4225;
wire n_3514;
wire n_3091;
wire n_4037;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_3859;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_3957;
wire n_3660;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_4308;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_4271;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3634;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_3788;
wire n_1377;
wire n_2473;
wire n_4096;
wire n_1583;
wire n_3520;
wire n_4404;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_974;
wire n_1036;
wire n_2599;
wire n_1831;
wire n_3626;
wire n_3733;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_3684;
wire n_1634;
wire n_3986;
wire n_2853;
wire n_1932;
wire n_3775;
wire n_1452;
wire n_1552;
wire n_1318;
wire n_4006;
wire n_1508;
wire n_2217;
wire n_3741;
wire n_3854;
wire n_1217;
wire n_3594;
wire n_2866;
wire n_3970;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_3966;
wire n_4293;
wire n_1189;
wire n_4008;
wire n_3300;
wire n_1713;
wire n_3621;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_4039;
wire n_4253;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_4122;
wire n_2622;
wire n_3232;
wire n_4250;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_3815;
wire n_4374;
wire n_1140;
wire n_1985;
wire n_4375;
wire n_4205;
wire n_1772;
wire n_2858;
wire n_3708;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3790;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_4403;
wire n_1421;
wire n_1203;
wire n_3640;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_4230;
wire n_859;
wire n_3849;
wire n_1109;
wire n_965;
wire n_4402;
wire n_2741;
wire n_2793;
wire n_4333;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_4070;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_4134;
wire n_1051;
wire n_4180;
wire n_4131;
wire n_1008;
wire n_2964;
wire n_3065;
wire n_2375;
wire n_4062;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_4330;
wire n_1656;
wire n_1207;
wire n_4040;
wire n_1735;
wire n_1076;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_1884;
wire n_2176;
wire n_3813;
wire n_1825;
wire n_2805;
wire n_4232;
wire n_1589;
wire n_2717;
wire n_4199;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_3757;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_4033;
wire n_3855;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3964;
wire n_3110;
wire n_1677;
wire n_1246;
wire n_1236;
wire n_3364;
wire n_4384;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_4231;
wire n_3188;
wire n_3037;
wire n_2780;
wire n_3787;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1477;
wire n_1184;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_4005;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_4323;
wire n_4407;
wire n_4184;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_4073;
wire n_1918;
wire n_2606;
wire n_3642;
wire n_2549;
wire n_4325;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_4113;
wire n_1229;
wire n_4337;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_3680;
wire n_1153;
wire n_3624;
wire n_1751;
wire n_2787;
wire n_3785;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_4292;
wire n_4187;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_3821;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_4261;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_3872;
wire n_1014;
wire n_3801;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_4063;
wire n_1464;
wire n_1566;
wire n_4362;
wire n_3568;
wire n_944;
wire n_3312;
wire n_4128;
wire n_4092;
wire n_3003;
wire n_4244;
wire n_1848;
wire n_4009;
wire n_2062;
wire n_2277;
wire n_3841;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_3932;
wire n_2888;
wire n_2339;
wire n_3614;
wire n_1334;
wire n_3879;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_2999;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_3331;
wire n_2590;
wire n_4414;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_4114;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_4347;
wire n_1852;
wire n_4191;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_3868;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_4209;
wire n_3554;
wire n_2481;
wire n_3692;
wire n_1064;
wire n_4409;
wire n_1408;
wire n_2832;
wire n_3913;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_3730;
wire n_2808;
wire n_2287;
wire n_3597;
wire n_3396;
wire n_4011;
wire n_4190;
wire n_2954;
wire n_4307;
wire n_3526;
wire n_2102;
wire n_4356;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_3558;
wire n_2142;
wire n_1548;
wire n_3703;
wire n_2977;
wire n_1682;
wire n_4151;
wire n_1608;
wire n_3776;
wire n_3599;
wire n_4170;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_4097;
wire n_1436;
wire n_3239;
wire n_4137;
wire n_2600;
wire n_1485;
wire n_1069;
wire n_2239;
wire n_4152;
wire n_1465;
wire n_3952;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_3826;
wire n_4365;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_3781;
wire n_4415;
wire n_1345;
wire n_4215;
wire n_4315;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_3578;
wire n_1628;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_3580;
wire n_2369;
wire n_3584;
wire n_3797;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_3470;
wire n_1395;
wire n_1115;
wire n_1729;
wire n_998;
wire n_2551;
wire n_3281;
wire n_2823;
wire n_3274;
wire n_4064;
wire n_4110;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_4379;
wire n_3397;
wire n_2934;
wire n_4145;
wire n_2807;
wire n_4047;
wire n_882;
wire n_4157;
wire n_942;
wire n_1627;
wire n_1431;
wire n_3956;
wire n_3880;
wire n_4042;
wire n_2525;
wire n_3829;
wire n_1864;
wire n_943;
wire n_4317;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_3587;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_3796;
wire n_2648;
wire n_2458;
wire n_4041;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_4297;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_4115;
wire n_2905;
wire n_3460;
wire n_3978;
wire n_3954;
wire n_2570;
wire n_4051;
wire n_4321;
wire n_3123;
wire n_4025;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2418;
wire n_2184;
wire n_1087;
wire n_3390;
wire n_3948;
wire n_3719;
wire n_1599;
wire n_1400;
wire n_1539;
wire n_1806;
wire n_2711;
wire n_3070;
wire n_2842;
wire n_3646;
wire n_3477;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_4416;
wire n_3074;
wire n_3897;
wire n_4077;
wire n_4024;
wire n_3020;
wire n_3142;
wire n_3975;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_4010;
wire n_4255;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_4059;
wire n_4130;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_3991;
wire n_4361;
wire n_3974;
wire n_1574;
wire n_2200;
wire n_1705;
wire n_3625;
wire n_2304;
wire n_4237;
wire n_1746;
wire n_1439;
wire n_2263;
wire n_2352;
wire n_2212;
wire n_2716;
wire n_3495;
wire n_863;
wire n_2185;
wire n_4141;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_3759;
wire n_4035;
wire n_2781;
wire n_4291;
wire n_3419;
wire n_3629;
wire n_2460;
wire n_2170;
wire n_3600;
wire n_1785;
wire n_4109;
wire n_1870;
wire n_2484;
wire n_3999;
wire n_4117;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_4087;
wire n_3167;
wire n_3687;
wire n_997;
wire n_4154;
wire n_2308;
wire n_3459;
wire n_3498;
wire n_2986;
wire n_3238;
wire n_1428;
wire n_2691;
wire n_4026;
wire n_4318;
wire n_2243;
wire n_2400;
wire n_3731;
wire n_3092;
wire n_3555;
wire n_4385;
wire n_2903;
wire n_891;
wire n_3659;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_4052;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_3682;
wire n_3434;
wire n_2463;
wire n_2654;
wire n_3840;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_4072;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_4245;
wire n_1512;
wire n_3672;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_3885;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_4100;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_3877;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_3936;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_3953;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_3834;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3656;
wire n_3257;
wire n_1048;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_3638;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_3816;
wire n_2450;
wire n_4195;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_3925;
wire n_4089;
wire n_4176;
wire n_1683;
wire n_1185;
wire n_4256;
wire n_3575;
wire n_4175;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_4278;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_3772;
wire n_2948;
wire n_916;
wire n_4322;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_4336;
wire n_3219;
wire n_2936;
wire n_895;
wire n_3955;
wire n_3867;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_4227;
wire n_2190;
wire n_1127;
wire n_932;
wire n_3657;
wire n_1972;
wire n_3080;
wire n_4030;
wire n_2772;
wire n_2778;
wire n_947;
wire n_1004;
wire n_4276;
wire n_831;
wire n_3929;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1845;
wire n_1104;
wire n_2205;
wire n_1011;
wire n_2875;
wire n_2684;
wire n_2524;
wire n_3835;
wire n_1437;
wire n_3284;
wire n_3723;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_3927;
wire n_4185;
wire n_2422;
wire n_3902;
wire n_4203;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_3564;
wire n_2385;
wire n_3095;
wire n_3864;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3695;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_4381;
wire n_1917;
wire n_4314;
wire n_1444;
wire n_4133;
wire n_920;
wire n_4316;
wire n_2442;
wire n_3985;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_4083;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_4020;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_4306;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_2896;
wire n_3064;
wire n_4228;
wire n_3314;
wire n_3747;
wire n_1349;
wire n_991;
wire n_1331;
wire n_961;
wire n_1223;
wire n_2127;
wire n_3735;
wire n_1323;
wire n_3891;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3228;
wire n_3028;
wire n_3710;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3706;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3588;
wire n_4003;
wire n_4254;
wire n_3420;
wire n_1432;
wire n_4192;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_4247;
wire n_4071;
wire n_4388;
wire n_996;
wire n_3632;
wire n_3914;
wire n_915;
wire n_2238;
wire n_3289;
wire n_1174;
wire n_1834;
wire n_1874;
wire n_3372;
wire n_3499;
wire n_4138;
wire n_3552;
wire n_4121;
wire n_3850;
wire n_2862;
wire n_3100;
wire n_4116;
wire n_4164;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3784;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_4118;
wire n_4142;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_3828;
wire n_1291;
wire n_2895;
wire n_3763;
wire n_1914;
wire n_3833;
wire n_4284;
wire n_1458;
wire n_1694;
wire n_4370;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_3673;
wire n_3990;
wire n_4066;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_4044;
wire n_1826;
wire n_1855;
wire n_4241;
wire n_1662;
wire n_2187;
wire n_2105;
wire n_3556;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3609;
wire n_4135;
wire n_3447;
wire n_3771;
wire n_2647;
wire n_1626;
wire n_3995;
wire n_4104;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3876;
wire n_3152;
wire n_4000;
wire n_3154;
wire n_4123;
wire n_2344;
wire n_3589;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_3616;
wire n_3908;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_3696;
wire n_4305;
wire n_2902;
wire n_4048;
wire n_4084;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3960;
wire n_4007;
wire n_3608;
wire n_4339;
wire n_4269;
wire n_4085;
wire n_3190;
wire n_1524;
wire n_1055;
wire n_3878;
wire n_4016;
wire n_2849;
wire n_2947;
wire n_4080;
wire n_1754;
wire n_4286;
wire n_3048;
wire n_3686;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_4028;
wire n_2210;
wire n_1517;
wire n_3940;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_3670;
wire n_1624;
wire n_1952;
wire n_2180;
wire n_3002;
wire n_3376;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_4289;
wire n_2617;
wire n_3585;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_1491;
wire n_1860;
wire n_4163;
wire n_2831;
wire n_1810;
wire n_1763;
wire n_923;
wire n_3778;
wire n_3912;
wire n_3818;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_2959;
wire n_1625;
wire n_3047;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_3993;
wire n_2120;
wire n_1037;
wire n_1899;
wire n_2031;
wire n_3669;
wire n_3427;
wire n_4001;
wire n_1289;
wire n_1348;
wire n_838;
wire n_2892;
wire n_1021;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_4099;
wire n_4377;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_3783;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_4264;
wire n_1942;
wire n_4326;
wire n_3666;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_1617;
wire n_1839;
wire n_3899;
wire n_3930;
wire n_1587;
wire n_2555;
wire n_2330;
wire n_2639;
wire n_4149;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_3712;
wire n_4101;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_4057;
wire n_2410;
wire n_3760;
wire n_4319;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_3736;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_4021;
wire n_1538;
wire n_2528;
wire n_3773;
wire n_4383;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_3717;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_2604;
wire n_3745;
wire n_3424;
wire n_3462;
wire n_4373;
wire n_2437;
wire n_2351;
wire n_3664;
wire n_2049;
wire n_1456;
wire n_3907;
wire n_1889;
wire n_3245;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3862;
wire n_3302;
wire n_1673;
wire n_4132;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_851;
wire n_993;
wire n_4202;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_4287;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2320;
wire n_2237;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_4300;
wire n_3921;
wire n_1800;
wire n_3277;
wire n_3746;
wire n_2758;
wire n_3480;
wire n_4417;
wire n_1494;
wire n_1550;
wire n_3906;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_4022;
wire n_4212;
wire n_1241;
wire n_3645;
wire n_4262;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_4019;
wire n_2736;
wire n_4320;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_3506;
wire n_2845;
wire n_2735;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_2984;
wire n_3162;
wire n_1906;
wire n_3004;
wire n_3886;
wire n_1647;
wire n_1901;
wire n_4357;
wire n_3096;
wire n_3333;
wire n_839;
wire n_3705;
wire n_4023;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_3276;
wire n_4366;
wire n_1006;
wire n_2956;
wire n_1415;
wire n_1238;
wire n_3959;
wire n_3743;
wire n_976;
wire n_1710;
wire n_4139;
wire n_3021;
wire n_1063;
wire n_4068;
wire n_4288;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_4340;
wire n_3825;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_3892;
wire n_1406;
wire n_1489;
wire n_3591;
wire n_1880;
wire n_1993;
wire n_3860;
wire n_2137;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_4034;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_3920;
wire n_1202;
wire n_3848;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_4082;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_3273;
wire n_4367;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_4282;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_4222;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_3734;
wire n_3637;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3650;
wire n_3327;
wire n_2265;
wire n_1114;
wire n_3513;
wire n_3709;
wire n_3011;
wire n_818;
wire n_1167;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3623;
wire n_3647;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_4029;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3619;
wire n_3349;
wire n_3928;
wire n_4043;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_4167;
wire n_3058;
wire n_3454;
wire n_4334;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_4143;
wire n_2272;
wire n_1956;
wire n_3574;
wire n_4410;
wire n_2608;
wire n_4270;
wire n_3384;
wire n_2983;
wire n_4273;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_3739;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_858;
wire n_1018;
wire n_2345;
wire n_1324;
wire n_4338;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3604;
wire n_1838;
wire n_3649;
wire n_833;
wire n_3540;
wire n_3824;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_4198;
wire n_1513;
wire n_3740;
wire n_4397;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_4181;
wire n_2161;
wire n_2191;
wire n_3611;
wire n_2329;
wire n_1788;
wire n_4186;
wire n_2348;
wire n_2093;
wire n_2675;
wire n_2417;
wire n_2576;
wire n_2043;
wire n_3601;
wire n_4344;
wire n_2366;
wire n_4229;
wire n_4294;
wire n_1621;
wire n_2338;
wire n_3571;
wire n_1919;
wire n_1342;
wire n_4351;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_4111;
wire n_4162;
wire n_4200;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_3962;
wire n_3875;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_3846;
wire n_4341;
wire n_4328;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_4127;
wire n_1688;
wire n_2973;
wire n_3651;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3059;
wire n_3085;
wire n_1242;
wire n_1119;
wire n_2229;
wire n_2810;
wire n_2867;
wire n_3871;
wire n_1085;
wire n_3027;
wire n_4076;
wire n_4189;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_4390;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_3994;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_3648;
wire n_2471;
wire n_1288;
wire n_4058;
wire n_1275;
wire n_985;
wire n_1165;
wire n_4148;
wire n_1622;
wire n_897;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_4081;
wire n_4391;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_4032;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_4268;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_3236;
wire n_3576;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_4265;
wire n_3062;
wire n_3806;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_1565;
wire n_1257;
wire n_3805;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_4260;
wire n_3391;
wire n_4017;
wire n_1547;
wire n_1542;
wire n_946;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_4178;
wire n_4324;
wire n_1097;
wire n_3354;
wire n_4069;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_4236;
wire n_3012;
wire n_4313;
wire n_4140;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_3561;
wire n_956;
wire n_4125;
wire n_3586;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_4242;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_3767;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_3942;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_4243;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3820;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_3697;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_4053;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_4279;
wire n_3937;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_4235;
wire n_3227;
wire n_1438;
wire n_3774;
wire n_3972;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2494;
wire n_2156;
wire n_4036;
wire n_2126;
wire n_1147;
wire n_3863;
wire n_1363;
wire n_3403;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1518;
wire n_1366;
wire n_4350;
wire n_4380;
wire n_1361;
wire n_1187;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_4281;
wire n_4345;
wire n_2411;
wire n_4332;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_3998;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_3866;
wire n_3761;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3803;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_3989;
wire n_2119;
wire n_1010;
wire n_3844;
wire n_883;
wire n_2207;
wire n_4210;
wire n_4049;
wire n_2044;
wire n_2542;
wire n_2091;
wire n_3918;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_4165;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_1635;
wire n_1572;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_3643;
wire n_2615;
wire n_3278;
wire n_2487;
wire n_2701;
wire n_3163;
wire n_2929;
wire n_3343;
wire n_3752;
wire n_4310;
wire n_3786;
wire n_4061;
wire n_2637;
wire n_1329;
wire n_2409;
wire n_2337;
wire n_4045;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_4405;
wire n_3118;
wire n_1369;
wire n_1297;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_3742;
wire n_3655;
wire n_3791;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_4091;
wire n_2323;
wire n_3532;
wire n_4257;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_2997;
wire n_967;
wire n_2561;
wire n_4263;
wire n_3725;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_4363;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_4196;
wire n_4335;
wire n_2371;
wire n_914;
wire n_4147;
wire n_3992;
wire n_3444;
wire n_1986;
wire n_3898;
wire n_4218;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_4301;
wire n_4107;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2429;
wire n_2408;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3581;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3547;
wire n_3423;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_3700;
wire n_4161;
wire n_2514;
wire n_2466;
wire n_3661;
wire n_4267;
wire n_4386;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_1299;
wire n_2942;
wire n_3947;
wire n_2096;
wire n_3663;
wire n_3562;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_3665;
wire n_2079;
wire n_4193;
wire n_2296;
wire n_4342;
wire n_3782;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_3831;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_3683;
wire n_3919;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_4302;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_4013;
wire n_1397;
wire n_1211;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_3794;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_3702;
wire n_3981;
wire n_1532;
wire n_4406;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3430;
wire n_3200;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1488;
wire n_1193;
wire n_849;
wire n_980;
wire n_2928;
wire n_3067;
wire n_2227;
wire n_2652;
wire n_3225;
wire n_1074;
wire n_3557;
wire n_3380;
wire n_3207;
wire n_3596;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3606;
wire n_3369;
wire n_3823;
wire n_4086;
wire n_3185;
wire n_2326;
wire n_3869;
wire n_1866;
wire n_3852;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_4112;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_4207;
wire n_960;
wire n_1022;
wire n_4412;
wire n_1760;
wire n_3737;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_4266;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_3286;
wire n_999;
wire n_2634;
wire n_2982;
wire n_4038;
wire n_1092;
wire n_3124;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_3636;
wire n_910;
wire n_2291;
wire n_3837;
wire n_4102;
wire n_3612;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_1385;
wire n_2927;
wire n_4274;
wire n_1062;
wire n_4395;
wire n_1230;
wire n_1516;
wire n_1027;
wire n_3893;
wire n_3622;
wire n_3857;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_4272;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2303;
wire n_2104;
wire n_949;
wire n_2148;
wire n_2653;
wire n_2618;
wire n_2357;
wire n_2855;
wire n_3938;
wire n_4354;
wire n_924;
wire n_2937;
wire n_3728;
wire n_3359;
wire n_4401;
wire n_3114;
wire n_2331;
wire n_4296;
wire n_3332;
wire n_3905;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_4413;
wire n_1757;
wire n_4088;
wire n_2136;
wire n_4309;
wire n_3617;
wire n_4027;
wire n_3602;
wire n_4298;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_3922;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_3894;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_1450;
wire n_2082;
wire n_2453;
wire n_2560;
wire n_2302;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_4208;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3052;
wire n_2802;
wire n_3189;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_2066;
wire n_1719;
wire n_1974;
wire n_1158;
wire n_2988;
wire n_3945;
wire n_1882;
wire n_4046;
wire n_4275;
wire n_2961;
wire n_2770;
wire n_2996;
wire n_2704;
wire n_3924;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_3689;
wire n_3582;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_4094;
wire n_3613;
wire n_1383;
wire n_990;
wire n_4108;
wire n_1968;
wire n_3675;
wire n_2057;
wire n_2609;
wire n_4018;
wire n_2378;
wire n_888;
wire n_2749;
wire n_3658;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3901;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_3715;
wire n_4194;
wire n_1059;
wire n_2969;
wire n_3713;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3889;
wire n_3325;
wire n_4299;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_3744;
wire n_1414;
wire n_2246;
wire n_2324;
wire n_2738;
wire n_3861;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_4150;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_3941;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_3933;
wire n_4188;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2619;
wire n_2917;
wire n_2726;
wire n_3873;
wire n_3738;
wire n_2073;
wire n_4093;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_4226;
wire n_1551;
wire n_3793;
wire n_4153;
wire n_1533;
wire n_1145;
wire n_2307;
wire n_2515;
wire n_3792;
wire n_3546;
wire n_1511;
wire n_4329;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3988;
wire n_2327;
wire n_3758;
wire n_3442;
wire n_4327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_4106;
wire n_4251;
wire n_4168;
wire n_1164;
wire n_2258;
wire n_3944;
wire n_3662;
wire n_3595;
wire n_1732;
wire n_3749;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_4396;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_3691;
wire n_2544;
wire n_856;
wire n_3193;
wire n_3635;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_4280;
wire n_2285;
wire n_3213;
wire n_3789;
wire n_1934;
wire n_4394;
wire n_1900;
wire n_2040;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_3934;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_4183;
wire n_1678;
wire n_1780;
wire n_1091;
wire n_2725;
wire n_3865;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_4220;
wire n_4075;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_3997;
wire n_3593;
wire n_2349;
wire n_2100;
wire n_1902;
wire n_2536;
wire n_3903;
wire n_2474;
wire n_3895;
wire n_1150;
wire n_1194;
wire n_1399;
wire n_3685;
wire n_3851;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_3768;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_4224;
wire n_970;
wire n_3654;
wire n_3980;
wire n_2430;
wire n_2673;
wire n_921;
wire n_2676;
wire n_3515;
wire n_3489;
wire n_4213;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3644;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_4387;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_3615;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_3677;
wire n_2657;
wire n_3935;
wire n_1186;
wire n_2065;
wire n_2901;
wire n_3180;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;
wire n_2658;

INVx1_ASAP7_75t_SL g815 ( 
.A(n_354),
.Y(n_815)
);

BUFx6f_ASAP7_75t_L g816 ( 
.A(n_508),
.Y(n_816)
);

CKINVDCx5p33_ASAP7_75t_R g817 ( 
.A(n_326),
.Y(n_817)
);

NOR2xp67_ASAP7_75t_L g818 ( 
.A(n_300),
.B(n_711),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_138),
.Y(n_819)
);

CKINVDCx5p33_ASAP7_75t_R g820 ( 
.A(n_23),
.Y(n_820)
);

BUFx10_ASAP7_75t_L g821 ( 
.A(n_59),
.Y(n_821)
);

INVx1_ASAP7_75t_L g822 ( 
.A(n_250),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_446),
.Y(n_823)
);

INVx1_ASAP7_75t_L g824 ( 
.A(n_636),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_380),
.Y(n_825)
);

BUFx6f_ASAP7_75t_L g826 ( 
.A(n_420),
.Y(n_826)
);

BUFx3_ASAP7_75t_L g827 ( 
.A(n_327),
.Y(n_827)
);

CKINVDCx20_ASAP7_75t_R g828 ( 
.A(n_525),
.Y(n_828)
);

INVx1_ASAP7_75t_L g829 ( 
.A(n_710),
.Y(n_829)
);

INVx2_ASAP7_75t_SL g830 ( 
.A(n_534),
.Y(n_830)
);

CKINVDCx16_ASAP7_75t_R g831 ( 
.A(n_64),
.Y(n_831)
);

INVx1_ASAP7_75t_SL g832 ( 
.A(n_111),
.Y(n_832)
);

INVx1_ASAP7_75t_L g833 ( 
.A(n_379),
.Y(n_833)
);

CKINVDCx5p33_ASAP7_75t_R g834 ( 
.A(n_525),
.Y(n_834)
);

NOR2xp67_ASAP7_75t_L g835 ( 
.A(n_469),
.B(n_592),
.Y(n_835)
);

CKINVDCx5p33_ASAP7_75t_R g836 ( 
.A(n_721),
.Y(n_836)
);

CKINVDCx5p33_ASAP7_75t_R g837 ( 
.A(n_697),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_697),
.Y(n_838)
);

CKINVDCx5p33_ASAP7_75t_R g839 ( 
.A(n_233),
.Y(n_839)
);

INVx1_ASAP7_75t_SL g840 ( 
.A(n_812),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_439),
.Y(n_841)
);

HB1xp67_ASAP7_75t_L g842 ( 
.A(n_594),
.Y(n_842)
);

INVx1_ASAP7_75t_SL g843 ( 
.A(n_743),
.Y(n_843)
);

CKINVDCx5p33_ASAP7_75t_R g844 ( 
.A(n_475),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_735),
.Y(n_845)
);

INVx2_ASAP7_75t_L g846 ( 
.A(n_691),
.Y(n_846)
);

CKINVDCx5p33_ASAP7_75t_R g847 ( 
.A(n_527),
.Y(n_847)
);

CKINVDCx5p33_ASAP7_75t_R g848 ( 
.A(n_291),
.Y(n_848)
);

INVx1_ASAP7_75t_SL g849 ( 
.A(n_148),
.Y(n_849)
);

CKINVDCx5p33_ASAP7_75t_R g850 ( 
.A(n_95),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_676),
.Y(n_851)
);

CKINVDCx5p33_ASAP7_75t_R g852 ( 
.A(n_62),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_550),
.Y(n_853)
);

CKINVDCx20_ASAP7_75t_R g854 ( 
.A(n_19),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_675),
.Y(n_855)
);

CKINVDCx5p33_ASAP7_75t_R g856 ( 
.A(n_706),
.Y(n_856)
);

INVx2_ASAP7_75t_SL g857 ( 
.A(n_680),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_209),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_356),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_61),
.Y(n_860)
);

BUFx2_ASAP7_75t_L g861 ( 
.A(n_96),
.Y(n_861)
);

INVx1_ASAP7_75t_L g862 ( 
.A(n_566),
.Y(n_862)
);

CKINVDCx5p33_ASAP7_75t_R g863 ( 
.A(n_192),
.Y(n_863)
);

INVx1_ASAP7_75t_L g864 ( 
.A(n_364),
.Y(n_864)
);

BUFx3_ASAP7_75t_L g865 ( 
.A(n_407),
.Y(n_865)
);

CKINVDCx5p33_ASAP7_75t_R g866 ( 
.A(n_45),
.Y(n_866)
);

CKINVDCx5p33_ASAP7_75t_R g867 ( 
.A(n_515),
.Y(n_867)
);

INVx1_ASAP7_75t_L g868 ( 
.A(n_694),
.Y(n_868)
);

INVx1_ASAP7_75t_L g869 ( 
.A(n_810),
.Y(n_869)
);

CKINVDCx5p33_ASAP7_75t_R g870 ( 
.A(n_216),
.Y(n_870)
);

BUFx3_ASAP7_75t_L g871 ( 
.A(n_671),
.Y(n_871)
);

CKINVDCx5p33_ASAP7_75t_R g872 ( 
.A(n_546),
.Y(n_872)
);

INVx1_ASAP7_75t_L g873 ( 
.A(n_750),
.Y(n_873)
);

INVx1_ASAP7_75t_L g874 ( 
.A(n_317),
.Y(n_874)
);

INVx1_ASAP7_75t_L g875 ( 
.A(n_70),
.Y(n_875)
);

CKINVDCx5p33_ASAP7_75t_R g876 ( 
.A(n_693),
.Y(n_876)
);

INVx1_ASAP7_75t_L g877 ( 
.A(n_96),
.Y(n_877)
);

CKINVDCx20_ASAP7_75t_R g878 ( 
.A(n_140),
.Y(n_878)
);

CKINVDCx20_ASAP7_75t_R g879 ( 
.A(n_480),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_313),
.Y(n_880)
);

CKINVDCx5p33_ASAP7_75t_R g881 ( 
.A(n_227),
.Y(n_881)
);

INVx2_ASAP7_75t_L g882 ( 
.A(n_496),
.Y(n_882)
);

INVx1_ASAP7_75t_L g883 ( 
.A(n_568),
.Y(n_883)
);

CKINVDCx20_ASAP7_75t_R g884 ( 
.A(n_567),
.Y(n_884)
);

INVx1_ASAP7_75t_L g885 ( 
.A(n_678),
.Y(n_885)
);

INVx1_ASAP7_75t_L g886 ( 
.A(n_167),
.Y(n_886)
);

INVx1_ASAP7_75t_L g887 ( 
.A(n_753),
.Y(n_887)
);

INVx1_ASAP7_75t_L g888 ( 
.A(n_715),
.Y(n_888)
);

INVx1_ASAP7_75t_L g889 ( 
.A(n_691),
.Y(n_889)
);

INVx1_ASAP7_75t_L g890 ( 
.A(n_462),
.Y(n_890)
);

BUFx3_ASAP7_75t_L g891 ( 
.A(n_604),
.Y(n_891)
);

BUFx2_ASAP7_75t_L g892 ( 
.A(n_667),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_686),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_395),
.Y(n_894)
);

NOR2xp67_ASAP7_75t_L g895 ( 
.A(n_622),
.B(n_102),
.Y(n_895)
);

INVx1_ASAP7_75t_L g896 ( 
.A(n_82),
.Y(n_896)
);

INVx1_ASAP7_75t_L g897 ( 
.A(n_3),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_0),
.Y(n_898)
);

INVxp67_ASAP7_75t_SL g899 ( 
.A(n_130),
.Y(n_899)
);

CKINVDCx5p33_ASAP7_75t_R g900 ( 
.A(n_807),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_191),
.Y(n_901)
);

INVx1_ASAP7_75t_L g902 ( 
.A(n_221),
.Y(n_902)
);

INVx1_ASAP7_75t_L g903 ( 
.A(n_797),
.Y(n_903)
);

CKINVDCx5p33_ASAP7_75t_R g904 ( 
.A(n_272),
.Y(n_904)
);

BUFx6f_ASAP7_75t_L g905 ( 
.A(n_677),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_771),
.Y(n_906)
);

INVx1_ASAP7_75t_L g907 ( 
.A(n_708),
.Y(n_907)
);

INVx1_ASAP7_75t_L g908 ( 
.A(n_198),
.Y(n_908)
);

CKINVDCx20_ASAP7_75t_R g909 ( 
.A(n_374),
.Y(n_909)
);

CKINVDCx5p33_ASAP7_75t_R g910 ( 
.A(n_375),
.Y(n_910)
);

INVx1_ASAP7_75t_L g911 ( 
.A(n_572),
.Y(n_911)
);

CKINVDCx11_ASAP7_75t_R g912 ( 
.A(n_437),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_22),
.Y(n_913)
);

CKINVDCx16_ASAP7_75t_R g914 ( 
.A(n_436),
.Y(n_914)
);

CKINVDCx5p33_ASAP7_75t_R g915 ( 
.A(n_459),
.Y(n_915)
);

INVx1_ASAP7_75t_L g916 ( 
.A(n_516),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_793),
.Y(n_917)
);

INVx1_ASAP7_75t_SL g918 ( 
.A(n_719),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_723),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_469),
.Y(n_920)
);

INVx1_ASAP7_75t_L g921 ( 
.A(n_518),
.Y(n_921)
);

CKINVDCx5p33_ASAP7_75t_R g922 ( 
.A(n_235),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_572),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_106),
.Y(n_924)
);

CKINVDCx5p33_ASAP7_75t_R g925 ( 
.A(n_614),
.Y(n_925)
);

INVx1_ASAP7_75t_L g926 ( 
.A(n_664),
.Y(n_926)
);

CKINVDCx5p33_ASAP7_75t_R g927 ( 
.A(n_155),
.Y(n_927)
);

CKINVDCx5p33_ASAP7_75t_R g928 ( 
.A(n_774),
.Y(n_928)
);

CKINVDCx5p33_ASAP7_75t_R g929 ( 
.A(n_726),
.Y(n_929)
);

INVx1_ASAP7_75t_SL g930 ( 
.A(n_178),
.Y(n_930)
);

INVx1_ASAP7_75t_L g931 ( 
.A(n_176),
.Y(n_931)
);

INVx1_ASAP7_75t_SL g932 ( 
.A(n_316),
.Y(n_932)
);

CKINVDCx5p33_ASAP7_75t_R g933 ( 
.A(n_23),
.Y(n_933)
);

BUFx3_ASAP7_75t_L g934 ( 
.A(n_803),
.Y(n_934)
);

CKINVDCx5p33_ASAP7_75t_R g935 ( 
.A(n_775),
.Y(n_935)
);

BUFx3_ASAP7_75t_L g936 ( 
.A(n_705),
.Y(n_936)
);

INVx1_ASAP7_75t_L g937 ( 
.A(n_707),
.Y(n_937)
);

CKINVDCx20_ASAP7_75t_R g938 ( 
.A(n_806),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_693),
.Y(n_939)
);

CKINVDCx5p33_ASAP7_75t_R g940 ( 
.A(n_440),
.Y(n_940)
);

BUFx6f_ASAP7_75t_L g941 ( 
.A(n_637),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_189),
.Y(n_942)
);

CKINVDCx20_ASAP7_75t_R g943 ( 
.A(n_321),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_620),
.Y(n_944)
);

BUFx3_ASAP7_75t_L g945 ( 
.A(n_73),
.Y(n_945)
);

CKINVDCx5p33_ASAP7_75t_R g946 ( 
.A(n_725),
.Y(n_946)
);

CKINVDCx5p33_ASAP7_75t_R g947 ( 
.A(n_390),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_118),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_105),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_143),
.Y(n_950)
);

INVx1_ASAP7_75t_L g951 ( 
.A(n_63),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_83),
.Y(n_952)
);

INVx1_ASAP7_75t_L g953 ( 
.A(n_741),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_809),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_227),
.Y(n_955)
);

INVx1_ASAP7_75t_L g956 ( 
.A(n_698),
.Y(n_956)
);

CKINVDCx20_ASAP7_75t_R g957 ( 
.A(n_411),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_551),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_686),
.Y(n_959)
);

CKINVDCx5p33_ASAP7_75t_R g960 ( 
.A(n_504),
.Y(n_960)
);

CKINVDCx20_ASAP7_75t_R g961 ( 
.A(n_397),
.Y(n_961)
);

INVx1_ASAP7_75t_L g962 ( 
.A(n_392),
.Y(n_962)
);

CKINVDCx5p33_ASAP7_75t_R g963 ( 
.A(n_81),
.Y(n_963)
);

INVx1_ASAP7_75t_SL g964 ( 
.A(n_727),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_578),
.Y(n_965)
);

BUFx10_ASAP7_75t_L g966 ( 
.A(n_523),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_709),
.Y(n_967)
);

CKINVDCx5p33_ASAP7_75t_R g968 ( 
.A(n_642),
.Y(n_968)
);

CKINVDCx20_ASAP7_75t_R g969 ( 
.A(n_69),
.Y(n_969)
);

INVx1_ASAP7_75t_L g970 ( 
.A(n_3),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_792),
.Y(n_971)
);

INVx1_ASAP7_75t_L g972 ( 
.A(n_547),
.Y(n_972)
);

BUFx6f_ASAP7_75t_L g973 ( 
.A(n_700),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_450),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_714),
.Y(n_975)
);

HB1xp67_ASAP7_75t_L g976 ( 
.A(n_233),
.Y(n_976)
);

INVx2_ASAP7_75t_L g977 ( 
.A(n_35),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_297),
.Y(n_978)
);

INVx1_ASAP7_75t_SL g979 ( 
.A(n_673),
.Y(n_979)
);

INVx1_ASAP7_75t_L g980 ( 
.A(n_91),
.Y(n_980)
);

INVx1_ASAP7_75t_L g981 ( 
.A(n_431),
.Y(n_981)
);

CKINVDCx5p33_ASAP7_75t_R g982 ( 
.A(n_680),
.Y(n_982)
);

CKINVDCx5p33_ASAP7_75t_R g983 ( 
.A(n_357),
.Y(n_983)
);

CKINVDCx20_ASAP7_75t_R g984 ( 
.A(n_661),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_135),
.Y(n_985)
);

BUFx2_ASAP7_75t_L g986 ( 
.A(n_188),
.Y(n_986)
);

CKINVDCx5p33_ASAP7_75t_R g987 ( 
.A(n_544),
.Y(n_987)
);

BUFx3_ASAP7_75t_L g988 ( 
.A(n_431),
.Y(n_988)
);

CKINVDCx14_ASAP7_75t_R g989 ( 
.A(n_733),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_699),
.Y(n_990)
);

INVx2_ASAP7_75t_SL g991 ( 
.A(n_213),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_56),
.Y(n_992)
);

INVx1_ASAP7_75t_L g993 ( 
.A(n_495),
.Y(n_993)
);

CKINVDCx5p33_ASAP7_75t_R g994 ( 
.A(n_768),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_378),
.Y(n_995)
);

INVx1_ASAP7_75t_L g996 ( 
.A(n_279),
.Y(n_996)
);

CKINVDCx5p33_ASAP7_75t_R g997 ( 
.A(n_151),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_273),
.Y(n_998)
);

CKINVDCx20_ASAP7_75t_R g999 ( 
.A(n_331),
.Y(n_999)
);

INVx1_ASAP7_75t_L g1000 ( 
.A(n_504),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_690),
.Y(n_1001)
);

CKINVDCx5p33_ASAP7_75t_R g1002 ( 
.A(n_30),
.Y(n_1002)
);

CKINVDCx5p33_ASAP7_75t_R g1003 ( 
.A(n_728),
.Y(n_1003)
);

CKINVDCx5p33_ASAP7_75t_R g1004 ( 
.A(n_498),
.Y(n_1004)
);

CKINVDCx5p33_ASAP7_75t_R g1005 ( 
.A(n_399),
.Y(n_1005)
);

INVx1_ASAP7_75t_L g1006 ( 
.A(n_712),
.Y(n_1006)
);

BUFx10_ASAP7_75t_L g1007 ( 
.A(n_272),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_412),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_393),
.Y(n_1009)
);

INVx3_ASAP7_75t_L g1010 ( 
.A(n_32),
.Y(n_1010)
);

CKINVDCx5p33_ASAP7_75t_R g1011 ( 
.A(n_169),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_221),
.Y(n_1012)
);

INVx1_ASAP7_75t_SL g1013 ( 
.A(n_385),
.Y(n_1013)
);

CKINVDCx20_ASAP7_75t_R g1014 ( 
.A(n_140),
.Y(n_1014)
);

CKINVDCx16_ASAP7_75t_R g1015 ( 
.A(n_747),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_713),
.Y(n_1016)
);

CKINVDCx5p33_ASAP7_75t_R g1017 ( 
.A(n_143),
.Y(n_1017)
);

INVx1_ASAP7_75t_L g1018 ( 
.A(n_732),
.Y(n_1018)
);

HB1xp67_ASAP7_75t_L g1019 ( 
.A(n_764),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_716),
.Y(n_1020)
);

INVx1_ASAP7_75t_L g1021 ( 
.A(n_263),
.Y(n_1021)
);

INVxp67_ASAP7_75t_L g1022 ( 
.A(n_317),
.Y(n_1022)
);

CKINVDCx20_ASAP7_75t_R g1023 ( 
.A(n_375),
.Y(n_1023)
);

CKINVDCx5p33_ASAP7_75t_R g1024 ( 
.A(n_194),
.Y(n_1024)
);

INVx1_ASAP7_75t_L g1025 ( 
.A(n_641),
.Y(n_1025)
);

INVx1_ASAP7_75t_L g1026 ( 
.A(n_286),
.Y(n_1026)
);

INVx1_ASAP7_75t_L g1027 ( 
.A(n_527),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_334),
.Y(n_1028)
);

CKINVDCx5p33_ASAP7_75t_R g1029 ( 
.A(n_668),
.Y(n_1029)
);

INVx1_ASAP7_75t_L g1030 ( 
.A(n_4),
.Y(n_1030)
);

CKINVDCx5p33_ASAP7_75t_R g1031 ( 
.A(n_36),
.Y(n_1031)
);

INVx1_ASAP7_75t_L g1032 ( 
.A(n_177),
.Y(n_1032)
);

INVx1_ASAP7_75t_L g1033 ( 
.A(n_43),
.Y(n_1033)
);

INVx1_ASAP7_75t_L g1034 ( 
.A(n_477),
.Y(n_1034)
);

CKINVDCx5p33_ASAP7_75t_R g1035 ( 
.A(n_318),
.Y(n_1035)
);

CKINVDCx5p33_ASAP7_75t_R g1036 ( 
.A(n_500),
.Y(n_1036)
);

INVx2_ASAP7_75t_L g1037 ( 
.A(n_224),
.Y(n_1037)
);

CKINVDCx20_ASAP7_75t_R g1038 ( 
.A(n_440),
.Y(n_1038)
);

INVx1_ASAP7_75t_L g1039 ( 
.A(n_429),
.Y(n_1039)
);

CKINVDCx20_ASAP7_75t_R g1040 ( 
.A(n_460),
.Y(n_1040)
);

INVx1_ASAP7_75t_SL g1041 ( 
.A(n_290),
.Y(n_1041)
);

INVx2_ASAP7_75t_L g1042 ( 
.A(n_625),
.Y(n_1042)
);

CKINVDCx20_ASAP7_75t_R g1043 ( 
.A(n_745),
.Y(n_1043)
);

INVx1_ASAP7_75t_L g1044 ( 
.A(n_223),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_186),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_672),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_626),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_271),
.Y(n_1048)
);

INVx2_ASAP7_75t_L g1049 ( 
.A(n_184),
.Y(n_1049)
);

CKINVDCx5p33_ASAP7_75t_R g1050 ( 
.A(n_717),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_44),
.Y(n_1051)
);

CKINVDCx5p33_ASAP7_75t_R g1052 ( 
.A(n_654),
.Y(n_1052)
);

CKINVDCx5p33_ASAP7_75t_R g1053 ( 
.A(n_419),
.Y(n_1053)
);

CKINVDCx20_ASAP7_75t_R g1054 ( 
.A(n_661),
.Y(n_1054)
);

CKINVDCx5p33_ASAP7_75t_R g1055 ( 
.A(n_674),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_359),
.Y(n_1056)
);

CKINVDCx5p33_ASAP7_75t_R g1057 ( 
.A(n_517),
.Y(n_1057)
);

CKINVDCx5p33_ASAP7_75t_R g1058 ( 
.A(n_178),
.Y(n_1058)
);

BUFx3_ASAP7_75t_L g1059 ( 
.A(n_682),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_47),
.Y(n_1060)
);

INVx2_ASAP7_75t_SL g1061 ( 
.A(n_264),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_720),
.Y(n_1062)
);

INVx1_ASAP7_75t_L g1063 ( 
.A(n_241),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_656),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_412),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_390),
.Y(n_1066)
);

CKINVDCx5p33_ASAP7_75t_R g1067 ( 
.A(n_117),
.Y(n_1067)
);

INVx1_ASAP7_75t_L g1068 ( 
.A(n_115),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_296),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_139),
.Y(n_1070)
);

INVx1_ASAP7_75t_L g1071 ( 
.A(n_428),
.Y(n_1071)
);

INVx1_ASAP7_75t_L g1072 ( 
.A(n_197),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_786),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_321),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_684),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_164),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_707),
.Y(n_1077)
);

INVx2_ASAP7_75t_L g1078 ( 
.A(n_335),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_20),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_300),
.Y(n_1080)
);

INVx1_ASAP7_75t_L g1081 ( 
.A(n_808),
.Y(n_1081)
);

CKINVDCx5p33_ASAP7_75t_R g1082 ( 
.A(n_512),
.Y(n_1082)
);

INVx2_ASAP7_75t_SL g1083 ( 
.A(n_405),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_396),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_314),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_791),
.Y(n_1086)
);

BUFx6f_ASAP7_75t_L g1087 ( 
.A(n_31),
.Y(n_1087)
);

CKINVDCx5p33_ASAP7_75t_R g1088 ( 
.A(n_694),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_408),
.Y(n_1089)
);

CKINVDCx16_ASAP7_75t_R g1090 ( 
.A(n_406),
.Y(n_1090)
);

INVx1_ASAP7_75t_L g1091 ( 
.A(n_532),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_703),
.Y(n_1092)
);

CKINVDCx5p33_ASAP7_75t_R g1093 ( 
.A(n_630),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_107),
.Y(n_1094)
);

BUFx10_ASAP7_75t_L g1095 ( 
.A(n_561),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_757),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_552),
.Y(n_1097)
);

CKINVDCx5p33_ASAP7_75t_R g1098 ( 
.A(n_545),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_695),
.Y(n_1099)
);

INVx1_ASAP7_75t_L g1100 ( 
.A(n_279),
.Y(n_1100)
);

INVx1_ASAP7_75t_L g1101 ( 
.A(n_696),
.Y(n_1101)
);

CKINVDCx5p33_ASAP7_75t_R g1102 ( 
.A(n_82),
.Y(n_1102)
);

CKINVDCx5p33_ASAP7_75t_R g1103 ( 
.A(n_355),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_701),
.Y(n_1104)
);

CKINVDCx20_ASAP7_75t_R g1105 ( 
.A(n_510),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_436),
.Y(n_1106)
);

INVx2_ASAP7_75t_SL g1107 ( 
.A(n_89),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_217),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_798),
.Y(n_1109)
);

CKINVDCx20_ASAP7_75t_R g1110 ( 
.A(n_58),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_218),
.Y(n_1111)
);

BUFx3_ASAP7_75t_L g1112 ( 
.A(n_668),
.Y(n_1112)
);

CKINVDCx5p33_ASAP7_75t_R g1113 ( 
.A(n_685),
.Y(n_1113)
);

HB1xp67_ASAP7_75t_L g1114 ( 
.A(n_516),
.Y(n_1114)
);

CKINVDCx5p33_ASAP7_75t_R g1115 ( 
.A(n_327),
.Y(n_1115)
);

CKINVDCx20_ASAP7_75t_R g1116 ( 
.A(n_11),
.Y(n_1116)
);

INVx1_ASAP7_75t_SL g1117 ( 
.A(n_471),
.Y(n_1117)
);

CKINVDCx5p33_ASAP7_75t_R g1118 ( 
.A(n_530),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_573),
.Y(n_1119)
);

INVx1_ASAP7_75t_L g1120 ( 
.A(n_308),
.Y(n_1120)
);

INVx1_ASAP7_75t_SL g1121 ( 
.A(n_536),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_142),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_562),
.Y(n_1123)
);

BUFx2_ASAP7_75t_L g1124 ( 
.A(n_243),
.Y(n_1124)
);

CKINVDCx5p33_ASAP7_75t_R g1125 ( 
.A(n_45),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_692),
.Y(n_1126)
);

CKINVDCx5p33_ASAP7_75t_R g1127 ( 
.A(n_704),
.Y(n_1127)
);

BUFx5_ASAP7_75t_L g1128 ( 
.A(n_612),
.Y(n_1128)
);

INVx2_ASAP7_75t_L g1129 ( 
.A(n_296),
.Y(n_1129)
);

INVx1_ASAP7_75t_L g1130 ( 
.A(n_502),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_422),
.Y(n_1131)
);

CKINVDCx20_ASAP7_75t_R g1132 ( 
.A(n_510),
.Y(n_1132)
);

CKINVDCx5p33_ASAP7_75t_R g1133 ( 
.A(n_71),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_687),
.Y(n_1134)
);

INVx1_ASAP7_75t_L g1135 ( 
.A(n_681),
.Y(n_1135)
);

CKINVDCx5p33_ASAP7_75t_R g1136 ( 
.A(n_389),
.Y(n_1136)
);

BUFx2_ASAP7_75t_L g1137 ( 
.A(n_190),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_526),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_156),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_93),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_134),
.Y(n_1141)
);

INVx1_ASAP7_75t_L g1142 ( 
.A(n_658),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_196),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_310),
.Y(n_1144)
);

CKINVDCx5p33_ASAP7_75t_R g1145 ( 
.A(n_704),
.Y(n_1145)
);

CKINVDCx5p33_ASAP7_75t_R g1146 ( 
.A(n_621),
.Y(n_1146)
);

INVx2_ASAP7_75t_L g1147 ( 
.A(n_716),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_614),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_4),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_456),
.Y(n_1150)
);

INVx1_ASAP7_75t_L g1151 ( 
.A(n_784),
.Y(n_1151)
);

INVx1_ASAP7_75t_L g1152 ( 
.A(n_433),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_376),
.Y(n_1153)
);

CKINVDCx5p33_ASAP7_75t_R g1154 ( 
.A(n_655),
.Y(n_1154)
);

INVx1_ASAP7_75t_L g1155 ( 
.A(n_523),
.Y(n_1155)
);

INVx1_ASAP7_75t_L g1156 ( 
.A(n_126),
.Y(n_1156)
);

CKINVDCx16_ASAP7_75t_R g1157 ( 
.A(n_121),
.Y(n_1157)
);

INVxp67_ASAP7_75t_SL g1158 ( 
.A(n_416),
.Y(n_1158)
);

CKINVDCx20_ASAP7_75t_R g1159 ( 
.A(n_161),
.Y(n_1159)
);

INVx2_ASAP7_75t_L g1160 ( 
.A(n_679),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_794),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_131),
.Y(n_1162)
);

CKINVDCx20_ASAP7_75t_R g1163 ( 
.A(n_139),
.Y(n_1163)
);

CKINVDCx16_ASAP7_75t_R g1164 ( 
.A(n_170),
.Y(n_1164)
);

CKINVDCx5p33_ASAP7_75t_R g1165 ( 
.A(n_720),
.Y(n_1165)
);

CKINVDCx20_ASAP7_75t_R g1166 ( 
.A(n_388),
.Y(n_1166)
);

CKINVDCx5p33_ASAP7_75t_R g1167 ( 
.A(n_226),
.Y(n_1167)
);

INVx1_ASAP7_75t_L g1168 ( 
.A(n_198),
.Y(n_1168)
);

CKINVDCx5p33_ASAP7_75t_R g1169 ( 
.A(n_288),
.Y(n_1169)
);

CKINVDCx5p33_ASAP7_75t_R g1170 ( 
.A(n_35),
.Y(n_1170)
);

INVx1_ASAP7_75t_L g1171 ( 
.A(n_724),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_671),
.Y(n_1172)
);

INVx1_ASAP7_75t_L g1173 ( 
.A(n_594),
.Y(n_1173)
);

BUFx2_ASAP7_75t_L g1174 ( 
.A(n_814),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_371),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_101),
.Y(n_1176)
);

INVx1_ASAP7_75t_L g1177 ( 
.A(n_722),
.Y(n_1177)
);

CKINVDCx14_ASAP7_75t_R g1178 ( 
.A(n_190),
.Y(n_1178)
);

INVx1_ASAP7_75t_L g1179 ( 
.A(n_252),
.Y(n_1179)
);

INVx1_ASAP7_75t_L g1180 ( 
.A(n_423),
.Y(n_1180)
);

CKINVDCx5p33_ASAP7_75t_R g1181 ( 
.A(n_151),
.Y(n_1181)
);

CKINVDCx20_ASAP7_75t_R g1182 ( 
.A(n_146),
.Y(n_1182)
);

CKINVDCx5p33_ASAP7_75t_R g1183 ( 
.A(n_674),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_349),
.Y(n_1184)
);

INVx1_ASAP7_75t_L g1185 ( 
.A(n_64),
.Y(n_1185)
);

CKINVDCx16_ASAP7_75t_R g1186 ( 
.A(n_150),
.Y(n_1186)
);

CKINVDCx16_ASAP7_75t_R g1187 ( 
.A(n_740),
.Y(n_1187)
);

INVx1_ASAP7_75t_L g1188 ( 
.A(n_41),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_189),
.Y(n_1189)
);

INVx1_ASAP7_75t_L g1190 ( 
.A(n_384),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_230),
.Y(n_1191)
);

BUFx2_ASAP7_75t_L g1192 ( 
.A(n_325),
.Y(n_1192)
);

CKINVDCx5p33_ASAP7_75t_R g1193 ( 
.A(n_730),
.Y(n_1193)
);

INVx1_ASAP7_75t_L g1194 ( 
.A(n_191),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_702),
.Y(n_1195)
);

CKINVDCx20_ASAP7_75t_R g1196 ( 
.A(n_370),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_664),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_93),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_669),
.Y(n_1199)
);

BUFx2_ASAP7_75t_L g1200 ( 
.A(n_314),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_407),
.Y(n_1201)
);

CKINVDCx5p33_ASAP7_75t_R g1202 ( 
.A(n_739),
.Y(n_1202)
);

INVx1_ASAP7_75t_L g1203 ( 
.A(n_324),
.Y(n_1203)
);

BUFx10_ASAP7_75t_L g1204 ( 
.A(n_663),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_425),
.Y(n_1205)
);

CKINVDCx5p33_ASAP7_75t_R g1206 ( 
.A(n_95),
.Y(n_1206)
);

CKINVDCx5p33_ASAP7_75t_R g1207 ( 
.A(n_89),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_598),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_446),
.Y(n_1209)
);

CKINVDCx20_ASAP7_75t_R g1210 ( 
.A(n_624),
.Y(n_1210)
);

INVx1_ASAP7_75t_L g1211 ( 
.A(n_9),
.Y(n_1211)
);

CKINVDCx5p33_ASAP7_75t_R g1212 ( 
.A(n_236),
.Y(n_1212)
);

CKINVDCx5p33_ASAP7_75t_R g1213 ( 
.A(n_127),
.Y(n_1213)
);

HB1xp67_ASAP7_75t_L g1214 ( 
.A(n_193),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_85),
.Y(n_1215)
);

BUFx2_ASAP7_75t_SL g1216 ( 
.A(n_770),
.Y(n_1216)
);

CKINVDCx20_ASAP7_75t_R g1217 ( 
.A(n_718),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_112),
.Y(n_1218)
);

CKINVDCx5p33_ASAP7_75t_R g1219 ( 
.A(n_767),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_494),
.Y(n_1220)
);

CKINVDCx20_ASAP7_75t_R g1221 ( 
.A(n_255),
.Y(n_1221)
);

INVx1_ASAP7_75t_SL g1222 ( 
.A(n_681),
.Y(n_1222)
);

CKINVDCx5p33_ASAP7_75t_R g1223 ( 
.A(n_666),
.Y(n_1223)
);

INVx1_ASAP7_75t_L g1224 ( 
.A(n_591),
.Y(n_1224)
);

CKINVDCx5p33_ASAP7_75t_R g1225 ( 
.A(n_447),
.Y(n_1225)
);

CKINVDCx5p33_ASAP7_75t_R g1226 ( 
.A(n_173),
.Y(n_1226)
);

INVx1_ASAP7_75t_L g1227 ( 
.A(n_512),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_204),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_81),
.Y(n_1229)
);

INVx1_ASAP7_75t_L g1230 ( 
.A(n_79),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_683),
.Y(n_1231)
);

CKINVDCx5p33_ASAP7_75t_R g1232 ( 
.A(n_290),
.Y(n_1232)
);

BUFx2_ASAP7_75t_L g1233 ( 
.A(n_406),
.Y(n_1233)
);

BUFx6f_ASAP7_75t_L g1234 ( 
.A(n_511),
.Y(n_1234)
);

CKINVDCx5p33_ASAP7_75t_R g1235 ( 
.A(n_736),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_796),
.Y(n_1236)
);

CKINVDCx5p33_ASAP7_75t_R g1237 ( 
.A(n_631),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_351),
.Y(n_1238)
);

BUFx2_ASAP7_75t_L g1239 ( 
.A(n_654),
.Y(n_1239)
);

INVx1_ASAP7_75t_L g1240 ( 
.A(n_204),
.Y(n_1240)
);

BUFx3_ASAP7_75t_L g1241 ( 
.A(n_638),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_381),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_128),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_182),
.Y(n_1244)
);

NOR2xp67_ASAP7_75t_L g1245 ( 
.A(n_629),
.B(n_726),
.Y(n_1245)
);

INVx1_ASAP7_75t_L g1246 ( 
.A(n_63),
.Y(n_1246)
);

INVx1_ASAP7_75t_L g1247 ( 
.A(n_124),
.Y(n_1247)
);

CKINVDCx5p33_ASAP7_75t_R g1248 ( 
.A(n_705),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_631),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_602),
.Y(n_1250)
);

CKINVDCx5p33_ASAP7_75t_R g1251 ( 
.A(n_613),
.Y(n_1251)
);

BUFx3_ASAP7_75t_L g1252 ( 
.A(n_155),
.Y(n_1252)
);

CKINVDCx20_ASAP7_75t_R g1253 ( 
.A(n_275),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_577),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_687),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_689),
.Y(n_1256)
);

CKINVDCx5p33_ASAP7_75t_R g1257 ( 
.A(n_688),
.Y(n_1257)
);

BUFx10_ASAP7_75t_L g1258 ( 
.A(n_199),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_488),
.Y(n_1259)
);

INVx1_ASAP7_75t_SL g1260 ( 
.A(n_685),
.Y(n_1260)
);

CKINVDCx5p33_ASAP7_75t_R g1261 ( 
.A(n_411),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_670),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_69),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_86),
.Y(n_1264)
);

AND2x2_ASAP7_75t_L g1265 ( 
.A(n_989),
.B(n_1178),
.Y(n_1265)
);

BUFx12f_ASAP7_75t_L g1266 ( 
.A(n_821),
.Y(n_1266)
);

INVx2_ASAP7_75t_L g1267 ( 
.A(n_1128),
.Y(n_1267)
);

INVx2_ASAP7_75t_L g1268 ( 
.A(n_1128),
.Y(n_1268)
);

AND2x4_ASAP7_75t_L g1269 ( 
.A(n_1010),
.B(n_830),
.Y(n_1269)
);

AND2x2_ASAP7_75t_L g1270 ( 
.A(n_989),
.B(n_0),
.Y(n_1270)
);

AND2x4_ASAP7_75t_L g1271 ( 
.A(n_1010),
.B(n_1),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_1010),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_1128),
.Y(n_1273)
);

HB1xp67_ASAP7_75t_L g1274 ( 
.A(n_842),
.Y(n_1274)
);

BUFx12f_ASAP7_75t_L g1275 ( 
.A(n_821),
.Y(n_1275)
);

INVx1_ASAP7_75t_L g1276 ( 
.A(n_1128),
.Y(n_1276)
);

AND2x2_ASAP7_75t_L g1277 ( 
.A(n_1178),
.B(n_1),
.Y(n_1277)
);

BUFx6f_ASAP7_75t_L g1278 ( 
.A(n_816),
.Y(n_1278)
);

BUFx6f_ASAP7_75t_L g1279 ( 
.A(n_816),
.Y(n_1279)
);

AND2x2_ASAP7_75t_L g1280 ( 
.A(n_861),
.B(n_2),
.Y(n_1280)
);

BUFx6f_ASAP7_75t_L g1281 ( 
.A(n_816),
.Y(n_1281)
);

INVx4_ASAP7_75t_L g1282 ( 
.A(n_1174),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_821),
.Y(n_1283)
);

HB1xp67_ASAP7_75t_L g1284 ( 
.A(n_976),
.Y(n_1284)
);

INVx1_ASAP7_75t_L g1285 ( 
.A(n_1019),
.Y(n_1285)
);

NAND2xp5_ASAP7_75t_L g1286 ( 
.A(n_892),
.B(n_5),
.Y(n_1286)
);

INVx1_ASAP7_75t_L g1287 ( 
.A(n_830),
.Y(n_1287)
);

NAND2xp5_ASAP7_75t_L g1288 ( 
.A(n_986),
.B(n_5),
.Y(n_1288)
);

INVx1_ASAP7_75t_L g1289 ( 
.A(n_1128),
.Y(n_1289)
);

BUFx3_ASAP7_75t_L g1290 ( 
.A(n_934),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_1128),
.Y(n_1291)
);

AND2x4_ASAP7_75t_L g1292 ( 
.A(n_857),
.B(n_2),
.Y(n_1292)
);

OAI21x1_ASAP7_75t_L g1293 ( 
.A1(n_869),
.A2(n_758),
.B(n_756),
.Y(n_1293)
);

INVx2_ASAP7_75t_L g1294 ( 
.A(n_1128),
.Y(n_1294)
);

OAI22x1_ASAP7_75t_L g1295 ( 
.A1(n_858),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1295)
);

INVx1_ASAP7_75t_L g1296 ( 
.A(n_846),
.Y(n_1296)
);

INVx2_ASAP7_75t_L g1297 ( 
.A(n_827),
.Y(n_1297)
);

BUFx12f_ASAP7_75t_L g1298 ( 
.A(n_966),
.Y(n_1298)
);

CKINVDCx5p33_ASAP7_75t_R g1299 ( 
.A(n_938),
.Y(n_1299)
);

INVx2_ASAP7_75t_L g1300 ( 
.A(n_827),
.Y(n_1300)
);

BUFx6f_ASAP7_75t_L g1301 ( 
.A(n_816),
.Y(n_1301)
);

AND2x6_ASAP7_75t_L g1302 ( 
.A(n_934),
.B(n_811),
.Y(n_1302)
);

INVx2_ASAP7_75t_L g1303 ( 
.A(n_865),
.Y(n_1303)
);

BUFx8_ASAP7_75t_SL g1304 ( 
.A(n_828),
.Y(n_1304)
);

INVx1_ASAP7_75t_L g1305 ( 
.A(n_846),
.Y(n_1305)
);

INVx1_ASAP7_75t_L g1306 ( 
.A(n_882),
.Y(n_1306)
);

INVx1_ASAP7_75t_L g1307 ( 
.A(n_882),
.Y(n_1307)
);

INVx1_ASAP7_75t_L g1308 ( 
.A(n_967),
.Y(n_1308)
);

OAI21x1_ASAP7_75t_L g1309 ( 
.A1(n_903),
.A2(n_760),
.B(n_759),
.Y(n_1309)
);

INVx2_ASAP7_75t_L g1310 ( 
.A(n_865),
.Y(n_1310)
);

OAI22x1_ASAP7_75t_L g1311 ( 
.A1(n_858),
.A2(n_8),
.B1(n_6),
.B2(n_7),
.Y(n_1311)
);

AND2x4_ASAP7_75t_L g1312 ( 
.A(n_857),
.B(n_9),
.Y(n_1312)
);

CKINVDCx5p33_ASAP7_75t_R g1313 ( 
.A(n_938),
.Y(n_1313)
);

INVx4_ASAP7_75t_L g1314 ( 
.A(n_900),
.Y(n_1314)
);

INVx3_ASAP7_75t_L g1315 ( 
.A(n_966),
.Y(n_1315)
);

OAI22x1_ASAP7_75t_R g1316 ( 
.A1(n_828),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1316)
);

INVx3_ASAP7_75t_L g1317 ( 
.A(n_966),
.Y(n_1317)
);

BUFx6f_ASAP7_75t_L g1318 ( 
.A(n_826),
.Y(n_1318)
);

INVx1_ASAP7_75t_L g1319 ( 
.A(n_991),
.Y(n_1319)
);

INVx2_ASAP7_75t_L g1320 ( 
.A(n_871),
.Y(n_1320)
);

BUFx6f_ASAP7_75t_L g1321 ( 
.A(n_826),
.Y(n_1321)
);

INVx3_ASAP7_75t_L g1322 ( 
.A(n_1007),
.Y(n_1322)
);

NAND2xp5_ASAP7_75t_L g1323 ( 
.A(n_1124),
.B(n_12),
.Y(n_1323)
);

BUFx8_ASAP7_75t_SL g1324 ( 
.A(n_854),
.Y(n_1324)
);

BUFx6f_ASAP7_75t_L g1325 ( 
.A(n_826),
.Y(n_1325)
);

BUFx2_ASAP7_75t_L g1326 ( 
.A(n_1137),
.Y(n_1326)
);

BUFx8_ASAP7_75t_SL g1327 ( 
.A(n_854),
.Y(n_1327)
);

BUFx3_ASAP7_75t_L g1328 ( 
.A(n_871),
.Y(n_1328)
);

AND2x6_ASAP7_75t_L g1329 ( 
.A(n_906),
.B(n_801),
.Y(n_1329)
);

INVx2_ASAP7_75t_L g1330 ( 
.A(n_891),
.Y(n_1330)
);

AOI22xp5_ASAP7_75t_SL g1331 ( 
.A1(n_878),
.A2(n_14),
.B1(n_10),
.B2(n_13),
.Y(n_1331)
);

AOI22xp5_ASAP7_75t_L g1332 ( 
.A1(n_991),
.A2(n_15),
.B1(n_13),
.B2(n_14),
.Y(n_1332)
);

BUFx6f_ASAP7_75t_L g1333 ( 
.A(n_905),
.Y(n_1333)
);

INVx2_ASAP7_75t_L g1334 ( 
.A(n_891),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_967),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_977),
.Y(n_1336)
);

BUFx12f_ASAP7_75t_L g1337 ( 
.A(n_1007),
.Y(n_1337)
);

INVx1_ASAP7_75t_L g1338 ( 
.A(n_1061),
.Y(n_1338)
);

INVx3_ASAP7_75t_L g1339 ( 
.A(n_1007),
.Y(n_1339)
);

OAI21x1_ASAP7_75t_L g1340 ( 
.A1(n_917),
.A2(n_762),
.B(n_761),
.Y(n_1340)
);

INVx4_ASAP7_75t_L g1341 ( 
.A(n_928),
.Y(n_1341)
);

INVx3_ASAP7_75t_L g1342 ( 
.A(n_1095),
.Y(n_1342)
);

INVx5_ASAP7_75t_L g1343 ( 
.A(n_905),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_905),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1061),
.Y(n_1345)
);

CKINVDCx5p33_ASAP7_75t_R g1346 ( 
.A(n_1161),
.Y(n_1346)
);

BUFx6f_ASAP7_75t_L g1347 ( 
.A(n_905),
.Y(n_1347)
);

BUFx6f_ASAP7_75t_L g1348 ( 
.A(n_941),
.Y(n_1348)
);

NOR2xp33_ASAP7_75t_L g1349 ( 
.A(n_954),
.B(n_15),
.Y(n_1349)
);

INVx2_ASAP7_75t_L g1350 ( 
.A(n_936),
.Y(n_1350)
);

BUFx3_ASAP7_75t_L g1351 ( 
.A(n_936),
.Y(n_1351)
);

INVx1_ASAP7_75t_L g1352 ( 
.A(n_1083),
.Y(n_1352)
);

INVx3_ASAP7_75t_L g1353 ( 
.A(n_1095),
.Y(n_1353)
);

OA21x2_ASAP7_75t_L g1354 ( 
.A1(n_1073),
.A2(n_765),
.B(n_763),
.Y(n_1354)
);

BUFx12f_ASAP7_75t_L g1355 ( 
.A(n_1095),
.Y(n_1355)
);

OAI21x1_ASAP7_75t_L g1356 ( 
.A1(n_1081),
.A2(n_769),
.B(n_766),
.Y(n_1356)
);

AND2x2_ASAP7_75t_L g1357 ( 
.A(n_1192),
.B(n_16),
.Y(n_1357)
);

BUFx6f_ASAP7_75t_L g1358 ( 
.A(n_941),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_1083),
.Y(n_1359)
);

NOR2xp33_ASAP7_75t_SL g1360 ( 
.A(n_935),
.B(n_788),
.Y(n_1360)
);

INVx2_ASAP7_75t_L g1361 ( 
.A(n_945),
.Y(n_1361)
);

BUFx6f_ASAP7_75t_L g1362 ( 
.A(n_941),
.Y(n_1362)
);

INVx1_ASAP7_75t_L g1363 ( 
.A(n_1037),
.Y(n_1363)
);

HB1xp67_ASAP7_75t_L g1364 ( 
.A(n_1114),
.Y(n_1364)
);

INVx3_ASAP7_75t_L g1365 ( 
.A(n_1204),
.Y(n_1365)
);

AND2x6_ASAP7_75t_L g1366 ( 
.A(n_1151),
.B(n_789),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_1161),
.Y(n_1367)
);

BUFx6f_ASAP7_75t_L g1368 ( 
.A(n_941),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_1042),
.Y(n_1369)
);

AOI22xp5_ASAP7_75t_L g1370 ( 
.A1(n_1107),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1370)
);

INVx2_ASAP7_75t_L g1371 ( 
.A(n_945),
.Y(n_1371)
);

BUFx6f_ASAP7_75t_L g1372 ( 
.A(n_973),
.Y(n_1372)
);

CKINVDCx5p33_ASAP7_75t_R g1373 ( 
.A(n_1299),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_1313),
.Y(n_1374)
);

AND2x2_ASAP7_75t_L g1375 ( 
.A(n_1326),
.B(n_1200),
.Y(n_1375)
);

INVx1_ASAP7_75t_L g1376 ( 
.A(n_1271),
.Y(n_1376)
);

CKINVDCx5p33_ASAP7_75t_R g1377 ( 
.A(n_1346),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1328),
.Y(n_1378)
);

INVx1_ASAP7_75t_L g1379 ( 
.A(n_1271),
.Y(n_1379)
);

INVx1_ASAP7_75t_L g1380 ( 
.A(n_1292),
.Y(n_1380)
);

INVx1_ASAP7_75t_L g1381 ( 
.A(n_1292),
.Y(n_1381)
);

CKINVDCx5p33_ASAP7_75t_R g1382 ( 
.A(n_1367),
.Y(n_1382)
);

NAND2xp5_ASAP7_75t_SL g1383 ( 
.A(n_1265),
.B(n_971),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1351),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_1304),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_1324),
.Y(n_1386)
);

BUFx6f_ASAP7_75t_L g1387 ( 
.A(n_1278),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_1327),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_1266),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_1312),
.Y(n_1390)
);

CKINVDCx5p33_ASAP7_75t_R g1391 ( 
.A(n_1275),
.Y(n_1391)
);

AND2x2_ASAP7_75t_L g1392 ( 
.A(n_1274),
.B(n_1233),
.Y(n_1392)
);

CKINVDCx5p33_ASAP7_75t_R g1393 ( 
.A(n_1298),
.Y(n_1393)
);

INVx2_ASAP7_75t_L g1394 ( 
.A(n_1297),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_1337),
.Y(n_1395)
);

INVx8_ASAP7_75t_L g1396 ( 
.A(n_1355),
.Y(n_1396)
);

BUFx10_ASAP7_75t_L g1397 ( 
.A(n_1269),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_L g1398 ( 
.A(n_1282),
.B(n_1239),
.Y(n_1398)
);

CKINVDCx20_ASAP7_75t_R g1399 ( 
.A(n_1284),
.Y(n_1399)
);

INVx2_ASAP7_75t_L g1400 ( 
.A(n_1300),
.Y(n_1400)
);

INVx2_ASAP7_75t_L g1401 ( 
.A(n_1303),
.Y(n_1401)
);

INVx3_ASAP7_75t_L g1402 ( 
.A(n_1269),
.Y(n_1402)
);

INVx2_ASAP7_75t_L g1403 ( 
.A(n_1310),
.Y(n_1403)
);

INVx2_ASAP7_75t_L g1404 ( 
.A(n_1320),
.Y(n_1404)
);

INVx2_ASAP7_75t_L g1405 ( 
.A(n_1330),
.Y(n_1405)
);

NOR2xp33_ASAP7_75t_R g1406 ( 
.A(n_1283),
.B(n_1315),
.Y(n_1406)
);

INVx1_ASAP7_75t_L g1407 ( 
.A(n_1287),
.Y(n_1407)
);

CKINVDCx20_ASAP7_75t_R g1408 ( 
.A(n_1364),
.Y(n_1408)
);

NOR2xp67_ASAP7_75t_L g1409 ( 
.A(n_1283),
.B(n_1214),
.Y(n_1409)
);

INVx1_ASAP7_75t_L g1410 ( 
.A(n_1319),
.Y(n_1410)
);

AND2x2_ASAP7_75t_L g1411 ( 
.A(n_1282),
.B(n_831),
.Y(n_1411)
);

NAND2xp33_ASAP7_75t_R g1412 ( 
.A(n_1315),
.B(n_859),
.Y(n_1412)
);

CKINVDCx5p33_ASAP7_75t_R g1413 ( 
.A(n_1314),
.Y(n_1413)
);

INVx1_ASAP7_75t_L g1414 ( 
.A(n_1338),
.Y(n_1414)
);

CKINVDCx20_ASAP7_75t_R g1415 ( 
.A(n_1270),
.Y(n_1415)
);

INVx1_ASAP7_75t_L g1416 ( 
.A(n_1345),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_1314),
.Y(n_1417)
);

NAND2xp5_ASAP7_75t_L g1418 ( 
.A(n_1341),
.B(n_859),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_1341),
.Y(n_1419)
);

CKINVDCx5p33_ASAP7_75t_R g1420 ( 
.A(n_1317),
.Y(n_1420)
);

NOR2xp33_ASAP7_75t_R g1421 ( 
.A(n_1317),
.B(n_914),
.Y(n_1421)
);

CKINVDCx5p33_ASAP7_75t_R g1422 ( 
.A(n_1322),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_1322),
.Y(n_1423)
);

INVx2_ASAP7_75t_L g1424 ( 
.A(n_1334),
.Y(n_1424)
);

AOI22xp5_ASAP7_75t_L g1425 ( 
.A1(n_1285),
.A2(n_1090),
.B1(n_1157),
.B2(n_1015),
.Y(n_1425)
);

CKINVDCx5p33_ASAP7_75t_R g1426 ( 
.A(n_1339),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_1352),
.Y(n_1427)
);

INVxp33_ASAP7_75t_SL g1428 ( 
.A(n_1277),
.Y(n_1428)
);

BUFx6f_ASAP7_75t_L g1429 ( 
.A(n_1278),
.Y(n_1429)
);

INVx2_ASAP7_75t_L g1430 ( 
.A(n_1350),
.Y(n_1430)
);

BUFx2_ASAP7_75t_L g1431 ( 
.A(n_1342),
.Y(n_1431)
);

INVx1_ASAP7_75t_L g1432 ( 
.A(n_1359),
.Y(n_1432)
);

CKINVDCx5p33_ASAP7_75t_R g1433 ( 
.A(n_1342),
.Y(n_1433)
);

CKINVDCx5p33_ASAP7_75t_R g1434 ( 
.A(n_1353),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_R g1435 ( 
.A(n_1353),
.B(n_1365),
.Y(n_1435)
);

BUFx3_ASAP7_75t_L g1436 ( 
.A(n_1290),
.Y(n_1436)
);

CKINVDCx20_ASAP7_75t_R g1437 ( 
.A(n_1316),
.Y(n_1437)
);

CKINVDCx5p33_ASAP7_75t_R g1438 ( 
.A(n_1365),
.Y(n_1438)
);

INVxp67_ASAP7_75t_SL g1439 ( 
.A(n_1272),
.Y(n_1439)
);

INVx2_ASAP7_75t_L g1440 ( 
.A(n_1361),
.Y(n_1440)
);

INVx2_ASAP7_75t_L g1441 ( 
.A(n_1371),
.Y(n_1441)
);

CKINVDCx5p33_ASAP7_75t_R g1442 ( 
.A(n_1280),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1272),
.Y(n_1443)
);

AND3x2_ASAP7_75t_L g1444 ( 
.A(n_1360),
.B(n_1158),
.C(n_899),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_1273),
.Y(n_1445)
);

CKINVDCx5p33_ASAP7_75t_R g1446 ( 
.A(n_1357),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_1331),
.Y(n_1447)
);

INVxp67_ASAP7_75t_SL g1448 ( 
.A(n_1286),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_1288),
.Y(n_1449)
);

NOR2xp33_ASAP7_75t_R g1450 ( 
.A(n_1329),
.B(n_1164),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_1323),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_R g1452 ( 
.A(n_1329),
.B(n_1186),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_1295),
.Y(n_1453)
);

NOR2xp33_ASAP7_75t_L g1454 ( 
.A(n_1296),
.B(n_1022),
.Y(n_1454)
);

BUFx10_ASAP7_75t_L g1455 ( 
.A(n_1349),
.Y(n_1455)
);

INVx1_ASAP7_75t_L g1456 ( 
.A(n_1273),
.Y(n_1456)
);

INVx1_ASAP7_75t_L g1457 ( 
.A(n_1276),
.Y(n_1457)
);

CKINVDCx20_ASAP7_75t_R g1458 ( 
.A(n_1332),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_1311),
.Y(n_1459)
);

CKINVDCx5p33_ASAP7_75t_R g1460 ( 
.A(n_1370),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_1296),
.Y(n_1461)
);

INVx1_ASAP7_75t_L g1462 ( 
.A(n_1289),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_1289),
.Y(n_1463)
);

OAI21x1_ASAP7_75t_L g1464 ( 
.A1(n_1293),
.A2(n_1049),
.B(n_1042),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_1305),
.Y(n_1465)
);

CKINVDCx5p33_ASAP7_75t_R g1466 ( 
.A(n_1305),
.Y(n_1466)
);

INVx1_ASAP7_75t_L g1467 ( 
.A(n_1267),
.Y(n_1467)
);

INVx1_ASAP7_75t_L g1468 ( 
.A(n_1268),
.Y(n_1468)
);

NAND2xp5_ASAP7_75t_SL g1469 ( 
.A(n_1291),
.B(n_994),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_1306),
.Y(n_1470)
);

NOR2xp33_ASAP7_75t_R g1471 ( 
.A(n_1329),
.B(n_1187),
.Y(n_1471)
);

NOR2xp33_ASAP7_75t_R g1472 ( 
.A(n_1329),
.B(n_912),
.Y(n_1472)
);

CKINVDCx20_ASAP7_75t_R g1473 ( 
.A(n_1306),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_1307),
.Y(n_1474)
);

INVx1_ASAP7_75t_L g1475 ( 
.A(n_1294),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_1307),
.Y(n_1476)
);

INVx1_ASAP7_75t_L g1477 ( 
.A(n_1308),
.Y(n_1477)
);

HB1xp67_ASAP7_75t_L g1478 ( 
.A(n_1335),
.Y(n_1478)
);

CKINVDCx20_ASAP7_75t_R g1479 ( 
.A(n_1336),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_1336),
.Y(n_1480)
);

NOR2xp33_ASAP7_75t_R g1481 ( 
.A(n_1366),
.B(n_912),
.Y(n_1481)
);

NOR2xp67_ASAP7_75t_L g1482 ( 
.A(n_1363),
.B(n_1369),
.Y(n_1482)
);

BUFx6f_ASAP7_75t_L g1483 ( 
.A(n_1278),
.Y(n_1483)
);

CKINVDCx20_ASAP7_75t_R g1484 ( 
.A(n_1354),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_1343),
.Y(n_1485)
);

XNOR2xp5_ASAP7_75t_L g1486 ( 
.A(n_1309),
.B(n_878),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_1343),
.Y(n_1487)
);

INVx2_ASAP7_75t_L g1488 ( 
.A(n_1279),
.Y(n_1488)
);

CKINVDCx16_ASAP7_75t_R g1489 ( 
.A(n_1302),
.Y(n_1489)
);

INVx2_ASAP7_75t_L g1490 ( 
.A(n_1279),
.Y(n_1490)
);

CKINVDCx20_ASAP7_75t_R g1491 ( 
.A(n_1354),
.Y(n_1491)
);

CKINVDCx5p33_ASAP7_75t_R g1492 ( 
.A(n_1302),
.Y(n_1492)
);

INVx3_ASAP7_75t_L g1493 ( 
.A(n_1340),
.Y(n_1493)
);

NOR2xp33_ASAP7_75t_R g1494 ( 
.A(n_1366),
.B(n_1086),
.Y(n_1494)
);

INVx2_ASAP7_75t_L g1495 ( 
.A(n_1279),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_1302),
.Y(n_1496)
);

CKINVDCx5p33_ASAP7_75t_R g1497 ( 
.A(n_1302),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_1366),
.Y(n_1498)
);

INVx1_ASAP7_75t_L g1499 ( 
.A(n_1356),
.Y(n_1499)
);

CKINVDCx5p33_ASAP7_75t_R g1500 ( 
.A(n_1281),
.Y(n_1500)
);

INVx2_ASAP7_75t_L g1501 ( 
.A(n_1281),
.Y(n_1501)
);

NOR2x1p5_ASAP7_75t_L g1502 ( 
.A(n_1281),
.B(n_860),
.Y(n_1502)
);

NOR2xp33_ASAP7_75t_R g1503 ( 
.A(n_1301),
.B(n_863),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_1301),
.Y(n_1504)
);

INVx2_ASAP7_75t_L g1505 ( 
.A(n_1301),
.Y(n_1505)
);

CKINVDCx16_ASAP7_75t_R g1506 ( 
.A(n_1318),
.Y(n_1506)
);

CKINVDCx5p33_ASAP7_75t_R g1507 ( 
.A(n_1318),
.Y(n_1507)
);

CKINVDCx5p33_ASAP7_75t_R g1508 ( 
.A(n_1318),
.Y(n_1508)
);

INVx1_ASAP7_75t_L g1509 ( 
.A(n_1321),
.Y(n_1509)
);

CKINVDCx5p33_ASAP7_75t_R g1510 ( 
.A(n_1321),
.Y(n_1510)
);

CKINVDCx5p33_ASAP7_75t_R g1511 ( 
.A(n_1321),
.Y(n_1511)
);

INVx2_ASAP7_75t_L g1512 ( 
.A(n_1325),
.Y(n_1512)
);

INVx3_ASAP7_75t_L g1513 ( 
.A(n_1325),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_1325),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_1333),
.Y(n_1515)
);

CKINVDCx20_ASAP7_75t_R g1516 ( 
.A(n_1333),
.Y(n_1516)
);

INVxp67_ASAP7_75t_L g1517 ( 
.A(n_1344),
.Y(n_1517)
);

INVx1_ASAP7_75t_L g1518 ( 
.A(n_1344),
.Y(n_1518)
);

CKINVDCx20_ASAP7_75t_R g1519 ( 
.A(n_1344),
.Y(n_1519)
);

INVx1_ASAP7_75t_L g1520 ( 
.A(n_1347),
.Y(n_1520)
);

CKINVDCx20_ASAP7_75t_R g1521 ( 
.A(n_1347),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_1347),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_1348),
.Y(n_1523)
);

INVx2_ASAP7_75t_L g1524 ( 
.A(n_1348),
.Y(n_1524)
);

INVx2_ASAP7_75t_L g1525 ( 
.A(n_1348),
.Y(n_1525)
);

INVx2_ASAP7_75t_L g1526 ( 
.A(n_1358),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_1358),
.Y(n_1527)
);

INVx1_ASAP7_75t_L g1528 ( 
.A(n_1358),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_1362),
.Y(n_1529)
);

CKINVDCx20_ASAP7_75t_R g1530 ( 
.A(n_1372),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_1372),
.Y(n_1531)
);

INVx3_ASAP7_75t_L g1532 ( 
.A(n_1362),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_1368),
.Y(n_1533)
);

AND2x2_ASAP7_75t_L g1534 ( 
.A(n_1368),
.B(n_1204),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1368),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1326),
.B(n_1204),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_1328),
.Y(n_1537)
);

CKINVDCx20_ASAP7_75t_R g1538 ( 
.A(n_1304),
.Y(n_1538)
);

HB1xp67_ASAP7_75t_L g1539 ( 
.A(n_1265),
.Y(n_1539)
);

CKINVDCx5p33_ASAP7_75t_R g1540 ( 
.A(n_1299),
.Y(n_1540)
);

CKINVDCx20_ASAP7_75t_R g1541 ( 
.A(n_1304),
.Y(n_1541)
);

CKINVDCx5p33_ASAP7_75t_R g1542 ( 
.A(n_1299),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_1299),
.Y(n_1543)
);

AO21x2_ASAP7_75t_L g1544 ( 
.A1(n_1293),
.A2(n_824),
.B(n_822),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_1299),
.Y(n_1545)
);

CKINVDCx5p33_ASAP7_75t_R g1546 ( 
.A(n_1299),
.Y(n_1546)
);

NAND2xp33_ASAP7_75t_R g1547 ( 
.A(n_1265),
.B(n_863),
.Y(n_1547)
);

CKINVDCx5p33_ASAP7_75t_R g1548 ( 
.A(n_1299),
.Y(n_1548)
);

CKINVDCx20_ASAP7_75t_R g1549 ( 
.A(n_1304),
.Y(n_1549)
);

CKINVDCx5p33_ASAP7_75t_R g1550 ( 
.A(n_1299),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_1299),
.Y(n_1551)
);

CKINVDCx20_ASAP7_75t_R g1552 ( 
.A(n_1304),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1328),
.Y(n_1553)
);

INVx1_ASAP7_75t_L g1554 ( 
.A(n_1402),
.Y(n_1554)
);

INVx2_ASAP7_75t_L g1555 ( 
.A(n_1394),
.Y(n_1555)
);

NAND3xp33_ASAP7_75t_L g1556 ( 
.A(n_1442),
.B(n_1056),
.C(n_866),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1448),
.B(n_1096),
.Y(n_1557)
);

INVx2_ASAP7_75t_L g1558 ( 
.A(n_1400),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_L g1559 ( 
.A(n_1448),
.B(n_1109),
.Y(n_1559)
);

NOR2xp33_ASAP7_75t_SL g1560 ( 
.A(n_1489),
.B(n_879),
.Y(n_1560)
);

NOR2xp33_ASAP7_75t_L g1561 ( 
.A(n_1402),
.B(n_840),
.Y(n_1561)
);

NAND2xp5_ASAP7_75t_SL g1562 ( 
.A(n_1450),
.B(n_1219),
.Y(n_1562)
);

NAND2xp5_ASAP7_75t_SL g1563 ( 
.A(n_1452),
.B(n_1236),
.Y(n_1563)
);

INVx2_ASAP7_75t_L g1564 ( 
.A(n_1401),
.Y(n_1564)
);

INVx2_ASAP7_75t_L g1565 ( 
.A(n_1403),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1478),
.Y(n_1566)
);

NAND2xp5_ASAP7_75t_L g1567 ( 
.A(n_1439),
.B(n_866),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1418),
.B(n_1216),
.Y(n_1568)
);

NOR2xp33_ASAP7_75t_SL g1569 ( 
.A(n_1396),
.B(n_879),
.Y(n_1569)
);

NAND2xp5_ASAP7_75t_SL g1570 ( 
.A(n_1471),
.B(n_973),
.Y(n_1570)
);

AO221x1_ASAP7_75t_L g1571 ( 
.A1(n_1399),
.A2(n_920),
.B1(n_943),
.B2(n_909),
.C(n_884),
.Y(n_1571)
);

NAND2xp5_ASAP7_75t_SL g1572 ( 
.A(n_1413),
.B(n_973),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_SL g1573 ( 
.A(n_1417),
.B(n_973),
.Y(n_1573)
);

NOR2xp33_ASAP7_75t_L g1574 ( 
.A(n_1431),
.B(n_817),
.Y(n_1574)
);

INVx1_ASAP7_75t_SL g1575 ( 
.A(n_1408),
.Y(n_1575)
);

INVx1_ASAP7_75t_L g1576 ( 
.A(n_1478),
.Y(n_1576)
);

INVx2_ASAP7_75t_L g1577 ( 
.A(n_1404),
.Y(n_1577)
);

INVx2_ASAP7_75t_L g1578 ( 
.A(n_1405),
.Y(n_1578)
);

AND2x2_ASAP7_75t_L g1579 ( 
.A(n_1392),
.B(n_1258),
.Y(n_1579)
);

BUFx3_ASAP7_75t_L g1580 ( 
.A(n_1396),
.Y(n_1580)
);

INVx2_ASAP7_75t_L g1581 ( 
.A(n_1424),
.Y(n_1581)
);

A2O1A1Ixp33_ASAP7_75t_L g1582 ( 
.A1(n_1380),
.A2(n_1059),
.B(n_1112),
.C(n_988),
.Y(n_1582)
);

NAND2xp5_ASAP7_75t_L g1583 ( 
.A(n_1461),
.B(n_1056),
.Y(n_1583)
);

NAND2xp5_ASAP7_75t_L g1584 ( 
.A(n_1465),
.B(n_1082),
.Y(n_1584)
);

INVx2_ASAP7_75t_L g1585 ( 
.A(n_1430),
.Y(n_1585)
);

NOR2xp33_ASAP7_75t_L g1586 ( 
.A(n_1397),
.B(n_819),
.Y(n_1586)
);

AND2x4_ASAP7_75t_L g1587 ( 
.A(n_1409),
.B(n_818),
.Y(n_1587)
);

NOR2xp33_ASAP7_75t_L g1588 ( 
.A(n_1397),
.B(n_820),
.Y(n_1588)
);

NAND2xp5_ASAP7_75t_L g1589 ( 
.A(n_1466),
.B(n_1082),
.Y(n_1589)
);

AOI22xp33_ASAP7_75t_L g1590 ( 
.A1(n_1381),
.A2(n_1059),
.B1(n_1112),
.B2(n_988),
.Y(n_1590)
);

INVx2_ASAP7_75t_SL g1591 ( 
.A(n_1396),
.Y(n_1591)
);

INVx1_ASAP7_75t_L g1592 ( 
.A(n_1407),
.Y(n_1592)
);

NAND2xp5_ASAP7_75t_L g1593 ( 
.A(n_1470),
.B(n_1085),
.Y(n_1593)
);

INVx1_ASAP7_75t_L g1594 ( 
.A(n_1410),
.Y(n_1594)
);

NOR2xp67_ASAP7_75t_L g1595 ( 
.A(n_1390),
.B(n_779),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1474),
.B(n_1085),
.Y(n_1596)
);

NAND2xp5_ASAP7_75t_L g1597 ( 
.A(n_1480),
.B(n_1232),
.Y(n_1597)
);

NOR2xp33_ASAP7_75t_L g1598 ( 
.A(n_1383),
.B(n_823),
.Y(n_1598)
);

BUFx6f_ASAP7_75t_L g1599 ( 
.A(n_1464),
.Y(n_1599)
);

NAND2xp5_ASAP7_75t_SL g1600 ( 
.A(n_1419),
.B(n_1472),
.Y(n_1600)
);

INVx3_ASAP7_75t_L g1601 ( 
.A(n_1534),
.Y(n_1601)
);

INVxp67_ASAP7_75t_SL g1602 ( 
.A(n_1473),
.Y(n_1602)
);

NAND2xp5_ASAP7_75t_SL g1603 ( 
.A(n_1481),
.B(n_1087),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1420),
.B(n_834),
.Y(n_1604)
);

BUFx6f_ASAP7_75t_L g1605 ( 
.A(n_1492),
.Y(n_1605)
);

INVx2_ASAP7_75t_L g1606 ( 
.A(n_1440),
.Y(n_1606)
);

BUFx2_ASAP7_75t_L g1607 ( 
.A(n_1479),
.Y(n_1607)
);

INVx8_ASAP7_75t_L g1608 ( 
.A(n_1422),
.Y(n_1608)
);

NOR2xp33_ASAP7_75t_L g1609 ( 
.A(n_1423),
.B(n_836),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_SL g1610 ( 
.A(n_1494),
.B(n_1087),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1426),
.B(n_837),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1414),
.Y(n_1612)
);

INVx1_ASAP7_75t_L g1613 ( 
.A(n_1416),
.Y(n_1613)
);

INVxp33_ASAP7_75t_L g1614 ( 
.A(n_1421),
.Y(n_1614)
);

NAND2xp5_ASAP7_75t_SL g1615 ( 
.A(n_1496),
.B(n_1087),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1398),
.B(n_1241),
.Y(n_1616)
);

NAND2xp5_ASAP7_75t_SL g1617 ( 
.A(n_1497),
.B(n_1087),
.Y(n_1617)
);

NOR2xp33_ASAP7_75t_L g1618 ( 
.A(n_1433),
.B(n_838),
.Y(n_1618)
);

NAND2xp5_ASAP7_75t_SL g1619 ( 
.A(n_1498),
.B(n_1234),
.Y(n_1619)
);

NOR2xp33_ASAP7_75t_L g1620 ( 
.A(n_1434),
.B(n_839),
.Y(n_1620)
);

NAND3xp33_ASAP7_75t_L g1621 ( 
.A(n_1446),
.B(n_847),
.C(n_844),
.Y(n_1621)
);

INVx2_ASAP7_75t_SL g1622 ( 
.A(n_1406),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1441),
.Y(n_1623)
);

NAND2xp5_ASAP7_75t_L g1624 ( 
.A(n_1376),
.B(n_1379),
.Y(n_1624)
);

INVx2_ASAP7_75t_SL g1625 ( 
.A(n_1435),
.Y(n_1625)
);

NOR2xp33_ASAP7_75t_L g1626 ( 
.A(n_1438),
.B(n_848),
.Y(n_1626)
);

INVx2_ASAP7_75t_L g1627 ( 
.A(n_1476),
.Y(n_1627)
);

NAND2xp5_ASAP7_75t_L g1628 ( 
.A(n_1449),
.B(n_1252),
.Y(n_1628)
);

INVx2_ASAP7_75t_L g1629 ( 
.A(n_1477),
.Y(n_1629)
);

INVx1_ASAP7_75t_L g1630 ( 
.A(n_1427),
.Y(n_1630)
);

INVx2_ASAP7_75t_SL g1631 ( 
.A(n_1502),
.Y(n_1631)
);

INVx2_ASAP7_75t_SL g1632 ( 
.A(n_1411),
.Y(n_1632)
);

INVx1_ASAP7_75t_SL g1633 ( 
.A(n_1415),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1432),
.Y(n_1634)
);

INVx2_ASAP7_75t_L g1635 ( 
.A(n_1378),
.Y(n_1635)
);

OR2x6_ASAP7_75t_L g1636 ( 
.A(n_1536),
.B(n_835),
.Y(n_1636)
);

INVx1_ASAP7_75t_L g1637 ( 
.A(n_1443),
.Y(n_1637)
);

NOR2xp33_ASAP7_75t_L g1638 ( 
.A(n_1455),
.B(n_850),
.Y(n_1638)
);

NAND2xp5_ASAP7_75t_L g1639 ( 
.A(n_1451),
.B(n_1252),
.Y(n_1639)
);

NAND2xp5_ASAP7_75t_L g1640 ( 
.A(n_1539),
.B(n_1428),
.Y(n_1640)
);

NOR2xp33_ASAP7_75t_L g1641 ( 
.A(n_1455),
.B(n_852),
.Y(n_1641)
);

INVx1_ASAP7_75t_SL g1642 ( 
.A(n_1373),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1482),
.Y(n_1643)
);

INVx2_ASAP7_75t_SL g1644 ( 
.A(n_1539),
.Y(n_1644)
);

INVx1_ASAP7_75t_L g1645 ( 
.A(n_1384),
.Y(n_1645)
);

INVx2_ASAP7_75t_SL g1646 ( 
.A(n_1375),
.Y(n_1646)
);

NOR2xp67_ASAP7_75t_L g1647 ( 
.A(n_1499),
.B(n_1486),
.Y(n_1647)
);

INVx1_ASAP7_75t_L g1648 ( 
.A(n_1537),
.Y(n_1648)
);

INVx2_ASAP7_75t_L g1649 ( 
.A(n_1553),
.Y(n_1649)
);

OR2x6_ASAP7_75t_L g1650 ( 
.A(n_1538),
.B(n_895),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1436),
.B(n_853),
.Y(n_1651)
);

AOI22xp5_ASAP7_75t_L g1652 ( 
.A1(n_1412),
.A2(n_1255),
.B1(n_1257),
.B2(n_1254),
.Y(n_1652)
);

NAND2xp5_ASAP7_75t_L g1653 ( 
.A(n_1454),
.B(n_855),
.Y(n_1653)
);

NOR2xp33_ASAP7_75t_L g1654 ( 
.A(n_1469),
.B(n_1454),
.Y(n_1654)
);

NOR2xp33_ASAP7_75t_L g1655 ( 
.A(n_1425),
.B(n_856),
.Y(n_1655)
);

NOR2xp33_ASAP7_75t_L g1656 ( 
.A(n_1389),
.B(n_867),
.Y(n_1656)
);

NOR2xp33_ASAP7_75t_L g1657 ( 
.A(n_1391),
.B(n_870),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1445),
.B(n_872),
.Y(n_1658)
);

AO221x1_ASAP7_75t_L g1659 ( 
.A1(n_1493),
.A2(n_920),
.B1(n_943),
.B2(n_909),
.C(n_884),
.Y(n_1659)
);

NOR3xp33_ASAP7_75t_L g1660 ( 
.A(n_1447),
.B(n_832),
.C(n_815),
.Y(n_1660)
);

NOR2xp67_ASAP7_75t_L g1661 ( 
.A(n_1493),
.B(n_780),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1456),
.B(n_876),
.Y(n_1662)
);

AOI22xp5_ASAP7_75t_L g1663 ( 
.A1(n_1460),
.A2(n_829),
.B1(n_833),
.B2(n_825),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1485),
.Y(n_1664)
);

BUFx5_ASAP7_75t_L g1665 ( 
.A(n_1467),
.Y(n_1665)
);

NAND2xp5_ASAP7_75t_SL g1666 ( 
.A(n_1506),
.B(n_1234),
.Y(n_1666)
);

NAND2xp5_ASAP7_75t_L g1667 ( 
.A(n_1457),
.B(n_881),
.Y(n_1667)
);

INVx1_ASAP7_75t_SL g1668 ( 
.A(n_1374),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1544),
.Y(n_1669)
);

NOR3xp33_ASAP7_75t_L g1670 ( 
.A(n_1453),
.B(n_849),
.C(n_843),
.Y(n_1670)
);

INVx1_ASAP7_75t_L g1671 ( 
.A(n_1487),
.Y(n_1671)
);

INVx8_ASAP7_75t_L g1672 ( 
.A(n_1393),
.Y(n_1672)
);

INVx2_ASAP7_75t_SL g1673 ( 
.A(n_1395),
.Y(n_1673)
);

BUFx6f_ASAP7_75t_L g1674 ( 
.A(n_1544),
.Y(n_1674)
);

NAND2xp5_ASAP7_75t_L g1675 ( 
.A(n_1462),
.B(n_1463),
.Y(n_1675)
);

NAND3xp33_ASAP7_75t_L g1676 ( 
.A(n_1547),
.B(n_894),
.C(n_893),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1377),
.B(n_898),
.Y(n_1677)
);

NOR2xp33_ASAP7_75t_L g1678 ( 
.A(n_1382),
.B(n_1540),
.Y(n_1678)
);

NAND2xp5_ASAP7_75t_L g1679 ( 
.A(n_1468),
.B(n_901),
.Y(n_1679)
);

INVx3_ASAP7_75t_L g1680 ( 
.A(n_1444),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1503),
.Y(n_1681)
);

HB1xp67_ASAP7_75t_L g1682 ( 
.A(n_1547),
.Y(n_1682)
);

INVx2_ASAP7_75t_L g1683 ( 
.A(n_1500),
.Y(n_1683)
);

INVxp67_ASAP7_75t_L g1684 ( 
.A(n_1542),
.Y(n_1684)
);

NAND3xp33_ASAP7_75t_L g1685 ( 
.A(n_1475),
.B(n_910),
.C(n_904),
.Y(n_1685)
);

INVx2_ASAP7_75t_SL g1686 ( 
.A(n_1444),
.Y(n_1686)
);

INVx1_ASAP7_75t_L g1687 ( 
.A(n_1516),
.Y(n_1687)
);

NAND2xp5_ASAP7_75t_L g1688 ( 
.A(n_1484),
.B(n_913),
.Y(n_1688)
);

NOR2xp33_ASAP7_75t_L g1689 ( 
.A(n_1543),
.B(n_915),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1519),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_SL g1691 ( 
.A(n_1545),
.B(n_1078),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1546),
.B(n_1078),
.Y(n_1692)
);

INVx4_ASAP7_75t_L g1693 ( 
.A(n_1504),
.Y(n_1693)
);

INVx2_ASAP7_75t_L g1694 ( 
.A(n_1507),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1508),
.Y(n_1695)
);

BUFx8_ASAP7_75t_L g1696 ( 
.A(n_1541),
.Y(n_1696)
);

NAND2xp5_ASAP7_75t_L g1697 ( 
.A(n_1491),
.B(n_919),
.Y(n_1697)
);

NAND2xp5_ASAP7_75t_L g1698 ( 
.A(n_1510),
.B(n_922),
.Y(n_1698)
);

NOR3xp33_ASAP7_75t_L g1699 ( 
.A(n_1459),
.B(n_930),
.C(n_918),
.Y(n_1699)
);

NOR2xp33_ASAP7_75t_L g1700 ( 
.A(n_1548),
.B(n_925),
.Y(n_1700)
);

INVx2_ASAP7_75t_L g1701 ( 
.A(n_1511),
.Y(n_1701)
);

NAND2xp5_ASAP7_75t_L g1702 ( 
.A(n_1514),
.B(n_927),
.Y(n_1702)
);

INVx2_ASAP7_75t_L g1703 ( 
.A(n_1515),
.Y(n_1703)
);

INVx2_ASAP7_75t_SL g1704 ( 
.A(n_1521),
.Y(n_1704)
);

NOR2xp67_ASAP7_75t_SL g1705 ( 
.A(n_1550),
.B(n_1261),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1530),
.Y(n_1706)
);

INVx5_ASAP7_75t_L g1707 ( 
.A(n_1513),
.Y(n_1707)
);

INVx2_ASAP7_75t_SL g1708 ( 
.A(n_1531),
.Y(n_1708)
);

AND2x2_ASAP7_75t_L g1709 ( 
.A(n_1551),
.B(n_1258),
.Y(n_1709)
);

CKINVDCx20_ASAP7_75t_R g1710 ( 
.A(n_1549),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1533),
.Y(n_1711)
);

INVx2_ASAP7_75t_L g1712 ( 
.A(n_1522),
.Y(n_1712)
);

AO221x1_ASAP7_75t_L g1713 ( 
.A1(n_1437),
.A2(n_969),
.B1(n_984),
.B2(n_961),
.C(n_957),
.Y(n_1713)
);

NOR2xp33_ASAP7_75t_L g1714 ( 
.A(n_1458),
.B(n_929),
.Y(n_1714)
);

NAND2xp33_ASAP7_75t_L g1715 ( 
.A(n_1523),
.B(n_933),
.Y(n_1715)
);

INVx2_ASAP7_75t_L g1716 ( 
.A(n_1527),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1529),
.B(n_939),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1517),
.B(n_940),
.Y(n_1718)
);

INVx2_ASAP7_75t_L g1719 ( 
.A(n_1517),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1532),
.B(n_942),
.Y(n_1720)
);

INVx2_ASAP7_75t_L g1721 ( 
.A(n_1532),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1385),
.B(n_946),
.Y(n_1722)
);

NOR3xp33_ASAP7_75t_L g1723 ( 
.A(n_1386),
.B(n_1388),
.C(n_964),
.Y(n_1723)
);

INVxp67_ASAP7_75t_L g1724 ( 
.A(n_1552),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1509),
.B(n_947),
.Y(n_1725)
);

INVxp33_ASAP7_75t_L g1726 ( 
.A(n_1387),
.Y(n_1726)
);

XOR2xp5_ASAP7_75t_L g1727 ( 
.A(n_1518),
.B(n_957),
.Y(n_1727)
);

NAND2xp5_ASAP7_75t_L g1728 ( 
.A(n_1520),
.B(n_949),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1528),
.B(n_950),
.Y(n_1729)
);

INVx1_ASAP7_75t_L g1730 ( 
.A(n_1535),
.Y(n_1730)
);

INVx1_ASAP7_75t_L g1731 ( 
.A(n_1488),
.Y(n_1731)
);

INVx2_ASAP7_75t_L g1732 ( 
.A(n_1490),
.Y(n_1732)
);

NAND2xp5_ASAP7_75t_L g1733 ( 
.A(n_1495),
.B(n_952),
.Y(n_1733)
);

XNOR2x2_ASAP7_75t_L g1734 ( 
.A(n_1501),
.B(n_932),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_L g1735 ( 
.A(n_1505),
.B(n_958),
.Y(n_1735)
);

NOR2xp33_ASAP7_75t_L g1736 ( 
.A(n_1526),
.B(n_960),
.Y(n_1736)
);

INVx2_ASAP7_75t_SL g1737 ( 
.A(n_1387),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_L g1738 ( 
.A(n_1512),
.B(n_963),
.Y(n_1738)
);

AND2x2_ASAP7_75t_L g1739 ( 
.A(n_1525),
.B(n_1258),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1524),
.B(n_968),
.Y(n_1740)
);

NOR2xp33_ASAP7_75t_L g1741 ( 
.A(n_1483),
.B(n_974),
.Y(n_1741)
);

NOR2xp67_ASAP7_75t_L g1742 ( 
.A(n_1387),
.B(n_781),
.Y(n_1742)
);

NOR3xp33_ASAP7_75t_L g1743 ( 
.A(n_1429),
.B(n_1013),
.C(n_979),
.Y(n_1743)
);

INVx1_ASAP7_75t_L g1744 ( 
.A(n_1429),
.Y(n_1744)
);

NAND2xp33_ASAP7_75t_L g1745 ( 
.A(n_1429),
.B(n_978),
.Y(n_1745)
);

OR2x2_ASAP7_75t_L g1746 ( 
.A(n_1429),
.B(n_1041),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1483),
.B(n_982),
.Y(n_1747)
);

INVx1_ASAP7_75t_L g1748 ( 
.A(n_1402),
.Y(n_1748)
);

NAND2xp5_ASAP7_75t_L g1749 ( 
.A(n_1448),
.B(n_983),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_L g1750 ( 
.A(n_1448),
.B(n_987),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_L g1751 ( 
.A(n_1448),
.B(n_990),
.Y(n_1751)
);

NOR2xp33_ASAP7_75t_L g1752 ( 
.A(n_1402),
.B(n_992),
.Y(n_1752)
);

AND2x2_ASAP7_75t_L g1753 ( 
.A(n_1392),
.B(n_997),
.Y(n_1753)
);

NOR3xp33_ASAP7_75t_L g1754 ( 
.A(n_1447),
.B(n_1121),
.C(n_1117),
.Y(n_1754)
);

INVx1_ASAP7_75t_L g1755 ( 
.A(n_1402),
.Y(n_1755)
);

BUFx8_ASAP7_75t_L g1756 ( 
.A(n_1411),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_SL g1757 ( 
.A(n_1450),
.B(n_1129),
.Y(n_1757)
);

INVx1_ASAP7_75t_L g1758 ( 
.A(n_1402),
.Y(n_1758)
);

INVx2_ASAP7_75t_L g1759 ( 
.A(n_1394),
.Y(n_1759)
);

NAND2xp5_ASAP7_75t_L g1760 ( 
.A(n_1448),
.B(n_1001),
.Y(n_1760)
);

NOR2xp33_ASAP7_75t_L g1761 ( 
.A(n_1402),
.B(n_1002),
.Y(n_1761)
);

NAND2xp5_ASAP7_75t_L g1762 ( 
.A(n_1448),
.B(n_1003),
.Y(n_1762)
);

INVx2_ASAP7_75t_SL g1763 ( 
.A(n_1397),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1402),
.B(n_1004),
.Y(n_1764)
);

INVxp67_ASAP7_75t_L g1765 ( 
.A(n_1412),
.Y(n_1765)
);

NAND2xp33_ASAP7_75t_L g1766 ( 
.A(n_1492),
.B(n_1005),
.Y(n_1766)
);

NAND2xp5_ASAP7_75t_SL g1767 ( 
.A(n_1450),
.B(n_1147),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1448),
.B(n_1008),
.Y(n_1768)
);

NOR2xp33_ASAP7_75t_L g1769 ( 
.A(n_1402),
.B(n_1009),
.Y(n_1769)
);

NOR2xp33_ASAP7_75t_L g1770 ( 
.A(n_1402),
.B(n_1011),
.Y(n_1770)
);

INVx2_ASAP7_75t_L g1771 ( 
.A(n_1394),
.Y(n_1771)
);

NAND2xp5_ASAP7_75t_L g1772 ( 
.A(n_1448),
.B(n_1016),
.Y(n_1772)
);

OR2x6_ASAP7_75t_L g1773 ( 
.A(n_1396),
.B(n_1245),
.Y(n_1773)
);

INVx1_ASAP7_75t_L g1774 ( 
.A(n_1402),
.Y(n_1774)
);

INVx1_ASAP7_75t_L g1775 ( 
.A(n_1402),
.Y(n_1775)
);

AOI22xp33_ASAP7_75t_L g1776 ( 
.A1(n_1448),
.A2(n_845),
.B1(n_851),
.B2(n_841),
.Y(n_1776)
);

INVx1_ASAP7_75t_L g1777 ( 
.A(n_1402),
.Y(n_1777)
);

INVx2_ASAP7_75t_SL g1778 ( 
.A(n_1397),
.Y(n_1778)
);

NAND2xp5_ASAP7_75t_SL g1779 ( 
.A(n_1450),
.B(n_1147),
.Y(n_1779)
);

INVx2_ASAP7_75t_L g1780 ( 
.A(n_1394),
.Y(n_1780)
);

NOR2xp33_ASAP7_75t_L g1781 ( 
.A(n_1402),
.B(n_1017),
.Y(n_1781)
);

NAND2xp5_ASAP7_75t_L g1782 ( 
.A(n_1448),
.B(n_1024),
.Y(n_1782)
);

NOR3xp33_ASAP7_75t_L g1783 ( 
.A(n_1447),
.B(n_1260),
.C(n_1222),
.Y(n_1783)
);

NAND2xp5_ASAP7_75t_L g1784 ( 
.A(n_1448),
.B(n_1028),
.Y(n_1784)
);

NOR2xp33_ASAP7_75t_L g1785 ( 
.A(n_1402),
.B(n_1029),
.Y(n_1785)
);

BUFx2_ASAP7_75t_SL g1786 ( 
.A(n_1399),
.Y(n_1786)
);

INVx1_ASAP7_75t_L g1787 ( 
.A(n_1402),
.Y(n_1787)
);

BUFx6f_ASAP7_75t_L g1788 ( 
.A(n_1464),
.Y(n_1788)
);

NOR2xp33_ASAP7_75t_L g1789 ( 
.A(n_1402),
.B(n_1031),
.Y(n_1789)
);

OR2x2_ASAP7_75t_L g1790 ( 
.A(n_1396),
.B(n_1251),
.Y(n_1790)
);

NAND2xp5_ASAP7_75t_SL g1791 ( 
.A(n_1450),
.B(n_1150),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1402),
.Y(n_1792)
);

INVx1_ASAP7_75t_L g1793 ( 
.A(n_1402),
.Y(n_1793)
);

NOR3xp33_ASAP7_75t_L g1794 ( 
.A(n_1447),
.B(n_1036),
.C(n_1035),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1402),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1448),
.B(n_1045),
.Y(n_1796)
);

NAND2xp5_ASAP7_75t_L g1797 ( 
.A(n_1448),
.B(n_1046),
.Y(n_1797)
);

INVx1_ASAP7_75t_L g1798 ( 
.A(n_1402),
.Y(n_1798)
);

NAND3xp33_ASAP7_75t_L g1799 ( 
.A(n_1442),
.B(n_1052),
.C(n_1050),
.Y(n_1799)
);

INVx2_ASAP7_75t_L g1800 ( 
.A(n_1394),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1394),
.Y(n_1801)
);

NOR3xp33_ASAP7_75t_L g1802 ( 
.A(n_1447),
.B(n_1055),
.C(n_1053),
.Y(n_1802)
);

INVx2_ASAP7_75t_L g1803 ( 
.A(n_1394),
.Y(n_1803)
);

OR2x6_ASAP7_75t_L g1804 ( 
.A(n_1786),
.B(n_1150),
.Y(n_1804)
);

NAND2xp5_ASAP7_75t_L g1805 ( 
.A(n_1566),
.B(n_1057),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1580),
.Y(n_1806)
);

INVx2_ASAP7_75t_SL g1807 ( 
.A(n_1591),
.Y(n_1807)
);

INVx2_ASAP7_75t_L g1808 ( 
.A(n_1665),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1576),
.B(n_1058),
.Y(n_1809)
);

NAND2xp5_ASAP7_75t_L g1810 ( 
.A(n_1567),
.B(n_1749),
.Y(n_1810)
);

BUFx4f_ASAP7_75t_L g1811 ( 
.A(n_1672),
.Y(n_1811)
);

INVx2_ASAP7_75t_L g1812 ( 
.A(n_1665),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1592),
.Y(n_1813)
);

INVx1_ASAP7_75t_L g1814 ( 
.A(n_1594),
.Y(n_1814)
);

AND2x4_ASAP7_75t_L g1815 ( 
.A(n_1763),
.B(n_862),
.Y(n_1815)
);

AOI21xp5_ASAP7_75t_L g1816 ( 
.A1(n_1675),
.A2(n_868),
.B(n_864),
.Y(n_1816)
);

INVx1_ASAP7_75t_L g1817 ( 
.A(n_1612),
.Y(n_1817)
);

INVx3_ASAP7_75t_L g1818 ( 
.A(n_1672),
.Y(n_1818)
);

AOI21xp5_ASAP7_75t_L g1819 ( 
.A1(n_1624),
.A2(n_874),
.B(n_873),
.Y(n_1819)
);

INVxp67_ASAP7_75t_L g1820 ( 
.A(n_1575),
.Y(n_1820)
);

INVx2_ASAP7_75t_SL g1821 ( 
.A(n_1608),
.Y(n_1821)
);

INVxp33_ASAP7_75t_SL g1822 ( 
.A(n_1569),
.Y(n_1822)
);

XOR2xp5_ASAP7_75t_L g1823 ( 
.A(n_1710),
.B(n_961),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1778),
.B(n_875),
.Y(n_1824)
);

INVx1_ASAP7_75t_L g1825 ( 
.A(n_1613),
.Y(n_1825)
);

INVx1_ASAP7_75t_L g1826 ( 
.A(n_1630),
.Y(n_1826)
);

INVx2_ASAP7_75t_SL g1827 ( 
.A(n_1608),
.Y(n_1827)
);

NAND2xp5_ASAP7_75t_L g1828 ( 
.A(n_1750),
.B(n_1060),
.Y(n_1828)
);

NAND2xp5_ASAP7_75t_SL g1829 ( 
.A(n_1665),
.B(n_1062),
.Y(n_1829)
);

NAND2xp5_ASAP7_75t_L g1830 ( 
.A(n_1751),
.B(n_1064),
.Y(n_1830)
);

BUFx4f_ASAP7_75t_L g1831 ( 
.A(n_1672),
.Y(n_1831)
);

OR2x6_ASAP7_75t_L g1832 ( 
.A(n_1608),
.B(n_1160),
.Y(n_1832)
);

INVx2_ASAP7_75t_L g1833 ( 
.A(n_1627),
.Y(n_1833)
);

BUFx3_ASAP7_75t_L g1834 ( 
.A(n_1696),
.Y(n_1834)
);

O2A1O1Ixp33_ASAP7_75t_L g1835 ( 
.A1(n_1640),
.A2(n_1646),
.B(n_1644),
.C(n_1632),
.Y(n_1835)
);

INVx2_ASAP7_75t_L g1836 ( 
.A(n_1629),
.Y(n_1836)
);

NOR2xp33_ASAP7_75t_R g1837 ( 
.A(n_1673),
.B(n_969),
.Y(n_1837)
);

NAND2xp5_ASAP7_75t_L g1838 ( 
.A(n_1760),
.B(n_1065),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1601),
.B(n_877),
.Y(n_1839)
);

BUFx3_ASAP7_75t_L g1840 ( 
.A(n_1696),
.Y(n_1840)
);

NAND2xp5_ASAP7_75t_L g1841 ( 
.A(n_1762),
.B(n_1066),
.Y(n_1841)
);

BUFx3_ASAP7_75t_L g1842 ( 
.A(n_1756),
.Y(n_1842)
);

AND2x4_ASAP7_75t_L g1843 ( 
.A(n_1601),
.B(n_880),
.Y(n_1843)
);

INVx2_ASAP7_75t_L g1844 ( 
.A(n_1554),
.Y(n_1844)
);

INVx2_ASAP7_75t_SL g1845 ( 
.A(n_1704),
.Y(n_1845)
);

AOI22xp33_ASAP7_75t_L g1846 ( 
.A1(n_1682),
.A2(n_999),
.B1(n_1014),
.B2(n_984),
.Y(n_1846)
);

NAND2xp5_ASAP7_75t_L g1847 ( 
.A(n_1768),
.B(n_1067),
.Y(n_1847)
);

INVx3_ASAP7_75t_L g1848 ( 
.A(n_1693),
.Y(n_1848)
);

NOR2xp33_ASAP7_75t_L g1849 ( 
.A(n_1614),
.B(n_999),
.Y(n_1849)
);

HB1xp67_ASAP7_75t_L g1850 ( 
.A(n_1607),
.Y(n_1850)
);

NOR2xp33_ASAP7_75t_L g1851 ( 
.A(n_1579),
.B(n_1014),
.Y(n_1851)
);

NOR2x1p5_ASAP7_75t_L g1852 ( 
.A(n_1602),
.B(n_1790),
.Y(n_1852)
);

AND2x2_ASAP7_75t_SL g1853 ( 
.A(n_1560),
.B(n_1023),
.Y(n_1853)
);

INVx2_ASAP7_75t_L g1854 ( 
.A(n_1748),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1772),
.B(n_1069),
.Y(n_1855)
);

AND2x4_ASAP7_75t_L g1856 ( 
.A(n_1622),
.B(n_883),
.Y(n_1856)
);

NAND2xp5_ASAP7_75t_L g1857 ( 
.A(n_1782),
.B(n_1070),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1756),
.Y(n_1858)
);

INVx1_ASAP7_75t_SL g1859 ( 
.A(n_1633),
.Y(n_1859)
);

INVx2_ASAP7_75t_SL g1860 ( 
.A(n_1708),
.Y(n_1860)
);

AND2x4_ASAP7_75t_L g1861 ( 
.A(n_1625),
.B(n_885),
.Y(n_1861)
);

NAND2xp5_ASAP7_75t_L g1862 ( 
.A(n_1784),
.B(n_1074),
.Y(n_1862)
);

AOI22xp33_ASAP7_75t_L g1863 ( 
.A1(n_1686),
.A2(n_1038),
.B1(n_1040),
.B2(n_1023),
.Y(n_1863)
);

INVx1_ASAP7_75t_L g1864 ( 
.A(n_1634),
.Y(n_1864)
);

INVx1_ASAP7_75t_L g1865 ( 
.A(n_1755),
.Y(n_1865)
);

INVx1_ASAP7_75t_L g1866 ( 
.A(n_1758),
.Y(n_1866)
);

NOR2xp33_ASAP7_75t_L g1867 ( 
.A(n_1753),
.B(n_1038),
.Y(n_1867)
);

NOR2x2_ASAP7_75t_L g1868 ( 
.A(n_1650),
.B(n_1253),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1774),
.Y(n_1869)
);

BUFx6f_ASAP7_75t_SL g1870 ( 
.A(n_1650),
.Y(n_1870)
);

NAND2x1p5_ASAP7_75t_L g1871 ( 
.A(n_1642),
.B(n_886),
.Y(n_1871)
);

AOI22xp5_ASAP7_75t_L g1872 ( 
.A1(n_1655),
.A2(n_1089),
.B1(n_1092),
.B2(n_1088),
.Y(n_1872)
);

AND2x4_ASAP7_75t_L g1873 ( 
.A(n_1631),
.B(n_887),
.Y(n_1873)
);

AOI22xp33_ASAP7_75t_L g1874 ( 
.A1(n_1680),
.A2(n_1043),
.B1(n_1054),
.B2(n_1040),
.Y(n_1874)
);

BUFx2_ASAP7_75t_L g1875 ( 
.A(n_1711),
.Y(n_1875)
);

AOI22xp5_ASAP7_75t_L g1876 ( 
.A1(n_1583),
.A2(n_1094),
.B1(n_1097),
.B2(n_1093),
.Y(n_1876)
);

INVx3_ASAP7_75t_L g1877 ( 
.A(n_1693),
.Y(n_1877)
);

INVx1_ASAP7_75t_L g1878 ( 
.A(n_1775),
.Y(n_1878)
);

INVx2_ASAP7_75t_L g1879 ( 
.A(n_1777),
.Y(n_1879)
);

AO22x1_ASAP7_75t_L g1880 ( 
.A1(n_1668),
.A2(n_1054),
.B1(n_1105),
.B2(n_1043),
.Y(n_1880)
);

AND2x2_ASAP7_75t_SL g1881 ( 
.A(n_1678),
.B(n_1105),
.Y(n_1881)
);

INVx2_ASAP7_75t_L g1882 ( 
.A(n_1787),
.Y(n_1882)
);

INVxp67_ASAP7_75t_L g1883 ( 
.A(n_1796),
.Y(n_1883)
);

INVx1_ASAP7_75t_L g1884 ( 
.A(n_1792),
.Y(n_1884)
);

INVx1_ASAP7_75t_L g1885 ( 
.A(n_1793),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1795),
.Y(n_1886)
);

NOR2xp33_ASAP7_75t_L g1887 ( 
.A(n_1638),
.B(n_1641),
.Y(n_1887)
);

BUFx2_ASAP7_75t_L g1888 ( 
.A(n_1684),
.Y(n_1888)
);

INVx2_ASAP7_75t_L g1889 ( 
.A(n_1798),
.Y(n_1889)
);

NAND2xp5_ASAP7_75t_L g1890 ( 
.A(n_1797),
.B(n_1098),
.Y(n_1890)
);

NOR2xp33_ASAP7_75t_SL g1891 ( 
.A(n_1724),
.B(n_1110),
.Y(n_1891)
);

INVx8_ASAP7_75t_L g1892 ( 
.A(n_1773),
.Y(n_1892)
);

INVx4_ASAP7_75t_L g1893 ( 
.A(n_1773),
.Y(n_1893)
);

NOR2xp33_ASAP7_75t_L g1894 ( 
.A(n_1584),
.B(n_1110),
.Y(n_1894)
);

HB1xp67_ASAP7_75t_L g1895 ( 
.A(n_1727),
.Y(n_1895)
);

OAI22xp5_ASAP7_75t_L g1896 ( 
.A1(n_1688),
.A2(n_1132),
.B1(n_1159),
.B2(n_1116),
.Y(n_1896)
);

INVx2_ASAP7_75t_L g1897 ( 
.A(n_1555),
.Y(n_1897)
);

INVx2_ASAP7_75t_L g1898 ( 
.A(n_1558),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1557),
.B(n_1102),
.Y(n_1899)
);

AOI22xp5_ASAP7_75t_L g1900 ( 
.A1(n_1589),
.A2(n_1104),
.B1(n_1111),
.B2(n_1103),
.Y(n_1900)
);

NOR2xp33_ASAP7_75t_L g1901 ( 
.A(n_1593),
.B(n_1116),
.Y(n_1901)
);

NAND2xp5_ASAP7_75t_L g1902 ( 
.A(n_1559),
.B(n_1113),
.Y(n_1902)
);

AND2x2_ASAP7_75t_L g1903 ( 
.A(n_1663),
.B(n_1132),
.Y(n_1903)
);

INVx1_ASAP7_75t_L g1904 ( 
.A(n_1637),
.Y(n_1904)
);

OR2x2_ASAP7_75t_L g1905 ( 
.A(n_1714),
.B(n_1115),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_SL g1906 ( 
.A(n_1670),
.B(n_1163),
.C(n_1159),
.Y(n_1906)
);

INVx2_ASAP7_75t_L g1907 ( 
.A(n_1564),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1596),
.B(n_1163),
.Y(n_1908)
);

BUFx6f_ASAP7_75t_L g1909 ( 
.A(n_1605),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_L g1910 ( 
.A(n_1654),
.B(n_1118),
.Y(n_1910)
);

OAI22xp5_ASAP7_75t_SL g1911 ( 
.A1(n_1663),
.A2(n_1182),
.B1(n_1196),
.B2(n_1166),
.Y(n_1911)
);

OR2x6_ASAP7_75t_L g1912 ( 
.A(n_1687),
.B(n_1160),
.Y(n_1912)
);

INVx2_ASAP7_75t_L g1913 ( 
.A(n_1565),
.Y(n_1913)
);

AOI22xp33_ASAP7_75t_L g1914 ( 
.A1(n_1765),
.A2(n_1182),
.B1(n_1196),
.B2(n_1166),
.Y(n_1914)
);

OAI22xp5_ASAP7_75t_L g1915 ( 
.A1(n_1697),
.A2(n_1217),
.B1(n_1221),
.B2(n_1210),
.Y(n_1915)
);

NOR2x2_ASAP7_75t_L g1916 ( 
.A(n_1636),
.B(n_1210),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1643),
.Y(n_1917)
);

INVx1_ASAP7_75t_L g1918 ( 
.A(n_1577),
.Y(n_1918)
);

INVx2_ASAP7_75t_L g1919 ( 
.A(n_1578),
.Y(n_1919)
);

NOR2xp67_ASAP7_75t_L g1920 ( 
.A(n_1556),
.B(n_17),
.Y(n_1920)
);

BUFx4f_ASAP7_75t_L g1921 ( 
.A(n_1690),
.Y(n_1921)
);

AND2x4_ASAP7_75t_L g1922 ( 
.A(n_1739),
.B(n_888),
.Y(n_1922)
);

INVx2_ASAP7_75t_L g1923 ( 
.A(n_1581),
.Y(n_1923)
);

AND2x4_ASAP7_75t_L g1924 ( 
.A(n_1600),
.B(n_889),
.Y(n_1924)
);

BUFx3_ASAP7_75t_L g1925 ( 
.A(n_1706),
.Y(n_1925)
);

INVx2_ASAP7_75t_SL g1926 ( 
.A(n_1709),
.Y(n_1926)
);

O2A1O1Ixp33_ASAP7_75t_L g1927 ( 
.A1(n_1582),
.A2(n_896),
.B(n_897),
.C(n_890),
.Y(n_1927)
);

INVx1_ASAP7_75t_L g1928 ( 
.A(n_1585),
.Y(n_1928)
);

INVx1_ASAP7_75t_L g1929 ( 
.A(n_1606),
.Y(n_1929)
);

NOR2xp33_ASAP7_75t_L g1930 ( 
.A(n_1597),
.B(n_1217),
.Y(n_1930)
);

INVx4_ASAP7_75t_L g1931 ( 
.A(n_1746),
.Y(n_1931)
);

AOI22xp5_ASAP7_75t_L g1932 ( 
.A1(n_1586),
.A2(n_1125),
.B1(n_1126),
.B2(n_1122),
.Y(n_1932)
);

OAI21xp5_ASAP7_75t_L g1933 ( 
.A1(n_1661),
.A2(n_907),
.B(n_902),
.Y(n_1933)
);

NOR2xp33_ASAP7_75t_L g1934 ( 
.A(n_1621),
.B(n_1221),
.Y(n_1934)
);

INVx2_ASAP7_75t_L g1935 ( 
.A(n_1623),
.Y(n_1935)
);

AND2x6_ASAP7_75t_L g1936 ( 
.A(n_1605),
.B(n_1208),
.Y(n_1936)
);

INVx1_ASAP7_75t_L g1937 ( 
.A(n_1759),
.Y(n_1937)
);

AO22x1_ASAP7_75t_L g1938 ( 
.A1(n_1723),
.A2(n_1253),
.B1(n_1133),
.B2(n_1134),
.Y(n_1938)
);

INVx1_ASAP7_75t_L g1939 ( 
.A(n_1771),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1776),
.B(n_1127),
.Y(n_1940)
);

NOR2x2_ASAP7_75t_L g1941 ( 
.A(n_1636),
.B(n_1208),
.Y(n_1941)
);

NOR2x2_ASAP7_75t_L g1942 ( 
.A(n_1571),
.B(n_1238),
.Y(n_1942)
);

BUFx3_ASAP7_75t_L g1943 ( 
.A(n_1645),
.Y(n_1943)
);

INVxp67_ASAP7_75t_L g1944 ( 
.A(n_1574),
.Y(n_1944)
);

INVx1_ASAP7_75t_SL g1945 ( 
.A(n_1628),
.Y(n_1945)
);

NOR2xp33_ASAP7_75t_L g1946 ( 
.A(n_1799),
.B(n_1136),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_L g1947 ( 
.A(n_1639),
.B(n_1658),
.Y(n_1947)
);

INVx5_ASAP7_75t_L g1948 ( 
.A(n_1605),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1662),
.B(n_1139),
.Y(n_1949)
);

A2O1A1Ixp33_ASAP7_75t_L g1950 ( 
.A1(n_1595),
.A2(n_911),
.B(n_916),
.C(n_908),
.Y(n_1950)
);

HB1xp67_ASAP7_75t_L g1951 ( 
.A(n_1677),
.Y(n_1951)
);

NAND2xp5_ASAP7_75t_SL g1952 ( 
.A(n_1588),
.B(n_1141),
.Y(n_1952)
);

NOR3xp33_ASAP7_75t_SL g1953 ( 
.A(n_1722),
.B(n_1145),
.C(n_1143),
.Y(n_1953)
);

NAND2xp33_ASAP7_75t_SL g1954 ( 
.A(n_1705),
.B(n_1249),
.Y(n_1954)
);

AND2x4_ASAP7_75t_L g1955 ( 
.A(n_1647),
.B(n_921),
.Y(n_1955)
);

INVx1_ASAP7_75t_L g1956 ( 
.A(n_1780),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1667),
.B(n_1146),
.Y(n_1957)
);

INVx2_ASAP7_75t_L g1958 ( 
.A(n_1800),
.Y(n_1958)
);

INVx2_ASAP7_75t_L g1959 ( 
.A(n_1801),
.Y(n_1959)
);

BUFx2_ASAP7_75t_L g1960 ( 
.A(n_1734),
.Y(n_1960)
);

AND2x4_ASAP7_75t_L g1961 ( 
.A(n_1647),
.B(n_923),
.Y(n_1961)
);

CKINVDCx20_ASAP7_75t_R g1962 ( 
.A(n_1652),
.Y(n_1962)
);

INVx1_ASAP7_75t_L g1963 ( 
.A(n_1803),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_L g1964 ( 
.A(n_1616),
.B(n_1148),
.Y(n_1964)
);

AND2x4_ASAP7_75t_L g1965 ( 
.A(n_1685),
.B(n_924),
.Y(n_1965)
);

NAND2xp5_ASAP7_75t_L g1966 ( 
.A(n_1653),
.B(n_1149),
.Y(n_1966)
);

AND2x2_ASAP7_75t_L g1967 ( 
.A(n_1689),
.B(n_1153),
.Y(n_1967)
);

NAND2xp33_ASAP7_75t_SL g1968 ( 
.A(n_1679),
.B(n_1154),
.Y(n_1968)
);

INVx2_ASAP7_75t_L g1969 ( 
.A(n_1664),
.Y(n_1969)
);

CKINVDCx5p33_ASAP7_75t_R g1970 ( 
.A(n_1656),
.Y(n_1970)
);

CKINVDCx5p33_ASAP7_75t_R g1971 ( 
.A(n_1657),
.Y(n_1971)
);

INVx1_ASAP7_75t_L g1972 ( 
.A(n_1671),
.Y(n_1972)
);

INVx1_ASAP7_75t_L g1973 ( 
.A(n_1648),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1599),
.A2(n_931),
.B(n_926),
.Y(n_1974)
);

AND2x2_ASAP7_75t_L g1975 ( 
.A(n_1700),
.B(n_1162),
.Y(n_1975)
);

OAI22xp5_ASAP7_75t_L g1976 ( 
.A1(n_1590),
.A2(n_944),
.B1(n_948),
.B2(n_937),
.Y(n_1976)
);

INVx1_ASAP7_75t_L g1977 ( 
.A(n_1635),
.Y(n_1977)
);

CKINVDCx5p33_ASAP7_75t_R g1978 ( 
.A(n_1604),
.Y(n_1978)
);

BUFx8_ASAP7_75t_L g1979 ( 
.A(n_1587),
.Y(n_1979)
);

INVx3_ASAP7_75t_L g1980 ( 
.A(n_1649),
.Y(n_1980)
);

XOR2xp5_ASAP7_75t_L g1981 ( 
.A(n_1676),
.B(n_1165),
.Y(n_1981)
);

O2A1O1Ixp33_ASAP7_75t_L g1982 ( 
.A1(n_1691),
.A2(n_953),
.B(n_955),
.C(n_951),
.Y(n_1982)
);

NOR2xp33_ASAP7_75t_L g1983 ( 
.A(n_1609),
.B(n_1167),
.Y(n_1983)
);

AND2x4_ASAP7_75t_L g1984 ( 
.A(n_1692),
.B(n_1651),
.Y(n_1984)
);

OR2x6_ASAP7_75t_L g1985 ( 
.A(n_1587),
.B(n_1757),
.Y(n_1985)
);

INVx1_ASAP7_75t_L g1986 ( 
.A(n_1733),
.Y(n_1986)
);

AND2x6_ASAP7_75t_L g1987 ( 
.A(n_1669),
.B(n_1238),
.Y(n_1987)
);

INVx1_ASAP7_75t_L g1988 ( 
.A(n_1735),
.Y(n_1988)
);

AOI22xp5_ASAP7_75t_L g1989 ( 
.A1(n_1752),
.A2(n_1170),
.B1(n_1175),
.B2(n_1169),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1738),
.Y(n_1990)
);

NOR2xp33_ASAP7_75t_R g1991 ( 
.A(n_1766),
.B(n_1176),
.Y(n_1991)
);

OR2x6_ASAP7_75t_L g1992 ( 
.A(n_1767),
.B(n_956),
.Y(n_1992)
);

AND2x4_ASAP7_75t_L g1993 ( 
.A(n_1562),
.B(n_959),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1568),
.B(n_1181),
.Y(n_1994)
);

AND2x2_ASAP7_75t_L g1995 ( 
.A(n_1611),
.B(n_1183),
.Y(n_1995)
);

BUFx6f_ASAP7_75t_L g1996 ( 
.A(n_1599),
.Y(n_1996)
);

INVxp33_ASAP7_75t_L g1997 ( 
.A(n_1794),
.Y(n_1997)
);

NAND2xp33_ASAP7_75t_L g1998 ( 
.A(n_1669),
.B(n_1674),
.Y(n_1998)
);

AND2x4_ASAP7_75t_L g1999 ( 
.A(n_1563),
.B(n_962),
.Y(n_1999)
);

NAND2xp33_ASAP7_75t_L g2000 ( 
.A(n_1669),
.B(n_1184),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1761),
.B(n_1189),
.Y(n_2001)
);

NOR2xp33_ASAP7_75t_L g2002 ( 
.A(n_1618),
.B(n_1191),
.Y(n_2002)
);

INVx1_ASAP7_75t_L g2003 ( 
.A(n_1720),
.Y(n_2003)
);

AND2x2_ASAP7_75t_SL g2004 ( 
.A(n_1802),
.B(n_965),
.Y(n_2004)
);

BUFx2_ASAP7_75t_L g2005 ( 
.A(n_1698),
.Y(n_2005)
);

INVx2_ASAP7_75t_L g2006 ( 
.A(n_1719),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_L g2007 ( 
.A(n_1764),
.B(n_1193),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1620),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_L g2009 ( 
.A(n_1769),
.B(n_1195),
.Y(n_2009)
);

AND2x2_ASAP7_75t_L g2010 ( 
.A(n_1626),
.B(n_1197),
.Y(n_2010)
);

INVx3_ASAP7_75t_L g2011 ( 
.A(n_1683),
.Y(n_2011)
);

INVx4_ASAP7_75t_L g2012 ( 
.A(n_1707),
.Y(n_2012)
);

NOR2xp67_ASAP7_75t_L g2013 ( 
.A(n_1598),
.B(n_18),
.Y(n_2013)
);

BUFx3_ASAP7_75t_L g2014 ( 
.A(n_1694),
.Y(n_2014)
);

NAND2xp5_ASAP7_75t_L g2015 ( 
.A(n_1770),
.B(n_1198),
.Y(n_2015)
);

INVx1_ASAP7_75t_L g2016 ( 
.A(n_1725),
.Y(n_2016)
);

AND2x6_ASAP7_75t_L g2017 ( 
.A(n_1674),
.B(n_970),
.Y(n_2017)
);

CKINVDCx5p33_ASAP7_75t_R g2018 ( 
.A(n_1717),
.Y(n_2018)
);

NAND2xp5_ASAP7_75t_L g2019 ( 
.A(n_1781),
.B(n_1199),
.Y(n_2019)
);

BUFx12f_ASAP7_75t_L g2020 ( 
.A(n_1713),
.Y(n_2020)
);

AND2x4_ASAP7_75t_L g2021 ( 
.A(n_1695),
.B(n_972),
.Y(n_2021)
);

CKINVDCx5p33_ASAP7_75t_R g2022 ( 
.A(n_1779),
.Y(n_2022)
);

OAI22xp33_ASAP7_75t_L g2023 ( 
.A1(n_1702),
.A2(n_1202),
.B1(n_1205),
.B2(n_1201),
.Y(n_2023)
);

INVx2_ASAP7_75t_L g2024 ( 
.A(n_1788),
.Y(n_2024)
);

NOR2x2_ASAP7_75t_L g2025 ( 
.A(n_1659),
.B(n_1244),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1785),
.B(n_1206),
.Y(n_2026)
);

AOI22xp5_ASAP7_75t_L g2027 ( 
.A1(n_1789),
.A2(n_1212),
.B1(n_1213),
.B2(n_1207),
.Y(n_2027)
);

INVx2_ASAP7_75t_SL g2028 ( 
.A(n_1701),
.Y(n_2028)
);

NOR2xp33_ASAP7_75t_L g2029 ( 
.A(n_1561),
.B(n_1791),
.Y(n_2029)
);

INVx2_ASAP7_75t_SL g2030 ( 
.A(n_1703),
.Y(n_2030)
);

INVx2_ASAP7_75t_SL g2031 ( 
.A(n_1712),
.Y(n_2031)
);

NOR2x1p5_ASAP7_75t_L g2032 ( 
.A(n_1681),
.B(n_1250),
.Y(n_2032)
);

AOI22xp33_ASAP7_75t_L g2033 ( 
.A1(n_1743),
.A2(n_980),
.B1(n_981),
.B2(n_975),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_L g2034 ( 
.A(n_1718),
.B(n_1218),
.Y(n_2034)
);

AND2x2_ASAP7_75t_L g2035 ( 
.A(n_1660),
.B(n_1220),
.Y(n_2035)
);

INVx5_ASAP7_75t_L g2036 ( 
.A(n_1716),
.Y(n_2036)
);

CKINVDCx16_ASAP7_75t_R g2037 ( 
.A(n_1741),
.Y(n_2037)
);

CKINVDCx5p33_ASAP7_75t_R g2038 ( 
.A(n_1666),
.Y(n_2038)
);

CKINVDCx5p33_ASAP7_75t_R g2039 ( 
.A(n_1603),
.Y(n_2039)
);

NOR2xp33_ASAP7_75t_L g2040 ( 
.A(n_1570),
.B(n_1223),
.Y(n_2040)
);

HB1xp67_ASAP7_75t_L g2041 ( 
.A(n_1754),
.Y(n_2041)
);

NOR2xp33_ASAP7_75t_L g2042 ( 
.A(n_1572),
.B(n_1225),
.Y(n_2042)
);

INVx1_ASAP7_75t_L g2043 ( 
.A(n_1728),
.Y(n_2043)
);

AND2x4_ASAP7_75t_L g2044 ( 
.A(n_1573),
.B(n_985),
.Y(n_2044)
);

NAND2xp5_ASAP7_75t_L g2045 ( 
.A(n_1715),
.B(n_1226),
.Y(n_2045)
);

INVx2_ASAP7_75t_L g2046 ( 
.A(n_1747),
.Y(n_2046)
);

BUFx2_ASAP7_75t_L g2047 ( 
.A(n_1729),
.Y(n_2047)
);

BUFx12f_ASAP7_75t_SL g2048 ( 
.A(n_1783),
.Y(n_2048)
);

NAND2xp33_ASAP7_75t_L g2049 ( 
.A(n_1726),
.B(n_1228),
.Y(n_2049)
);

AND3x1_ASAP7_75t_L g2050 ( 
.A(n_1699),
.B(n_995),
.C(n_993),
.Y(n_2050)
);

AOI22xp33_ASAP7_75t_L g2051 ( 
.A1(n_1610),
.A2(n_998),
.B1(n_1000),
.B2(n_996),
.Y(n_2051)
);

AND2x4_ASAP7_75t_L g2052 ( 
.A(n_1619),
.B(n_1006),
.Y(n_2052)
);

INVx1_ASAP7_75t_L g2053 ( 
.A(n_1736),
.Y(n_2053)
);

AOI22xp33_ASAP7_75t_L g2054 ( 
.A1(n_1740),
.A2(n_1018),
.B1(n_1020),
.B2(n_1012),
.Y(n_2054)
);

NOR2xp33_ASAP7_75t_R g2055 ( 
.A(n_1745),
.B(n_1229),
.Y(n_2055)
);

AND2x4_ASAP7_75t_L g2056 ( 
.A(n_1615),
.B(n_1021),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1617),
.B(n_1231),
.Y(n_2057)
);

HB1xp67_ASAP7_75t_L g2058 ( 
.A(n_1661),
.Y(n_2058)
);

NOR2xp33_ASAP7_75t_L g2059 ( 
.A(n_1730),
.B(n_1235),
.Y(n_2059)
);

INVx1_ASAP7_75t_L g2060 ( 
.A(n_1707),
.Y(n_2060)
);

INVx1_ASAP7_75t_L g2061 ( 
.A(n_1731),
.Y(n_2061)
);

O2A1O1Ixp5_ASAP7_75t_L g2062 ( 
.A1(n_1744),
.A2(n_1026),
.B(n_1027),
.C(n_1025),
.Y(n_2062)
);

OR2x2_ASAP7_75t_L g2063 ( 
.A(n_1721),
.B(n_1237),
.Y(n_2063)
);

INVx1_ASAP7_75t_L g2064 ( 
.A(n_1732),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1737),
.B(n_1248),
.Y(n_2065)
);

BUFx6f_ASAP7_75t_L g2066 ( 
.A(n_1742),
.Y(n_2066)
);

NAND2xp5_ASAP7_75t_L g2067 ( 
.A(n_1566),
.B(n_1259),
.Y(n_2067)
);

BUFx6f_ASAP7_75t_L g2068 ( 
.A(n_1605),
.Y(n_2068)
);

INVx1_ASAP7_75t_L g2069 ( 
.A(n_1592),
.Y(n_2069)
);

BUFx2_ASAP7_75t_L g2070 ( 
.A(n_1575),
.Y(n_2070)
);

INVx1_ASAP7_75t_L g2071 ( 
.A(n_1592),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_L g2072 ( 
.A(n_1566),
.B(n_1262),
.Y(n_2072)
);

INVxp67_ASAP7_75t_L g2073 ( 
.A(n_1786),
.Y(n_2073)
);

CKINVDCx5p33_ASAP7_75t_R g2074 ( 
.A(n_1786),
.Y(n_2074)
);

CKINVDCx20_ASAP7_75t_R g2075 ( 
.A(n_1710),
.Y(n_2075)
);

AND2x4_ASAP7_75t_L g2076 ( 
.A(n_1580),
.B(n_1030),
.Y(n_2076)
);

HB1xp67_ASAP7_75t_L g2077 ( 
.A(n_1575),
.Y(n_2077)
);

AOI22xp5_ASAP7_75t_L g2078 ( 
.A1(n_1632),
.A2(n_1263),
.B1(n_1033),
.B2(n_1034),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1665),
.B(n_1032),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1566),
.B(n_1039),
.Y(n_2080)
);

NOR2xp33_ASAP7_75t_L g2081 ( 
.A(n_1632),
.B(n_1227),
.Y(n_2081)
);

AND2x2_ASAP7_75t_L g2082 ( 
.A(n_1644),
.B(n_1044),
.Y(n_2082)
);

NAND2xp5_ASAP7_75t_L g2083 ( 
.A(n_1566),
.B(n_1047),
.Y(n_2083)
);

HB1xp67_ASAP7_75t_L g2084 ( 
.A(n_1575),
.Y(n_2084)
);

NAND2x1p5_ASAP7_75t_L g2085 ( 
.A(n_1580),
.B(n_1048),
.Y(n_2085)
);

BUFx6f_ASAP7_75t_L g2086 ( 
.A(n_1605),
.Y(n_2086)
);

INVx1_ASAP7_75t_L g2087 ( 
.A(n_1592),
.Y(n_2087)
);

INVx2_ASAP7_75t_SL g2088 ( 
.A(n_1580),
.Y(n_2088)
);

NOR3xp33_ASAP7_75t_SL g2089 ( 
.A(n_1714),
.B(n_1063),
.C(n_1051),
.Y(n_2089)
);

NOR3xp33_ASAP7_75t_L g2090 ( 
.A(n_1906),
.B(n_1264),
.C(n_1256),
.Y(n_2090)
);

INVx3_ASAP7_75t_L g2091 ( 
.A(n_1909),
.Y(n_2091)
);

NOR2xp33_ASAP7_75t_L g2092 ( 
.A(n_1851),
.B(n_1867),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_L g2093 ( 
.A(n_1883),
.B(n_1068),
.Y(n_2093)
);

AND2x4_ASAP7_75t_L g2094 ( 
.A(n_1984),
.B(n_1071),
.Y(n_2094)
);

OAI22xp5_ASAP7_75t_L g2095 ( 
.A1(n_1810),
.A2(n_1945),
.B1(n_1947),
.B2(n_1904),
.Y(n_2095)
);

CKINVDCx16_ASAP7_75t_R g2096 ( 
.A(n_1837),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1894),
.B(n_1190),
.Y(n_2097)
);

BUFx2_ASAP7_75t_L g2098 ( 
.A(n_2070),
.Y(n_2098)
);

INVx1_ASAP7_75t_L g2099 ( 
.A(n_1813),
.Y(n_2099)
);

AND2x4_ASAP7_75t_L g2100 ( 
.A(n_1984),
.B(n_1072),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1871),
.B(n_1075),
.Y(n_2101)
);

AOI21xp5_ASAP7_75t_L g2102 ( 
.A1(n_1998),
.A2(n_1077),
.B(n_1076),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1814),
.B(n_1215),
.Y(n_2103)
);

AND2x2_ASAP7_75t_L g2104 ( 
.A(n_1903),
.B(n_1224),
.Y(n_2104)
);

INVx1_ASAP7_75t_L g2105 ( 
.A(n_1817),
.Y(n_2105)
);

INVx1_ASAP7_75t_L g2106 ( 
.A(n_1825),
.Y(n_2106)
);

OAI21xp5_ASAP7_75t_L g2107 ( 
.A1(n_1974),
.A2(n_1080),
.B(n_1079),
.Y(n_2107)
);

O2A1O1Ixp33_ASAP7_75t_L g2108 ( 
.A1(n_1927),
.A2(n_1091),
.B(n_1099),
.C(n_1084),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1888),
.B(n_1100),
.Y(n_2109)
);

BUFx2_ASAP7_75t_L g2110 ( 
.A(n_2077),
.Y(n_2110)
);

AOI21xp5_ASAP7_75t_L g2111 ( 
.A1(n_1933),
.A2(n_1106),
.B(n_1101),
.Y(n_2111)
);

INVx2_ASAP7_75t_L g2112 ( 
.A(n_1826),
.Y(n_2112)
);

OR2x2_ASAP7_75t_L g2113 ( 
.A(n_1896),
.B(n_1108),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1864),
.B(n_1188),
.Y(n_2114)
);

NOR2xp33_ASAP7_75t_L g2115 ( 
.A(n_1901),
.B(n_1194),
.Y(n_2115)
);

AND2x4_ASAP7_75t_L g2116 ( 
.A(n_2003),
.B(n_1119),
.Y(n_2116)
);

OAI21xp33_ASAP7_75t_L g2117 ( 
.A1(n_1891),
.A2(n_1123),
.B(n_1120),
.Y(n_2117)
);

A2O1A1Ixp33_ASAP7_75t_L g2118 ( 
.A1(n_2016),
.A2(n_1131),
.B(n_1135),
.C(n_1130),
.Y(n_2118)
);

BUFx2_ASAP7_75t_L g2119 ( 
.A(n_2084),
.Y(n_2119)
);

INVx1_ASAP7_75t_L g2120 ( 
.A(n_2069),
.Y(n_2120)
);

BUFx3_ASAP7_75t_L g2121 ( 
.A(n_1834),
.Y(n_2121)
);

NOR2xp33_ASAP7_75t_SL g2122 ( 
.A(n_1811),
.B(n_1138),
.Y(n_2122)
);

NAND2xp5_ASAP7_75t_L g2123 ( 
.A(n_2071),
.B(n_1246),
.Y(n_2123)
);

INVx1_ASAP7_75t_SL g2124 ( 
.A(n_1859),
.Y(n_2124)
);

NOR2xp33_ASAP7_75t_R g2125 ( 
.A(n_2075),
.B(n_19),
.Y(n_2125)
);

INVx2_ASAP7_75t_L g2126 ( 
.A(n_2087),
.Y(n_2126)
);

NOR2xp67_ASAP7_75t_SL g2127 ( 
.A(n_1842),
.B(n_1140),
.Y(n_2127)
);

INVx4_ASAP7_75t_L g2128 ( 
.A(n_1831),
.Y(n_2128)
);

OAI21xp33_ASAP7_75t_SL g2129 ( 
.A1(n_2013),
.A2(n_1144),
.B(n_1142),
.Y(n_2129)
);

BUFx12f_ASAP7_75t_L g2130 ( 
.A(n_2074),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1972),
.Y(n_2131)
);

OAI22xp5_ASAP7_75t_L g2132 ( 
.A1(n_1833),
.A2(n_1836),
.B1(n_1944),
.B2(n_1943),
.Y(n_2132)
);

NOR2xp33_ASAP7_75t_L g2133 ( 
.A(n_1908),
.B(n_1173),
.Y(n_2133)
);

INVx3_ASAP7_75t_L g2134 ( 
.A(n_1909),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1819),
.B(n_1185),
.Y(n_2135)
);

NAND2x1_ASAP7_75t_L g2136 ( 
.A(n_2017),
.B(n_1152),
.Y(n_2136)
);

NOR3xp33_ASAP7_75t_SL g2137 ( 
.A(n_1970),
.B(n_1156),
.C(n_1155),
.Y(n_2137)
);

INVx1_ASAP7_75t_L g2138 ( 
.A(n_1969),
.Y(n_2138)
);

INVx1_ASAP7_75t_L g2139 ( 
.A(n_1973),
.Y(n_2139)
);

INVx1_ASAP7_75t_L g2140 ( 
.A(n_1839),
.Y(n_2140)
);

NOR2xp33_ASAP7_75t_R g2141 ( 
.A(n_1840),
.B(n_20),
.Y(n_2141)
);

OAI22xp5_ASAP7_75t_L g2142 ( 
.A1(n_1931),
.A2(n_1171),
.B1(n_1172),
.B2(n_1168),
.Y(n_2142)
);

INVx2_ASAP7_75t_L g2143 ( 
.A(n_1844),
.Y(n_2143)
);

A2O1A1Ixp33_ASAP7_75t_L g2144 ( 
.A1(n_2043),
.A2(n_2062),
.B(n_2029),
.C(n_1816),
.Y(n_2144)
);

INVx3_ASAP7_75t_L g2145 ( 
.A(n_2068),
.Y(n_2145)
);

INVx2_ASAP7_75t_L g2146 ( 
.A(n_1854),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_L g2147 ( 
.A(n_2082),
.B(n_1177),
.Y(n_2147)
);

OR2x2_ASAP7_75t_L g2148 ( 
.A(n_1915),
.B(n_1179),
.Y(n_2148)
);

INVx2_ASAP7_75t_L g2149 ( 
.A(n_1879),
.Y(n_2149)
);

AO22x1_ASAP7_75t_L g2150 ( 
.A1(n_1822),
.A2(n_1203),
.B1(n_1209),
.B2(n_1180),
.Y(n_2150)
);

OAI22xp5_ASAP7_75t_L g2151 ( 
.A1(n_2008),
.A2(n_1230),
.B1(n_1240),
.B2(n_1211),
.Y(n_2151)
);

A2O1A1Ixp33_ASAP7_75t_L g2152 ( 
.A1(n_1950),
.A2(n_1243),
.B(n_1247),
.C(n_1242),
.Y(n_2152)
);

NAND3xp33_ASAP7_75t_L g2153 ( 
.A(n_2089),
.B(n_2002),
.C(n_1983),
.Y(n_2153)
);

INVx1_ASAP7_75t_L g2154 ( 
.A(n_1839),
.Y(n_2154)
);

O2A1O1Ixp33_ASAP7_75t_L g2155 ( 
.A1(n_1976),
.A2(n_1982),
.B(n_1910),
.C(n_2041),
.Y(n_2155)
);

NOR2xp33_ASAP7_75t_L g2156 ( 
.A(n_1930),
.B(n_21),
.Y(n_2156)
);

NAND2xp5_ASAP7_75t_SL g2157 ( 
.A(n_1853),
.B(n_21),
.Y(n_2157)
);

NOR2xp33_ASAP7_75t_L g2158 ( 
.A(n_1820),
.B(n_24),
.Y(n_2158)
);

INVx4_ASAP7_75t_L g2159 ( 
.A(n_1948),
.Y(n_2159)
);

NOR2xp33_ASAP7_75t_L g2160 ( 
.A(n_1926),
.B(n_24),
.Y(n_2160)
);

HB1xp67_ASAP7_75t_L g2161 ( 
.A(n_1850),
.Y(n_2161)
);

BUFx10_ASAP7_75t_L g2162 ( 
.A(n_1832),
.Y(n_2162)
);

OR2x2_ASAP7_75t_L g2163 ( 
.A(n_1880),
.B(n_25),
.Y(n_2163)
);

INVx3_ASAP7_75t_L g2164 ( 
.A(n_2068),
.Y(n_2164)
);

OAI22xp5_ASAP7_75t_L g2165 ( 
.A1(n_1832),
.A2(n_1951),
.B1(n_2083),
.B2(n_2080),
.Y(n_2165)
);

OAI21xp5_ASAP7_75t_L g2166 ( 
.A1(n_1986),
.A2(n_1990),
.B(n_1988),
.Y(n_2166)
);

INVxp67_ASAP7_75t_L g2167 ( 
.A(n_1823),
.Y(n_2167)
);

NAND2xp5_ASAP7_75t_L g2168 ( 
.A(n_2021),
.B(n_26),
.Y(n_2168)
);

AOI21xp5_ASAP7_75t_L g2169 ( 
.A1(n_2079),
.A2(n_773),
.B(n_772),
.Y(n_2169)
);

AND2x2_ASAP7_75t_L g2170 ( 
.A(n_1881),
.B(n_26),
.Y(n_2170)
);

INVx2_ASAP7_75t_L g2171 ( 
.A(n_1882),
.Y(n_2171)
);

AND2x2_ASAP7_75t_L g2172 ( 
.A(n_2085),
.B(n_27),
.Y(n_2172)
);

AOI21xp5_ASAP7_75t_L g2173 ( 
.A1(n_1996),
.A2(n_777),
.B(n_776),
.Y(n_2173)
);

INVx1_ASAP7_75t_L g2174 ( 
.A(n_1843),
.Y(n_2174)
);

O2A1O1Ixp33_ASAP7_75t_L g2175 ( 
.A1(n_2053),
.A2(n_29),
.B(n_27),
.C(n_28),
.Y(n_2175)
);

NAND2xp5_ASAP7_75t_L g2176 ( 
.A(n_2021),
.B(n_28),
.Y(n_2176)
);

AOI21xp5_ASAP7_75t_L g2177 ( 
.A1(n_1996),
.A2(n_782),
.B(n_778),
.Y(n_2177)
);

NOR2xp33_ASAP7_75t_L g2178 ( 
.A(n_1905),
.B(n_29),
.Y(n_2178)
);

A2O1A1Ixp33_ASAP7_75t_L g2179 ( 
.A1(n_2046),
.A2(n_33),
.B(n_30),
.C(n_31),
.Y(n_2179)
);

NAND2xp5_ASAP7_75t_SL g2180 ( 
.A(n_1991),
.B(n_33),
.Y(n_2180)
);

CKINVDCx5p33_ASAP7_75t_R g2181 ( 
.A(n_1870),
.Y(n_2181)
);

NAND2xp5_ASAP7_75t_SL g2182 ( 
.A(n_1815),
.B(n_34),
.Y(n_2182)
);

AOI21xp5_ASAP7_75t_L g2183 ( 
.A1(n_1899),
.A2(n_785),
.B(n_783),
.Y(n_2183)
);

OAI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1918),
.A2(n_790),
.B(n_787),
.Y(n_2184)
);

AND2x2_ASAP7_75t_L g2185 ( 
.A(n_1815),
.B(n_34),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_1808),
.A2(n_799),
.B(n_795),
.Y(n_2186)
);

BUFx6f_ASAP7_75t_L g2187 ( 
.A(n_2068),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_1902),
.A2(n_802),
.B(n_800),
.Y(n_2188)
);

O2A1O1Ixp33_ASAP7_75t_L g2189 ( 
.A1(n_1835),
.A2(n_39),
.B(n_37),
.C(n_38),
.Y(n_2189)
);

INVx1_ASAP7_75t_L g2190 ( 
.A(n_1843),
.Y(n_2190)
);

BUFx4f_ASAP7_75t_L g2191 ( 
.A(n_1892),
.Y(n_2191)
);

OAI21xp33_ASAP7_75t_SL g2192 ( 
.A1(n_1928),
.A2(n_38),
.B(n_39),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_SL g2193 ( 
.A(n_1824),
.B(n_40),
.Y(n_2193)
);

INVx3_ASAP7_75t_L g2194 ( 
.A(n_2086),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1922),
.B(n_40),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1889),
.Y(n_2196)
);

NAND2xp5_ASAP7_75t_L g2197 ( 
.A(n_1922),
.B(n_41),
.Y(n_2197)
);

NAND2x2_ASAP7_75t_L g2198 ( 
.A(n_1858),
.B(n_42),
.Y(n_2198)
);

O2A1O1Ixp33_ASAP7_75t_L g2199 ( 
.A1(n_1940),
.A2(n_44),
.B(n_42),
.C(n_43),
.Y(n_2199)
);

OAI22xp5_ASAP7_75t_L g2200 ( 
.A1(n_1929),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2200)
);

AND2x2_ASAP7_75t_SL g2201 ( 
.A(n_1874),
.B(n_46),
.Y(n_2201)
);

AOI21x1_ASAP7_75t_L g2202 ( 
.A1(n_1829),
.A2(n_805),
.B(n_804),
.Y(n_2202)
);

AND2x2_ASAP7_75t_L g2203 ( 
.A(n_1824),
.B(n_48),
.Y(n_2203)
);

INVx1_ASAP7_75t_L g2204 ( 
.A(n_1937),
.Y(n_2204)
);

O2A1O1Ixp33_ASAP7_75t_L g2205 ( 
.A1(n_1966),
.A2(n_1960),
.B(n_1828),
.C(n_1830),
.Y(n_2205)
);

INVx2_ASAP7_75t_SL g2206 ( 
.A(n_1818),
.Y(n_2206)
);

INVxp67_ASAP7_75t_L g2207 ( 
.A(n_1911),
.Y(n_2207)
);

A2O1A1Ixp33_ASAP7_75t_L g2208 ( 
.A1(n_2081),
.A2(n_51),
.B(n_49),
.C(n_50),
.Y(n_2208)
);

AOI33xp33_ASAP7_75t_L g2209 ( 
.A1(n_2054),
.A2(n_51),
.A3(n_53),
.B1(n_49),
.B2(n_50),
.B3(n_52),
.Y(n_2209)
);

AND2x2_ASAP7_75t_L g2210 ( 
.A(n_2005),
.B(n_1852),
.Y(n_2210)
);

AOI22xp33_ASAP7_75t_L g2211 ( 
.A1(n_1934),
.A2(n_54),
.B1(n_52),
.B2(n_53),
.Y(n_2211)
);

A2O1A1Ixp33_ASAP7_75t_L g2212 ( 
.A1(n_1920),
.A2(n_56),
.B(n_54),
.C(n_55),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1939),
.Y(n_2213)
);

NAND2xp5_ASAP7_75t_L g2214 ( 
.A(n_2047),
.B(n_57),
.Y(n_2214)
);

INVx4_ASAP7_75t_L g2215 ( 
.A(n_1948),
.Y(n_2215)
);

AOI22xp33_ASAP7_75t_L g2216 ( 
.A1(n_1962),
.A2(n_61),
.B1(n_59),
.B2(n_60),
.Y(n_2216)
);

INVx1_ASAP7_75t_L g2217 ( 
.A(n_1956),
.Y(n_2217)
);

INVx1_ASAP7_75t_L g2218 ( 
.A(n_1963),
.Y(n_2218)
);

AND2x2_ASAP7_75t_L g2219 ( 
.A(n_1863),
.B(n_60),
.Y(n_2219)
);

INVx1_ASAP7_75t_L g2220 ( 
.A(n_2006),
.Y(n_2220)
);

INVx4_ASAP7_75t_L g2221 ( 
.A(n_1948),
.Y(n_2221)
);

NAND2xp5_ASAP7_75t_L g2222 ( 
.A(n_1838),
.B(n_65),
.Y(n_2222)
);

INVx1_ASAP7_75t_L g2223 ( 
.A(n_1865),
.Y(n_2223)
);

AOI21xp5_ASAP7_75t_L g2224 ( 
.A1(n_1841),
.A2(n_813),
.B(n_65),
.Y(n_2224)
);

BUFx12f_ASAP7_75t_L g2225 ( 
.A(n_1804),
.Y(n_2225)
);

OAI22xp5_ASAP7_75t_L g2226 ( 
.A1(n_1847),
.A2(n_68),
.B1(n_66),
.B2(n_67),
.Y(n_2226)
);

INVx4_ASAP7_75t_L g2227 ( 
.A(n_2086),
.Y(n_2227)
);

NAND2xp5_ASAP7_75t_L g2228 ( 
.A(n_1855),
.B(n_68),
.Y(n_2228)
);

INVxp67_ASAP7_75t_L g2229 ( 
.A(n_1804),
.Y(n_2229)
);

INVx2_ASAP7_75t_L g2230 ( 
.A(n_1897),
.Y(n_2230)
);

NAND2xp5_ASAP7_75t_L g2231 ( 
.A(n_1857),
.B(n_70),
.Y(n_2231)
);

AND2x2_ASAP7_75t_L g2232 ( 
.A(n_1967),
.B(n_71),
.Y(n_2232)
);

AOI21x1_ASAP7_75t_L g2233 ( 
.A1(n_2061),
.A2(n_72),
.B(n_74),
.Y(n_2233)
);

INVx2_ASAP7_75t_SL g2234 ( 
.A(n_1821),
.Y(n_2234)
);

INVx3_ASAP7_75t_L g2235 ( 
.A(n_2012),
.Y(n_2235)
);

AND2x4_ASAP7_75t_L g2236 ( 
.A(n_1827),
.B(n_72),
.Y(n_2236)
);

NOR2xp33_ASAP7_75t_L g2237 ( 
.A(n_1849),
.B(n_739),
.Y(n_2237)
);

AND2x6_ASAP7_75t_L g2238 ( 
.A(n_1812),
.B(n_74),
.Y(n_2238)
);

OAI22xp5_ASAP7_75t_L g2239 ( 
.A1(n_1862),
.A2(n_77),
.B1(n_75),
.B2(n_76),
.Y(n_2239)
);

NAND2xp5_ASAP7_75t_SL g2240 ( 
.A(n_1807),
.B(n_76),
.Y(n_2240)
);

OAI221xp5_ASAP7_75t_L g2241 ( 
.A1(n_1846),
.A2(n_80),
.B1(n_78),
.B2(n_79),
.C(n_83),
.Y(n_2241)
);

INVx2_ASAP7_75t_L g2242 ( 
.A(n_1898),
.Y(n_2242)
);

INVx2_ASAP7_75t_L g2243 ( 
.A(n_1907),
.Y(n_2243)
);

NAND2xp5_ASAP7_75t_L g2244 ( 
.A(n_1890),
.B(n_84),
.Y(n_2244)
);

HB1xp67_ASAP7_75t_L g2245 ( 
.A(n_1875),
.Y(n_2245)
);

BUFx6f_ASAP7_75t_L g2246 ( 
.A(n_2017),
.Y(n_2246)
);

BUFx2_ASAP7_75t_L g2247 ( 
.A(n_2017),
.Y(n_2247)
);

OR2x2_ASAP7_75t_L g2248 ( 
.A(n_1914),
.B(n_87),
.Y(n_2248)
);

AND2x2_ASAP7_75t_L g2249 ( 
.A(n_1975),
.B(n_88),
.Y(n_2249)
);

NAND2xp5_ASAP7_75t_L g2250 ( 
.A(n_1955),
.B(n_90),
.Y(n_2250)
);

INVx3_ASAP7_75t_L g2251 ( 
.A(n_2012),
.Y(n_2251)
);

O2A1O1Ixp33_ASAP7_75t_L g2252 ( 
.A1(n_2001),
.A2(n_97),
.B(n_92),
.C(n_94),
.Y(n_2252)
);

NAND2xp5_ASAP7_75t_L g2253 ( 
.A(n_1955),
.B(n_97),
.Y(n_2253)
);

NAND2xp5_ASAP7_75t_L g2254 ( 
.A(n_1961),
.B(n_98),
.Y(n_2254)
);

NAND2xp5_ASAP7_75t_L g2255 ( 
.A(n_1961),
.B(n_98),
.Y(n_2255)
);

AND2x2_ASAP7_75t_L g2256 ( 
.A(n_2035),
.B(n_99),
.Y(n_2256)
);

AND2x2_ASAP7_75t_L g2257 ( 
.A(n_1995),
.B(n_99),
.Y(n_2257)
);

AOI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_1949),
.A2(n_100),
.B(n_101),
.Y(n_2258)
);

NAND2xp5_ASAP7_75t_L g2259 ( 
.A(n_1805),
.B(n_100),
.Y(n_2259)
);

A2O1A1Ixp33_ASAP7_75t_L g2260 ( 
.A1(n_1965),
.A2(n_104),
.B(n_102),
.C(n_103),
.Y(n_2260)
);

INVx1_ASAP7_75t_L g2261 ( 
.A(n_1866),
.Y(n_2261)
);

NOR2xp33_ASAP7_75t_L g2262 ( 
.A(n_1997),
.B(n_751),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_1809),
.B(n_105),
.Y(n_2263)
);

NAND2xp5_ASAP7_75t_L g2264 ( 
.A(n_2067),
.B(n_106),
.Y(n_2264)
);

AND2x4_ASAP7_75t_L g2265 ( 
.A(n_2032),
.B(n_107),
.Y(n_2265)
);

AOI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_1957),
.A2(n_108),
.B(n_109),
.Y(n_2266)
);

NAND2xp5_ASAP7_75t_SL g2267 ( 
.A(n_2023),
.B(n_108),
.Y(n_2267)
);

BUFx6f_ASAP7_75t_L g2268 ( 
.A(n_2017),
.Y(n_2268)
);

AOI21xp5_ASAP7_75t_L g2269 ( 
.A1(n_1994),
.A2(n_109),
.B(n_110),
.Y(n_2269)
);

NOR2xp33_ASAP7_75t_L g2270 ( 
.A(n_2073),
.B(n_110),
.Y(n_2270)
);

NAND2xp5_ASAP7_75t_L g2271 ( 
.A(n_2072),
.B(n_111),
.Y(n_2271)
);

NAND3xp33_ASAP7_75t_SL g2272 ( 
.A(n_2018),
.B(n_742),
.C(n_740),
.Y(n_2272)
);

AOI21xp5_ASAP7_75t_L g2273 ( 
.A1(n_2034),
.A2(n_112),
.B(n_113),
.Y(n_2273)
);

OR2x2_ASAP7_75t_L g2274 ( 
.A(n_1895),
.B(n_113),
.Y(n_2274)
);

OAI22x1_ASAP7_75t_L g2275 ( 
.A1(n_1916),
.A2(n_117),
.B1(n_114),
.B2(n_116),
.Y(n_2275)
);

NOR2xp33_ASAP7_75t_SL g2276 ( 
.A(n_1893),
.B(n_116),
.Y(n_2276)
);

BUFx4f_ASAP7_75t_L g2277 ( 
.A(n_1892),
.Y(n_2277)
);

INVx1_ASAP7_75t_SL g2278 ( 
.A(n_2076),
.Y(n_2278)
);

NOR3xp33_ASAP7_75t_SL g2279 ( 
.A(n_1971),
.B(n_119),
.C(n_120),
.Y(n_2279)
);

INVx2_ASAP7_75t_L g2280 ( 
.A(n_1913),
.Y(n_2280)
);

AND2x2_ASAP7_75t_L g2281 ( 
.A(n_2010),
.B(n_120),
.Y(n_2281)
);

INVxp67_ASAP7_75t_L g2282 ( 
.A(n_1912),
.Y(n_2282)
);

AOI22xp5_ASAP7_75t_L g2283 ( 
.A1(n_1978),
.A2(n_123),
.B1(n_121),
.B2(n_122),
.Y(n_2283)
);

HB1xp67_ASAP7_75t_L g2284 ( 
.A(n_1912),
.Y(n_2284)
);

OR2x6_ASAP7_75t_L g2285 ( 
.A(n_2088),
.B(n_122),
.Y(n_2285)
);

AOI22xp5_ASAP7_75t_L g2286 ( 
.A1(n_2004),
.A2(n_125),
.B1(n_123),
.B2(n_124),
.Y(n_2286)
);

INVx2_ASAP7_75t_L g2287 ( 
.A(n_1919),
.Y(n_2287)
);

OR2x6_ASAP7_75t_L g2288 ( 
.A(n_1938),
.B(n_125),
.Y(n_2288)
);

O2A1O1Ixp5_ASAP7_75t_SL g2289 ( 
.A1(n_1917),
.A2(n_128),
.B(n_126),
.C(n_127),
.Y(n_2289)
);

BUFx8_ASAP7_75t_L g2290 ( 
.A(n_1845),
.Y(n_2290)
);

INVx5_ASAP7_75t_L g2291 ( 
.A(n_1987),
.Y(n_2291)
);

NAND2xp5_ASAP7_75t_L g2292 ( 
.A(n_1965),
.B(n_1993),
.Y(n_2292)
);

HB1xp67_ASAP7_75t_L g2293 ( 
.A(n_2076),
.Y(n_2293)
);

NAND2xp5_ASAP7_75t_L g2294 ( 
.A(n_1993),
.B(n_129),
.Y(n_2294)
);

BUFx6f_ASAP7_75t_L g2295 ( 
.A(n_1987),
.Y(n_2295)
);

NOR2xp33_ASAP7_75t_L g2296 ( 
.A(n_1925),
.B(n_747),
.Y(n_2296)
);

NAND2xp5_ASAP7_75t_SL g2297 ( 
.A(n_1921),
.B(n_130),
.Y(n_2297)
);

NAND3xp33_ASAP7_75t_SL g2298 ( 
.A(n_1953),
.B(n_751),
.C(n_749),
.Y(n_2298)
);

INVx1_ASAP7_75t_L g2299 ( 
.A(n_1869),
.Y(n_2299)
);

CKINVDCx12_ASAP7_75t_R g2300 ( 
.A(n_1985),
.Y(n_2300)
);

AOI22xp5_ASAP7_75t_L g2301 ( 
.A1(n_2050),
.A2(n_135),
.B1(n_132),
.B2(n_133),
.Y(n_2301)
);

INVx2_ASAP7_75t_L g2302 ( 
.A(n_1923),
.Y(n_2302)
);

INVx2_ASAP7_75t_SL g2303 ( 
.A(n_1979),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_1878),
.Y(n_2304)
);

OAI22xp5_ASAP7_75t_L g2305 ( 
.A1(n_2063),
.A2(n_137),
.B1(n_132),
.B2(n_136),
.Y(n_2305)
);

NOR2xp33_ASAP7_75t_L g2306 ( 
.A(n_1860),
.B(n_2022),
.Y(n_2306)
);

INVx2_ASAP7_75t_L g2307 ( 
.A(n_1935),
.Y(n_2307)
);

INVx4_ASAP7_75t_SL g2308 ( 
.A(n_1936),
.Y(n_2308)
);

HB1xp67_ASAP7_75t_L g2309 ( 
.A(n_1806),
.Y(n_2309)
);

CKINVDCx16_ASAP7_75t_R g2310 ( 
.A(n_2055),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_1958),
.Y(n_2311)
);

BUFx4f_ASAP7_75t_SL g2312 ( 
.A(n_1979),
.Y(n_2312)
);

BUFx2_ASAP7_75t_L g2313 ( 
.A(n_1987),
.Y(n_2313)
);

AND2x2_ASAP7_75t_L g2314 ( 
.A(n_1856),
.B(n_138),
.Y(n_2314)
);

OAI22xp5_ASAP7_75t_L g2315 ( 
.A1(n_2007),
.A2(n_145),
.B1(n_141),
.B2(n_144),
.Y(n_2315)
);

BUFx12f_ASAP7_75t_L g2316 ( 
.A(n_2020),
.Y(n_2316)
);

NAND2xp5_ASAP7_75t_L g2317 ( 
.A(n_1999),
.B(n_1964),
.Y(n_2317)
);

INVx2_ASAP7_75t_L g2318 ( 
.A(n_1959),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_SL g2319 ( 
.A(n_1954),
.B(n_146),
.Y(n_2319)
);

NAND2xp33_ASAP7_75t_L g2320 ( 
.A(n_1987),
.B(n_1936),
.Y(n_2320)
);

AOI22xp5_ASAP7_75t_L g2321 ( 
.A1(n_1856),
.A2(n_1861),
.B1(n_1872),
.B2(n_1876),
.Y(n_2321)
);

AOI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2009),
.A2(n_147),
.B(n_148),
.Y(n_2322)
);

INVx4_ASAP7_75t_L g2323 ( 
.A(n_1936),
.Y(n_2323)
);

NOR3xp33_ASAP7_75t_L g2324 ( 
.A(n_2037),
.B(n_147),
.C(n_149),
.Y(n_2324)
);

NAND3xp33_ASAP7_75t_SL g2325 ( 
.A(n_2033),
.B(n_1932),
.C(n_2015),
.Y(n_2325)
);

BUFx2_ASAP7_75t_L g2326 ( 
.A(n_1936),
.Y(n_2326)
);

AOI21xp5_ASAP7_75t_L g2327 ( 
.A1(n_2019),
.A2(n_152),
.B(n_153),
.Y(n_2327)
);

BUFx3_ASAP7_75t_L g2328 ( 
.A(n_2036),
.Y(n_2328)
);

AOI21xp5_ASAP7_75t_L g2329 ( 
.A1(n_2026),
.A2(n_154),
.B(n_156),
.Y(n_2329)
);

OR2x6_ASAP7_75t_SL g2330 ( 
.A(n_1868),
.B(n_154),
.Y(n_2330)
);

CKINVDCx16_ASAP7_75t_R g2331 ( 
.A(n_1981),
.Y(n_2331)
);

NAND2xp5_ASAP7_75t_L g2332 ( 
.A(n_1999),
.B(n_157),
.Y(n_2332)
);

OAI21xp5_ASAP7_75t_L g2333 ( 
.A1(n_1884),
.A2(n_157),
.B(n_158),
.Y(n_2333)
);

INVx1_ASAP7_75t_L g2334 ( 
.A(n_1885),
.Y(n_2334)
);

OAI21xp5_ASAP7_75t_L g2335 ( 
.A1(n_1886),
.A2(n_158),
.B(n_159),
.Y(n_2335)
);

AND2x2_ASAP7_75t_L g2336 ( 
.A(n_1861),
.B(n_159),
.Y(n_2336)
);

NAND2xp5_ASAP7_75t_L g2337 ( 
.A(n_2078),
.B(n_160),
.Y(n_2337)
);

NAND2xp5_ASAP7_75t_L g2338 ( 
.A(n_2014),
.B(n_160),
.Y(n_2338)
);

INVx1_ASAP7_75t_L g2339 ( 
.A(n_1977),
.Y(n_2339)
);

NOR2xp33_ASAP7_75t_L g2340 ( 
.A(n_1985),
.B(n_737),
.Y(n_2340)
);

OR2x2_ASAP7_75t_L g2341 ( 
.A(n_1900),
.B(n_161),
.Y(n_2341)
);

NOR2xp33_ASAP7_75t_L g2342 ( 
.A(n_1952),
.B(n_738),
.Y(n_2342)
);

CKINVDCx5p33_ASAP7_75t_R g2343 ( 
.A(n_2048),
.Y(n_2343)
);

BUFx6f_ASAP7_75t_L g2344 ( 
.A(n_1848),
.Y(n_2344)
);

AND3x1_ASAP7_75t_SL g2345 ( 
.A(n_1941),
.B(n_162),
.C(n_163),
.Y(n_2345)
);

BUFx3_ASAP7_75t_L g2346 ( 
.A(n_2036),
.Y(n_2346)
);

OAI22xp5_ASAP7_75t_L g2347 ( 
.A1(n_1992),
.A2(n_164),
.B1(n_162),
.B2(n_163),
.Y(n_2347)
);

BUFx6f_ASAP7_75t_L g2348 ( 
.A(n_1877),
.Y(n_2348)
);

NAND2xp5_ASAP7_75t_SL g2349 ( 
.A(n_2036),
.B(n_165),
.Y(n_2349)
);

NAND2x1p5_ASAP7_75t_L g2350 ( 
.A(n_2011),
.B(n_166),
.Y(n_2350)
);

INVx5_ASAP7_75t_L g2351 ( 
.A(n_1980),
.Y(n_2351)
);

OAI22xp5_ASAP7_75t_L g2352 ( 
.A1(n_1992),
.A2(n_167),
.B1(n_165),
.B2(n_166),
.Y(n_2352)
);

INVx2_ASAP7_75t_L g2353 ( 
.A(n_2064),
.Y(n_2353)
);

NOR2xp33_ASAP7_75t_SL g2354 ( 
.A(n_2038),
.B(n_168),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2059),
.A2(n_171),
.B(n_169),
.C(n_170),
.Y(n_2355)
);

A2O1A1Ixp33_ASAP7_75t_L g2356 ( 
.A1(n_1968),
.A2(n_173),
.B(n_171),
.C(n_172),
.Y(n_2356)
);

NOR2xp33_ASAP7_75t_L g2357 ( 
.A(n_2028),
.B(n_172),
.Y(n_2357)
);

OAI22xp5_ASAP7_75t_L g2358 ( 
.A1(n_2030),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2358)
);

AOI33xp33_ASAP7_75t_L g2359 ( 
.A1(n_1873),
.A2(n_177),
.A3(n_180),
.B1(n_174),
.B2(n_175),
.B3(n_179),
.Y(n_2359)
);

OAI21xp33_ASAP7_75t_L g2360 ( 
.A1(n_1989),
.A2(n_179),
.B(n_180),
.Y(n_2360)
);

NAND2xp5_ASAP7_75t_L g2361 ( 
.A(n_2031),
.B(n_181),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2044),
.Y(n_2362)
);

AND2x4_ASAP7_75t_L g2363 ( 
.A(n_1924),
.B(n_182),
.Y(n_2363)
);

INVx1_ASAP7_75t_L g2364 ( 
.A(n_2044),
.Y(n_2364)
);

OAI22xp5_ASAP7_75t_L g2365 ( 
.A1(n_2027),
.A2(n_186),
.B1(n_183),
.B2(n_185),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1946),
.B(n_185),
.Y(n_2366)
);

NOR2xp33_ASAP7_75t_L g2367 ( 
.A(n_2045),
.B(n_753),
.Y(n_2367)
);

NAND2xp5_ASAP7_75t_L g2368 ( 
.A(n_1924),
.B(n_187),
.Y(n_2368)
);

NOR2xp33_ASAP7_75t_L g2369 ( 
.A(n_1873),
.B(n_754),
.Y(n_2369)
);

AOI21xp5_ASAP7_75t_L g2370 ( 
.A1(n_2065),
.A2(n_187),
.B(n_188),
.Y(n_2370)
);

AOI22xp33_ASAP7_75t_L g2371 ( 
.A1(n_2052),
.A2(n_195),
.B1(n_193),
.B2(n_194),
.Y(n_2371)
);

BUFx2_ASAP7_75t_L g2372 ( 
.A(n_2025),
.Y(n_2372)
);

INVx3_ASAP7_75t_L g2373 ( 
.A(n_2060),
.Y(n_2373)
);

BUFx8_ASAP7_75t_L g2374 ( 
.A(n_2052),
.Y(n_2374)
);

INVx1_ASAP7_75t_SL g2375 ( 
.A(n_2049),
.Y(n_2375)
);

INVx1_ASAP7_75t_L g2376 ( 
.A(n_2056),
.Y(n_2376)
);

AOI22xp5_ASAP7_75t_L g2377 ( 
.A1(n_2056),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_2377)
);

NOR2xp33_ASAP7_75t_L g2378 ( 
.A(n_2057),
.B(n_738),
.Y(n_2378)
);

A2O1A1Ixp33_ASAP7_75t_SL g2379 ( 
.A1(n_2040),
.A2(n_743),
.B(n_744),
.C(n_742),
.Y(n_2379)
);

NAND2xp5_ASAP7_75t_L g2380 ( 
.A(n_2042),
.B(n_200),
.Y(n_2380)
);

AOI22xp33_ASAP7_75t_L g2381 ( 
.A1(n_2051),
.A2(n_203),
.B1(n_201),
.B2(n_202),
.Y(n_2381)
);

O2A1O1Ixp33_ASAP7_75t_L g2382 ( 
.A1(n_2000),
.A2(n_205),
.B(n_201),
.C(n_203),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2039),
.B(n_205),
.Y(n_2383)
);

AOI21xp5_ASAP7_75t_L g2384 ( 
.A1(n_2066),
.A2(n_206),
.B(n_207),
.Y(n_2384)
);

NOR2xp33_ASAP7_75t_R g2385 ( 
.A(n_2066),
.B(n_755),
.Y(n_2385)
);

NAND2xp5_ASAP7_75t_L g2386 ( 
.A(n_1942),
.B(n_208),
.Y(n_2386)
);

AOI22xp5_ASAP7_75t_L g2387 ( 
.A1(n_1896),
.A2(n_211),
.B1(n_209),
.B2(n_210),
.Y(n_2387)
);

AO32x1_ASAP7_75t_L g2388 ( 
.A1(n_2024),
.A2(n_212),
.A3(n_210),
.B1(n_211),
.B2(n_213),
.Y(n_2388)
);

NAND2xp5_ASAP7_75t_L g2389 ( 
.A(n_1883),
.B(n_212),
.Y(n_2389)
);

INVx1_ASAP7_75t_L g2390 ( 
.A(n_1813),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_1813),
.Y(n_2391)
);

NAND2xp5_ASAP7_75t_SL g2392 ( 
.A(n_1871),
.B(n_214),
.Y(n_2392)
);

OAI22xp5_ASAP7_75t_L g2393 ( 
.A1(n_1883),
.A2(n_216),
.B1(n_214),
.B2(n_215),
.Y(n_2393)
);

OAI21xp33_ASAP7_75t_SL g2394 ( 
.A1(n_1933),
.A2(n_215),
.B(n_217),
.Y(n_2394)
);

NOR2xp33_ASAP7_75t_R g2395 ( 
.A(n_2075),
.B(n_748),
.Y(n_2395)
);

OAI22x1_ASAP7_75t_L g2396 ( 
.A1(n_1871),
.A2(n_222),
.B1(n_219),
.B2(n_220),
.Y(n_2396)
);

NAND2xp5_ASAP7_75t_L g2397 ( 
.A(n_1883),
.B(n_219),
.Y(n_2397)
);

HB1xp67_ASAP7_75t_L g2398 ( 
.A(n_2077),
.Y(n_2398)
);

BUFx2_ASAP7_75t_L g2399 ( 
.A(n_2070),
.Y(n_2399)
);

NOR2xp33_ASAP7_75t_L g2400 ( 
.A(n_1851),
.B(n_754),
.Y(n_2400)
);

AO21x1_ASAP7_75t_L g2401 ( 
.A1(n_1933),
.A2(n_220),
.B(n_222),
.Y(n_2401)
);

INVx1_ASAP7_75t_L g2402 ( 
.A(n_1813),
.Y(n_2402)
);

NAND2xp5_ASAP7_75t_L g2403 ( 
.A(n_1883),
.B(n_223),
.Y(n_2403)
);

INVx2_ASAP7_75t_L g2404 ( 
.A(n_1904),
.Y(n_2404)
);

INVx2_ASAP7_75t_SL g2405 ( 
.A(n_1811),
.Y(n_2405)
);

NAND2xp5_ASAP7_75t_SL g2406 ( 
.A(n_1871),
.B(n_224),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_1883),
.B(n_225),
.Y(n_2407)
);

NOR2xp33_ASAP7_75t_L g2408 ( 
.A(n_1851),
.B(n_731),
.Y(n_2408)
);

NAND2xp5_ASAP7_75t_L g2409 ( 
.A(n_1883),
.B(n_228),
.Y(n_2409)
);

INVx2_ASAP7_75t_SL g2410 ( 
.A(n_1811),
.Y(n_2410)
);

NAND3xp33_ASAP7_75t_L g2411 ( 
.A(n_1887),
.B(n_229),
.C(n_230),
.Y(n_2411)
);

OAI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_1883),
.A2(n_234),
.B1(n_231),
.B2(n_232),
.Y(n_2412)
);

A2O1A1Ixp33_ASAP7_75t_L g2413 ( 
.A1(n_1810),
.A2(n_235),
.B(n_232),
.C(n_234),
.Y(n_2413)
);

HB1xp67_ASAP7_75t_L g2414 ( 
.A(n_2077),
.Y(n_2414)
);

BUFx6f_ASAP7_75t_L g2415 ( 
.A(n_1996),
.Y(n_2415)
);

INVx1_ASAP7_75t_L g2416 ( 
.A(n_1813),
.Y(n_2416)
);

INVx2_ASAP7_75t_L g2417 ( 
.A(n_1904),
.Y(n_2417)
);

INVx5_ASAP7_75t_L g2418 ( 
.A(n_2017),
.Y(n_2418)
);

INVx3_ASAP7_75t_SL g2419 ( 
.A(n_2074),
.Y(n_2419)
);

INVx1_ASAP7_75t_L g2420 ( 
.A(n_1813),
.Y(n_2420)
);

INVx1_ASAP7_75t_L g2421 ( 
.A(n_1813),
.Y(n_2421)
);

OR2x2_ASAP7_75t_SL g2422 ( 
.A(n_1906),
.B(n_237),
.Y(n_2422)
);

INVx3_ASAP7_75t_L g2423 ( 
.A(n_1909),
.Y(n_2423)
);

AND2x2_ASAP7_75t_L g2424 ( 
.A(n_1903),
.B(n_237),
.Y(n_2424)
);

O2A1O1Ixp5_ASAP7_75t_L g2425 ( 
.A1(n_1887),
.A2(n_240),
.B(n_238),
.C(n_239),
.Y(n_2425)
);

NAND2xp5_ASAP7_75t_SL g2426 ( 
.A(n_1871),
.B(n_240),
.Y(n_2426)
);

INVx3_ASAP7_75t_L g2427 ( 
.A(n_1909),
.Y(n_2427)
);

INVx3_ASAP7_75t_L g2428 ( 
.A(n_1909),
.Y(n_2428)
);

OR2x2_ASAP7_75t_L g2429 ( 
.A(n_1903),
.B(n_241),
.Y(n_2429)
);

BUFx6f_ASAP7_75t_L g2430 ( 
.A(n_1996),
.Y(n_2430)
);

NOR2xp33_ASAP7_75t_L g2431 ( 
.A(n_1851),
.B(n_729),
.Y(n_2431)
);

O2A1O1Ixp33_ASAP7_75t_L g2432 ( 
.A1(n_1810),
.A2(n_244),
.B(n_242),
.C(n_243),
.Y(n_2432)
);

INVx1_ASAP7_75t_L g2433 ( 
.A(n_1813),
.Y(n_2433)
);

INVx1_ASAP7_75t_L g2434 ( 
.A(n_1813),
.Y(n_2434)
);

NOR2xp33_ASAP7_75t_L g2435 ( 
.A(n_1851),
.B(n_733),
.Y(n_2435)
);

NOR2xp33_ASAP7_75t_L g2436 ( 
.A(n_1851),
.B(n_734),
.Y(n_2436)
);

AO21x1_ASAP7_75t_L g2437 ( 
.A1(n_1933),
.A2(n_245),
.B(n_246),
.Y(n_2437)
);

NAND2xp5_ASAP7_75t_L g2438 ( 
.A(n_1883),
.B(n_247),
.Y(n_2438)
);

NAND2xp5_ASAP7_75t_L g2439 ( 
.A(n_1883),
.B(n_248),
.Y(n_2439)
);

NAND2x1p5_ASAP7_75t_L g2440 ( 
.A(n_1811),
.B(n_250),
.Y(n_2440)
);

NAND2xp5_ASAP7_75t_R g2441 ( 
.A(n_1903),
.B(n_249),
.Y(n_2441)
);

A2O1A1Ixp33_ASAP7_75t_SL g2442 ( 
.A1(n_1887),
.A2(n_746),
.B(n_748),
.C(n_745),
.Y(n_2442)
);

BUFx12f_ASAP7_75t_L g2443 ( 
.A(n_2074),
.Y(n_2443)
);

A2O1A1Ixp33_ASAP7_75t_L g2444 ( 
.A1(n_1810),
.A2(n_252),
.B(n_249),
.C(n_251),
.Y(n_2444)
);

NAND2xp5_ASAP7_75t_L g2445 ( 
.A(n_1883),
.B(n_251),
.Y(n_2445)
);

OAI22xp5_ASAP7_75t_L g2446 ( 
.A1(n_1883),
.A2(n_255),
.B1(n_253),
.B2(n_254),
.Y(n_2446)
);

NAND2xp5_ASAP7_75t_L g2447 ( 
.A(n_1883),
.B(n_253),
.Y(n_2447)
);

INVx2_ASAP7_75t_L g2448 ( 
.A(n_1904),
.Y(n_2448)
);

INVxp67_ASAP7_75t_SL g2449 ( 
.A(n_1896),
.Y(n_2449)
);

AOI22xp33_ASAP7_75t_SL g2450 ( 
.A1(n_1853),
.A2(n_257),
.B1(n_254),
.B2(n_256),
.Y(n_2450)
);

BUFx6f_ASAP7_75t_L g2451 ( 
.A(n_1996),
.Y(n_2451)
);

AOI21xp5_ASAP7_75t_L g2452 ( 
.A1(n_1810),
.A2(n_256),
.B(n_257),
.Y(n_2452)
);

INVx1_ASAP7_75t_L g2453 ( 
.A(n_1813),
.Y(n_2453)
);

INVx1_ASAP7_75t_L g2454 ( 
.A(n_1813),
.Y(n_2454)
);

BUFx6f_ASAP7_75t_L g2455 ( 
.A(n_1996),
.Y(n_2455)
);

NAND2xp5_ASAP7_75t_SL g2456 ( 
.A(n_1871),
.B(n_258),
.Y(n_2456)
);

NAND2xp5_ASAP7_75t_SL g2457 ( 
.A(n_1871),
.B(n_259),
.Y(n_2457)
);

NAND2xp5_ASAP7_75t_L g2458 ( 
.A(n_1883),
.B(n_260),
.Y(n_2458)
);

NAND2xp5_ASAP7_75t_L g2459 ( 
.A(n_1883),
.B(n_260),
.Y(n_2459)
);

BUFx12f_ASAP7_75t_L g2460 ( 
.A(n_2074),
.Y(n_2460)
);

NOR2xp33_ASAP7_75t_L g2461 ( 
.A(n_1851),
.B(n_261),
.Y(n_2461)
);

OAI22xp5_ASAP7_75t_L g2462 ( 
.A1(n_1883),
.A2(n_263),
.B1(n_261),
.B2(n_262),
.Y(n_2462)
);

NOR2x1_ASAP7_75t_L g2463 ( 
.A(n_1810),
.B(n_262),
.Y(n_2463)
);

INVx1_ASAP7_75t_L g2464 ( 
.A(n_1813),
.Y(n_2464)
);

OR2x6_ASAP7_75t_L g2465 ( 
.A(n_1834),
.B(n_264),
.Y(n_2465)
);

NAND2x1p5_ASAP7_75t_L g2466 ( 
.A(n_1811),
.B(n_265),
.Y(n_2466)
);

NAND2xp5_ASAP7_75t_L g2467 ( 
.A(n_1883),
.B(n_265),
.Y(n_2467)
);

OAI22xp5_ASAP7_75t_L g2468 ( 
.A1(n_1883),
.A2(n_268),
.B1(n_266),
.B2(n_267),
.Y(n_2468)
);

NAND2xp33_ASAP7_75t_L g2469 ( 
.A(n_2017),
.B(n_268),
.Y(n_2469)
);

NOR2xp33_ASAP7_75t_L g2470 ( 
.A(n_1851),
.B(n_269),
.Y(n_2470)
);

OR2x2_ASAP7_75t_L g2471 ( 
.A(n_1903),
.B(n_269),
.Y(n_2471)
);

NAND2xp5_ASAP7_75t_SL g2472 ( 
.A(n_1871),
.B(n_270),
.Y(n_2472)
);

BUFx2_ASAP7_75t_L g2473 ( 
.A(n_2070),
.Y(n_2473)
);

A2O1A1Ixp33_ASAP7_75t_SL g2474 ( 
.A1(n_1887),
.A2(n_275),
.B(n_273),
.C(n_274),
.Y(n_2474)
);

INVx1_ASAP7_75t_L g2475 ( 
.A(n_1813),
.Y(n_2475)
);

AND2x2_ASAP7_75t_SL g2476 ( 
.A(n_1853),
.B(n_274),
.Y(n_2476)
);

BUFx2_ASAP7_75t_L g2477 ( 
.A(n_2070),
.Y(n_2477)
);

NAND2x1p5_ASAP7_75t_L g2478 ( 
.A(n_1811),
.B(n_276),
.Y(n_2478)
);

OAI22x1_ASAP7_75t_L g2479 ( 
.A1(n_1871),
.A2(n_278),
.B1(n_276),
.B2(n_277),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_1883),
.B(n_277),
.Y(n_2480)
);

INVx1_ASAP7_75t_L g2481 ( 
.A(n_1813),
.Y(n_2481)
);

NOR2x1_ASAP7_75t_SL g2482 ( 
.A(n_1832),
.B(n_278),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_1837),
.Y(n_2483)
);

OAI22xp5_ASAP7_75t_L g2484 ( 
.A1(n_1883),
.A2(n_282),
.B1(n_280),
.B2(n_281),
.Y(n_2484)
);

AOI21xp5_ASAP7_75t_L g2485 ( 
.A1(n_1810),
.A2(n_280),
.B(n_281),
.Y(n_2485)
);

NAND2xp5_ASAP7_75t_L g2486 ( 
.A(n_1883),
.B(n_282),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_1813),
.Y(n_2487)
);

BUFx6f_ASAP7_75t_L g2488 ( 
.A(n_1996),
.Y(n_2488)
);

BUFx12f_ASAP7_75t_L g2489 ( 
.A(n_2074),
.Y(n_2489)
);

INVx1_ASAP7_75t_SL g2490 ( 
.A(n_2070),
.Y(n_2490)
);

A2O1A1Ixp33_ASAP7_75t_L g2491 ( 
.A1(n_1810),
.A2(n_285),
.B(n_283),
.C(n_284),
.Y(n_2491)
);

INVx2_ASAP7_75t_L g2492 ( 
.A(n_1904),
.Y(n_2492)
);

NAND2xp5_ASAP7_75t_SL g2493 ( 
.A(n_1871),
.B(n_283),
.Y(n_2493)
);

INVx2_ASAP7_75t_L g2494 ( 
.A(n_1904),
.Y(n_2494)
);

OAI22xp5_ASAP7_75t_L g2495 ( 
.A1(n_1883),
.A2(n_286),
.B1(n_284),
.B2(n_285),
.Y(n_2495)
);

NOR2xp33_ASAP7_75t_L g2496 ( 
.A(n_1851),
.B(n_287),
.Y(n_2496)
);

AOI22xp5_ASAP7_75t_L g2497 ( 
.A1(n_1810),
.A2(n_289),
.B1(n_287),
.B2(n_288),
.Y(n_2497)
);

NAND2x1p5_ASAP7_75t_L g2498 ( 
.A(n_1811),
.B(n_289),
.Y(n_2498)
);

AOI21xp5_ASAP7_75t_L g2499 ( 
.A1(n_1810),
.A2(n_291),
.B(n_292),
.Y(n_2499)
);

AOI21xp5_ASAP7_75t_L g2500 ( 
.A1(n_1810),
.A2(n_292),
.B(n_293),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1813),
.Y(n_2501)
);

INVx2_ASAP7_75t_L g2502 ( 
.A(n_1904),
.Y(n_2502)
);

AO32x1_ASAP7_75t_L g2503 ( 
.A1(n_2024),
.A2(n_755),
.A3(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_2503)
);

AOI22xp5_ASAP7_75t_L g2504 ( 
.A1(n_1896),
.A2(n_298),
.B1(n_294),
.B2(n_295),
.Y(n_2504)
);

CKINVDCx20_ASAP7_75t_R g2505 ( 
.A(n_2075),
.Y(n_2505)
);

NOR3xp33_ASAP7_75t_SL g2506 ( 
.A(n_1906),
.B(n_299),
.C(n_301),
.Y(n_2506)
);

AOI22xp5_ASAP7_75t_L g2507 ( 
.A1(n_1896),
.A2(n_302),
.B1(n_299),
.B2(n_301),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_1813),
.Y(n_2508)
);

INVx1_ASAP7_75t_L g2509 ( 
.A(n_1813),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_1813),
.Y(n_2510)
);

AND2x2_ASAP7_75t_L g2511 ( 
.A(n_1903),
.B(n_303),
.Y(n_2511)
);

INVx1_ASAP7_75t_L g2512 ( 
.A(n_1813),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_1813),
.Y(n_2513)
);

OAI21x1_ASAP7_75t_SL g2514 ( 
.A1(n_1933),
.A2(n_304),
.B(n_305),
.Y(n_2514)
);

INVx3_ASAP7_75t_L g2515 ( 
.A(n_1909),
.Y(n_2515)
);

INVx1_ASAP7_75t_L g2516 ( 
.A(n_1813),
.Y(n_2516)
);

NOR2xp33_ASAP7_75t_L g2517 ( 
.A(n_1851),
.B(n_304),
.Y(n_2517)
);

NAND2xp5_ASAP7_75t_SL g2518 ( 
.A(n_1871),
.B(n_305),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_1903),
.B(n_306),
.Y(n_2519)
);

INVx1_ASAP7_75t_SL g2520 ( 
.A(n_2070),
.Y(n_2520)
);

INVx1_ASAP7_75t_SL g2521 ( 
.A(n_2070),
.Y(n_2521)
);

NAND2xp5_ASAP7_75t_L g2522 ( 
.A(n_1883),
.B(n_307),
.Y(n_2522)
);

INVx2_ASAP7_75t_L g2523 ( 
.A(n_1904),
.Y(n_2523)
);

NAND2xp5_ASAP7_75t_L g2524 ( 
.A(n_1883),
.B(n_308),
.Y(n_2524)
);

OAI22xp5_ASAP7_75t_L g2525 ( 
.A1(n_1883),
.A2(n_311),
.B1(n_309),
.B2(n_310),
.Y(n_2525)
);

CKINVDCx5p33_ASAP7_75t_R g2526 ( 
.A(n_1837),
.Y(n_2526)
);

AO31x2_ASAP7_75t_L g2527 ( 
.A1(n_1950),
.A2(n_312),
.A3(n_309),
.B(n_311),
.Y(n_2527)
);

O2A1O1Ixp33_ASAP7_75t_L g2528 ( 
.A1(n_1810),
.A2(n_315),
.B(n_312),
.C(n_313),
.Y(n_2528)
);

NAND2xp5_ASAP7_75t_SL g2529 ( 
.A(n_1871),
.B(n_315),
.Y(n_2529)
);

NAND3xp33_ASAP7_75t_SL g2530 ( 
.A(n_1837),
.B(n_316),
.C(n_318),
.Y(n_2530)
);

NAND2xp5_ASAP7_75t_SL g2531 ( 
.A(n_1871),
.B(n_319),
.Y(n_2531)
);

AOI22xp5_ASAP7_75t_L g2532 ( 
.A1(n_1896),
.A2(n_322),
.B1(n_319),
.B2(n_320),
.Y(n_2532)
);

BUFx6f_ASAP7_75t_L g2533 ( 
.A(n_1996),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_SL g2534 ( 
.A(n_1871),
.B(n_320),
.Y(n_2534)
);

OAI22xp5_ASAP7_75t_L g2535 ( 
.A1(n_1883),
.A2(n_324),
.B1(n_322),
.B2(n_323),
.Y(n_2535)
);

AOI21x1_ASAP7_75t_L g2536 ( 
.A1(n_2058),
.A2(n_323),
.B(n_325),
.Y(n_2536)
);

AO32x2_ASAP7_75t_L g2537 ( 
.A1(n_1976),
.A2(n_329),
.A3(n_326),
.B1(n_328),
.B2(n_330),
.Y(n_2537)
);

INVx3_ASAP7_75t_L g2538 ( 
.A(n_1909),
.Y(n_2538)
);

INVx1_ASAP7_75t_L g2539 ( 
.A(n_1813),
.Y(n_2539)
);

HB1xp67_ASAP7_75t_L g2540 ( 
.A(n_2077),
.Y(n_2540)
);

NAND2xp5_ASAP7_75t_L g2541 ( 
.A(n_1883),
.B(n_332),
.Y(n_2541)
);

INVx2_ASAP7_75t_L g2542 ( 
.A(n_1904),
.Y(n_2542)
);

NAND2xp5_ASAP7_75t_L g2543 ( 
.A(n_1883),
.B(n_332),
.Y(n_2543)
);

AND2x6_ASAP7_75t_L g2544 ( 
.A(n_1909),
.B(n_333),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_1813),
.Y(n_2545)
);

OAI22x1_ASAP7_75t_L g2546 ( 
.A1(n_1871),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2546)
);

NAND2xp5_ASAP7_75t_L g2547 ( 
.A(n_1883),
.B(n_336),
.Y(n_2547)
);

INVx2_ASAP7_75t_SL g2548 ( 
.A(n_1811),
.Y(n_2548)
);

INVx2_ASAP7_75t_L g2549 ( 
.A(n_1904),
.Y(n_2549)
);

NOR2xp67_ASAP7_75t_SL g2550 ( 
.A(n_1888),
.B(n_336),
.Y(n_2550)
);

NOR2xp33_ASAP7_75t_L g2551 ( 
.A(n_1851),
.B(n_337),
.Y(n_2551)
);

NOR2xp67_ASAP7_75t_L g2552 ( 
.A(n_1948),
.B(n_752),
.Y(n_2552)
);

BUFx6f_ASAP7_75t_L g2553 ( 
.A(n_1996),
.Y(n_2553)
);

NAND2xp5_ASAP7_75t_L g2554 ( 
.A(n_1883),
.B(n_337),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_1904),
.Y(n_2555)
);

NOR2x1_ASAP7_75t_L g2556 ( 
.A(n_1810),
.B(n_338),
.Y(n_2556)
);

INVx2_ASAP7_75t_L g2557 ( 
.A(n_1904),
.Y(n_2557)
);

AOI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_1810),
.A2(n_341),
.B1(n_339),
.B2(n_340),
.Y(n_2558)
);

NOR2xp33_ASAP7_75t_L g2559 ( 
.A(n_1851),
.B(n_341),
.Y(n_2559)
);

OR2x2_ASAP7_75t_L g2560 ( 
.A(n_1903),
.B(n_342),
.Y(n_2560)
);

A2O1A1Ixp33_ASAP7_75t_L g2561 ( 
.A1(n_1810),
.A2(n_344),
.B(n_342),
.C(n_343),
.Y(n_2561)
);

AO221x2_ASAP7_75t_L g2562 ( 
.A1(n_1911),
.A2(n_345),
.B1(n_343),
.B2(n_344),
.C(n_346),
.Y(n_2562)
);

NAND2xp5_ASAP7_75t_L g2563 ( 
.A(n_1883),
.B(n_347),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_1813),
.Y(n_2564)
);

AND2x4_ASAP7_75t_L g2565 ( 
.A(n_1984),
.B(n_348),
.Y(n_2565)
);

NAND2xp5_ASAP7_75t_SL g2566 ( 
.A(n_1871),
.B(n_348),
.Y(n_2566)
);

INVx5_ASAP7_75t_L g2567 ( 
.A(n_2544),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2112),
.Y(n_2568)
);

INVx3_ASAP7_75t_L g2569 ( 
.A(n_2159),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2424),
.B(n_349),
.Y(n_2570)
);

BUFx2_ASAP7_75t_SL g2571 ( 
.A(n_2128),
.Y(n_2571)
);

INVx8_ASAP7_75t_L g2572 ( 
.A(n_2544),
.Y(n_2572)
);

INVx1_ASAP7_75t_L g2573 ( 
.A(n_2126),
.Y(n_2573)
);

BUFx6f_ASAP7_75t_L g2574 ( 
.A(n_2187),
.Y(n_2574)
);

AND2x4_ASAP7_75t_L g2575 ( 
.A(n_2166),
.B(n_350),
.Y(n_2575)
);

INVx5_ASAP7_75t_SL g2576 ( 
.A(n_2465),
.Y(n_2576)
);

INVx6_ASAP7_75t_SL g2577 ( 
.A(n_2465),
.Y(n_2577)
);

CKINVDCx20_ASAP7_75t_R g2578 ( 
.A(n_2312),
.Y(n_2578)
);

OAI21x1_ASAP7_75t_L g2579 ( 
.A1(n_2186),
.A2(n_352),
.B(n_353),
.Y(n_2579)
);

AND2x2_ASAP7_75t_L g2580 ( 
.A(n_2511),
.B(n_352),
.Y(n_2580)
);

INVx1_ASAP7_75t_L g2581 ( 
.A(n_2404),
.Y(n_2581)
);

INVx3_ASAP7_75t_L g2582 ( 
.A(n_2159),
.Y(n_2582)
);

INVx1_ASAP7_75t_L g2583 ( 
.A(n_2417),
.Y(n_2583)
);

INVx2_ASAP7_75t_L g2584 ( 
.A(n_2448),
.Y(n_2584)
);

INVxp67_ASAP7_75t_SL g2585 ( 
.A(n_2320),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2492),
.Y(n_2586)
);

BUFx12f_ASAP7_75t_L g2587 ( 
.A(n_2303),
.Y(n_2587)
);

NOR2x1_ASAP7_75t_SL g2588 ( 
.A(n_2418),
.B(n_353),
.Y(n_2588)
);

INVx1_ASAP7_75t_SL g2589 ( 
.A(n_2124),
.Y(n_2589)
);

OAI21x1_ASAP7_75t_L g2590 ( 
.A1(n_2202),
.A2(n_357),
.B(n_358),
.Y(n_2590)
);

INVx6_ASAP7_75t_L g2591 ( 
.A(n_2290),
.Y(n_2591)
);

INVx6_ASAP7_75t_L g2592 ( 
.A(n_2290),
.Y(n_2592)
);

INVx2_ASAP7_75t_L g2593 ( 
.A(n_2494),
.Y(n_2593)
);

INVx2_ASAP7_75t_L g2594 ( 
.A(n_2502),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2523),
.Y(n_2595)
);

AO21x2_ASAP7_75t_L g2596 ( 
.A1(n_2514),
.A2(n_358),
.B(n_359),
.Y(n_2596)
);

INVx3_ASAP7_75t_L g2597 ( 
.A(n_2215),
.Y(n_2597)
);

AND2x4_ASAP7_75t_L g2598 ( 
.A(n_2128),
.B(n_360),
.Y(n_2598)
);

NAND2xp5_ASAP7_75t_L g2599 ( 
.A(n_2095),
.B(n_361),
.Y(n_2599)
);

INVx1_ASAP7_75t_L g2600 ( 
.A(n_2542),
.Y(n_2600)
);

INVx1_ASAP7_75t_L g2601 ( 
.A(n_2549),
.Y(n_2601)
);

BUFx5_ASAP7_75t_L g2602 ( 
.A(n_2544),
.Y(n_2602)
);

INVx1_ASAP7_75t_L g2603 ( 
.A(n_2555),
.Y(n_2603)
);

NAND2x1p5_ASAP7_75t_L g2604 ( 
.A(n_2418),
.B(n_362),
.Y(n_2604)
);

NAND2x1p5_ASAP7_75t_L g2605 ( 
.A(n_2418),
.B(n_2215),
.Y(n_2605)
);

AND2x2_ASAP7_75t_L g2606 ( 
.A(n_2519),
.B(n_362),
.Y(n_2606)
);

OR2x2_ASAP7_75t_L g2607 ( 
.A(n_2429),
.B(n_2471),
.Y(n_2607)
);

NOR2x1_ASAP7_75t_SL g2608 ( 
.A(n_2323),
.B(n_363),
.Y(n_2608)
);

INVx3_ASAP7_75t_L g2609 ( 
.A(n_2221),
.Y(n_2609)
);

NAND2x1p5_ASAP7_75t_L g2610 ( 
.A(n_2221),
.B(n_365),
.Y(n_2610)
);

HB1xp67_ASAP7_75t_L g2611 ( 
.A(n_2246),
.Y(n_2611)
);

CKINVDCx20_ASAP7_75t_R g2612 ( 
.A(n_2505),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2557),
.Y(n_2613)
);

OA21x2_ASAP7_75t_L g2614 ( 
.A1(n_2184),
.A2(n_365),
.B(n_366),
.Y(n_2614)
);

BUFx12f_ASAP7_75t_L g2615 ( 
.A(n_2181),
.Y(n_2615)
);

OAI21x1_ASAP7_75t_L g2616 ( 
.A1(n_2173),
.A2(n_366),
.B(n_367),
.Y(n_2616)
);

BUFx3_ASAP7_75t_L g2617 ( 
.A(n_2121),
.Y(n_2617)
);

BUFx12f_ASAP7_75t_L g2618 ( 
.A(n_2130),
.Y(n_2618)
);

NOR2xp33_ASAP7_75t_L g2619 ( 
.A(n_2092),
.B(n_2449),
.Y(n_2619)
);

OAI21x1_ASAP7_75t_SL g2620 ( 
.A1(n_2323),
.A2(n_367),
.B(n_368),
.Y(n_2620)
);

INVx1_ASAP7_75t_L g2621 ( 
.A(n_2099),
.Y(n_2621)
);

NAND2xp5_ASAP7_75t_L g2622 ( 
.A(n_2105),
.B(n_368),
.Y(n_2622)
);

OR3x4_ASAP7_75t_SL g2623 ( 
.A(n_2330),
.B(n_369),
.C(n_370),
.Y(n_2623)
);

INVx2_ASAP7_75t_L g2624 ( 
.A(n_2353),
.Y(n_2624)
);

NAND2xp5_ASAP7_75t_L g2625 ( 
.A(n_2106),
.B(n_369),
.Y(n_2625)
);

CKINVDCx20_ASAP7_75t_R g2626 ( 
.A(n_2310),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2120),
.Y(n_2627)
);

OA21x2_ASAP7_75t_L g2628 ( 
.A1(n_2425),
.A2(n_371),
.B(n_372),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2131),
.Y(n_2629)
);

AO21x2_ASAP7_75t_L g2630 ( 
.A1(n_2442),
.A2(n_372),
.B(n_373),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2390),
.Y(n_2631)
);

HB1xp67_ASAP7_75t_L g2632 ( 
.A(n_2246),
.Y(n_2632)
);

HB1xp67_ASAP7_75t_L g2633 ( 
.A(n_2246),
.Y(n_2633)
);

INVx2_ASAP7_75t_L g2634 ( 
.A(n_2391),
.Y(n_2634)
);

OAI21x1_ASAP7_75t_L g2635 ( 
.A1(n_2177),
.A2(n_377),
.B(n_378),
.Y(n_2635)
);

OAI21x1_ASAP7_75t_L g2636 ( 
.A1(n_2091),
.A2(n_377),
.B(n_379),
.Y(n_2636)
);

INVx1_ASAP7_75t_L g2637 ( 
.A(n_2402),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2416),
.B(n_380),
.Y(n_2638)
);

CKINVDCx5p33_ASAP7_75t_R g2639 ( 
.A(n_2191),
.Y(n_2639)
);

CKINVDCx20_ASAP7_75t_R g2640 ( 
.A(n_2096),
.Y(n_2640)
);

INVx1_ASAP7_75t_L g2641 ( 
.A(n_2420),
.Y(n_2641)
);

INVx1_ASAP7_75t_L g2642 ( 
.A(n_2421),
.Y(n_2642)
);

INVx3_ASAP7_75t_L g2643 ( 
.A(n_2268),
.Y(n_2643)
);

HB1xp67_ASAP7_75t_L g2644 ( 
.A(n_2268),
.Y(n_2644)
);

INVx4_ASAP7_75t_L g2645 ( 
.A(n_2191),
.Y(n_2645)
);

AND2x4_ASAP7_75t_L g2646 ( 
.A(n_2308),
.B(n_382),
.Y(n_2646)
);

BUFx2_ASAP7_75t_L g2647 ( 
.A(n_2098),
.Y(n_2647)
);

INVxp67_ASAP7_75t_SL g2648 ( 
.A(n_2268),
.Y(n_2648)
);

INVx5_ASAP7_75t_L g2649 ( 
.A(n_2544),
.Y(n_2649)
);

BUFx2_ASAP7_75t_R g2650 ( 
.A(n_2483),
.Y(n_2650)
);

INVx2_ASAP7_75t_L g2651 ( 
.A(n_2433),
.Y(n_2651)
);

BUFx2_ASAP7_75t_SL g2652 ( 
.A(n_2405),
.Y(n_2652)
);

BUFx3_ASAP7_75t_L g2653 ( 
.A(n_2277),
.Y(n_2653)
);

INVx3_ASAP7_75t_L g2654 ( 
.A(n_2227),
.Y(n_2654)
);

INVx1_ASAP7_75t_L g2655 ( 
.A(n_2434),
.Y(n_2655)
);

HB1xp67_ASAP7_75t_L g2656 ( 
.A(n_2291),
.Y(n_2656)
);

OA21x2_ASAP7_75t_L g2657 ( 
.A1(n_2333),
.A2(n_2335),
.B(n_2188),
.Y(n_2657)
);

BUFx3_ASAP7_75t_L g2658 ( 
.A(n_2277),
.Y(n_2658)
);

INVx1_ASAP7_75t_L g2659 ( 
.A(n_2453),
.Y(n_2659)
);

AO21x2_ASAP7_75t_L g2660 ( 
.A1(n_2474),
.A2(n_383),
.B(n_384),
.Y(n_2660)
);

AO21x2_ASAP7_75t_L g2661 ( 
.A1(n_2144),
.A2(n_383),
.B(n_385),
.Y(n_2661)
);

AND2x2_ASAP7_75t_L g2662 ( 
.A(n_2476),
.B(n_386),
.Y(n_2662)
);

AND2x2_ASAP7_75t_L g2663 ( 
.A(n_2201),
.B(n_386),
.Y(n_2663)
);

OAI21x1_ASAP7_75t_L g2664 ( 
.A1(n_2134),
.A2(n_387),
.B(n_388),
.Y(n_2664)
);

INVx2_ASAP7_75t_SL g2665 ( 
.A(n_2374),
.Y(n_2665)
);

AO21x2_ASAP7_75t_L g2666 ( 
.A1(n_2401),
.A2(n_387),
.B(n_389),
.Y(n_2666)
);

CKINVDCx5p33_ASAP7_75t_R g2667 ( 
.A(n_2316),
.Y(n_2667)
);

INVxp67_ASAP7_75t_SL g2668 ( 
.A(n_2295),
.Y(n_2668)
);

OR2x6_ASAP7_75t_L g2669 ( 
.A(n_2225),
.B(n_391),
.Y(n_2669)
);

BUFx12f_ASAP7_75t_L g2670 ( 
.A(n_2443),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2454),
.Y(n_2671)
);

CKINVDCx16_ASAP7_75t_R g2672 ( 
.A(n_2122),
.Y(n_2672)
);

BUFx8_ASAP7_75t_SL g2673 ( 
.A(n_2460),
.Y(n_2673)
);

OR2x6_ASAP7_75t_L g2674 ( 
.A(n_2285),
.B(n_393),
.Y(n_2674)
);

OAI21xp5_ASAP7_75t_L g2675 ( 
.A1(n_2289),
.A2(n_394),
.B(n_395),
.Y(n_2675)
);

OAI21xp5_ASAP7_75t_L g2676 ( 
.A1(n_2152),
.A2(n_394),
.B(n_397),
.Y(n_2676)
);

INVx1_ASAP7_75t_L g2677 ( 
.A(n_2464),
.Y(n_2677)
);

INVxp67_ASAP7_75t_L g2678 ( 
.A(n_2398),
.Y(n_2678)
);

INVx2_ASAP7_75t_L g2679 ( 
.A(n_2475),
.Y(n_2679)
);

OAI21x1_ASAP7_75t_L g2680 ( 
.A1(n_2145),
.A2(n_2194),
.B(n_2164),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2481),
.Y(n_2681)
);

INVx2_ASAP7_75t_SL g2682 ( 
.A(n_2374),
.Y(n_2682)
);

NAND2x1p5_ASAP7_75t_L g2683 ( 
.A(n_2291),
.B(n_398),
.Y(n_2683)
);

AO21x2_ASAP7_75t_L g2684 ( 
.A1(n_2437),
.A2(n_399),
.B(n_400),
.Y(n_2684)
);

NAND2xp5_ASAP7_75t_L g2685 ( 
.A(n_2487),
.B(n_400),
.Y(n_2685)
);

INVx3_ASAP7_75t_SL g2686 ( 
.A(n_2419),
.Y(n_2686)
);

AO21x2_ASAP7_75t_L g2687 ( 
.A1(n_2379),
.A2(n_401),
.B(n_402),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2501),
.Y(n_2688)
);

BUFx3_ASAP7_75t_L g2689 ( 
.A(n_2399),
.Y(n_2689)
);

OAI21x1_ASAP7_75t_L g2690 ( 
.A1(n_2423),
.A2(n_401),
.B(n_402),
.Y(n_2690)
);

INVx2_ASAP7_75t_L g2691 ( 
.A(n_2508),
.Y(n_2691)
);

AND2x6_ASAP7_75t_L g2692 ( 
.A(n_2295),
.B(n_752),
.Y(n_2692)
);

AND2x4_ASAP7_75t_L g2693 ( 
.A(n_2308),
.B(n_403),
.Y(n_2693)
);

INVx1_ASAP7_75t_L g2694 ( 
.A(n_2509),
.Y(n_2694)
);

BUFx2_ASAP7_75t_L g2695 ( 
.A(n_2473),
.Y(n_2695)
);

OAI21x1_ASAP7_75t_L g2696 ( 
.A1(n_2423),
.A2(n_403),
.B(n_404),
.Y(n_2696)
);

BUFx2_ASAP7_75t_L g2697 ( 
.A(n_2477),
.Y(n_2697)
);

INVx2_ASAP7_75t_L g2698 ( 
.A(n_2510),
.Y(n_2698)
);

OAI21x1_ASAP7_75t_L g2699 ( 
.A1(n_2427),
.A2(n_2515),
.B(n_2428),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2512),
.Y(n_2700)
);

OAI21x1_ASAP7_75t_L g2701 ( 
.A1(n_2427),
.A2(n_404),
.B(n_405),
.Y(n_2701)
);

AND2x4_ASAP7_75t_L g2702 ( 
.A(n_2565),
.B(n_408),
.Y(n_2702)
);

BUFx3_ASAP7_75t_L g2703 ( 
.A(n_2489),
.Y(n_2703)
);

OR3x4_ASAP7_75t_SL g2704 ( 
.A(n_2562),
.B(n_409),
.C(n_410),
.Y(n_2704)
);

AND2x4_ASAP7_75t_L g2705 ( 
.A(n_2565),
.B(n_409),
.Y(n_2705)
);

AO21x2_ASAP7_75t_L g2706 ( 
.A1(n_2102),
.A2(n_410),
.B(n_413),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2513),
.Y(n_2707)
);

CKINVDCx14_ASAP7_75t_R g2708 ( 
.A(n_2125),
.Y(n_2708)
);

NAND2xp5_ASAP7_75t_SL g2709 ( 
.A(n_2291),
.B(n_414),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2516),
.Y(n_2710)
);

INVx3_ASAP7_75t_L g2711 ( 
.A(n_2227),
.Y(n_2711)
);

NAND2x1p5_ASAP7_75t_L g2712 ( 
.A(n_2247),
.B(n_415),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2539),
.Y(n_2713)
);

INVx2_ASAP7_75t_SL g2714 ( 
.A(n_2162),
.Y(n_2714)
);

AO21x2_ASAP7_75t_L g2715 ( 
.A1(n_2233),
.A2(n_415),
.B(n_416),
.Y(n_2715)
);

NAND2x1p5_ASAP7_75t_L g2716 ( 
.A(n_2295),
.B(n_417),
.Y(n_2716)
);

NAND2x1p5_ASAP7_75t_L g2717 ( 
.A(n_2326),
.B(n_417),
.Y(n_2717)
);

AOI21xp5_ASAP7_75t_L g2718 ( 
.A1(n_2205),
.A2(n_418),
.B(n_419),
.Y(n_2718)
);

AO21x2_ASAP7_75t_L g2719 ( 
.A1(n_2536),
.A2(n_418),
.B(n_420),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2104),
.B(n_421),
.Y(n_2720)
);

BUFx4f_ASAP7_75t_L g2721 ( 
.A(n_2288),
.Y(n_2721)
);

AND2x2_ASAP7_75t_L g2722 ( 
.A(n_2560),
.B(n_421),
.Y(n_2722)
);

HB1xp67_ASAP7_75t_L g2723 ( 
.A(n_2236),
.Y(n_2723)
);

HB1xp67_ASAP7_75t_L g2724 ( 
.A(n_2236),
.Y(n_2724)
);

INVx1_ASAP7_75t_L g2725 ( 
.A(n_2545),
.Y(n_2725)
);

INVx8_ASAP7_75t_L g2726 ( 
.A(n_2285),
.Y(n_2726)
);

BUFx12f_ASAP7_75t_L g2727 ( 
.A(n_2526),
.Y(n_2727)
);

INVx8_ASAP7_75t_L g2728 ( 
.A(n_2288),
.Y(n_2728)
);

BUFx3_ASAP7_75t_L g2729 ( 
.A(n_2328),
.Y(n_2729)
);

BUFx3_ASAP7_75t_L g2730 ( 
.A(n_2346),
.Y(n_2730)
);

INVx1_ASAP7_75t_L g2731 ( 
.A(n_2564),
.Y(n_2731)
);

AND2x2_ASAP7_75t_SL g2732 ( 
.A(n_2469),
.B(n_746),
.Y(n_2732)
);

CKINVDCx20_ASAP7_75t_R g2733 ( 
.A(n_2395),
.Y(n_2733)
);

INVx4_ASAP7_75t_L g2734 ( 
.A(n_2162),
.Y(n_2734)
);

AO21x2_ASAP7_75t_L g2735 ( 
.A1(n_2224),
.A2(n_424),
.B(n_425),
.Y(n_2735)
);

INVx1_ASAP7_75t_L g2736 ( 
.A(n_2138),
.Y(n_2736)
);

CKINVDCx5p33_ASAP7_75t_R g2737 ( 
.A(n_2141),
.Y(n_2737)
);

INVx1_ASAP7_75t_L g2738 ( 
.A(n_2139),
.Y(n_2738)
);

AND2x2_ASAP7_75t_L g2739 ( 
.A(n_2363),
.B(n_426),
.Y(n_2739)
);

OR2x6_ASAP7_75t_L g2740 ( 
.A(n_2363),
.B(n_427),
.Y(n_2740)
);

INVx1_ASAP7_75t_SL g2741 ( 
.A(n_2490),
.Y(n_2741)
);

BUFx10_ASAP7_75t_L g2742 ( 
.A(n_2410),
.Y(n_2742)
);

INVx2_ASAP7_75t_SL g2743 ( 
.A(n_2548),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2207),
.B(n_430),
.Y(n_2744)
);

INVx2_ASAP7_75t_L g2745 ( 
.A(n_2143),
.Y(n_2745)
);

OAI21x1_ASAP7_75t_L g2746 ( 
.A1(n_2538),
.A2(n_430),
.B(n_432),
.Y(n_2746)
);

OAI21x1_ASAP7_75t_L g2747 ( 
.A1(n_2183),
.A2(n_432),
.B(n_433),
.Y(n_2747)
);

INVx1_ASAP7_75t_L g2748 ( 
.A(n_2204),
.Y(n_2748)
);

BUFx3_ASAP7_75t_L g2749 ( 
.A(n_2110),
.Y(n_2749)
);

NOR2xp33_ASAP7_75t_L g2750 ( 
.A(n_2321),
.B(n_434),
.Y(n_2750)
);

OAI21x1_ASAP7_75t_L g2751 ( 
.A1(n_2169),
.A2(n_2556),
.B(n_2463),
.Y(n_2751)
);

AND2x4_ASAP7_75t_L g2752 ( 
.A(n_2235),
.B(n_435),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2146),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2213),
.Y(n_2754)
);

NOR2xp67_ASAP7_75t_SL g2755 ( 
.A(n_2331),
.B(n_435),
.Y(n_2755)
);

INVx2_ASAP7_75t_L g2756 ( 
.A(n_2149),
.Y(n_2756)
);

HB1xp67_ASAP7_75t_L g2757 ( 
.A(n_2119),
.Y(n_2757)
);

BUFx3_ASAP7_75t_L g2758 ( 
.A(n_2520),
.Y(n_2758)
);

BUFx4f_ASAP7_75t_SL g2759 ( 
.A(n_2521),
.Y(n_2759)
);

INVx3_ASAP7_75t_L g2760 ( 
.A(n_2235),
.Y(n_2760)
);

BUFx3_ASAP7_75t_L g2761 ( 
.A(n_2414),
.Y(n_2761)
);

INVx3_ASAP7_75t_L g2762 ( 
.A(n_2251),
.Y(n_2762)
);

OAI21x1_ASAP7_75t_L g2763 ( 
.A1(n_2463),
.A2(n_437),
.B(n_438),
.Y(n_2763)
);

INVx3_ASAP7_75t_L g2764 ( 
.A(n_2251),
.Y(n_2764)
);

NOR2xp33_ASAP7_75t_L g2765 ( 
.A(n_2292),
.B(n_439),
.Y(n_2765)
);

AOI22x1_ASAP7_75t_L g2766 ( 
.A1(n_2322),
.A2(n_443),
.B1(n_441),
.B2(n_442),
.Y(n_2766)
);

CKINVDCx16_ASAP7_75t_R g2767 ( 
.A(n_2276),
.Y(n_2767)
);

INVx1_ASAP7_75t_L g2768 ( 
.A(n_2217),
.Y(n_2768)
);

INVx6_ASAP7_75t_L g2769 ( 
.A(n_2351),
.Y(n_2769)
);

OAI21x1_ASAP7_75t_L g2770 ( 
.A1(n_2556),
.A2(n_441),
.B(n_442),
.Y(n_2770)
);

BUFx3_ASAP7_75t_L g2771 ( 
.A(n_2540),
.Y(n_2771)
);

BUFx3_ASAP7_75t_L g2772 ( 
.A(n_2245),
.Y(n_2772)
);

BUFx3_ASAP7_75t_L g2773 ( 
.A(n_2234),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2171),
.Y(n_2774)
);

AO21x1_ASAP7_75t_L g2775 ( 
.A1(n_2382),
.A2(n_443),
.B(n_444),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2161),
.Y(n_2776)
);

AO21x2_ASAP7_75t_L g2777 ( 
.A1(n_2107),
.A2(n_444),
.B(n_445),
.Y(n_2777)
);

CKINVDCx6p67_ASAP7_75t_R g2778 ( 
.A(n_2275),
.Y(n_2778)
);

INVx2_ASAP7_75t_SL g2779 ( 
.A(n_2351),
.Y(n_2779)
);

CKINVDCx20_ASAP7_75t_R g2780 ( 
.A(n_2343),
.Y(n_2780)
);

AOI22x1_ASAP7_75t_L g2781 ( 
.A1(n_2327),
.A2(n_448),
.B1(n_445),
.B2(n_447),
.Y(n_2781)
);

AND2x4_ASAP7_75t_L g2782 ( 
.A(n_2223),
.B(n_449),
.Y(n_2782)
);

NAND2x1p5_ASAP7_75t_L g2783 ( 
.A(n_2136),
.B(n_450),
.Y(n_2783)
);

INVx3_ASAP7_75t_SL g2784 ( 
.A(n_2278),
.Y(n_2784)
);

BUFx5_ASAP7_75t_L g2785 ( 
.A(n_2238),
.Y(n_2785)
);

NAND2xp5_ASAP7_75t_L g2786 ( 
.A(n_2261),
.B(n_451),
.Y(n_2786)
);

INVx1_ASAP7_75t_L g2787 ( 
.A(n_2218),
.Y(n_2787)
);

BUFx3_ASAP7_75t_L g2788 ( 
.A(n_2372),
.Y(n_2788)
);

BUFx2_ASAP7_75t_R g2789 ( 
.A(n_2157),
.Y(n_2789)
);

INVx5_ASAP7_75t_SL g2790 ( 
.A(n_2265),
.Y(n_2790)
);

OR2x6_ASAP7_75t_L g2791 ( 
.A(n_2440),
.B(n_452),
.Y(n_2791)
);

BUFx3_ASAP7_75t_L g2792 ( 
.A(n_2309),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2339),
.Y(n_2793)
);

AND2x4_ASAP7_75t_L g2794 ( 
.A(n_2299),
.B(n_453),
.Y(n_2794)
);

OAI21x1_ASAP7_75t_L g2795 ( 
.A1(n_2373),
.A2(n_453),
.B(n_454),
.Y(n_2795)
);

INVx2_ASAP7_75t_SL g2796 ( 
.A(n_2351),
.Y(n_2796)
);

AOI21x1_ASAP7_75t_L g2797 ( 
.A1(n_2313),
.A2(n_454),
.B(n_455),
.Y(n_2797)
);

AND2x2_ASAP7_75t_L g2798 ( 
.A(n_2210),
.B(n_455),
.Y(n_2798)
);

NOR2xp33_ASAP7_75t_L g2799 ( 
.A(n_2165),
.B(n_456),
.Y(n_2799)
);

INVx1_ASAP7_75t_L g2800 ( 
.A(n_2304),
.Y(n_2800)
);

NAND2x1p5_ASAP7_75t_L g2801 ( 
.A(n_2415),
.B(n_457),
.Y(n_2801)
);

NOR2xp33_ASAP7_75t_L g2802 ( 
.A(n_2317),
.B(n_457),
.Y(n_2802)
);

BUFx12f_ASAP7_75t_L g2803 ( 
.A(n_2466),
.Y(n_2803)
);

BUFx2_ASAP7_75t_SL g2804 ( 
.A(n_2552),
.Y(n_2804)
);

BUFx3_ASAP7_75t_L g2805 ( 
.A(n_2344),
.Y(n_2805)
);

INVx2_ASAP7_75t_L g2806 ( 
.A(n_2196),
.Y(n_2806)
);

BUFx3_ASAP7_75t_L g2807 ( 
.A(n_2344),
.Y(n_2807)
);

AO21x2_ASAP7_75t_L g2808 ( 
.A1(n_2222),
.A2(n_458),
.B(n_460),
.Y(n_2808)
);

BUFx2_ASAP7_75t_SL g2809 ( 
.A(n_2552),
.Y(n_2809)
);

OAI21x1_ASAP7_75t_L g2810 ( 
.A1(n_2373),
.A2(n_461),
.B(n_462),
.Y(n_2810)
);

BUFx2_ASAP7_75t_L g2811 ( 
.A(n_2229),
.Y(n_2811)
);

AO21x2_ASAP7_75t_L g2812 ( 
.A1(n_2228),
.A2(n_461),
.B(n_463),
.Y(n_2812)
);

AOI22x1_ASAP7_75t_L g2813 ( 
.A1(n_2329),
.A2(n_465),
.B1(n_463),
.B2(n_464),
.Y(n_2813)
);

AND2x4_ASAP7_75t_L g2814 ( 
.A(n_2334),
.B(n_464),
.Y(n_2814)
);

AO21x2_ASAP7_75t_L g2815 ( 
.A1(n_2231),
.A2(n_465),
.B(n_466),
.Y(n_2815)
);

BUFx3_ASAP7_75t_L g2816 ( 
.A(n_2344),
.Y(n_2816)
);

AND2x4_ASAP7_75t_L g2817 ( 
.A(n_2362),
.B(n_466),
.Y(n_2817)
);

INVx2_ASAP7_75t_L g2818 ( 
.A(n_2220),
.Y(n_2818)
);

BUFx2_ASAP7_75t_L g2819 ( 
.A(n_2284),
.Y(n_2819)
);

OAI21x1_ASAP7_75t_SL g2820 ( 
.A1(n_2482),
.A2(n_467),
.B(n_468),
.Y(n_2820)
);

INVx5_ASAP7_75t_L g2821 ( 
.A(n_2238),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2359),
.Y(n_2822)
);

INVx2_ASAP7_75t_L g2823 ( 
.A(n_2230),
.Y(n_2823)
);

CKINVDCx20_ASAP7_75t_R g2824 ( 
.A(n_2385),
.Y(n_2824)
);

AO21x2_ASAP7_75t_L g2825 ( 
.A1(n_2244),
.A2(n_467),
.B(n_468),
.Y(n_2825)
);

INVxp67_ASAP7_75t_SL g2826 ( 
.A(n_2430),
.Y(n_2826)
);

OAI21x1_ASAP7_75t_L g2827 ( 
.A1(n_2384),
.A2(n_470),
.B(n_471),
.Y(n_2827)
);

HB1xp67_ASAP7_75t_L g2828 ( 
.A(n_2293),
.Y(n_2828)
);

OAI21xp5_ASAP7_75t_L g2829 ( 
.A1(n_2118),
.A2(n_470),
.B(n_472),
.Y(n_2829)
);

CKINVDCx11_ASAP7_75t_R g2830 ( 
.A(n_2198),
.Y(n_2830)
);

BUFx2_ASAP7_75t_SL g2831 ( 
.A(n_2238),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2209),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2219),
.B(n_472),
.Y(n_2833)
);

AO21x2_ASAP7_75t_L g2834 ( 
.A1(n_2111),
.A2(n_473),
.B(n_474),
.Y(n_2834)
);

INVx1_ASAP7_75t_SL g2835 ( 
.A(n_2172),
.Y(n_2835)
);

INVx1_ASAP7_75t_L g2836 ( 
.A(n_2441),
.Y(n_2836)
);

OAI21x1_ASAP7_75t_L g2837 ( 
.A1(n_2349),
.A2(n_475),
.B(n_476),
.Y(n_2837)
);

BUFx5_ASAP7_75t_L g2838 ( 
.A(n_2238),
.Y(n_2838)
);

INVx8_ASAP7_75t_L g2839 ( 
.A(n_2348),
.Y(n_2839)
);

NAND2x1p5_ASAP7_75t_L g2840 ( 
.A(n_2451),
.B(n_478),
.Y(n_2840)
);

HB1xp67_ASAP7_75t_L g2841 ( 
.A(n_2132),
.Y(n_2841)
);

INVx3_ASAP7_75t_L g2842 ( 
.A(n_2348),
.Y(n_2842)
);

BUFx3_ASAP7_75t_L g2843 ( 
.A(n_2348),
.Y(n_2843)
);

NOR2xp33_ASAP7_75t_L g2844 ( 
.A(n_2325),
.B(n_478),
.Y(n_2844)
);

OAI21x1_ASAP7_75t_SL g2845 ( 
.A1(n_2377),
.A2(n_2301),
.B(n_2497),
.Y(n_2845)
);

AO21x2_ASAP7_75t_L g2846 ( 
.A1(n_2411),
.A2(n_479),
.B(n_481),
.Y(n_2846)
);

AO21x2_ASAP7_75t_L g2847 ( 
.A1(n_2366),
.A2(n_481),
.B(n_482),
.Y(n_2847)
);

BUFx2_ASAP7_75t_L g2848 ( 
.A(n_2282),
.Y(n_2848)
);

AOI22x1_ASAP7_75t_L g2849 ( 
.A1(n_2452),
.A2(n_484),
.B1(n_482),
.B2(n_483),
.Y(n_2849)
);

OAI21xp5_ASAP7_75t_L g2850 ( 
.A1(n_2394),
.A2(n_484),
.B(n_485),
.Y(n_2850)
);

INVx2_ASAP7_75t_L g2851 ( 
.A(n_2242),
.Y(n_2851)
);

AOI21xp5_ASAP7_75t_L g2852 ( 
.A1(n_2155),
.A2(n_486),
.B(n_487),
.Y(n_2852)
);

INVx8_ASAP7_75t_L g2853 ( 
.A(n_2265),
.Y(n_2853)
);

BUFx3_ASAP7_75t_L g2854 ( 
.A(n_2206),
.Y(n_2854)
);

NAND2x1p5_ASAP7_75t_L g2855 ( 
.A(n_2451),
.B(n_487),
.Y(n_2855)
);

BUFx2_ASAP7_75t_L g2856 ( 
.A(n_2478),
.Y(n_2856)
);

INVx1_ASAP7_75t_L g2857 ( 
.A(n_2140),
.Y(n_2857)
);

INVx2_ASAP7_75t_L g2858 ( 
.A(n_2243),
.Y(n_2858)
);

NOR2xp33_ASAP7_75t_L g2859 ( 
.A(n_2153),
.B(n_488),
.Y(n_2859)
);

BUFx2_ASAP7_75t_R g2860 ( 
.A(n_2386),
.Y(n_2860)
);

NAND2xp5_ASAP7_75t_L g2861 ( 
.A(n_2280),
.B(n_2287),
.Y(n_2861)
);

BUFx6f_ASAP7_75t_L g2862 ( 
.A(n_2455),
.Y(n_2862)
);

AO21x2_ASAP7_75t_L g2863 ( 
.A1(n_2485),
.A2(n_489),
.B(n_490),
.Y(n_2863)
);

INVx3_ASAP7_75t_L g2864 ( 
.A(n_2455),
.Y(n_2864)
);

INVx3_ASAP7_75t_L g2865 ( 
.A(n_2488),
.Y(n_2865)
);

INVx8_ASAP7_75t_L g2866 ( 
.A(n_2185),
.Y(n_2866)
);

INVx1_ASAP7_75t_SL g2867 ( 
.A(n_2203),
.Y(n_2867)
);

INVx2_ASAP7_75t_L g2868 ( 
.A(n_2302),
.Y(n_2868)
);

AO21x2_ASAP7_75t_L g2869 ( 
.A1(n_2499),
.A2(n_491),
.B(n_492),
.Y(n_2869)
);

BUFx3_ASAP7_75t_L g2870 ( 
.A(n_2498),
.Y(n_2870)
);

INVx1_ASAP7_75t_L g2871 ( 
.A(n_2154),
.Y(n_2871)
);

OAI21xp5_ASAP7_75t_L g2872 ( 
.A1(n_2394),
.A2(n_491),
.B(n_492),
.Y(n_2872)
);

AO21x2_ASAP7_75t_L g2873 ( 
.A1(n_2500),
.A2(n_493),
.B(n_494),
.Y(n_2873)
);

CKINVDCx5p33_ASAP7_75t_R g2874 ( 
.A(n_2300),
.Y(n_2874)
);

BUFx3_ASAP7_75t_L g2875 ( 
.A(n_2350),
.Y(n_2875)
);

CKINVDCx20_ASAP7_75t_R g2876 ( 
.A(n_2345),
.Y(n_2876)
);

CKINVDCx16_ASAP7_75t_R g2877 ( 
.A(n_2354),
.Y(n_2877)
);

CKINVDCx14_ASAP7_75t_R g2878 ( 
.A(n_2530),
.Y(n_2878)
);

BUFx12f_ASAP7_75t_L g2879 ( 
.A(n_2274),
.Y(n_2879)
);

BUFx5_ASAP7_75t_L g2880 ( 
.A(n_2364),
.Y(n_2880)
);

AOI22xp33_ASAP7_75t_L g2881 ( 
.A1(n_2562),
.A2(n_496),
.B1(n_493),
.B2(n_495),
.Y(n_2881)
);

HB1xp67_ASAP7_75t_L g2882 ( 
.A(n_2174),
.Y(n_2882)
);

INVx1_ASAP7_75t_L g2883 ( 
.A(n_2190),
.Y(n_2883)
);

INVx2_ASAP7_75t_L g2884 ( 
.A(n_2307),
.Y(n_2884)
);

OAI21x1_ASAP7_75t_SL g2885 ( 
.A1(n_2377),
.A2(n_497),
.B(n_499),
.Y(n_2885)
);

NAND2x1p5_ASAP7_75t_L g2886 ( 
.A(n_2533),
.B(n_499),
.Y(n_2886)
);

INVx1_ASAP7_75t_L g2887 ( 
.A(n_2376),
.Y(n_2887)
);

INVx1_ASAP7_75t_L g2888 ( 
.A(n_2497),
.Y(n_2888)
);

INVx1_ASAP7_75t_L g2889 ( 
.A(n_2558),
.Y(n_2889)
);

OA21x2_ASAP7_75t_L g2890 ( 
.A1(n_2360),
.A2(n_500),
.B(n_501),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2311),
.B(n_501),
.Y(n_2891)
);

INVx1_ASAP7_75t_L g2892 ( 
.A(n_2558),
.Y(n_2892)
);

INVx2_ASAP7_75t_L g2893 ( 
.A(n_2318),
.Y(n_2893)
);

NOR2xp33_ASAP7_75t_L g2894 ( 
.A(n_2097),
.B(n_502),
.Y(n_2894)
);

NOR2xp33_ASAP7_75t_L g2895 ( 
.A(n_2115),
.B(n_2133),
.Y(n_2895)
);

INVx8_ASAP7_75t_L g2896 ( 
.A(n_2116),
.Y(n_2896)
);

BUFx3_ASAP7_75t_L g2897 ( 
.A(n_2306),
.Y(n_2897)
);

AND2x4_ASAP7_75t_L g2898 ( 
.A(n_2101),
.B(n_503),
.Y(n_2898)
);

BUFx3_ASAP7_75t_L g2899 ( 
.A(n_2383),
.Y(n_2899)
);

BUFx12f_ASAP7_75t_L g2900 ( 
.A(n_2163),
.Y(n_2900)
);

BUFx3_ASAP7_75t_L g2901 ( 
.A(n_2116),
.Y(n_2901)
);

INVxp67_ASAP7_75t_SL g2902 ( 
.A(n_2553),
.Y(n_2902)
);

AO21x2_ASAP7_75t_L g2903 ( 
.A1(n_2259),
.A2(n_505),
.B(n_506),
.Y(n_2903)
);

AOI22x1_ASAP7_75t_L g2904 ( 
.A1(n_2258),
.A2(n_508),
.B1(n_506),
.B2(n_507),
.Y(n_2904)
);

NAND2x1p5_ASAP7_75t_L g2905 ( 
.A(n_2553),
.B(n_507),
.Y(n_2905)
);

INVx8_ASAP7_75t_L g2906 ( 
.A(n_2553),
.Y(n_2906)
);

AOI22x1_ASAP7_75t_L g2907 ( 
.A1(n_2266),
.A2(n_513),
.B1(n_509),
.B2(n_511),
.Y(n_2907)
);

BUFx6f_ASAP7_75t_L g2908 ( 
.A(n_2338),
.Y(n_2908)
);

AOI22x1_ASAP7_75t_L g2909 ( 
.A1(n_2273),
.A2(n_514),
.B1(n_509),
.B2(n_513),
.Y(n_2909)
);

INVx2_ASAP7_75t_SL g2910 ( 
.A(n_2314),
.Y(n_2910)
);

BUFx3_ASAP7_75t_L g2911 ( 
.A(n_2094),
.Y(n_2911)
);

CKINVDCx12_ASAP7_75t_R g2912 ( 
.A(n_2170),
.Y(n_2912)
);

INVx1_ASAP7_75t_L g2913 ( 
.A(n_2168),
.Y(n_2913)
);

BUFx6f_ASAP7_75t_L g2914 ( 
.A(n_2094),
.Y(n_2914)
);

INVx1_ASAP7_75t_L g2915 ( 
.A(n_2176),
.Y(n_2915)
);

BUFx2_ASAP7_75t_L g2916 ( 
.A(n_2336),
.Y(n_2916)
);

INVx1_ASAP7_75t_L g2917 ( 
.A(n_2248),
.Y(n_2917)
);

NAND2x1p5_ASAP7_75t_L g2918 ( 
.A(n_2127),
.B(n_518),
.Y(n_2918)
);

BUFx2_ASAP7_75t_L g2919 ( 
.A(n_2167),
.Y(n_2919)
);

INVx1_ASAP7_75t_L g2920 ( 
.A(n_2195),
.Y(n_2920)
);

INVx8_ASAP7_75t_L g2921 ( 
.A(n_2100),
.Y(n_2921)
);

AO21x2_ASAP7_75t_L g2922 ( 
.A1(n_2263),
.A2(n_519),
.B(n_520),
.Y(n_2922)
);

AO21x2_ASAP7_75t_L g2923 ( 
.A1(n_2264),
.A2(n_519),
.B(n_520),
.Y(n_2923)
);

AO21x2_ASAP7_75t_L g2924 ( 
.A1(n_2271),
.A2(n_521),
.B(n_522),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2137),
.B(n_521),
.Y(n_2925)
);

BUFx2_ASAP7_75t_R g2926 ( 
.A(n_2180),
.Y(n_2926)
);

INVx2_ASAP7_75t_L g2927 ( 
.A(n_2527),
.Y(n_2927)
);

OAI22xp33_ASAP7_75t_L g2928 ( 
.A1(n_2301),
.A2(n_528),
.B1(n_524),
.B2(n_526),
.Y(n_2928)
);

AO21x2_ASAP7_75t_L g2929 ( 
.A1(n_2413),
.A2(n_529),
.B(n_530),
.Y(n_2929)
);

INVx1_ASAP7_75t_L g2930 ( 
.A(n_2197),
.Y(n_2930)
);

CKINVDCx20_ASAP7_75t_R g2931 ( 
.A(n_2109),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2527),
.Y(n_2932)
);

INVx1_ASAP7_75t_L g2933 ( 
.A(n_2527),
.Y(n_2933)
);

NAND3xp33_ASAP7_75t_L g2934 ( 
.A(n_2279),
.B(n_529),
.C(n_531),
.Y(n_2934)
);

INVx2_ASAP7_75t_SL g2935 ( 
.A(n_2341),
.Y(n_2935)
);

NAND2x1p5_ASAP7_75t_L g2936 ( 
.A(n_2550),
.B(n_532),
.Y(n_2936)
);

AOI21x1_ASAP7_75t_L g2937 ( 
.A1(n_2380),
.A2(n_533),
.B(n_534),
.Y(n_2937)
);

NAND2xp5_ASAP7_75t_L g2938 ( 
.A(n_2103),
.B(n_533),
.Y(n_2938)
);

NAND2x1_ASAP7_75t_L g2939 ( 
.A(n_2232),
.B(n_535),
.Y(n_2939)
);

INVx1_ASAP7_75t_L g2940 ( 
.A(n_2294),
.Y(n_2940)
);

INVx1_ASAP7_75t_L g2941 ( 
.A(n_2332),
.Y(n_2941)
);

BUFx6f_ASAP7_75t_SL g2942 ( 
.A(n_2100),
.Y(n_2942)
);

INVx4_ASAP7_75t_L g2943 ( 
.A(n_2256),
.Y(n_2943)
);

BUFx6f_ASAP7_75t_L g2944 ( 
.A(n_2361),
.Y(n_2944)
);

OA21x2_ASAP7_75t_L g2945 ( 
.A1(n_2444),
.A2(n_537),
.B(n_538),
.Y(n_2945)
);

NAND2xp5_ASAP7_75t_L g2946 ( 
.A(n_2114),
.B(n_2123),
.Y(n_2946)
);

OA21x2_ASAP7_75t_L g2947 ( 
.A1(n_2491),
.A2(n_537),
.B(n_538),
.Y(n_2947)
);

INVx6_ASAP7_75t_L g2948 ( 
.A(n_2249),
.Y(n_2948)
);

BUFx2_ASAP7_75t_L g2949 ( 
.A(n_2375),
.Y(n_2949)
);

BUFx6f_ASAP7_75t_L g2950 ( 
.A(n_2368),
.Y(n_2950)
);

CKINVDCx8_ASAP7_75t_R g2951 ( 
.A(n_2340),
.Y(n_2951)
);

AO21x2_ASAP7_75t_L g2952 ( 
.A1(n_2561),
.A2(n_539),
.B(n_540),
.Y(n_2952)
);

HB1xp67_ASAP7_75t_L g2953 ( 
.A(n_2182),
.Y(n_2953)
);

INVx6_ASAP7_75t_L g2954 ( 
.A(n_2257),
.Y(n_2954)
);

AND2x4_ASAP7_75t_L g2955 ( 
.A(n_2281),
.B(n_541),
.Y(n_2955)
);

OR2x6_ASAP7_75t_L g2956 ( 
.A(n_2193),
.B(n_542),
.Y(n_2956)
);

INVx3_ASAP7_75t_L g2957 ( 
.A(n_2250),
.Y(n_2957)
);

OAI21x1_ASAP7_75t_L g2958 ( 
.A1(n_2432),
.A2(n_543),
.B(n_544),
.Y(n_2958)
);

CKINVDCx14_ASAP7_75t_R g2959 ( 
.A(n_2298),
.Y(n_2959)
);

INVx6_ASAP7_75t_L g2960 ( 
.A(n_2113),
.Y(n_2960)
);

INVx5_ASAP7_75t_L g2961 ( 
.A(n_2192),
.Y(n_2961)
);

INVx2_ASAP7_75t_L g2962 ( 
.A(n_2537),
.Y(n_2962)
);

INVx1_ASAP7_75t_SL g2963 ( 
.A(n_2214),
.Y(n_2963)
);

INVx1_ASAP7_75t_L g2964 ( 
.A(n_2305),
.Y(n_2964)
);

OR2x2_ASAP7_75t_L g2965 ( 
.A(n_2148),
.B(n_2093),
.Y(n_2965)
);

OAI21x1_ASAP7_75t_L g2966 ( 
.A1(n_2528),
.A2(n_543),
.B(n_545),
.Y(n_2966)
);

INVx2_ASAP7_75t_L g2967 ( 
.A(n_2537),
.Y(n_2967)
);

INVx4_ASAP7_75t_L g2968 ( 
.A(n_2396),
.Y(n_2968)
);

INVx3_ASAP7_75t_L g2969 ( 
.A(n_2253),
.Y(n_2969)
);

INVx2_ASAP7_75t_L g2970 ( 
.A(n_2135),
.Y(n_2970)
);

BUFx6f_ASAP7_75t_L g2971 ( 
.A(n_2254),
.Y(n_2971)
);

NAND2xp5_ASAP7_75t_L g2972 ( 
.A(n_2178),
.B(n_548),
.Y(n_2972)
);

AOI22x1_ASAP7_75t_L g2973 ( 
.A1(n_2269),
.A2(n_550),
.B1(n_548),
.B2(n_549),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2393),
.Y(n_2974)
);

NOR2xp67_ASAP7_75t_L g2975 ( 
.A(n_2129),
.B(n_553),
.Y(n_2975)
);

AND2x2_ASAP7_75t_L g2976 ( 
.A(n_2090),
.B(n_554),
.Y(n_2976)
);

INVx3_ASAP7_75t_L g2977 ( 
.A(n_2255),
.Y(n_2977)
);

INVx1_ASAP7_75t_L g2978 ( 
.A(n_2412),
.Y(n_2978)
);

BUFx6f_ASAP7_75t_L g2979 ( 
.A(n_2319),
.Y(n_2979)
);

BUFx12f_ASAP7_75t_L g2980 ( 
.A(n_2422),
.Y(n_2980)
);

CKINVDCx5p33_ASAP7_75t_R g2981 ( 
.A(n_2578),
.Y(n_2981)
);

INVx4_ASAP7_75t_L g2982 ( 
.A(n_2591),
.Y(n_2982)
);

OAI22xp33_ASAP7_75t_L g2983 ( 
.A1(n_2740),
.A2(n_2286),
.B1(n_2283),
.B2(n_2387),
.Y(n_2983)
);

INVx6_ASAP7_75t_L g2984 ( 
.A(n_2591),
.Y(n_2984)
);

INVx2_ASAP7_75t_L g2985 ( 
.A(n_2584),
.Y(n_2985)
);

HB1xp67_ASAP7_75t_L g2986 ( 
.A(n_2757),
.Y(n_2986)
);

INVx2_ASAP7_75t_L g2987 ( 
.A(n_2586),
.Y(n_2987)
);

INVx1_ASAP7_75t_L g2988 ( 
.A(n_2621),
.Y(n_2988)
);

INVx3_ASAP7_75t_SL g2989 ( 
.A(n_2591),
.Y(n_2989)
);

INVx1_ASAP7_75t_L g2990 ( 
.A(n_2627),
.Y(n_2990)
);

INVx2_ASAP7_75t_L g2991 ( 
.A(n_2593),
.Y(n_2991)
);

OAI22xp5_ASAP7_75t_L g2992 ( 
.A1(n_2740),
.A2(n_2450),
.B1(n_2507),
.B2(n_2504),
.Y(n_2992)
);

INVx6_ASAP7_75t_L g2993 ( 
.A(n_2592),
.Y(n_2993)
);

NAND2x1p5_ASAP7_75t_L g2994 ( 
.A(n_2567),
.B(n_2392),
.Y(n_2994)
);

INVx2_ASAP7_75t_L g2995 ( 
.A(n_2594),
.Y(n_2995)
);

AND2x2_ASAP7_75t_L g2996 ( 
.A(n_2960),
.B(n_2506),
.Y(n_2996)
);

NAND2x1p5_ASAP7_75t_L g2997 ( 
.A(n_2567),
.B(n_2406),
.Y(n_2997)
);

OAI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_2740),
.A2(n_2532),
.B1(n_2546),
.B2(n_2479),
.Y(n_2998)
);

INVx2_ASAP7_75t_L g2999 ( 
.A(n_2624),
.Y(n_2999)
);

BUFx2_ASAP7_75t_L g3000 ( 
.A(n_2759),
.Y(n_3000)
);

INVx1_ASAP7_75t_L g3001 ( 
.A(n_2631),
.Y(n_3001)
);

AOI22xp33_ASAP7_75t_L g3002 ( 
.A1(n_2895),
.A2(n_2400),
.B1(n_2431),
.B2(n_2408),
.Y(n_3002)
);

INVx2_ASAP7_75t_L g3003 ( 
.A(n_2629),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2637),
.Y(n_3004)
);

AOI22xp33_ASAP7_75t_L g3005 ( 
.A1(n_2895),
.A2(n_2845),
.B1(n_2960),
.B2(n_2721),
.Y(n_3005)
);

INVx1_ASAP7_75t_L g3006 ( 
.A(n_2641),
.Y(n_3006)
);

AND2x4_ASAP7_75t_L g3007 ( 
.A(n_2567),
.B(n_2370),
.Y(n_3007)
);

INVx2_ASAP7_75t_L g3008 ( 
.A(n_2634),
.Y(n_3008)
);

BUFx6f_ASAP7_75t_SL g3009 ( 
.A(n_2653),
.Y(n_3009)
);

INVx1_ASAP7_75t_L g3010 ( 
.A(n_2642),
.Y(n_3010)
);

INVx1_ASAP7_75t_L g3011 ( 
.A(n_2655),
.Y(n_3011)
);

INVx2_ASAP7_75t_L g3012 ( 
.A(n_2651),
.Y(n_3012)
);

OAI21xp5_ASAP7_75t_L g3013 ( 
.A1(n_2852),
.A2(n_2832),
.B(n_2619),
.Y(n_3013)
);

AOI22xp33_ASAP7_75t_L g3014 ( 
.A1(n_2960),
.A2(n_2721),
.B1(n_2750),
.B2(n_2619),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2592),
.Y(n_3015)
);

OAI21x1_ASAP7_75t_SL g3016 ( 
.A1(n_2850),
.A2(n_2872),
.B(n_2608),
.Y(n_3016)
);

INVx1_ASAP7_75t_L g3017 ( 
.A(n_2659),
.Y(n_3017)
);

CKINVDCx5p33_ASAP7_75t_R g3018 ( 
.A(n_2673),
.Y(n_3018)
);

OAI21xp5_ASAP7_75t_SL g3019 ( 
.A1(n_2881),
.A2(n_2272),
.B(n_2216),
.Y(n_3019)
);

INVx2_ASAP7_75t_L g3020 ( 
.A(n_2679),
.Y(n_3020)
);

INVx1_ASAP7_75t_L g3021 ( 
.A(n_2671),
.Y(n_3021)
);

BUFx3_ASAP7_75t_L g3022 ( 
.A(n_2592),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2888),
.B(n_2156),
.Y(n_3023)
);

INVx2_ASAP7_75t_L g3024 ( 
.A(n_2681),
.Y(n_3024)
);

INVx6_ASAP7_75t_L g3025 ( 
.A(n_2645),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2677),
.Y(n_3026)
);

OAI22xp5_ASAP7_75t_L g3027 ( 
.A1(n_2732),
.A2(n_2241),
.B1(n_2371),
.B2(n_2260),
.Y(n_3027)
);

NAND2x1p5_ASAP7_75t_L g3028 ( 
.A(n_2567),
.B(n_2426),
.Y(n_3028)
);

INVx4_ASAP7_75t_L g3029 ( 
.A(n_2572),
.Y(n_3029)
);

INVx2_ASAP7_75t_L g3030 ( 
.A(n_2691),
.Y(n_3030)
);

INVx2_ASAP7_75t_L g3031 ( 
.A(n_2698),
.Y(n_3031)
);

INVx2_ASAP7_75t_L g3032 ( 
.A(n_2818),
.Y(n_3032)
);

CKINVDCx11_ASAP7_75t_R g3033 ( 
.A(n_2618),
.Y(n_3033)
);

BUFx3_ASAP7_75t_L g3034 ( 
.A(n_2686),
.Y(n_3034)
);

INVx1_ASAP7_75t_L g3035 ( 
.A(n_2688),
.Y(n_3035)
);

INVx2_ASAP7_75t_L g3036 ( 
.A(n_2568),
.Y(n_3036)
);

BUFx3_ASAP7_75t_L g3037 ( 
.A(n_2686),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2694),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2700),
.Y(n_3039)
);

AOI22xp33_ASAP7_75t_L g3040 ( 
.A1(n_2750),
.A2(n_2436),
.B1(n_2461),
.B2(n_2435),
.Y(n_3040)
);

AND2x4_ASAP7_75t_L g3041 ( 
.A(n_2649),
.B(n_2240),
.Y(n_3041)
);

INVx1_ASAP7_75t_SL g3042 ( 
.A(n_2589),
.Y(n_3042)
);

OAI21x1_ASAP7_75t_L g3043 ( 
.A1(n_2751),
.A2(n_2199),
.B(n_2252),
.Y(n_3043)
);

INVxp33_ASAP7_75t_L g3044 ( 
.A(n_2757),
.Y(n_3044)
);

INVx2_ASAP7_75t_L g3045 ( 
.A(n_2573),
.Y(n_3045)
);

AOI22xp33_ASAP7_75t_L g3046 ( 
.A1(n_2935),
.A2(n_2496),
.B1(n_2517),
.B2(n_2470),
.Y(n_3046)
);

INVx4_ASAP7_75t_L g3047 ( 
.A(n_2572),
.Y(n_3047)
);

HB1xp67_ASAP7_75t_SL g3048 ( 
.A(n_2602),
.Y(n_3048)
);

AOI22xp33_ASAP7_75t_L g3049 ( 
.A1(n_2889),
.A2(n_2559),
.B1(n_2551),
.B2(n_2324),
.Y(n_3049)
);

INVx6_ASAP7_75t_L g3050 ( 
.A(n_2645),
.Y(n_3050)
);

INVx2_ASAP7_75t_L g3051 ( 
.A(n_2581),
.Y(n_3051)
);

INVx8_ASAP7_75t_L g3052 ( 
.A(n_2572),
.Y(n_3052)
);

CKINVDCx5p33_ASAP7_75t_R g3053 ( 
.A(n_2673),
.Y(n_3053)
);

INVx2_ASAP7_75t_L g3054 ( 
.A(n_2583),
.Y(n_3054)
);

INVx2_ASAP7_75t_L g3055 ( 
.A(n_2595),
.Y(n_3055)
);

AO21x1_ASAP7_75t_L g3056 ( 
.A1(n_2850),
.A2(n_2200),
.B(n_2347),
.Y(n_3056)
);

OA21x2_ASAP7_75t_L g3057 ( 
.A1(n_2932),
.A2(n_2933),
.B(n_2927),
.Y(n_3057)
);

AOI22xp5_ASAP7_75t_L g3058 ( 
.A1(n_2892),
.A2(n_2262),
.B1(n_2365),
.B2(n_2117),
.Y(n_3058)
);

INVx2_ASAP7_75t_L g3059 ( 
.A(n_2600),
.Y(n_3059)
);

INVx2_ASAP7_75t_L g3060 ( 
.A(n_2601),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2707),
.Y(n_3061)
);

INVx2_ASAP7_75t_L g3062 ( 
.A(n_2603),
.Y(n_3062)
);

OAI22xp5_ASAP7_75t_L g3063 ( 
.A1(n_2575),
.A2(n_2211),
.B1(n_2208),
.B2(n_2355),
.Y(n_3063)
);

INVx3_ASAP7_75t_L g3064 ( 
.A(n_2605),
.Y(n_3064)
);

HB1xp67_ASAP7_75t_L g3065 ( 
.A(n_2761),
.Y(n_3065)
);

INVx4_ASAP7_75t_L g3066 ( 
.A(n_2639),
.Y(n_3066)
);

BUFx3_ASAP7_75t_L g3067 ( 
.A(n_2617),
.Y(n_3067)
);

INVx4_ASAP7_75t_L g3068 ( 
.A(n_2649),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2710),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2713),
.Y(n_3070)
);

INVx1_ASAP7_75t_SL g3071 ( 
.A(n_2589),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2725),
.Y(n_3072)
);

BUFx2_ASAP7_75t_L g3073 ( 
.A(n_2759),
.Y(n_3073)
);

AND2x2_ASAP7_75t_L g3074 ( 
.A(n_2835),
.B(n_2369),
.Y(n_3074)
);

INVx4_ASAP7_75t_L g3075 ( 
.A(n_2649),
.Y(n_3075)
);

AND2x2_ASAP7_75t_L g3076 ( 
.A(n_2835),
.B(n_2720),
.Y(n_3076)
);

INVx2_ASAP7_75t_L g3077 ( 
.A(n_2613),
.Y(n_3077)
);

OAI21xp5_ASAP7_75t_L g3078 ( 
.A1(n_2852),
.A2(n_2189),
.B(n_2108),
.Y(n_3078)
);

INVx2_ASAP7_75t_L g3079 ( 
.A(n_2745),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2917),
.B(n_2378),
.Y(n_3080)
);

INVx1_ASAP7_75t_L g3081 ( 
.A(n_2731),
.Y(n_3081)
);

AOI22xp33_ASAP7_75t_L g3082 ( 
.A1(n_2728),
.A2(n_2237),
.B1(n_2457),
.B2(n_2456),
.Y(n_3082)
);

AOI22xp33_ASAP7_75t_SL g3083 ( 
.A1(n_2728),
.A2(n_2352),
.B1(n_2462),
.B2(n_2446),
.Y(n_3083)
);

CKINVDCx5p33_ASAP7_75t_R g3084 ( 
.A(n_2612),
.Y(n_3084)
);

INVx1_ASAP7_75t_SL g3085 ( 
.A(n_2784),
.Y(n_3085)
);

BUFx2_ASAP7_75t_L g3086 ( 
.A(n_2577),
.Y(n_3086)
);

BUFx2_ASAP7_75t_L g3087 ( 
.A(n_2577),
.Y(n_3087)
);

OAI22xp5_ASAP7_75t_L g3088 ( 
.A1(n_2575),
.A2(n_2493),
.B1(n_2518),
.B2(n_2472),
.Y(n_3088)
);

NAND2x1p5_ASAP7_75t_L g3089 ( 
.A(n_2649),
.B(n_2529),
.Y(n_3089)
);

AOI22xp33_ASAP7_75t_SL g3090 ( 
.A1(n_2728),
.A2(n_2468),
.B1(n_2495),
.B2(n_2484),
.Y(n_3090)
);

INVx2_ASAP7_75t_SL g3091 ( 
.A(n_2658),
.Y(n_3091)
);

INVx6_ASAP7_75t_L g3092 ( 
.A(n_2587),
.Y(n_3092)
);

INVx5_ASAP7_75t_L g3093 ( 
.A(n_2674),
.Y(n_3093)
);

AOI22xp33_ASAP7_75t_L g3094 ( 
.A1(n_2876),
.A2(n_2531),
.B1(n_2566),
.B2(n_2534),
.Y(n_3094)
);

INVx2_ASAP7_75t_L g3095 ( 
.A(n_2753),
.Y(n_3095)
);

INVx4_ASAP7_75t_L g3096 ( 
.A(n_2674),
.Y(n_3096)
);

BUFx2_ASAP7_75t_R g3097 ( 
.A(n_2667),
.Y(n_3097)
);

INVx3_ASAP7_75t_L g3098 ( 
.A(n_2605),
.Y(n_3098)
);

BUFx8_ASAP7_75t_L g3099 ( 
.A(n_2670),
.Y(n_3099)
);

BUFx2_ASAP7_75t_R g3100 ( 
.A(n_2874),
.Y(n_3100)
);

INVx3_ASAP7_75t_L g3101 ( 
.A(n_2821),
.Y(n_3101)
);

INVx1_ASAP7_75t_L g3102 ( 
.A(n_2738),
.Y(n_3102)
);

INVx1_ASAP7_75t_L g3103 ( 
.A(n_2800),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2748),
.Y(n_3104)
);

INVx2_ASAP7_75t_L g3105 ( 
.A(n_2756),
.Y(n_3105)
);

INVx1_ASAP7_75t_L g3106 ( 
.A(n_2754),
.Y(n_3106)
);

INVx1_ASAP7_75t_SL g3107 ( 
.A(n_2784),
.Y(n_3107)
);

AOI22xp33_ASAP7_75t_L g3108 ( 
.A1(n_2876),
.A2(n_2267),
.B1(n_2367),
.B2(n_2342),
.Y(n_3108)
);

INVx2_ASAP7_75t_SL g3109 ( 
.A(n_2726),
.Y(n_3109)
);

AOI22xp33_ASAP7_75t_L g3110 ( 
.A1(n_2799),
.A2(n_2296),
.B1(n_2158),
.B2(n_2160),
.Y(n_3110)
);

NAND2xp5_ASAP7_75t_L g3111 ( 
.A(n_2822),
.B(n_2389),
.Y(n_3111)
);

INVx1_ASAP7_75t_L g3112 ( 
.A(n_2768),
.Y(n_3112)
);

INVx2_ASAP7_75t_L g3113 ( 
.A(n_2774),
.Y(n_3113)
);

INVx2_ASAP7_75t_L g3114 ( 
.A(n_2806),
.Y(n_3114)
);

INVxp67_ASAP7_75t_SL g3115 ( 
.A(n_2841),
.Y(n_3115)
);

INVx2_ASAP7_75t_L g3116 ( 
.A(n_2736),
.Y(n_3116)
);

INVx2_ASAP7_75t_L g3117 ( 
.A(n_2823),
.Y(n_3117)
);

AOI22xp33_ASAP7_75t_L g3118 ( 
.A1(n_2799),
.A2(n_2357),
.B1(n_2337),
.B2(n_2297),
.Y(n_3118)
);

AO21x2_ASAP7_75t_L g3119 ( 
.A1(n_2675),
.A2(n_2179),
.B(n_2212),
.Y(n_3119)
);

BUFx12f_ASAP7_75t_L g3120 ( 
.A(n_2615),
.Y(n_3120)
);

BUFx12f_ASAP7_75t_SL g3121 ( 
.A(n_2669),
.Y(n_3121)
);

INVx3_ASAP7_75t_L g3122 ( 
.A(n_2821),
.Y(n_3122)
);

BUFx3_ASAP7_75t_L g3123 ( 
.A(n_2729),
.Y(n_3123)
);

AOI22xp33_ASAP7_75t_L g3124 ( 
.A1(n_2894),
.A2(n_2270),
.B1(n_2226),
.B2(n_2239),
.Y(n_3124)
);

AOI22xp33_ASAP7_75t_L g3125 ( 
.A1(n_2894),
.A2(n_2535),
.B1(n_2525),
.B2(n_2315),
.Y(n_3125)
);

OAI22xp5_ASAP7_75t_L g3126 ( 
.A1(n_2674),
.A2(n_2961),
.B1(n_2705),
.B2(n_2702),
.Y(n_3126)
);

INVx1_ASAP7_75t_L g3127 ( 
.A(n_2787),
.Y(n_3127)
);

CKINVDCx6p67_ASAP7_75t_R g3128 ( 
.A(n_2803),
.Y(n_3128)
);

NOR2xp33_ASAP7_75t_L g3129 ( 
.A(n_2931),
.B(n_2150),
.Y(n_3129)
);

BUFx3_ASAP7_75t_L g3130 ( 
.A(n_2730),
.Y(n_3130)
);

OR2x6_ASAP7_75t_L g3131 ( 
.A(n_2726),
.B(n_2175),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2793),
.Y(n_3132)
);

NAND2x1p5_ASAP7_75t_L g3133 ( 
.A(n_2821),
.B(n_2563),
.Y(n_3133)
);

BUFx6f_ASAP7_75t_L g3134 ( 
.A(n_2906),
.Y(n_3134)
);

AOI22xp33_ASAP7_75t_SL g3135 ( 
.A1(n_2726),
.A2(n_2358),
.B1(n_2403),
.B2(n_2397),
.Y(n_3135)
);

INVx2_ASAP7_75t_L g3136 ( 
.A(n_2851),
.Y(n_3136)
);

HB1xp67_ASAP7_75t_L g3137 ( 
.A(n_2771),
.Y(n_3137)
);

OAI21x1_ASAP7_75t_L g3138 ( 
.A1(n_2680),
.A2(n_2409),
.B(n_2407),
.Y(n_3138)
);

HB1xp67_ASAP7_75t_L g3139 ( 
.A(n_2776),
.Y(n_3139)
);

INVx1_ASAP7_75t_L g3140 ( 
.A(n_2622),
.Y(n_3140)
);

INVx2_ASAP7_75t_L g3141 ( 
.A(n_2858),
.Y(n_3141)
);

INVx1_ASAP7_75t_L g3142 ( 
.A(n_2622),
.Y(n_3142)
);

INVx2_ASAP7_75t_L g3143 ( 
.A(n_2868),
.Y(n_3143)
);

INVx2_ASAP7_75t_L g3144 ( 
.A(n_2884),
.Y(n_3144)
);

NAND2xp5_ASAP7_75t_L g3145 ( 
.A(n_2964),
.B(n_2438),
.Y(n_3145)
);

HB1xp67_ASAP7_75t_L g3146 ( 
.A(n_2749),
.Y(n_3146)
);

INVx5_ASAP7_75t_L g3147 ( 
.A(n_2692),
.Y(n_3147)
);

INVx1_ASAP7_75t_SL g3148 ( 
.A(n_2741),
.Y(n_3148)
);

INVx2_ASAP7_75t_SL g3149 ( 
.A(n_2742),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2625),
.Y(n_3150)
);

INVx2_ASAP7_75t_L g3151 ( 
.A(n_2893),
.Y(n_3151)
);

NOR2x1_ASAP7_75t_R g3152 ( 
.A(n_2737),
.B(n_2439),
.Y(n_3152)
);

INVx1_ASAP7_75t_L g3153 ( 
.A(n_2625),
.Y(n_3153)
);

INVx2_ASAP7_75t_L g3154 ( 
.A(n_2861),
.Y(n_3154)
);

NAND2xp5_ASAP7_75t_L g3155 ( 
.A(n_2974),
.B(n_2445),
.Y(n_3155)
);

AOI22xp33_ASAP7_75t_L g3156 ( 
.A1(n_2980),
.A2(n_2778),
.B1(n_2878),
.B2(n_2900),
.Y(n_3156)
);

BUFx3_ASAP7_75t_L g3157 ( 
.A(n_2772),
.Y(n_3157)
);

INVx2_ASAP7_75t_SL g3158 ( 
.A(n_2742),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_2861),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2638),
.Y(n_3160)
);

HB1xp67_ASAP7_75t_L g3161 ( 
.A(n_2758),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_2638),
.Y(n_3162)
);

OAI22xp5_ASAP7_75t_L g3163 ( 
.A1(n_2961),
.A2(n_2705),
.B1(n_2702),
.B2(n_2723),
.Y(n_3163)
);

BUFx3_ASAP7_75t_L g3164 ( 
.A(n_2689),
.Y(n_3164)
);

INVx1_ASAP7_75t_L g3165 ( 
.A(n_2685),
.Y(n_3165)
);

AOI22xp33_ASAP7_75t_L g3166 ( 
.A1(n_2878),
.A2(n_2447),
.B1(n_2459),
.B2(n_2458),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2685),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2786),
.Y(n_3168)
);

AOI22xp33_ASAP7_75t_L g3169 ( 
.A1(n_2978),
.A2(n_2467),
.B1(n_2486),
.B2(n_2480),
.Y(n_3169)
);

INVx1_ASAP7_75t_SL g3170 ( 
.A(n_2741),
.Y(n_3170)
);

INVx2_ASAP7_75t_L g3171 ( 
.A(n_2795),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_2739),
.B(n_2151),
.Y(n_3172)
);

NAND2x1p5_ASAP7_75t_L g3173 ( 
.A(n_2821),
.B(n_2554),
.Y(n_3173)
);

NAND2xp5_ASAP7_75t_L g3174 ( 
.A(n_2970),
.B(n_2522),
.Y(n_3174)
);

CKINVDCx11_ASAP7_75t_R g3175 ( 
.A(n_2780),
.Y(n_3175)
);

INVxp67_ASAP7_75t_L g3176 ( 
.A(n_2723),
.Y(n_3176)
);

HB1xp67_ASAP7_75t_SL g3177 ( 
.A(n_2602),
.Y(n_3177)
);

HB1xp67_ASAP7_75t_L g3178 ( 
.A(n_2647),
.Y(n_3178)
);

BUFx2_ASAP7_75t_R g3179 ( 
.A(n_2703),
.Y(n_3179)
);

NOR2xp33_ASAP7_75t_L g3180 ( 
.A(n_2931),
.B(n_2142),
.Y(n_3180)
);

BUFx2_ASAP7_75t_R g3181 ( 
.A(n_2571),
.Y(n_3181)
);

INVx1_ASAP7_75t_L g3182 ( 
.A(n_2786),
.Y(n_3182)
);

INVx2_ASAP7_75t_L g3183 ( 
.A(n_2810),
.Y(n_3183)
);

BUFx6f_ASAP7_75t_L g3184 ( 
.A(n_2906),
.Y(n_3184)
);

INVx3_ASAP7_75t_L g3185 ( 
.A(n_2906),
.Y(n_3185)
);

INVx2_ASAP7_75t_L g3186 ( 
.A(n_2887),
.Y(n_3186)
);

OAI22xp33_ASAP7_75t_L g3187 ( 
.A1(n_2672),
.A2(n_2541),
.B1(n_2543),
.B2(n_2524),
.Y(n_3187)
);

BUFx3_ASAP7_75t_L g3188 ( 
.A(n_2792),
.Y(n_3188)
);

INVx1_ASAP7_75t_L g3189 ( 
.A(n_2857),
.Y(n_3189)
);

INVx1_ASAP7_75t_L g3190 ( 
.A(n_2871),
.Y(n_3190)
);

INVx2_ASAP7_75t_L g3191 ( 
.A(n_2883),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2636),
.Y(n_3192)
);

BUFx2_ASAP7_75t_SL g3193 ( 
.A(n_2665),
.Y(n_3193)
);

INVx1_ASAP7_75t_L g3194 ( 
.A(n_2782),
.Y(n_3194)
);

NOR2xp33_ASAP7_75t_L g3195 ( 
.A(n_2943),
.B(n_2547),
.Y(n_3195)
);

AND2x2_ASAP7_75t_L g3196 ( 
.A(n_2867),
.B(n_2147),
.Y(n_3196)
);

HB1xp67_ASAP7_75t_L g3197 ( 
.A(n_2961),
.Y(n_3197)
);

AO21x1_ASAP7_75t_L g3198 ( 
.A1(n_2968),
.A2(n_2503),
.B(n_2388),
.Y(n_3198)
);

INVx1_ASAP7_75t_L g3199 ( 
.A(n_2782),
.Y(n_3199)
);

AOI22xp33_ASAP7_75t_L g3200 ( 
.A1(n_2956),
.A2(n_2381),
.B1(n_2356),
.B2(n_2503),
.Y(n_3200)
);

AND2x2_ASAP7_75t_L g3201 ( 
.A(n_2867),
.B(n_554),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_2794),
.Y(n_3202)
);

INVx1_ASAP7_75t_L g3203 ( 
.A(n_2794),
.Y(n_3203)
);

INVx1_ASAP7_75t_L g3204 ( 
.A(n_2814),
.Y(n_3204)
);

CKINVDCx5p33_ASAP7_75t_R g3205 ( 
.A(n_2708),
.Y(n_3205)
);

INVx1_ASAP7_75t_L g3206 ( 
.A(n_2814),
.Y(n_3206)
);

INVx2_ASAP7_75t_SL g3207 ( 
.A(n_2853),
.Y(n_3207)
);

OAI22xp5_ASAP7_75t_L g3208 ( 
.A1(n_2961),
.A2(n_2724),
.B1(n_2881),
.B2(n_2975),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_2916),
.B(n_555),
.Y(n_3209)
);

AOI22xp33_ASAP7_75t_L g3210 ( 
.A1(n_2956),
.A2(n_557),
.B1(n_555),
.B2(n_556),
.Y(n_3210)
);

INVx2_ASAP7_75t_L g3211 ( 
.A(n_2664),
.Y(n_3211)
);

INVx3_ASAP7_75t_L g3212 ( 
.A(n_2569),
.Y(n_3212)
);

INVx3_ASAP7_75t_L g3213 ( 
.A(n_2569),
.Y(n_3213)
);

CKINVDCx6p67_ASAP7_75t_R g3214 ( 
.A(n_2669),
.Y(n_3214)
);

INVx5_ASAP7_75t_L g3215 ( 
.A(n_2692),
.Y(n_3215)
);

BUFx2_ASAP7_75t_R g3216 ( 
.A(n_2951),
.Y(n_3216)
);

INVx3_ASAP7_75t_L g3217 ( 
.A(n_2582),
.Y(n_3217)
);

NOR2xp33_ASAP7_75t_L g3218 ( 
.A(n_2943),
.B(n_556),
.Y(n_3218)
);

HB1xp67_ASAP7_75t_L g3219 ( 
.A(n_2695),
.Y(n_3219)
);

INVx1_ASAP7_75t_L g3220 ( 
.A(n_2817),
.Y(n_3220)
);

AOI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_2956),
.A2(n_559),
.B1(n_557),
.B2(n_558),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_2817),
.Y(n_3222)
);

OAI21x1_ASAP7_75t_L g3223 ( 
.A1(n_2699),
.A2(n_558),
.B(n_559),
.Y(n_3223)
);

AOI22xp5_ASAP7_75t_L g3224 ( 
.A1(n_2928),
.A2(n_562),
.B1(n_560),
.B2(n_561),
.Y(n_3224)
);

AND2x4_ASAP7_75t_L g3225 ( 
.A(n_2582),
.B(n_560),
.Y(n_3225)
);

HB1xp67_ASAP7_75t_L g3226 ( 
.A(n_2697),
.Y(n_3226)
);

BUFx6f_ASAP7_75t_L g3227 ( 
.A(n_2574),
.Y(n_3227)
);

AOI22xp33_ASAP7_75t_L g3228 ( 
.A1(n_2968),
.A2(n_565),
.B1(n_563),
.B2(n_564),
.Y(n_3228)
);

INVx2_ASAP7_75t_L g3229 ( 
.A(n_2690),
.Y(n_3229)
);

INVx1_ASAP7_75t_SL g3230 ( 
.A(n_2831),
.Y(n_3230)
);

INVx3_ASAP7_75t_L g3231 ( 
.A(n_2597),
.Y(n_3231)
);

AND2x2_ASAP7_75t_L g3232 ( 
.A(n_2722),
.B(n_563),
.Y(n_3232)
);

CKINVDCx20_ASAP7_75t_R g3233 ( 
.A(n_2626),
.Y(n_3233)
);

HB1xp67_ASAP7_75t_L g3234 ( 
.A(n_2678),
.Y(n_3234)
);

INVx1_ASAP7_75t_L g3235 ( 
.A(n_2891),
.Y(n_3235)
);

BUFx2_ASAP7_75t_L g3236 ( 
.A(n_2896),
.Y(n_3236)
);

BUFx3_ASAP7_75t_L g3237 ( 
.A(n_2682),
.Y(n_3237)
);

INVx3_ASAP7_75t_L g3238 ( 
.A(n_2597),
.Y(n_3238)
);

AOI22xp33_ASAP7_75t_SL g3239 ( 
.A1(n_2877),
.A2(n_566),
.B1(n_564),
.B2(n_565),
.Y(n_3239)
);

INVx2_ASAP7_75t_L g3240 ( 
.A(n_2696),
.Y(n_3240)
);

AOI22xp33_ASAP7_75t_SL g3241 ( 
.A1(n_2663),
.A2(n_569),
.B1(n_567),
.B2(n_568),
.Y(n_3241)
);

INVx1_ASAP7_75t_L g3242 ( 
.A(n_2891),
.Y(n_3242)
);

AOI22xp33_ASAP7_75t_L g3243 ( 
.A1(n_2959),
.A2(n_571),
.B1(n_569),
.B2(n_570),
.Y(n_3243)
);

INVx3_ASAP7_75t_L g3244 ( 
.A(n_2609),
.Y(n_3244)
);

INVx2_ASAP7_75t_L g3245 ( 
.A(n_2701),
.Y(n_3245)
);

BUFx2_ASAP7_75t_SL g3246 ( 
.A(n_2626),
.Y(n_3246)
);

OAI22xp5_ASAP7_75t_L g3247 ( 
.A1(n_2724),
.A2(n_573),
.B1(n_570),
.B2(n_571),
.Y(n_3247)
);

BUFx3_ASAP7_75t_L g3248 ( 
.A(n_2773),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_L g3249 ( 
.A1(n_2959),
.A2(n_576),
.B1(n_574),
.B2(n_575),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_2965),
.B(n_574),
.Y(n_3250)
);

BUFx2_ASAP7_75t_L g3251 ( 
.A(n_2896),
.Y(n_3251)
);

NAND2xp5_ASAP7_75t_L g3252 ( 
.A(n_2841),
.B(n_577),
.Y(n_3252)
);

AND2x2_ASAP7_75t_L g3253 ( 
.A(n_2607),
.B(n_579),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_2752),
.Y(n_3254)
);

OAI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_2844),
.A2(n_579),
.B(n_580),
.Y(n_3255)
);

AO21x2_ASAP7_75t_L g3256 ( 
.A1(n_2675),
.A2(n_580),
.B(n_581),
.Y(n_3256)
);

INVx2_ASAP7_75t_SL g3257 ( 
.A(n_2853),
.Y(n_3257)
);

INVx1_ASAP7_75t_L g3258 ( 
.A(n_2752),
.Y(n_3258)
);

CKINVDCx20_ASAP7_75t_R g3259 ( 
.A(n_2733),
.Y(n_3259)
);

NAND2xp5_ASAP7_75t_L g3260 ( 
.A(n_2940),
.B(n_581),
.Y(n_3260)
);

INVx1_ASAP7_75t_L g3261 ( 
.A(n_2882),
.Y(n_3261)
);

INVx3_ASAP7_75t_L g3262 ( 
.A(n_2609),
.Y(n_3262)
);

INVx2_ASAP7_75t_SL g3263 ( 
.A(n_2853),
.Y(n_3263)
);

INVx3_ASAP7_75t_L g3264 ( 
.A(n_2839),
.Y(n_3264)
);

HB1xp67_ASAP7_75t_L g3265 ( 
.A(n_2678),
.Y(n_3265)
);

BUFx8_ASAP7_75t_L g3266 ( 
.A(n_2942),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_2882),
.Y(n_3267)
);

AOI21x1_ASAP7_75t_L g3268 ( 
.A1(n_2718),
.A2(n_582),
.B(n_583),
.Y(n_3268)
);

NOR2xp33_ASAP7_75t_L g3269 ( 
.A(n_2942),
.B(n_582),
.Y(n_3269)
);

OAI21xp5_ASAP7_75t_L g3270 ( 
.A1(n_2844),
.A2(n_583),
.B(n_584),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_L g3271 ( 
.A(n_2879),
.B(n_584),
.Y(n_3271)
);

OAI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_2946),
.A2(n_585),
.B(n_586),
.Y(n_3272)
);

INVx2_ASAP7_75t_SL g3273 ( 
.A(n_2839),
.Y(n_3273)
);

CKINVDCx20_ASAP7_75t_R g3274 ( 
.A(n_2824),
.Y(n_3274)
);

AOI22xp33_ASAP7_75t_L g3275 ( 
.A1(n_2953),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_2836),
.Y(n_3276)
);

AOI22xp33_ASAP7_75t_SL g3277 ( 
.A1(n_2767),
.A2(n_589),
.B1(n_587),
.B2(n_588),
.Y(n_3277)
);

AO21x1_ASAP7_75t_L g3278 ( 
.A1(n_2928),
.A2(n_590),
.B(n_591),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_2599),
.Y(n_3279)
);

INVx2_ASAP7_75t_L g3280 ( 
.A(n_2746),
.Y(n_3280)
);

INVxp33_ASAP7_75t_L g3281 ( 
.A(n_2856),
.Y(n_3281)
);

AOI21x1_ASAP7_75t_L g3282 ( 
.A1(n_2718),
.A2(n_590),
.B(n_592),
.Y(n_3282)
);

OAI22xp5_ASAP7_75t_L g3283 ( 
.A1(n_2975),
.A2(n_596),
.B1(n_593),
.B2(n_595),
.Y(n_3283)
);

AOI21x1_ASAP7_75t_L g3284 ( 
.A1(n_2657),
.A2(n_595),
.B(n_596),
.Y(n_3284)
);

OAI22xp33_ASAP7_75t_L g3285 ( 
.A1(n_2791),
.A2(n_599),
.B1(n_597),
.B2(n_598),
.Y(n_3285)
);

INVx6_ASAP7_75t_L g3286 ( 
.A(n_2734),
.Y(n_3286)
);

INVx1_ASAP7_75t_L g3287 ( 
.A(n_2599),
.Y(n_3287)
);

INVx2_ASAP7_75t_SL g3288 ( 
.A(n_2839),
.Y(n_3288)
);

OA21x2_ASAP7_75t_L g3289 ( 
.A1(n_2962),
.A2(n_597),
.B(n_599),
.Y(n_3289)
);

INVx1_ASAP7_75t_L g3290 ( 
.A(n_2610),
.Y(n_3290)
);

BUFx2_ASAP7_75t_L g3291 ( 
.A(n_2896),
.Y(n_3291)
);

BUFx3_ASAP7_75t_L g3292 ( 
.A(n_2854),
.Y(n_3292)
);

CKINVDCx20_ASAP7_75t_R g3293 ( 
.A(n_2708),
.Y(n_3293)
);

INVx3_ASAP7_75t_L g3294 ( 
.A(n_2654),
.Y(n_3294)
);

AND2x2_ASAP7_75t_L g3295 ( 
.A(n_2662),
.B(n_600),
.Y(n_3295)
);

INVx1_ASAP7_75t_L g3296 ( 
.A(n_2610),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_2712),
.Y(n_3297)
);

AOI22xp33_ASAP7_75t_SL g3298 ( 
.A1(n_2576),
.A2(n_2790),
.B1(n_2921),
.B2(n_2885),
.Y(n_3298)
);

INVx1_ASAP7_75t_L g3299 ( 
.A(n_2712),
.Y(n_3299)
);

INVx2_ASAP7_75t_L g3300 ( 
.A(n_2967),
.Y(n_3300)
);

BUFx2_ASAP7_75t_R g3301 ( 
.A(n_2788),
.Y(n_3301)
);

BUFx4f_ASAP7_75t_SL g3302 ( 
.A(n_2727),
.Y(n_3302)
);

AOI22xp33_ASAP7_75t_SL g3303 ( 
.A1(n_2576),
.A2(n_600),
.B1(n_601),
.B2(n_602),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_2808),
.Y(n_3304)
);

AOI22xp33_ASAP7_75t_L g3305 ( 
.A1(n_2953),
.A2(n_601),
.B1(n_603),
.B2(n_604),
.Y(n_3305)
);

NAND2x1p5_ASAP7_75t_L g3306 ( 
.A(n_2734),
.B(n_603),
.Y(n_3306)
);

NAND2x1p5_ASAP7_75t_L g3307 ( 
.A(n_2870),
.B(n_605),
.Y(n_3307)
);

NAND2x1p5_ASAP7_75t_L g3308 ( 
.A(n_2875),
.B(n_605),
.Y(n_3308)
);

BUFx2_ASAP7_75t_L g3309 ( 
.A(n_2921),
.Y(n_3309)
);

BUFx2_ASAP7_75t_R g3310 ( 
.A(n_2897),
.Y(n_3310)
);

OAI21x1_ASAP7_75t_SL g3311 ( 
.A1(n_2588),
.A2(n_606),
.B(n_607),
.Y(n_3311)
);

NAND2xp5_ASAP7_75t_L g3312 ( 
.A(n_2941),
.B(n_606),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_2808),
.Y(n_3313)
);

INVx2_ASAP7_75t_SL g3314 ( 
.A(n_2921),
.Y(n_3314)
);

AOI22xp33_ASAP7_75t_SL g3315 ( 
.A1(n_2576),
.A2(n_607),
.B1(n_608),
.B2(n_609),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_2812),
.Y(n_3316)
);

AND2x2_ASAP7_75t_L g3317 ( 
.A(n_2570),
.B(n_608),
.Y(n_3317)
);

INVx1_ASAP7_75t_L g3318 ( 
.A(n_2812),
.Y(n_3318)
);

CKINVDCx6p67_ASAP7_75t_R g3319 ( 
.A(n_2669),
.Y(n_3319)
);

NAND2xp5_ASAP7_75t_L g3320 ( 
.A(n_2913),
.B(n_610),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_2815),
.Y(n_3321)
);

OAI21x1_ASAP7_75t_L g3322 ( 
.A1(n_2579),
.A2(n_611),
.B(n_612),
.Y(n_3322)
);

AOI22xp33_ASAP7_75t_L g3323 ( 
.A1(n_2934),
.A2(n_615),
.B1(n_616),
.B2(n_617),
.Y(n_3323)
);

INVx1_ASAP7_75t_L g3324 ( 
.A(n_2815),
.Y(n_3324)
);

INVx1_ASAP7_75t_L g3325 ( 
.A(n_2825),
.Y(n_3325)
);

INVx1_ASAP7_75t_L g3326 ( 
.A(n_2825),
.Y(n_3326)
);

OAI22xp33_ASAP7_75t_L g3327 ( 
.A1(n_2791),
.A2(n_615),
.B1(n_616),
.B2(n_617),
.Y(n_3327)
);

INVx1_ASAP7_75t_L g3328 ( 
.A(n_2903),
.Y(n_3328)
);

AND2x4_ASAP7_75t_L g3329 ( 
.A(n_2760),
.B(n_2762),
.Y(n_3329)
);

AOI22xp33_ASAP7_75t_SL g3330 ( 
.A1(n_2790),
.A2(n_618),
.B1(n_619),
.B2(n_620),
.Y(n_3330)
);

AOI22xp33_ASAP7_75t_SL g3331 ( 
.A1(n_2790),
.A2(n_618),
.B1(n_622),
.B2(n_623),
.Y(n_3331)
);

AOI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_2934),
.A2(n_623),
.B1(n_624),
.B2(n_625),
.Y(n_3332)
);

OAI21x1_ASAP7_75t_L g3333 ( 
.A1(n_2590),
.A2(n_626),
.B(n_627),
.Y(n_3333)
);

AOI22xp33_ASAP7_75t_SL g3334 ( 
.A1(n_2692),
.A2(n_627),
.B1(n_628),
.B2(n_629),
.Y(n_3334)
);

INVx1_ASAP7_75t_L g3335 ( 
.A(n_2903),
.Y(n_3335)
);

INVx2_ASAP7_75t_SL g3336 ( 
.A(n_2769),
.Y(n_3336)
);

BUFx4f_ASAP7_75t_SL g3337 ( 
.A(n_2640),
.Y(n_3337)
);

BUFx2_ASAP7_75t_SL g3338 ( 
.A(n_2640),
.Y(n_3338)
);

INVx1_ASAP7_75t_L g3339 ( 
.A(n_2922),
.Y(n_3339)
);

BUFx6f_ASAP7_75t_L g3340 ( 
.A(n_2574),
.Y(n_3340)
);

INVx1_ASAP7_75t_L g3341 ( 
.A(n_2922),
.Y(n_3341)
);

AND2x4_ASAP7_75t_L g3342 ( 
.A(n_2760),
.B(n_628),
.Y(n_3342)
);

BUFx8_ASAP7_75t_L g3343 ( 
.A(n_2919),
.Y(n_3343)
);

INVx1_ASAP7_75t_L g3344 ( 
.A(n_2923),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_2923),
.Y(n_3345)
);

INVx2_ASAP7_75t_L g3346 ( 
.A(n_2763),
.Y(n_3346)
);

BUFx8_ASAP7_75t_L g3347 ( 
.A(n_2598),
.Y(n_3347)
);

INVx3_ASAP7_75t_L g3348 ( 
.A(n_2654),
.Y(n_3348)
);

INVx1_ASAP7_75t_L g3349 ( 
.A(n_2924),
.Y(n_3349)
);

HB1xp67_ASAP7_75t_L g3350 ( 
.A(n_2826),
.Y(n_3350)
);

HB1xp67_ASAP7_75t_L g3351 ( 
.A(n_2901),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_2924),
.Y(n_3352)
);

INVx6_ASAP7_75t_L g3353 ( 
.A(n_2769),
.Y(n_3353)
);

CKINVDCx20_ASAP7_75t_R g3354 ( 
.A(n_2830),
.Y(n_3354)
);

AOI21xp5_ASAP7_75t_L g3355 ( 
.A1(n_2585),
.A2(n_630),
.B(n_632),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_2580),
.B(n_632),
.Y(n_3356)
);

HB1xp67_ASAP7_75t_L g3357 ( 
.A(n_2826),
.Y(n_3357)
);

BUFx2_ASAP7_75t_L g3358 ( 
.A(n_2911),
.Y(n_3358)
);

AO21x2_ASAP7_75t_L g3359 ( 
.A1(n_2661),
.A2(n_633),
.B(n_634),
.Y(n_3359)
);

INVx2_ASAP7_75t_L g3360 ( 
.A(n_2770),
.Y(n_3360)
);

BUFx5_ASAP7_75t_L g3361 ( 
.A(n_3290),
.Y(n_3361)
);

CKINVDCx16_ASAP7_75t_R g3362 ( 
.A(n_3233),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3196),
.B(n_2828),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_2988),
.Y(n_3364)
);

INVx1_ASAP7_75t_L g3365 ( 
.A(n_2990),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3076),
.B(n_2798),
.Y(n_3366)
);

NOR3xp33_ASAP7_75t_SL g3367 ( 
.A(n_3018),
.B(n_2859),
.C(n_2623),
.Y(n_3367)
);

INVx1_ASAP7_75t_L g3368 ( 
.A(n_3001),
.Y(n_3368)
);

NOR2xp33_ASAP7_75t_R g3369 ( 
.A(n_3128),
.B(n_2830),
.Y(n_3369)
);

AOI22xp33_ASAP7_75t_L g3370 ( 
.A1(n_2992),
.A2(n_2791),
.B1(n_2925),
.B2(n_2859),
.Y(n_3370)
);

INVx2_ASAP7_75t_L g3371 ( 
.A(n_3032),
.Y(n_3371)
);

NAND2xp5_ASAP7_75t_L g3372 ( 
.A(n_3004),
.B(n_2828),
.Y(n_3372)
);

INVx3_ASAP7_75t_L g3373 ( 
.A(n_3286),
.Y(n_3373)
);

CKINVDCx20_ASAP7_75t_R g3374 ( 
.A(n_3099),
.Y(n_3374)
);

AOI22xp33_ASAP7_75t_L g3375 ( 
.A1(n_2992),
.A2(n_2954),
.B1(n_2948),
.B2(n_2976),
.Y(n_3375)
);

OR2x2_ASAP7_75t_L g3376 ( 
.A(n_3148),
.B(n_2819),
.Y(n_3376)
);

INVx1_ASAP7_75t_L g3377 ( 
.A(n_3006),
.Y(n_3377)
);

AND2x2_ASAP7_75t_L g3378 ( 
.A(n_3253),
.B(n_2955),
.Y(n_3378)
);

AOI22xp33_ASAP7_75t_L g3379 ( 
.A1(n_3083),
.A2(n_2954),
.B1(n_2948),
.B2(n_2955),
.Y(n_3379)
);

HB1xp67_ASAP7_75t_L g3380 ( 
.A(n_3139),
.Y(n_3380)
);

INVxp67_ASAP7_75t_L g3381 ( 
.A(n_3065),
.Y(n_3381)
);

CKINVDCx5p33_ASAP7_75t_R g3382 ( 
.A(n_3099),
.Y(n_3382)
);

INVx1_ASAP7_75t_L g3383 ( 
.A(n_3010),
.Y(n_3383)
);

HB1xp67_ASAP7_75t_L g3384 ( 
.A(n_2986),
.Y(n_3384)
);

AND2x2_ASAP7_75t_L g3385 ( 
.A(n_3295),
.B(n_2744),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3317),
.B(n_2606),
.Y(n_3386)
);

HB1xp67_ASAP7_75t_L g3387 ( 
.A(n_3137),
.Y(n_3387)
);

OR2x2_ASAP7_75t_L g3388 ( 
.A(n_3148),
.B(n_2949),
.Y(n_3388)
);

OR2x6_ASAP7_75t_L g3389 ( 
.A(n_3052),
.B(n_2918),
.Y(n_3389)
);

INVx2_ASAP7_75t_L g3390 ( 
.A(n_2985),
.Y(n_3390)
);

AND2x4_ASAP7_75t_L g3391 ( 
.A(n_3147),
.B(n_2646),
.Y(n_3391)
);

OAI21xp5_ASAP7_75t_SL g3392 ( 
.A1(n_3126),
.A2(n_2918),
.B(n_2936),
.Y(n_3392)
);

OR2x2_ASAP7_75t_L g3393 ( 
.A(n_3170),
.B(n_3042),
.Y(n_3393)
);

NAND2xp33_ASAP7_75t_R g3394 ( 
.A(n_3000),
.B(n_2598),
.Y(n_3394)
);

INVx4_ASAP7_75t_L g3395 ( 
.A(n_2989),
.Y(n_3395)
);

AND2x2_ASAP7_75t_L g3396 ( 
.A(n_3356),
.B(n_2914),
.Y(n_3396)
);

INVx2_ASAP7_75t_L g3397 ( 
.A(n_2987),
.Y(n_3397)
);

AND2x2_ASAP7_75t_L g3398 ( 
.A(n_3250),
.B(n_2914),
.Y(n_3398)
);

INVx4_ASAP7_75t_L g3399 ( 
.A(n_3092),
.Y(n_3399)
);

AND2x2_ASAP7_75t_L g3400 ( 
.A(n_3232),
.B(n_2914),
.Y(n_3400)
);

INVx2_ASAP7_75t_SL g3401 ( 
.A(n_3092),
.Y(n_3401)
);

INVx2_ASAP7_75t_L g3402 ( 
.A(n_2991),
.Y(n_3402)
);

NOR2xp33_ASAP7_75t_R g3403 ( 
.A(n_3121),
.B(n_2912),
.Y(n_3403)
);

INVxp67_ASAP7_75t_L g3404 ( 
.A(n_3146),
.Y(n_3404)
);

BUFx3_ASAP7_75t_L g3405 ( 
.A(n_3123),
.Y(n_3405)
);

AND2x2_ASAP7_75t_L g3406 ( 
.A(n_3209),
.B(n_2833),
.Y(n_3406)
);

BUFx6f_ASAP7_75t_L g3407 ( 
.A(n_3134),
.Y(n_3407)
);

INVx1_ASAP7_75t_L g3408 ( 
.A(n_3011),
.Y(n_3408)
);

CKINVDCx5p33_ASAP7_75t_R g3409 ( 
.A(n_3033),
.Y(n_3409)
);

BUFx2_ASAP7_75t_L g3410 ( 
.A(n_3350),
.Y(n_3410)
);

INVx2_ASAP7_75t_L g3411 ( 
.A(n_2995),
.Y(n_3411)
);

INVx1_ASAP7_75t_L g3412 ( 
.A(n_3017),
.Y(n_3412)
);

INVx1_ASAP7_75t_L g3413 ( 
.A(n_3021),
.Y(n_3413)
);

INVx2_ASAP7_75t_L g3414 ( 
.A(n_2999),
.Y(n_3414)
);

NAND2xp5_ASAP7_75t_L g3415 ( 
.A(n_3026),
.B(n_2963),
.Y(n_3415)
);

INVx2_ASAP7_75t_L g3416 ( 
.A(n_3079),
.Y(n_3416)
);

INVx2_ASAP7_75t_L g3417 ( 
.A(n_3095),
.Y(n_3417)
);

AND2x4_ASAP7_75t_L g3418 ( 
.A(n_3147),
.B(n_2646),
.Y(n_3418)
);

AND2x4_ASAP7_75t_L g3419 ( 
.A(n_3147),
.B(n_2693),
.Y(n_3419)
);

BUFx3_ASAP7_75t_L g3420 ( 
.A(n_3130),
.Y(n_3420)
);

NAND2xp5_ASAP7_75t_L g3421 ( 
.A(n_3035),
.B(n_2963),
.Y(n_3421)
);

AOI222xp33_ASAP7_75t_L g3422 ( 
.A1(n_2998),
.A2(n_2755),
.B1(n_2829),
.B2(n_2676),
.C1(n_2946),
.C2(n_2920),
.Y(n_3422)
);

NAND2xp33_ASAP7_75t_R g3423 ( 
.A(n_3073),
.B(n_3053),
.Y(n_3423)
);

BUFx6f_ASAP7_75t_L g3424 ( 
.A(n_3134),
.Y(n_3424)
);

BUFx10_ASAP7_75t_L g3425 ( 
.A(n_2981),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3074),
.B(n_2899),
.Y(n_3426)
);

AND2x2_ASAP7_75t_L g3427 ( 
.A(n_3201),
.B(n_2910),
.Y(n_3427)
);

NAND2xp33_ASAP7_75t_R g3428 ( 
.A(n_3236),
.B(n_2693),
.Y(n_3428)
);

CKINVDCx16_ASAP7_75t_R g3429 ( 
.A(n_3274),
.Y(n_3429)
);

NOR3xp33_ASAP7_75t_SL g3430 ( 
.A(n_3205),
.B(n_2623),
.C(n_2829),
.Y(n_3430)
);

INVxp67_ASAP7_75t_L g3431 ( 
.A(n_3188),
.Y(n_3431)
);

INVx2_ASAP7_75t_L g3432 ( 
.A(n_3105),
.Y(n_3432)
);

AO31x2_ASAP7_75t_L g3433 ( 
.A1(n_3198),
.A2(n_2775),
.A3(n_2915),
.B(n_2802),
.Y(n_3433)
);

OR2x6_ASAP7_75t_L g3434 ( 
.A(n_3052),
.B(n_2866),
.Y(n_3434)
);

HB1xp67_ASAP7_75t_SL g3435 ( 
.A(n_3181),
.Y(n_3435)
);

INVx3_ASAP7_75t_SL g3436 ( 
.A(n_3084),
.Y(n_3436)
);

CKINVDCx16_ASAP7_75t_R g3437 ( 
.A(n_3293),
.Y(n_3437)
);

CKINVDCx8_ASAP7_75t_R g3438 ( 
.A(n_3193),
.Y(n_3438)
);

NOR2xp33_ASAP7_75t_R g3439 ( 
.A(n_3266),
.B(n_2866),
.Y(n_3439)
);

AND2x2_ASAP7_75t_L g3440 ( 
.A(n_3172),
.B(n_2898),
.Y(n_3440)
);

AND2x4_ASAP7_75t_L g3441 ( 
.A(n_3215),
.B(n_2711),
.Y(n_3441)
);

CKINVDCx5p33_ASAP7_75t_R g3442 ( 
.A(n_3175),
.Y(n_3442)
);

NAND2xp5_ASAP7_75t_L g3443 ( 
.A(n_3038),
.B(n_2930),
.Y(n_3443)
);

BUFx4f_ASAP7_75t_SL g3444 ( 
.A(n_3120),
.Y(n_3444)
);

OR2x6_ASAP7_75t_L g3445 ( 
.A(n_3052),
.B(n_2866),
.Y(n_3445)
);

INVx1_ASAP7_75t_L g3446 ( 
.A(n_3039),
.Y(n_3446)
);

OAI22xp33_ASAP7_75t_L g3447 ( 
.A1(n_3214),
.A2(n_2717),
.B1(n_2936),
.B2(n_2604),
.Y(n_3447)
);

A2O1A1Ixp33_ASAP7_75t_L g3448 ( 
.A1(n_3126),
.A2(n_3019),
.B(n_3218),
.C(n_3224),
.Y(n_3448)
);

AOI22xp33_ASAP7_75t_L g3449 ( 
.A1(n_3083),
.A2(n_2948),
.B1(n_2954),
.B2(n_2898),
.Y(n_3449)
);

NOR2xp33_ASAP7_75t_R g3450 ( 
.A(n_3266),
.B(n_2692),
.Y(n_3450)
);

AND2x2_ASAP7_75t_L g3451 ( 
.A(n_3157),
.B(n_2811),
.Y(n_3451)
);

BUFx6f_ASAP7_75t_L g3452 ( 
.A(n_3134),
.Y(n_3452)
);

INVx3_ASAP7_75t_L g3453 ( 
.A(n_3286),
.Y(n_3453)
);

OAI21xp5_ASAP7_75t_L g3454 ( 
.A1(n_3002),
.A2(n_2966),
.B(n_2958),
.Y(n_3454)
);

AOI22xp33_ASAP7_75t_L g3455 ( 
.A1(n_2983),
.A2(n_2950),
.B1(n_2676),
.B2(n_2971),
.Y(n_3455)
);

AND2x2_ASAP7_75t_L g3456 ( 
.A(n_3042),
.B(n_2848),
.Y(n_3456)
);

AO31x2_ASAP7_75t_L g3457 ( 
.A1(n_3171),
.A2(n_2802),
.A3(n_2972),
.B(n_2938),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3061),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3069),
.Y(n_3459)
);

OAI22xp5_ASAP7_75t_L g3460 ( 
.A1(n_3005),
.A2(n_2717),
.B1(n_2604),
.B2(n_2683),
.Y(n_3460)
);

INVx3_ASAP7_75t_L g3461 ( 
.A(n_2982),
.Y(n_3461)
);

BUFx6f_ASAP7_75t_L g3462 ( 
.A(n_3184),
.Y(n_3462)
);

AOI22xp33_ASAP7_75t_SL g3463 ( 
.A1(n_3096),
.A2(n_2602),
.B1(n_2838),
.B2(n_2785),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3070),
.Y(n_3464)
);

NAND2xp5_ASAP7_75t_SL g3465 ( 
.A(n_3093),
.B(n_3096),
.Y(n_3465)
);

INVx1_ASAP7_75t_L g3466 ( 
.A(n_3072),
.Y(n_3466)
);

INVx1_ASAP7_75t_L g3467 ( 
.A(n_3081),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3071),
.B(n_2805),
.Y(n_3468)
);

AND2x2_ASAP7_75t_L g3469 ( 
.A(n_3071),
.B(n_2807),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_SL g3470 ( 
.A(n_3093),
.B(n_2602),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_R g3471 ( 
.A(n_3347),
.B(n_2602),
.Y(n_3471)
);

INVx2_ASAP7_75t_L g3472 ( 
.A(n_3113),
.Y(n_3472)
);

NAND2xp33_ASAP7_75t_R g3473 ( 
.A(n_3251),
.B(n_2614),
.Y(n_3473)
);

CKINVDCx20_ASAP7_75t_R g3474 ( 
.A(n_3302),
.Y(n_3474)
);

CKINVDCx5p33_ASAP7_75t_R g3475 ( 
.A(n_3097),
.Y(n_3475)
);

AOI22xp33_ASAP7_75t_L g3476 ( 
.A1(n_3090),
.A2(n_2996),
.B1(n_3014),
.B2(n_3027),
.Y(n_3476)
);

NAND2xp5_ASAP7_75t_L g3477 ( 
.A(n_3102),
.B(n_2765),
.Y(n_3477)
);

OAI22xp5_ASAP7_75t_L g3478 ( 
.A1(n_3224),
.A2(n_2683),
.B1(n_2783),
.B2(n_2789),
.Y(n_3478)
);

NAND2xp33_ASAP7_75t_R g3479 ( 
.A(n_3291),
.B(n_2890),
.Y(n_3479)
);

CKINVDCx5p33_ASAP7_75t_R g3480 ( 
.A(n_3097),
.Y(n_3480)
);

NAND2xp5_ASAP7_75t_L g3481 ( 
.A(n_3103),
.B(n_2765),
.Y(n_3481)
);

OR2x6_ASAP7_75t_L g3482 ( 
.A(n_3029),
.B(n_2652),
.Y(n_3482)
);

BUFx6f_ASAP7_75t_L g3483 ( 
.A(n_3184),
.Y(n_3483)
);

INVx1_ASAP7_75t_SL g3484 ( 
.A(n_3181),
.Y(n_3484)
);

BUFx3_ASAP7_75t_L g3485 ( 
.A(n_3067),
.Y(n_3485)
);

INVx2_ASAP7_75t_L g3486 ( 
.A(n_3114),
.Y(n_3486)
);

OR2x2_ASAP7_75t_L g3487 ( 
.A(n_3170),
.B(n_2816),
.Y(n_3487)
);

NAND2xp5_ASAP7_75t_L g3488 ( 
.A(n_3104),
.B(n_2957),
.Y(n_3488)
);

CKINVDCx8_ASAP7_75t_R g3489 ( 
.A(n_3246),
.Y(n_3489)
);

CKINVDCx16_ASAP7_75t_R g3490 ( 
.A(n_3259),
.Y(n_3490)
);

BUFx3_ASAP7_75t_L g3491 ( 
.A(n_3034),
.Y(n_3491)
);

INVx1_ASAP7_75t_L g3492 ( 
.A(n_3106),
.Y(n_3492)
);

AO31x2_ASAP7_75t_L g3493 ( 
.A1(n_3183),
.A2(n_2972),
.A3(n_2938),
.B(n_2661),
.Y(n_3493)
);

OR2x6_ASAP7_75t_L g3494 ( 
.A(n_3029),
.B(n_2783),
.Y(n_3494)
);

NOR3xp33_ASAP7_75t_SL g3495 ( 
.A(n_3285),
.B(n_2709),
.C(n_2704),
.Y(n_3495)
);

CKINVDCx5p33_ASAP7_75t_R g3496 ( 
.A(n_3354),
.Y(n_3496)
);

AND2x2_ASAP7_75t_L g3497 ( 
.A(n_3164),
.B(n_2843),
.Y(n_3497)
);

AND2x2_ASAP7_75t_L g3498 ( 
.A(n_3036),
.B(n_2779),
.Y(n_3498)
);

NOR3xp33_ASAP7_75t_SL g3499 ( 
.A(n_3327),
.B(n_2709),
.C(n_2704),
.Y(n_3499)
);

NAND2xp5_ASAP7_75t_L g3500 ( 
.A(n_3112),
.B(n_2957),
.Y(n_3500)
);

AOI22xp33_ASAP7_75t_L g3501 ( 
.A1(n_3090),
.A2(n_2950),
.B1(n_2971),
.B2(n_2969),
.Y(n_3501)
);

OAI22xp5_ASAP7_75t_L g3502 ( 
.A1(n_3093),
.A2(n_2789),
.B1(n_2926),
.B2(n_2716),
.Y(n_3502)
);

AND2x2_ASAP7_75t_L g3503 ( 
.A(n_3045),
.B(n_2796),
.Y(n_3503)
);

AND2x2_ASAP7_75t_L g3504 ( 
.A(n_3051),
.B(n_633),
.Y(n_3504)
);

AOI22xp33_ASAP7_75t_L g3505 ( 
.A1(n_3027),
.A2(n_2950),
.B1(n_2971),
.B2(n_2969),
.Y(n_3505)
);

HB1xp67_ASAP7_75t_L g3506 ( 
.A(n_3234),
.Y(n_3506)
);

INVx2_ASAP7_75t_L g3507 ( 
.A(n_3117),
.Y(n_3507)
);

BUFx3_ASAP7_75t_L g3508 ( 
.A(n_3037),
.Y(n_3508)
);

NAND2xp33_ASAP7_75t_R g3509 ( 
.A(n_3309),
.B(n_3129),
.Y(n_3509)
);

NOR3xp33_ASAP7_75t_SL g3510 ( 
.A(n_3187),
.B(n_2650),
.C(n_2860),
.Y(n_3510)
);

NAND2xp5_ASAP7_75t_L g3511 ( 
.A(n_3127),
.B(n_2977),
.Y(n_3511)
);

AOI22xp33_ASAP7_75t_L g3512 ( 
.A1(n_3056),
.A2(n_2977),
.B1(n_2820),
.B2(n_2766),
.Y(n_3512)
);

CKINVDCx5p33_ASAP7_75t_R g3513 ( 
.A(n_3319),
.Y(n_3513)
);

INVx2_ASAP7_75t_SL g3514 ( 
.A(n_2984),
.Y(n_3514)
);

INVx2_ASAP7_75t_L g3515 ( 
.A(n_3136),
.Y(n_3515)
);

AND2x2_ASAP7_75t_L g3516 ( 
.A(n_3054),
.B(n_634),
.Y(n_3516)
);

CKINVDCx16_ASAP7_75t_R g3517 ( 
.A(n_3009),
.Y(n_3517)
);

AND2x2_ASAP7_75t_L g3518 ( 
.A(n_3055),
.B(n_635),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3132),
.Y(n_3519)
);

NOR2xp33_ASAP7_75t_R g3520 ( 
.A(n_3347),
.B(n_2785),
.Y(n_3520)
);

NAND2xp5_ASAP7_75t_L g3521 ( 
.A(n_3080),
.B(n_2847),
.Y(n_3521)
);

NAND3xp33_ASAP7_75t_L g3522 ( 
.A(n_3166),
.B(n_2813),
.C(n_2781),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3116),
.Y(n_3523)
);

AND2x2_ASAP7_75t_L g3524 ( 
.A(n_3059),
.B(n_635),
.Y(n_3524)
);

NAND2xp33_ASAP7_75t_R g3525 ( 
.A(n_3086),
.B(n_2945),
.Y(n_3525)
);

NOR2xp33_ASAP7_75t_L g3526 ( 
.A(n_3180),
.B(n_2860),
.Y(n_3526)
);

INVx2_ASAP7_75t_L g3527 ( 
.A(n_3141),
.Y(n_3527)
);

BUFx3_ASAP7_75t_L g3528 ( 
.A(n_3292),
.Y(n_3528)
);

OR2x2_ASAP7_75t_L g3529 ( 
.A(n_3265),
.B(n_2714),
.Y(n_3529)
);

AND2x2_ASAP7_75t_L g3530 ( 
.A(n_3060),
.B(n_636),
.Y(n_3530)
);

NOR2xp33_ASAP7_75t_R g3531 ( 
.A(n_3337),
.B(n_2785),
.Y(n_3531)
);

CKINVDCx8_ASAP7_75t_R g3532 ( 
.A(n_3338),
.Y(n_3532)
);

INVx1_ASAP7_75t_L g3533 ( 
.A(n_3189),
.Y(n_3533)
);

INVx8_ASAP7_75t_L g3534 ( 
.A(n_3009),
.Y(n_3534)
);

BUFx8_ASAP7_75t_SL g3535 ( 
.A(n_3087),
.Y(n_3535)
);

AND2x4_ASAP7_75t_L g3536 ( 
.A(n_3215),
.B(n_2711),
.Y(n_3536)
);

OAI21xp33_ASAP7_75t_L g3537 ( 
.A1(n_3277),
.A2(n_2926),
.B(n_2939),
.Y(n_3537)
);

CKINVDCx5p33_ASAP7_75t_R g3538 ( 
.A(n_3179),
.Y(n_3538)
);

INVx2_ASAP7_75t_L g3539 ( 
.A(n_3143),
.Y(n_3539)
);

CKINVDCx5p33_ASAP7_75t_R g3540 ( 
.A(n_3179),
.Y(n_3540)
);

OAI22xp5_ASAP7_75t_L g3541 ( 
.A1(n_3163),
.A2(n_2716),
.B1(n_2840),
.B2(n_2801),
.Y(n_3541)
);

NOR2xp33_ASAP7_75t_R g3542 ( 
.A(n_3064),
.B(n_2785),
.Y(n_3542)
);

NOR2x1_ASAP7_75t_L g3543 ( 
.A(n_2982),
.B(n_2834),
.Y(n_3543)
);

HB1xp67_ASAP7_75t_L g3544 ( 
.A(n_3178),
.Y(n_3544)
);

AOI22xp33_ASAP7_75t_L g3545 ( 
.A1(n_3040),
.A2(n_2907),
.B1(n_2909),
.B2(n_2904),
.Y(n_3545)
);

XNOR2x1_ASAP7_75t_L g3546 ( 
.A(n_3237),
.B(n_637),
.Y(n_3546)
);

BUFx2_ASAP7_75t_L g3547 ( 
.A(n_3064),
.Y(n_3547)
);

INVx2_ASAP7_75t_L g3548 ( 
.A(n_3144),
.Y(n_3548)
);

HB1xp67_ASAP7_75t_L g3549 ( 
.A(n_3219),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3190),
.Y(n_3550)
);

AND2x2_ASAP7_75t_L g3551 ( 
.A(n_3062),
.B(n_638),
.Y(n_3551)
);

OR2x2_ASAP7_75t_L g3552 ( 
.A(n_3226),
.B(n_2842),
.Y(n_3552)
);

AND2x2_ASAP7_75t_L g3553 ( 
.A(n_3077),
.B(n_3003),
.Y(n_3553)
);

INVx2_ASAP7_75t_L g3554 ( 
.A(n_3151),
.Y(n_3554)
);

NOR3xp33_ASAP7_75t_SL g3555 ( 
.A(n_3019),
.B(n_2650),
.C(n_2648),
.Y(n_3555)
);

OR2x6_ASAP7_75t_L g3556 ( 
.A(n_3047),
.B(n_2769),
.Y(n_3556)
);

OR2x2_ASAP7_75t_SL g3557 ( 
.A(n_2984),
.B(n_2656),
.Y(n_3557)
);

HB1xp67_ASAP7_75t_L g3558 ( 
.A(n_3350),
.Y(n_3558)
);

OAI21x1_ASAP7_75t_SL g3559 ( 
.A1(n_3016),
.A2(n_2620),
.B(n_2797),
.Y(n_3559)
);

CKINVDCx5p33_ASAP7_75t_R g3560 ( 
.A(n_3100),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3080),
.B(n_2847),
.Y(n_3561)
);

BUFx4f_ASAP7_75t_L g3562 ( 
.A(n_2993),
.Y(n_3562)
);

CKINVDCx11_ASAP7_75t_R g3563 ( 
.A(n_3015),
.Y(n_3563)
);

INVx3_ASAP7_75t_L g3564 ( 
.A(n_3184),
.Y(n_3564)
);

INVx1_ASAP7_75t_L g3565 ( 
.A(n_3186),
.Y(n_3565)
);

INVx1_ASAP7_75t_L g3566 ( 
.A(n_3191),
.Y(n_3566)
);

OR2x6_ASAP7_75t_L g3567 ( 
.A(n_3047),
.B(n_2804),
.Y(n_3567)
);

AND2x4_ASAP7_75t_SL g3568 ( 
.A(n_3066),
.B(n_2842),
.Y(n_3568)
);

AO31x2_ASAP7_75t_L g3569 ( 
.A1(n_3192),
.A2(n_2838),
.A3(n_2785),
.B(n_2630),
.Y(n_3569)
);

INVx1_ASAP7_75t_L g3570 ( 
.A(n_3008),
.Y(n_3570)
);

AND2x2_ASAP7_75t_L g3571 ( 
.A(n_3012),
.B(n_639),
.Y(n_3571)
);

HB1xp67_ASAP7_75t_L g3572 ( 
.A(n_3357),
.Y(n_3572)
);

INVx1_ASAP7_75t_L g3573 ( 
.A(n_3020),
.Y(n_3573)
);

BUFx10_ASAP7_75t_L g3574 ( 
.A(n_2993),
.Y(n_3574)
);

NOR2xp33_ASAP7_75t_L g3575 ( 
.A(n_3281),
.B(n_2743),
.Y(n_3575)
);

A2O1A1Ixp33_ASAP7_75t_L g3576 ( 
.A1(n_3255),
.A2(n_3270),
.B(n_3272),
.C(n_3163),
.Y(n_3576)
);

BUFx4f_ASAP7_75t_L g3577 ( 
.A(n_3306),
.Y(n_3577)
);

INVx1_ASAP7_75t_L g3578 ( 
.A(n_3024),
.Y(n_3578)
);

AO32x1_ASAP7_75t_L g3579 ( 
.A1(n_3208),
.A2(n_2838),
.A3(n_2684),
.B1(n_2666),
.B2(n_2596),
.Y(n_3579)
);

OR2x6_ASAP7_75t_L g3580 ( 
.A(n_3314),
.B(n_2809),
.Y(n_3580)
);

BUFx6f_ASAP7_75t_L g3581 ( 
.A(n_3248),
.Y(n_3581)
);

NOR2xp33_ASAP7_75t_R g3582 ( 
.A(n_3098),
.B(n_2838),
.Y(n_3582)
);

OAI21xp5_ASAP7_75t_SL g3583 ( 
.A1(n_3277),
.A2(n_2840),
.B(n_2801),
.Y(n_3583)
);

CKINVDCx16_ASAP7_75t_R g3584 ( 
.A(n_3022),
.Y(n_3584)
);

AOI22xp5_ASAP7_75t_L g3585 ( 
.A1(n_3049),
.A2(n_2929),
.B1(n_2952),
.B2(n_2880),
.Y(n_3585)
);

CKINVDCx5p33_ASAP7_75t_R g3586 ( 
.A(n_3100),
.Y(n_3586)
);

AND2x2_ASAP7_75t_SL g3587 ( 
.A(n_3156),
.B(n_2656),
.Y(n_3587)
);

AND2x2_ASAP7_75t_L g3588 ( 
.A(n_3030),
.B(n_639),
.Y(n_3588)
);

NAND2xp33_ASAP7_75t_L g3589 ( 
.A(n_3215),
.B(n_2838),
.Y(n_3589)
);

INVx1_ASAP7_75t_L g3590 ( 
.A(n_3031),
.Y(n_3590)
);

AND2x2_ASAP7_75t_L g3591 ( 
.A(n_3044),
.B(n_640),
.Y(n_3591)
);

OAI22xp5_ASAP7_75t_L g3592 ( 
.A1(n_3241),
.A2(n_2855),
.B1(n_2905),
.B2(n_2886),
.Y(n_3592)
);

NAND2xp33_ASAP7_75t_SL g3593 ( 
.A(n_3296),
.B(n_2596),
.Y(n_3593)
);

INVx2_ASAP7_75t_L g3594 ( 
.A(n_3154),
.Y(n_3594)
);

AND2x2_ASAP7_75t_L g3595 ( 
.A(n_3241),
.B(n_640),
.Y(n_3595)
);

AND2x4_ASAP7_75t_L g3596 ( 
.A(n_3098),
.B(n_2648),
.Y(n_3596)
);

AND2x2_ASAP7_75t_L g3597 ( 
.A(n_3225),
.B(n_641),
.Y(n_3597)
);

AND2x2_ASAP7_75t_L g3598 ( 
.A(n_3225),
.B(n_3161),
.Y(n_3598)
);

BUFx3_ASAP7_75t_L g3599 ( 
.A(n_3343),
.Y(n_3599)
);

AND2x2_ASAP7_75t_L g3600 ( 
.A(n_3085),
.B(n_642),
.Y(n_3600)
);

AOI22xp33_ASAP7_75t_L g3601 ( 
.A1(n_3278),
.A2(n_2849),
.B1(n_2973),
.B2(n_2944),
.Y(n_3601)
);

INVx1_ASAP7_75t_L g3602 ( 
.A(n_3261),
.Y(n_3602)
);

AOI22xp33_ASAP7_75t_L g3603 ( 
.A1(n_3131),
.A2(n_2944),
.B1(n_2908),
.B2(n_2979),
.Y(n_3603)
);

AO31x2_ASAP7_75t_L g3604 ( 
.A1(n_3211),
.A2(n_2660),
.A3(n_2687),
.B(n_2715),
.Y(n_3604)
);

BUFx2_ASAP7_75t_L g3605 ( 
.A(n_3358),
.Y(n_3605)
);

INVx2_ASAP7_75t_L g3606 ( 
.A(n_3159),
.Y(n_3606)
);

INVx1_ASAP7_75t_L g3607 ( 
.A(n_3267),
.Y(n_3607)
);

CKINVDCx5p33_ASAP7_75t_R g3608 ( 
.A(n_3343),
.Y(n_3608)
);

HB1xp67_ASAP7_75t_L g3609 ( 
.A(n_3357),
.Y(n_3609)
);

NAND2xp33_ASAP7_75t_SL g3610 ( 
.A(n_3068),
.B(n_2777),
.Y(n_3610)
);

HB1xp67_ASAP7_75t_L g3611 ( 
.A(n_3351),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3260),
.Y(n_3612)
);

AND2x2_ASAP7_75t_L g3613 ( 
.A(n_3085),
.B(n_643),
.Y(n_3613)
);

BUFx4f_ASAP7_75t_L g3614 ( 
.A(n_3306),
.Y(n_3614)
);

OR2x2_ASAP7_75t_L g3615 ( 
.A(n_3107),
.B(n_2762),
.Y(n_3615)
);

CKINVDCx5p33_ASAP7_75t_R g3616 ( 
.A(n_3216),
.Y(n_3616)
);

CKINVDCx16_ASAP7_75t_R g3617 ( 
.A(n_3066),
.Y(n_3617)
);

NAND2xp5_ASAP7_75t_L g3618 ( 
.A(n_3279),
.B(n_2834),
.Y(n_3618)
);

BUFx3_ASAP7_75t_L g3619 ( 
.A(n_3149),
.Y(n_3619)
);

INVx4_ASAP7_75t_R g3620 ( 
.A(n_3048),
.Y(n_3620)
);

INVx3_ASAP7_75t_L g3621 ( 
.A(n_3025),
.Y(n_3621)
);

BUFx2_ASAP7_75t_L g3622 ( 
.A(n_3197),
.Y(n_3622)
);

NAND2xp33_ASAP7_75t_R g3623 ( 
.A(n_3269),
.B(n_2945),
.Y(n_3623)
);

OR2x6_ASAP7_75t_L g3624 ( 
.A(n_3307),
.B(n_2855),
.Y(n_3624)
);

CKINVDCx5p33_ASAP7_75t_R g3625 ( 
.A(n_3216),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3289),
.Y(n_3626)
);

INVx2_ASAP7_75t_L g3627 ( 
.A(n_3289),
.Y(n_3627)
);

HB1xp67_ASAP7_75t_L g3628 ( 
.A(n_3176),
.Y(n_3628)
);

INVx1_ASAP7_75t_L g3629 ( 
.A(n_3260),
.Y(n_3629)
);

NAND2xp33_ASAP7_75t_R g3630 ( 
.A(n_3185),
.B(n_2947),
.Y(n_3630)
);

AND2x4_ASAP7_75t_L g3631 ( 
.A(n_3294),
.B(n_2611),
.Y(n_3631)
);

AOI22xp33_ASAP7_75t_SL g3632 ( 
.A1(n_3297),
.A2(n_2905),
.B1(n_2886),
.B2(n_2947),
.Y(n_3632)
);

BUFx3_ASAP7_75t_L g3633 ( 
.A(n_3158),
.Y(n_3633)
);

CKINVDCx16_ASAP7_75t_R g3634 ( 
.A(n_3109),
.Y(n_3634)
);

NAND2xp5_ASAP7_75t_L g3635 ( 
.A(n_3287),
.B(n_2929),
.Y(n_3635)
);

INVx8_ASAP7_75t_L g3636 ( 
.A(n_3185),
.Y(n_3636)
);

AND2x2_ASAP7_75t_L g3637 ( 
.A(n_3107),
.B(n_643),
.Y(n_3637)
);

AND2x2_ASAP7_75t_L g3638 ( 
.A(n_3239),
.B(n_644),
.Y(n_3638)
);

OR2x2_ASAP7_75t_L g3639 ( 
.A(n_3176),
.B(n_2764),
.Y(n_3639)
);

NOR3xp33_ASAP7_75t_SL g3640 ( 
.A(n_3271),
.B(n_2668),
.C(n_2585),
.Y(n_3640)
);

CKINVDCx8_ASAP7_75t_R g3641 ( 
.A(n_3342),
.Y(n_3641)
);

CKINVDCx5p33_ASAP7_75t_R g3642 ( 
.A(n_3301),
.Y(n_3642)
);

OR2x2_ASAP7_75t_L g3643 ( 
.A(n_3252),
.B(n_2764),
.Y(n_3643)
);

AND2x2_ASAP7_75t_L g3644 ( 
.A(n_3239),
.B(n_644),
.Y(n_3644)
);

AND2x4_ASAP7_75t_L g3645 ( 
.A(n_3294),
.B(n_2611),
.Y(n_3645)
);

INVx1_ASAP7_75t_L g3646 ( 
.A(n_3312),
.Y(n_3646)
);

AND2x2_ASAP7_75t_L g3647 ( 
.A(n_3303),
.B(n_645),
.Y(n_3647)
);

AND2x2_ASAP7_75t_L g3648 ( 
.A(n_3303),
.B(n_3315),
.Y(n_3648)
);

AOI22xp33_ASAP7_75t_L g3649 ( 
.A1(n_3131),
.A2(n_2944),
.B1(n_2908),
.B2(n_2979),
.Y(n_3649)
);

INVx1_ASAP7_75t_L g3650 ( 
.A(n_3312),
.Y(n_3650)
);

INVx2_ASAP7_75t_L g3651 ( 
.A(n_3300),
.Y(n_3651)
);

AOI22xp33_ASAP7_75t_L g3652 ( 
.A1(n_3131),
.A2(n_2908),
.B1(n_2979),
.B2(n_2952),
.Y(n_3652)
);

O2A1O1Ixp33_ASAP7_75t_L g3653 ( 
.A1(n_3023),
.A2(n_2846),
.B(n_2869),
.C(n_2863),
.Y(n_3653)
);

AND2x2_ASAP7_75t_L g3654 ( 
.A(n_3315),
.B(n_645),
.Y(n_3654)
);

AOI22xp5_ASAP7_75t_L g3655 ( 
.A1(n_3058),
.A2(n_2880),
.B1(n_2706),
.B2(n_2863),
.Y(n_3655)
);

HB1xp67_ASAP7_75t_L g3656 ( 
.A(n_3194),
.Y(n_3656)
);

NOR2xp33_ASAP7_75t_R g3657 ( 
.A(n_3207),
.B(n_2864),
.Y(n_3657)
);

NAND2xp5_ASAP7_75t_L g3658 ( 
.A(n_3023),
.B(n_2777),
.Y(n_3658)
);

OAI222xp33_ASAP7_75t_L g3659 ( 
.A1(n_3334),
.A2(n_2937),
.B1(n_2632),
.B2(n_2633),
.C1(n_2644),
.C2(n_2668),
.Y(n_3659)
);

CKINVDCx20_ASAP7_75t_R g3660 ( 
.A(n_3091),
.Y(n_3660)
);

INVx2_ASAP7_75t_L g3661 ( 
.A(n_3223),
.Y(n_3661)
);

BUFx6f_ASAP7_75t_L g3662 ( 
.A(n_3257),
.Y(n_3662)
);

INVx1_ASAP7_75t_L g3663 ( 
.A(n_3320),
.Y(n_3663)
);

AND2x4_ASAP7_75t_L g3664 ( 
.A(n_3348),
.B(n_3212),
.Y(n_3664)
);

INVx1_ASAP7_75t_L g3665 ( 
.A(n_3320),
.Y(n_3665)
);

INVx1_ASAP7_75t_L g3666 ( 
.A(n_3252),
.Y(n_3666)
);

AND2x2_ASAP7_75t_L g3667 ( 
.A(n_3330),
.B(n_646),
.Y(n_3667)
);

NAND2xp5_ASAP7_75t_L g3668 ( 
.A(n_3140),
.B(n_2706),
.Y(n_3668)
);

NAND2xp33_ASAP7_75t_R g3669 ( 
.A(n_3264),
.B(n_2628),
.Y(n_3669)
);

INVx2_ASAP7_75t_L g3670 ( 
.A(n_3322),
.Y(n_3670)
);

AND2x2_ASAP7_75t_L g3671 ( 
.A(n_3330),
.B(n_646),
.Y(n_3671)
);

AND2x4_ASAP7_75t_SL g3672 ( 
.A(n_3263),
.B(n_2632),
.Y(n_3672)
);

INVx3_ASAP7_75t_L g3673 ( 
.A(n_3025),
.Y(n_3673)
);

BUFx2_ASAP7_75t_L g3674 ( 
.A(n_3197),
.Y(n_3674)
);

AND2x2_ASAP7_75t_L g3675 ( 
.A(n_3331),
.B(n_647),
.Y(n_3675)
);

NAND2xp5_ASAP7_75t_L g3676 ( 
.A(n_3142),
.B(n_3150),
.Y(n_3676)
);

CKINVDCx16_ASAP7_75t_R g3677 ( 
.A(n_3048),
.Y(n_3677)
);

OR2x2_ASAP7_75t_L g3678 ( 
.A(n_3254),
.B(n_2633),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3276),
.Y(n_3679)
);

NAND2xp5_ASAP7_75t_L g3680 ( 
.A(n_3153),
.B(n_2869),
.Y(n_3680)
);

INVx2_ASAP7_75t_SL g3681 ( 
.A(n_3050),
.Y(n_3681)
);

AND2x2_ASAP7_75t_L g3682 ( 
.A(n_3331),
.B(n_647),
.Y(n_3682)
);

INVx1_ASAP7_75t_L g3683 ( 
.A(n_3199),
.Y(n_3683)
);

CKINVDCx5p33_ASAP7_75t_R g3684 ( 
.A(n_3301),
.Y(n_3684)
);

CKINVDCx5p33_ASAP7_75t_R g3685 ( 
.A(n_3310),
.Y(n_3685)
);

INVx1_ASAP7_75t_L g3686 ( 
.A(n_3202),
.Y(n_3686)
);

BUFx3_ASAP7_75t_L g3687 ( 
.A(n_3050),
.Y(n_3687)
);

HB1xp67_ASAP7_75t_L g3688 ( 
.A(n_3203),
.Y(n_3688)
);

NAND4xp25_ASAP7_75t_L g3689 ( 
.A(n_3243),
.B(n_3249),
.C(n_3046),
.D(n_3108),
.Y(n_3689)
);

INVx4_ASAP7_75t_SL g3690 ( 
.A(n_3353),
.Y(n_3690)
);

OR2x2_ASAP7_75t_L g3691 ( 
.A(n_3258),
.B(n_2644),
.Y(n_3691)
);

NOR3xp33_ASAP7_75t_SL g3692 ( 
.A(n_3247),
.B(n_2902),
.C(n_2873),
.Y(n_3692)
);

NAND2xp33_ASAP7_75t_R g3693 ( 
.A(n_3264),
.B(n_648),
.Y(n_3693)
);

INVxp33_ASAP7_75t_L g3694 ( 
.A(n_3152),
.Y(n_3694)
);

CKINVDCx5p33_ASAP7_75t_R g3695 ( 
.A(n_3310),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_L g3696 ( 
.A(n_3152),
.B(n_2643),
.Y(n_3696)
);

NAND2xp33_ASAP7_75t_R g3697 ( 
.A(n_3342),
.B(n_648),
.Y(n_3697)
);

AND2x4_ASAP7_75t_SL g3698 ( 
.A(n_3273),
.B(n_3288),
.Y(n_3698)
);

CKINVDCx16_ASAP7_75t_R g3699 ( 
.A(n_3177),
.Y(n_3699)
);

INVx2_ASAP7_75t_L g3700 ( 
.A(n_3390),
.Y(n_3700)
);

AND2x2_ASAP7_75t_L g3701 ( 
.A(n_3366),
.B(n_3204),
.Y(n_3701)
);

INVx1_ASAP7_75t_L g3702 ( 
.A(n_3651),
.Y(n_3702)
);

INVx1_ASAP7_75t_L g3703 ( 
.A(n_3680),
.Y(n_3703)
);

INVx1_ASAP7_75t_L g3704 ( 
.A(n_3668),
.Y(n_3704)
);

INVx1_ASAP7_75t_L g3705 ( 
.A(n_3618),
.Y(n_3705)
);

INVx1_ASAP7_75t_L g3706 ( 
.A(n_3635),
.Y(n_3706)
);

AND2x2_ASAP7_75t_L g3707 ( 
.A(n_3440),
.B(n_3206),
.Y(n_3707)
);

O2A1O1Ixp5_ASAP7_75t_L g3708 ( 
.A1(n_3577),
.A2(n_3283),
.B(n_3270),
.C(n_3255),
.Y(n_3708)
);

INVx2_ASAP7_75t_L g3709 ( 
.A(n_3397),
.Y(n_3709)
);

INVx2_ASAP7_75t_L g3710 ( 
.A(n_3402),
.Y(n_3710)
);

BUFx2_ASAP7_75t_L g3711 ( 
.A(n_3557),
.Y(n_3711)
);

AND2x2_ASAP7_75t_L g3712 ( 
.A(n_3456),
.B(n_3220),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3602),
.Y(n_3713)
);

HB1xp67_ASAP7_75t_L g3714 ( 
.A(n_3558),
.Y(n_3714)
);

INVx1_ASAP7_75t_L g3715 ( 
.A(n_3607),
.Y(n_3715)
);

INVx2_ASAP7_75t_L g3716 ( 
.A(n_3411),
.Y(n_3716)
);

INVx2_ASAP7_75t_L g3717 ( 
.A(n_3414),
.Y(n_3717)
);

INVx2_ASAP7_75t_L g3718 ( 
.A(n_3416),
.Y(n_3718)
);

BUFx12f_ASAP7_75t_L g3719 ( 
.A(n_3382),
.Y(n_3719)
);

INVx1_ASAP7_75t_L g3720 ( 
.A(n_3364),
.Y(n_3720)
);

NOR2xp33_ASAP7_75t_L g3721 ( 
.A(n_3634),
.B(n_3307),
.Y(n_3721)
);

INVx1_ASAP7_75t_L g3722 ( 
.A(n_3365),
.Y(n_3722)
);

INVx2_ASAP7_75t_L g3723 ( 
.A(n_3417),
.Y(n_3723)
);

INVx1_ASAP7_75t_L g3724 ( 
.A(n_3368),
.Y(n_3724)
);

INVx1_ASAP7_75t_L g3725 ( 
.A(n_3377),
.Y(n_3725)
);

INVx2_ASAP7_75t_L g3726 ( 
.A(n_3432),
.Y(n_3726)
);

OAI22xp5_ASAP7_75t_L g3727 ( 
.A1(n_3641),
.A2(n_3298),
.B1(n_3210),
.B2(n_3221),
.Y(n_3727)
);

NAND2xp5_ASAP7_75t_L g3728 ( 
.A(n_3363),
.B(n_3553),
.Y(n_3728)
);

AND2x2_ASAP7_75t_L g3729 ( 
.A(n_3426),
.B(n_3386),
.Y(n_3729)
);

HB1xp67_ASAP7_75t_L g3730 ( 
.A(n_3572),
.Y(n_3730)
);

INVx3_ASAP7_75t_L g3731 ( 
.A(n_3677),
.Y(n_3731)
);

AND2x2_ASAP7_75t_L g3732 ( 
.A(n_3387),
.B(n_3222),
.Y(n_3732)
);

INVx1_ASAP7_75t_L g3733 ( 
.A(n_3383),
.Y(n_3733)
);

HB1xp67_ASAP7_75t_L g3734 ( 
.A(n_3609),
.Y(n_3734)
);

OR2x2_ASAP7_75t_L g3735 ( 
.A(n_3384),
.B(n_3115),
.Y(n_3735)
);

BUFx2_ASAP7_75t_L g3736 ( 
.A(n_3699),
.Y(n_3736)
);

INVx1_ASAP7_75t_L g3737 ( 
.A(n_3408),
.Y(n_3737)
);

INVx1_ASAP7_75t_L g3738 ( 
.A(n_3412),
.Y(n_3738)
);

BUFx2_ASAP7_75t_SL g3739 ( 
.A(n_3438),
.Y(n_3739)
);

BUFx3_ASAP7_75t_L g3740 ( 
.A(n_3405),
.Y(n_3740)
);

INVx2_ASAP7_75t_L g3741 ( 
.A(n_3472),
.Y(n_3741)
);

AND2x2_ASAP7_75t_L g3742 ( 
.A(n_3406),
.B(n_3348),
.Y(n_3742)
);

NAND2xp5_ASAP7_75t_L g3743 ( 
.A(n_3523),
.B(n_3160),
.Y(n_3743)
);

AND2x2_ASAP7_75t_L g3744 ( 
.A(n_3378),
.B(n_3212),
.Y(n_3744)
);

INVx2_ASAP7_75t_SL g3745 ( 
.A(n_3534),
.Y(n_3745)
);

INVx1_ASAP7_75t_L g3746 ( 
.A(n_3413),
.Y(n_3746)
);

AOI22xp33_ASAP7_75t_L g3747 ( 
.A1(n_3648),
.A2(n_3063),
.B1(n_3135),
.B2(n_3078),
.Y(n_3747)
);

INVx1_ASAP7_75t_L g3748 ( 
.A(n_3446),
.Y(n_3748)
);

INVx2_ASAP7_75t_L g3749 ( 
.A(n_3486),
.Y(n_3749)
);

INVx1_ASAP7_75t_L g3750 ( 
.A(n_3458),
.Y(n_3750)
);

HB1xp67_ASAP7_75t_L g3751 ( 
.A(n_3410),
.Y(n_3751)
);

OR2x2_ASAP7_75t_L g3752 ( 
.A(n_3506),
.B(n_3115),
.Y(n_3752)
);

INVx1_ASAP7_75t_L g3753 ( 
.A(n_3459),
.Y(n_3753)
);

INVx1_ASAP7_75t_L g3754 ( 
.A(n_3464),
.Y(n_3754)
);

INVx1_ASAP7_75t_L g3755 ( 
.A(n_3466),
.Y(n_3755)
);

INVx1_ASAP7_75t_L g3756 ( 
.A(n_3467),
.Y(n_3756)
);

AND2x2_ASAP7_75t_L g3757 ( 
.A(n_3598),
.B(n_3213),
.Y(n_3757)
);

INVxp67_ASAP7_75t_L g3758 ( 
.A(n_3611),
.Y(n_3758)
);

INVx2_ASAP7_75t_L g3759 ( 
.A(n_3507),
.Y(n_3759)
);

INVx3_ASAP7_75t_L g3760 ( 
.A(n_3391),
.Y(n_3760)
);

INVx2_ASAP7_75t_L g3761 ( 
.A(n_3515),
.Y(n_3761)
);

AND2x2_ASAP7_75t_L g3762 ( 
.A(n_3396),
.B(n_3213),
.Y(n_3762)
);

INVx2_ASAP7_75t_L g3763 ( 
.A(n_3527),
.Y(n_3763)
);

INVx2_ASAP7_75t_L g3764 ( 
.A(n_3539),
.Y(n_3764)
);

OR2x2_ASAP7_75t_L g3765 ( 
.A(n_3380),
.B(n_3162),
.Y(n_3765)
);

OR2x6_ASAP7_75t_L g3766 ( 
.A(n_3482),
.B(n_3308),
.Y(n_3766)
);

INVxp67_ASAP7_75t_SL g3767 ( 
.A(n_3410),
.Y(n_3767)
);

INVx2_ASAP7_75t_L g3768 ( 
.A(n_3548),
.Y(n_3768)
);

INVx1_ASAP7_75t_L g3769 ( 
.A(n_3492),
.Y(n_3769)
);

INVx1_ASAP7_75t_L g3770 ( 
.A(n_3519),
.Y(n_3770)
);

BUFx6f_ASAP7_75t_L g3771 ( 
.A(n_3407),
.Y(n_3771)
);

AND2x2_ASAP7_75t_L g3772 ( 
.A(n_3498),
.B(n_3217),
.Y(n_3772)
);

INVx1_ASAP7_75t_L g3773 ( 
.A(n_3533),
.Y(n_3773)
);

OR2x2_ASAP7_75t_L g3774 ( 
.A(n_3393),
.B(n_3165),
.Y(n_3774)
);

AND2x4_ASAP7_75t_L g3775 ( 
.A(n_3622),
.B(n_3230),
.Y(n_3775)
);

HB1xp67_ASAP7_75t_L g3776 ( 
.A(n_3544),
.Y(n_3776)
);

INVx1_ASAP7_75t_L g3777 ( 
.A(n_3550),
.Y(n_3777)
);

HB1xp67_ASAP7_75t_L g3778 ( 
.A(n_3549),
.Y(n_3778)
);

BUFx3_ASAP7_75t_L g3779 ( 
.A(n_3420),
.Y(n_3779)
);

AND2x2_ASAP7_75t_L g3780 ( 
.A(n_3503),
.B(n_3217),
.Y(n_3780)
);

HB1xp67_ASAP7_75t_L g3781 ( 
.A(n_3628),
.Y(n_3781)
);

AND2x2_ASAP7_75t_L g3782 ( 
.A(n_3400),
.B(n_3231),
.Y(n_3782)
);

NOR2xp33_ASAP7_75t_L g3783 ( 
.A(n_3694),
.B(n_3308),
.Y(n_3783)
);

OR2x2_ASAP7_75t_L g3784 ( 
.A(n_3388),
.B(n_3167),
.Y(n_3784)
);

INVx2_ASAP7_75t_L g3785 ( 
.A(n_3554),
.Y(n_3785)
);

AND2x2_ASAP7_75t_L g3786 ( 
.A(n_3398),
.B(n_3231),
.Y(n_3786)
);

AND2x2_ASAP7_75t_L g3787 ( 
.A(n_3468),
.B(n_3238),
.Y(n_3787)
);

AND2x2_ASAP7_75t_L g3788 ( 
.A(n_3469),
.B(n_3238),
.Y(n_3788)
);

NAND2xp5_ASAP7_75t_L g3789 ( 
.A(n_3565),
.B(n_3168),
.Y(n_3789)
);

BUFx2_ASAP7_75t_L g3790 ( 
.A(n_3657),
.Y(n_3790)
);

INVx1_ASAP7_75t_L g3791 ( 
.A(n_3626),
.Y(n_3791)
);

AND2x2_ASAP7_75t_L g3792 ( 
.A(n_3605),
.B(n_3244),
.Y(n_3792)
);

AND2x2_ASAP7_75t_L g3793 ( 
.A(n_3427),
.B(n_3244),
.Y(n_3793)
);

INVx1_ASAP7_75t_L g3794 ( 
.A(n_3627),
.Y(n_3794)
);

NOR2x1_ASAP7_75t_SL g3795 ( 
.A(n_3392),
.B(n_3068),
.Y(n_3795)
);

NOR4xp25_ASAP7_75t_SL g3796 ( 
.A(n_3697),
.B(n_3394),
.C(n_3428),
.D(n_3693),
.Y(n_3796)
);

INVx1_ASAP7_75t_L g3797 ( 
.A(n_3658),
.Y(n_3797)
);

AND2x2_ASAP7_75t_L g3798 ( 
.A(n_3385),
.B(n_3262),
.Y(n_3798)
);

CKINVDCx20_ASAP7_75t_R g3799 ( 
.A(n_3374),
.Y(n_3799)
);

INVx1_ASAP7_75t_L g3800 ( 
.A(n_3594),
.Y(n_3800)
);

AND2x2_ASAP7_75t_L g3801 ( 
.A(n_3679),
.B(n_3262),
.Y(n_3801)
);

OR2x2_ASAP7_75t_L g3802 ( 
.A(n_3376),
.B(n_3182),
.Y(n_3802)
);

INVx2_ASAP7_75t_L g3803 ( 
.A(n_3371),
.Y(n_3803)
);

BUFx3_ASAP7_75t_L g3804 ( 
.A(n_3485),
.Y(n_3804)
);

INVx2_ASAP7_75t_L g3805 ( 
.A(n_3606),
.Y(n_3805)
);

OR2x2_ASAP7_75t_L g3806 ( 
.A(n_3381),
.B(n_3304),
.Y(n_3806)
);

HB1xp67_ASAP7_75t_L g3807 ( 
.A(n_3622),
.Y(n_3807)
);

HB1xp67_ASAP7_75t_L g3808 ( 
.A(n_3674),
.Y(n_3808)
);

AND2x4_ASAP7_75t_L g3809 ( 
.A(n_3674),
.B(n_3230),
.Y(n_3809)
);

BUFx2_ASAP7_75t_L g3810 ( 
.A(n_3520),
.Y(n_3810)
);

AND2x2_ASAP7_75t_L g3811 ( 
.A(n_3404),
.B(n_3299),
.Y(n_3811)
);

NAND2xp5_ASAP7_75t_L g3812 ( 
.A(n_3566),
.B(n_3235),
.Y(n_3812)
);

OR2x2_ASAP7_75t_L g3813 ( 
.A(n_3372),
.B(n_3313),
.Y(n_3813)
);

INVx2_ASAP7_75t_L g3814 ( 
.A(n_3570),
.Y(n_3814)
);

AND2x4_ASAP7_75t_L g3815 ( 
.A(n_3391),
.B(n_3101),
.Y(n_3815)
);

AND2x2_ASAP7_75t_L g3816 ( 
.A(n_3451),
.B(n_3329),
.Y(n_3816)
);

INVx2_ASAP7_75t_SL g3817 ( 
.A(n_3534),
.Y(n_3817)
);

INVx2_ASAP7_75t_L g3818 ( 
.A(n_3573),
.Y(n_3818)
);

AND2x2_ASAP7_75t_L g3819 ( 
.A(n_3497),
.B(n_3329),
.Y(n_3819)
);

INVx1_ASAP7_75t_L g3820 ( 
.A(n_3521),
.Y(n_3820)
);

INVx1_ASAP7_75t_L g3821 ( 
.A(n_3561),
.Y(n_3821)
);

BUFx2_ASAP7_75t_L g3822 ( 
.A(n_3482),
.Y(n_3822)
);

NAND2xp5_ASAP7_75t_L g3823 ( 
.A(n_3666),
.B(n_3242),
.Y(n_3823)
);

NAND2xp5_ASAP7_75t_L g3824 ( 
.A(n_3578),
.B(n_3145),
.Y(n_3824)
);

AND2x2_ASAP7_75t_L g3825 ( 
.A(n_3590),
.B(n_3336),
.Y(n_3825)
);

HB1xp67_ASAP7_75t_L g3826 ( 
.A(n_3487),
.Y(n_3826)
);

AND2x4_ASAP7_75t_L g3827 ( 
.A(n_3418),
.B(n_3101),
.Y(n_3827)
);

INVx2_ASAP7_75t_L g3828 ( 
.A(n_3683),
.Y(n_3828)
);

NAND2xp33_ASAP7_75t_SL g3829 ( 
.A(n_3450),
.B(n_3075),
.Y(n_3829)
);

AND2x2_ASAP7_75t_L g3830 ( 
.A(n_3552),
.B(n_3316),
.Y(n_3830)
);

BUFx3_ASAP7_75t_L g3831 ( 
.A(n_3660),
.Y(n_3831)
);

AND2x4_ASAP7_75t_L g3832 ( 
.A(n_3418),
.B(n_3122),
.Y(n_3832)
);

AND2x2_ASAP7_75t_L g3833 ( 
.A(n_3597),
.B(n_3318),
.Y(n_3833)
);

INVx1_ASAP7_75t_SL g3834 ( 
.A(n_3563),
.Y(n_3834)
);

NAND2xp5_ASAP7_75t_L g3835 ( 
.A(n_3612),
.B(n_3629),
.Y(n_3835)
);

AOI21xp5_ASAP7_75t_L g3836 ( 
.A1(n_3541),
.A2(n_3013),
.B(n_3088),
.Y(n_3836)
);

INVx1_ASAP7_75t_L g3837 ( 
.A(n_3415),
.Y(n_3837)
);

HB1xp67_ASAP7_75t_L g3838 ( 
.A(n_3615),
.Y(n_3838)
);

HB1xp67_ASAP7_75t_L g3839 ( 
.A(n_3529),
.Y(n_3839)
);

INVx2_ASAP7_75t_L g3840 ( 
.A(n_3686),
.Y(n_3840)
);

INVx1_ASAP7_75t_L g3841 ( 
.A(n_3421),
.Y(n_3841)
);

INVx1_ASAP7_75t_L g3842 ( 
.A(n_3676),
.Y(n_3842)
);

INVx1_ASAP7_75t_L g3843 ( 
.A(n_3488),
.Y(n_3843)
);

AND2x4_ASAP7_75t_L g3844 ( 
.A(n_3419),
.B(n_3122),
.Y(n_3844)
);

AND2x4_ASAP7_75t_L g3845 ( 
.A(n_3419),
.B(n_3555),
.Y(n_3845)
);

HB1xp67_ASAP7_75t_L g3846 ( 
.A(n_3547),
.Y(n_3846)
);

AND2x2_ASAP7_75t_L g3847 ( 
.A(n_3600),
.B(n_3321),
.Y(n_3847)
);

AND2x2_ASAP7_75t_L g3848 ( 
.A(n_3613),
.B(n_3324),
.Y(n_3848)
);

AOI22xp5_ASAP7_75t_L g3849 ( 
.A1(n_3422),
.A2(n_3058),
.B1(n_3110),
.B2(n_3195),
.Y(n_3849)
);

HB1xp67_ASAP7_75t_L g3850 ( 
.A(n_3656),
.Y(n_3850)
);

INVx2_ASAP7_75t_SL g3851 ( 
.A(n_3491),
.Y(n_3851)
);

INVx2_ASAP7_75t_R g3852 ( 
.A(n_3508),
.Y(n_3852)
);

AND2x2_ASAP7_75t_L g3853 ( 
.A(n_3637),
.B(n_3325),
.Y(n_3853)
);

INVx1_ASAP7_75t_L g3854 ( 
.A(n_3500),
.Y(n_3854)
);

INVx2_ASAP7_75t_L g3855 ( 
.A(n_3511),
.Y(n_3855)
);

AND2x2_ASAP7_75t_L g3856 ( 
.A(n_3476),
.B(n_3326),
.Y(n_3856)
);

OR2x2_ASAP7_75t_L g3857 ( 
.A(n_3584),
.B(n_3328),
.Y(n_3857)
);

AND2x2_ASAP7_75t_L g3858 ( 
.A(n_3688),
.B(n_3591),
.Y(n_3858)
);

INVx3_ASAP7_75t_L g3859 ( 
.A(n_3441),
.Y(n_3859)
);

INVx1_ASAP7_75t_L g3860 ( 
.A(n_3670),
.Y(n_3860)
);

NAND2xp5_ASAP7_75t_L g3861 ( 
.A(n_3646),
.B(n_3145),
.Y(n_3861)
);

OR2x2_ASAP7_75t_L g3862 ( 
.A(n_3431),
.B(n_3335),
.Y(n_3862)
);

INVx2_ASAP7_75t_L g3863 ( 
.A(n_3678),
.Y(n_3863)
);

AOI21xp5_ASAP7_75t_L g3864 ( 
.A1(n_3589),
.A2(n_3013),
.B(n_3088),
.Y(n_3864)
);

INVx1_ASAP7_75t_L g3865 ( 
.A(n_3443),
.Y(n_3865)
);

INVx2_ASAP7_75t_L g3866 ( 
.A(n_3691),
.Y(n_3866)
);

INVx2_ASAP7_75t_L g3867 ( 
.A(n_3361),
.Y(n_3867)
);

BUFx3_ASAP7_75t_L g3868 ( 
.A(n_3528),
.Y(n_3868)
);

INVx3_ASAP7_75t_L g3869 ( 
.A(n_3441),
.Y(n_3869)
);

INVxp67_ASAP7_75t_L g3870 ( 
.A(n_3619),
.Y(n_3870)
);

AOI221xp5_ASAP7_75t_L g3871 ( 
.A1(n_3370),
.A2(n_3247),
.B1(n_3283),
.B2(n_3155),
.C(n_3272),
.Y(n_3871)
);

INVx2_ASAP7_75t_L g3872 ( 
.A(n_3361),
.Y(n_3872)
);

BUFx2_ASAP7_75t_L g3873 ( 
.A(n_3471),
.Y(n_3873)
);

AND2x2_ASAP7_75t_L g3874 ( 
.A(n_3375),
.B(n_3339),
.Y(n_3874)
);

INVx2_ASAP7_75t_L g3875 ( 
.A(n_3361),
.Y(n_3875)
);

INVx1_ASAP7_75t_L g3876 ( 
.A(n_3650),
.Y(n_3876)
);

INVx1_ASAP7_75t_L g3877 ( 
.A(n_3663),
.Y(n_3877)
);

INVx3_ASAP7_75t_L g3878 ( 
.A(n_3536),
.Y(n_3878)
);

OR2x2_ASAP7_75t_L g3879 ( 
.A(n_3643),
.B(n_3341),
.Y(n_3879)
);

BUFx3_ASAP7_75t_L g3880 ( 
.A(n_3581),
.Y(n_3880)
);

HB1xp67_ASAP7_75t_L g3881 ( 
.A(n_3639),
.Y(n_3881)
);

HB1xp67_ASAP7_75t_L g3882 ( 
.A(n_3664),
.Y(n_3882)
);

INVx3_ASAP7_75t_L g3883 ( 
.A(n_3536),
.Y(n_3883)
);

OR2x2_ASAP7_75t_L g3884 ( 
.A(n_3665),
.B(n_3344),
.Y(n_3884)
);

INVx3_ASAP7_75t_L g3885 ( 
.A(n_3664),
.Y(n_3885)
);

INVx2_ASAP7_75t_L g3886 ( 
.A(n_3361),
.Y(n_3886)
);

BUFx2_ASAP7_75t_L g3887 ( 
.A(n_3531),
.Y(n_3887)
);

OR2x2_ASAP7_75t_L g3888 ( 
.A(n_3617),
.B(n_3345),
.Y(n_3888)
);

OR2x2_ASAP7_75t_L g3889 ( 
.A(n_3633),
.B(n_3349),
.Y(n_3889)
);

HB1xp67_ASAP7_75t_L g3890 ( 
.A(n_3631),
.Y(n_3890)
);

INVx2_ASAP7_75t_L g3891 ( 
.A(n_3596),
.Y(n_3891)
);

NAND2xp5_ASAP7_75t_L g3892 ( 
.A(n_3477),
.B(n_3155),
.Y(n_3892)
);

OR2x6_ASAP7_75t_L g3893 ( 
.A(n_3567),
.B(n_3075),
.Y(n_3893)
);

INVx2_ASAP7_75t_SL g3894 ( 
.A(n_3581),
.Y(n_3894)
);

INVx2_ASAP7_75t_L g3895 ( 
.A(n_3596),
.Y(n_3895)
);

OAI22xp5_ASAP7_75t_L g3896 ( 
.A1(n_3379),
.A2(n_3298),
.B1(n_3135),
.B2(n_3094),
.Y(n_3896)
);

AND2x4_ASAP7_75t_L g3897 ( 
.A(n_3465),
.B(n_3352),
.Y(n_3897)
);

INVx2_ASAP7_75t_L g3898 ( 
.A(n_3631),
.Y(n_3898)
);

AND2x2_ASAP7_75t_L g3899 ( 
.A(n_3645),
.B(n_3359),
.Y(n_3899)
);

OR2x2_ASAP7_75t_L g3900 ( 
.A(n_3481),
.B(n_3174),
.Y(n_3900)
);

AND2x2_ASAP7_75t_L g3901 ( 
.A(n_3645),
.B(n_3359),
.Y(n_3901)
);

INVx1_ASAP7_75t_L g3902 ( 
.A(n_3661),
.Y(n_3902)
);

AND2x2_ASAP7_75t_L g3903 ( 
.A(n_3504),
.B(n_3346),
.Y(n_3903)
);

INVx1_ASAP7_75t_L g3904 ( 
.A(n_3569),
.Y(n_3904)
);

BUFx2_ASAP7_75t_L g3905 ( 
.A(n_3580),
.Y(n_3905)
);

AND2x2_ASAP7_75t_L g3906 ( 
.A(n_3516),
.B(n_3518),
.Y(n_3906)
);

INVxp67_ASAP7_75t_SL g3907 ( 
.A(n_3543),
.Y(n_3907)
);

AND2x2_ASAP7_75t_L g3908 ( 
.A(n_3524),
.B(n_3360),
.Y(n_3908)
);

INVx2_ASAP7_75t_L g3909 ( 
.A(n_3571),
.Y(n_3909)
);

INVx1_ASAP7_75t_L g3910 ( 
.A(n_3569),
.Y(n_3910)
);

INVx1_ASAP7_75t_L g3911 ( 
.A(n_3569),
.Y(n_3911)
);

OR2x2_ASAP7_75t_L g3912 ( 
.A(n_3484),
.B(n_3174),
.Y(n_3912)
);

OA21x2_ASAP7_75t_L g3913 ( 
.A1(n_3692),
.A2(n_3240),
.B(n_3229),
.Y(n_3913)
);

INVx1_ASAP7_75t_L g3914 ( 
.A(n_3604),
.Y(n_3914)
);

INVx3_ASAP7_75t_L g3915 ( 
.A(n_3567),
.Y(n_3915)
);

BUFx2_ASAP7_75t_L g3916 ( 
.A(n_3580),
.Y(n_3916)
);

OR2x2_ASAP7_75t_L g3917 ( 
.A(n_3362),
.B(n_3057),
.Y(n_3917)
);

NAND2xp5_ASAP7_75t_L g3918 ( 
.A(n_3448),
.B(n_3111),
.Y(n_3918)
);

INVxp67_ASAP7_75t_SL g3919 ( 
.A(n_3669),
.Y(n_3919)
);

OR2x2_ASAP7_75t_SL g3920 ( 
.A(n_3517),
.B(n_3353),
.Y(n_3920)
);

AND2x2_ASAP7_75t_L g3921 ( 
.A(n_3530),
.B(n_2719),
.Y(n_3921)
);

BUFx3_ASAP7_75t_L g3922 ( 
.A(n_3474),
.Y(n_3922)
);

INVx1_ASAP7_75t_L g3923 ( 
.A(n_3604),
.Y(n_3923)
);

OR2x2_ASAP7_75t_L g3924 ( 
.A(n_3551),
.B(n_3057),
.Y(n_3924)
);

OR2x2_ASAP7_75t_L g3925 ( 
.A(n_3728),
.B(n_3457),
.Y(n_3925)
);

AND2x2_ASAP7_75t_L g3926 ( 
.A(n_3826),
.B(n_3729),
.Y(n_3926)
);

INVx2_ASAP7_75t_L g3927 ( 
.A(n_3700),
.Y(n_3927)
);

INVx1_ASAP7_75t_L g3928 ( 
.A(n_3720),
.Y(n_3928)
);

AND2x2_ASAP7_75t_L g3929 ( 
.A(n_3816),
.B(n_3501),
.Y(n_3929)
);

NOR2xp67_ASAP7_75t_L g3930 ( 
.A(n_3915),
.B(n_3583),
.Y(n_3930)
);

AND2x2_ASAP7_75t_L g3931 ( 
.A(n_3858),
.B(n_3587),
.Y(n_3931)
);

AND2x2_ASAP7_75t_L g3932 ( 
.A(n_3742),
.B(n_3449),
.Y(n_3932)
);

INVx1_ASAP7_75t_L g3933 ( 
.A(n_3720),
.Y(n_3933)
);

OR2x2_ASAP7_75t_L g3934 ( 
.A(n_3838),
.B(n_3457),
.Y(n_3934)
);

INVx1_ASAP7_75t_L g3935 ( 
.A(n_3722),
.Y(n_3935)
);

AOI22xp33_ASAP7_75t_L g3936 ( 
.A1(n_3747),
.A2(n_3689),
.B1(n_3478),
.B2(n_3537),
.Y(n_3936)
);

AOI22xp33_ASAP7_75t_L g3937 ( 
.A1(n_3896),
.A2(n_3638),
.B1(n_3644),
.B2(n_3595),
.Y(n_3937)
);

AND2x2_ASAP7_75t_L g3938 ( 
.A(n_3798),
.B(n_3652),
.Y(n_3938)
);

AND2x2_ASAP7_75t_L g3939 ( 
.A(n_3757),
.B(n_3603),
.Y(n_3939)
);

INVx1_ASAP7_75t_L g3940 ( 
.A(n_3722),
.Y(n_3940)
);

OR2x2_ASAP7_75t_L g3941 ( 
.A(n_3714),
.B(n_3457),
.Y(n_3941)
);

NAND2xp5_ASAP7_75t_L g3942 ( 
.A(n_3820),
.B(n_3655),
.Y(n_3942)
);

INVx1_ASAP7_75t_L g3943 ( 
.A(n_3724),
.Y(n_3943)
);

OR2x2_ASAP7_75t_L g3944 ( 
.A(n_3730),
.B(n_3395),
.Y(n_3944)
);

INVx1_ASAP7_75t_L g3945 ( 
.A(n_3724),
.Y(n_3945)
);

AND2x2_ASAP7_75t_L g3946 ( 
.A(n_3833),
.B(n_3649),
.Y(n_3946)
);

HB1xp67_ASAP7_75t_L g3947 ( 
.A(n_3734),
.Y(n_3947)
);

NAND2xp5_ASAP7_75t_L g3948 ( 
.A(n_3820),
.B(n_3585),
.Y(n_3948)
);

INVx2_ASAP7_75t_L g3949 ( 
.A(n_3709),
.Y(n_3949)
);

AND2x2_ASAP7_75t_L g3950 ( 
.A(n_3787),
.B(n_3788),
.Y(n_3950)
);

INVxp67_ASAP7_75t_L g3951 ( 
.A(n_3740),
.Y(n_3951)
);

INVx1_ASAP7_75t_L g3952 ( 
.A(n_3725),
.Y(n_3952)
);

AOI221xp5_ASAP7_75t_L g3953 ( 
.A1(n_3918),
.A2(n_3430),
.B1(n_3576),
.B2(n_3510),
.C(n_3367),
.Y(n_3953)
);

OR2x2_ASAP7_75t_L g3954 ( 
.A(n_3781),
.B(n_3599),
.Y(n_3954)
);

INVx1_ASAP7_75t_L g3955 ( 
.A(n_3725),
.Y(n_3955)
);

INVx1_ASAP7_75t_L g3956 ( 
.A(n_3748),
.Y(n_3956)
);

OR2x2_ASAP7_75t_L g3957 ( 
.A(n_3776),
.B(n_3461),
.Y(n_3957)
);

NAND2xp5_ASAP7_75t_L g3958 ( 
.A(n_3821),
.B(n_3653),
.Y(n_3958)
);

AOI21xp33_ASAP7_75t_L g3959 ( 
.A1(n_3708),
.A2(n_3623),
.B(n_3525),
.Y(n_3959)
);

INVx2_ASAP7_75t_L g3960 ( 
.A(n_3710),
.Y(n_3960)
);

HB1xp67_ASAP7_75t_L g3961 ( 
.A(n_3850),
.Y(n_3961)
);

OR2x2_ASAP7_75t_L g3962 ( 
.A(n_3778),
.B(n_3437),
.Y(n_3962)
);

AND2x2_ASAP7_75t_L g3963 ( 
.A(n_3744),
.B(n_3505),
.Y(n_3963)
);

INVx2_ASAP7_75t_L g3964 ( 
.A(n_3716),
.Y(n_3964)
);

INVx1_ASAP7_75t_L g3965 ( 
.A(n_3748),
.Y(n_3965)
);

OR2x2_ASAP7_75t_L g3966 ( 
.A(n_3752),
.B(n_3735),
.Y(n_3966)
);

OAI21xp5_ASAP7_75t_SL g3967 ( 
.A1(n_3810),
.A2(n_3447),
.B(n_3502),
.Y(n_3967)
);

INVx1_ASAP7_75t_L g3968 ( 
.A(n_3750),
.Y(n_3968)
);

NAND2xp5_ASAP7_75t_L g3969 ( 
.A(n_3821),
.B(n_3433),
.Y(n_3969)
);

OR2x2_ASAP7_75t_L g3970 ( 
.A(n_3917),
.B(n_3546),
.Y(n_3970)
);

AND2x4_ASAP7_75t_L g3971 ( 
.A(n_3795),
.B(n_3640),
.Y(n_3971)
);

INVx2_ASAP7_75t_L g3972 ( 
.A(n_3717),
.Y(n_3972)
);

INVx1_ASAP7_75t_L g3973 ( 
.A(n_3750),
.Y(n_3973)
);

AND2x2_ASAP7_75t_L g3974 ( 
.A(n_3793),
.B(n_3514),
.Y(n_3974)
);

NAND2xp5_ASAP7_75t_L g3975 ( 
.A(n_3797),
.B(n_3703),
.Y(n_3975)
);

NAND2xp5_ASAP7_75t_L g3976 ( 
.A(n_3797),
.B(n_3703),
.Y(n_3976)
);

BUFx2_ASAP7_75t_L g3977 ( 
.A(n_3920),
.Y(n_3977)
);

AND2x4_ASAP7_75t_L g3978 ( 
.A(n_3795),
.B(n_3687),
.Y(n_3978)
);

INVx2_ASAP7_75t_L g3979 ( 
.A(n_3718),
.Y(n_3979)
);

INVx2_ASAP7_75t_L g3980 ( 
.A(n_3723),
.Y(n_3980)
);

AND2x2_ASAP7_75t_SL g3981 ( 
.A(n_3873),
.B(n_3614),
.Y(n_3981)
);

NOR2xp33_ASAP7_75t_L g3982 ( 
.A(n_3894),
.B(n_3399),
.Y(n_3982)
);

AND2x2_ASAP7_75t_L g3983 ( 
.A(n_3712),
.B(n_3575),
.Y(n_3983)
);

INVx1_ASAP7_75t_L g3984 ( 
.A(n_3713),
.Y(n_3984)
);

AND2x2_ASAP7_75t_L g3985 ( 
.A(n_3890),
.B(n_3373),
.Y(n_3985)
);

AND2x2_ASAP7_75t_L g3986 ( 
.A(n_3786),
.B(n_3762),
.Y(n_3986)
);

AND2x2_ASAP7_75t_L g3987 ( 
.A(n_3782),
.B(n_3453),
.Y(n_3987)
);

AND2x4_ASAP7_75t_L g3988 ( 
.A(n_3919),
.B(n_3494),
.Y(n_3988)
);

INVxp67_ASAP7_75t_SL g3989 ( 
.A(n_3807),
.Y(n_3989)
);

HB1xp67_ASAP7_75t_L g3990 ( 
.A(n_3808),
.Y(n_3990)
);

INVx1_ASAP7_75t_L g3991 ( 
.A(n_3713),
.Y(n_3991)
);

INVx1_ASAP7_75t_L g3992 ( 
.A(n_3715),
.Y(n_3992)
);

AND2x2_ASAP7_75t_L g3993 ( 
.A(n_3701),
.B(n_3681),
.Y(n_3993)
);

NOR2xp67_ASAP7_75t_L g3994 ( 
.A(n_3915),
.B(n_3460),
.Y(n_3994)
);

INVx1_ASAP7_75t_L g3995 ( 
.A(n_3715),
.Y(n_3995)
);

NAND2xp5_ASAP7_75t_L g3996 ( 
.A(n_3704),
.B(n_3433),
.Y(n_3996)
);

INVx2_ASAP7_75t_L g3997 ( 
.A(n_3726),
.Y(n_3997)
);

INVx3_ASAP7_75t_L g3998 ( 
.A(n_3775),
.Y(n_3998)
);

NAND2xp5_ASAP7_75t_L g3999 ( 
.A(n_3704),
.B(n_3433),
.Y(n_3999)
);

BUFx3_ASAP7_75t_L g4000 ( 
.A(n_3779),
.Y(n_4000)
);

AND2x2_ASAP7_75t_L g4001 ( 
.A(n_3881),
.B(n_3455),
.Y(n_4001)
);

INVx2_ASAP7_75t_L g4002 ( 
.A(n_3741),
.Y(n_4002)
);

NAND2xp5_ASAP7_75t_SL g4003 ( 
.A(n_3790),
.B(n_3711),
.Y(n_4003)
);

AND2x2_ASAP7_75t_L g4004 ( 
.A(n_3847),
.B(n_3696),
.Y(n_4004)
);

NAND2xp5_ASAP7_75t_L g4005 ( 
.A(n_3705),
.B(n_3493),
.Y(n_4005)
);

NAND2xp5_ASAP7_75t_L g4006 ( 
.A(n_3705),
.B(n_3493),
.Y(n_4006)
);

NAND2xp5_ASAP7_75t_L g4007 ( 
.A(n_3706),
.B(n_3493),
.Y(n_4007)
);

INVx2_ASAP7_75t_L g4008 ( 
.A(n_3749),
.Y(n_4008)
);

INVxp67_ASAP7_75t_SL g4009 ( 
.A(n_3751),
.Y(n_4009)
);

AND2x2_ASAP7_75t_L g4010 ( 
.A(n_3848),
.B(n_3642),
.Y(n_4010)
);

INVx1_ASAP7_75t_L g4011 ( 
.A(n_3733),
.Y(n_4011)
);

INVx1_ASAP7_75t_L g4012 ( 
.A(n_3737),
.Y(n_4012)
);

OR2x2_ASAP7_75t_L g4013 ( 
.A(n_3863),
.B(n_3429),
.Y(n_4013)
);

AND2x2_ASAP7_75t_L g4014 ( 
.A(n_3853),
.B(n_3684),
.Y(n_4014)
);

BUFx2_ASAP7_75t_L g4015 ( 
.A(n_3822),
.Y(n_4015)
);

HB1xp67_ASAP7_75t_SL g4016 ( 
.A(n_3739),
.Y(n_4016)
);

AND2x2_ASAP7_75t_L g4017 ( 
.A(n_3819),
.B(n_3662),
.Y(n_4017)
);

INVx1_ASAP7_75t_L g4018 ( 
.A(n_3738),
.Y(n_4018)
);

INVx1_ASAP7_75t_L g4019 ( 
.A(n_3746),
.Y(n_4019)
);

INVx2_ASAP7_75t_L g4020 ( 
.A(n_3759),
.Y(n_4020)
);

INVx1_ASAP7_75t_L g4021 ( 
.A(n_3753),
.Y(n_4021)
);

AND2x2_ASAP7_75t_L g4022 ( 
.A(n_3811),
.B(n_3662),
.Y(n_4022)
);

INVx2_ASAP7_75t_L g4023 ( 
.A(n_3761),
.Y(n_4023)
);

AND2x2_ASAP7_75t_L g4024 ( 
.A(n_3792),
.B(n_3672),
.Y(n_4024)
);

AND2x4_ASAP7_75t_L g4025 ( 
.A(n_3775),
.B(n_3494),
.Y(n_4025)
);

INVx1_ASAP7_75t_L g4026 ( 
.A(n_3754),
.Y(n_4026)
);

HB1xp67_ASAP7_75t_L g4027 ( 
.A(n_3846),
.Y(n_4027)
);

BUFx2_ASAP7_75t_L g4028 ( 
.A(n_3905),
.Y(n_4028)
);

INVx1_ASAP7_75t_L g4029 ( 
.A(n_3755),
.Y(n_4029)
);

AND2x4_ASAP7_75t_L g4030 ( 
.A(n_3809),
.B(n_3470),
.Y(n_4030)
);

OAI221xp5_ASAP7_75t_SL g4031 ( 
.A1(n_3849),
.A2(n_3766),
.B1(n_3871),
.B2(n_3836),
.C(n_3916),
.Y(n_4031)
);

NAND2xp5_ASAP7_75t_L g4032 ( 
.A(n_3958),
.B(n_3706),
.Y(n_4032)
);

NOR3xp33_ASAP7_75t_L g4033 ( 
.A(n_4031),
.B(n_3727),
.C(n_3490),
.Y(n_4033)
);

AND2x2_ASAP7_75t_L g4034 ( 
.A(n_3950),
.B(n_3882),
.Y(n_4034)
);

INVx1_ASAP7_75t_L g4035 ( 
.A(n_3975),
.Y(n_4035)
);

NAND2xp5_ASAP7_75t_L g4036 ( 
.A(n_3958),
.B(n_3876),
.Y(n_4036)
);

INVx1_ASAP7_75t_L g4037 ( 
.A(n_3975),
.Y(n_4037)
);

INVx2_ASAP7_75t_L g4038 ( 
.A(n_3961),
.Y(n_4038)
);

OR2x2_ASAP7_75t_L g4039 ( 
.A(n_3966),
.B(n_3813),
.Y(n_4039)
);

AND2x2_ASAP7_75t_L g4040 ( 
.A(n_3986),
.B(n_4004),
.Y(n_4040)
);

AND2x2_ASAP7_75t_L g4041 ( 
.A(n_3926),
.B(n_3839),
.Y(n_4041)
);

INVx1_ASAP7_75t_L g4042 ( 
.A(n_3976),
.Y(n_4042)
);

OR2x2_ASAP7_75t_L g4043 ( 
.A(n_3925),
.B(n_3866),
.Y(n_4043)
);

AND2x2_ASAP7_75t_L g4044 ( 
.A(n_4028),
.B(n_3758),
.Y(n_4044)
);

AND2x2_ASAP7_75t_L g4045 ( 
.A(n_4015),
.B(n_3736),
.Y(n_4045)
);

AND2x2_ASAP7_75t_L g4046 ( 
.A(n_4027),
.B(n_3898),
.Y(n_4046)
);

INVx1_ASAP7_75t_L g4047 ( 
.A(n_3976),
.Y(n_4047)
);

AND2x2_ASAP7_75t_L g4048 ( 
.A(n_3938),
.B(n_3947),
.Y(n_4048)
);

INVx1_ASAP7_75t_L g4049 ( 
.A(n_4011),
.Y(n_4049)
);

NOR2x1p5_ASAP7_75t_L g4050 ( 
.A(n_4000),
.B(n_3731),
.Y(n_4050)
);

AND2x2_ASAP7_75t_L g4051 ( 
.A(n_3931),
.B(n_3731),
.Y(n_4051)
);

OR2x2_ASAP7_75t_L g4052 ( 
.A(n_3990),
.B(n_3924),
.Y(n_4052)
);

HB1xp67_ASAP7_75t_L g4053 ( 
.A(n_3989),
.Y(n_4053)
);

NOR2x1_ASAP7_75t_L g4054 ( 
.A(n_3967),
.B(n_3804),
.Y(n_4054)
);

AND2x2_ASAP7_75t_L g4055 ( 
.A(n_4022),
.B(n_3885),
.Y(n_4055)
);

AND2x2_ASAP7_75t_L g4056 ( 
.A(n_3946),
.B(n_3885),
.Y(n_4056)
);

AND2x2_ASAP7_75t_L g4057 ( 
.A(n_3983),
.B(n_3939),
.Y(n_4057)
);

NAND2xp5_ASAP7_75t_L g4058 ( 
.A(n_3969),
.B(n_3877),
.Y(n_4058)
);

AND2x2_ASAP7_75t_L g4059 ( 
.A(n_3985),
.B(n_3857),
.Y(n_4059)
);

INVx1_ASAP7_75t_L g4060 ( 
.A(n_4012),
.Y(n_4060)
);

OR2x2_ASAP7_75t_L g4061 ( 
.A(n_4009),
.B(n_3806),
.Y(n_4061)
);

NAND2xp33_ASAP7_75t_R g4062 ( 
.A(n_3971),
.B(n_3796),
.Y(n_4062)
);

AND2x2_ASAP7_75t_L g4063 ( 
.A(n_3987),
.B(n_3888),
.Y(n_4063)
);

INVx1_ASAP7_75t_L g4064 ( 
.A(n_4018),
.Y(n_4064)
);

AND2x2_ASAP7_75t_L g4065 ( 
.A(n_3998),
.B(n_3809),
.Y(n_4065)
);

AND2x2_ASAP7_75t_L g4066 ( 
.A(n_3998),
.B(n_3899),
.Y(n_4066)
);

INVx1_ASAP7_75t_L g4067 ( 
.A(n_4019),
.Y(n_4067)
);

OR2x2_ASAP7_75t_L g4068 ( 
.A(n_3934),
.B(n_3879),
.Y(n_4068)
);

INVx1_ASAP7_75t_L g4069 ( 
.A(n_4021),
.Y(n_4069)
);

AND2x2_ASAP7_75t_L g4070 ( 
.A(n_3974),
.B(n_3901),
.Y(n_4070)
);

BUFx2_ASAP7_75t_L g4071 ( 
.A(n_3978),
.Y(n_4071)
);

AND2x2_ASAP7_75t_L g4072 ( 
.A(n_4010),
.B(n_3891),
.Y(n_4072)
);

AND2x2_ASAP7_75t_L g4073 ( 
.A(n_4014),
.B(n_3895),
.Y(n_4073)
);

INVx2_ASAP7_75t_L g4074 ( 
.A(n_3927),
.Y(n_4074)
);

INVx1_ASAP7_75t_L g4075 ( 
.A(n_4026),
.Y(n_4075)
);

INVx1_ASAP7_75t_L g4076 ( 
.A(n_4029),
.Y(n_4076)
);

AND2x2_ASAP7_75t_L g4077 ( 
.A(n_4017),
.B(n_3767),
.Y(n_4077)
);

INVx1_ASAP7_75t_L g4078 ( 
.A(n_3928),
.Y(n_4078)
);

NAND2xp5_ASAP7_75t_L g4079 ( 
.A(n_3969),
.B(n_3837),
.Y(n_4079)
);

NAND2xp5_ASAP7_75t_L g4080 ( 
.A(n_3996),
.B(n_3841),
.Y(n_4080)
);

INVx1_ASAP7_75t_L g4081 ( 
.A(n_3933),
.Y(n_4081)
);

NAND2xp5_ASAP7_75t_SL g4082 ( 
.A(n_3981),
.B(n_3845),
.Y(n_4082)
);

NAND2xp5_ASAP7_75t_L g4083 ( 
.A(n_3996),
.B(n_3999),
.Y(n_4083)
);

AND2x2_ASAP7_75t_L g4084 ( 
.A(n_3929),
.B(n_3830),
.Y(n_4084)
);

INVx2_ASAP7_75t_SL g4085 ( 
.A(n_3954),
.Y(n_4085)
);

OR2x2_ASAP7_75t_L g4086 ( 
.A(n_3941),
.B(n_3949),
.Y(n_4086)
);

OR2x2_ASAP7_75t_L g4087 ( 
.A(n_3960),
.B(n_3765),
.Y(n_4087)
);

AND2x4_ASAP7_75t_L g4088 ( 
.A(n_3988),
.B(n_3897),
.Y(n_4088)
);

NOR2xp33_ASAP7_75t_L g4089 ( 
.A(n_3967),
.B(n_3912),
.Y(n_4089)
);

AND2x2_ASAP7_75t_L g4090 ( 
.A(n_3993),
.B(n_3732),
.Y(n_4090)
);

AND2x2_ASAP7_75t_L g4091 ( 
.A(n_3963),
.B(n_3707),
.Y(n_4091)
);

OR2x2_ASAP7_75t_L g4092 ( 
.A(n_3964),
.B(n_3774),
.Y(n_4092)
);

INVx1_ASAP7_75t_L g4093 ( 
.A(n_3935),
.Y(n_4093)
);

INVx1_ASAP7_75t_L g4094 ( 
.A(n_3940),
.Y(n_4094)
);

INVx3_ASAP7_75t_L g4095 ( 
.A(n_3978),
.Y(n_4095)
);

INVx2_ASAP7_75t_L g4096 ( 
.A(n_3972),
.Y(n_4096)
);

INVx1_ASAP7_75t_SL g4097 ( 
.A(n_3944),
.Y(n_4097)
);

HB1xp67_ASAP7_75t_L g4098 ( 
.A(n_3979),
.Y(n_4098)
);

AND2x2_ASAP7_75t_L g4099 ( 
.A(n_4001),
.B(n_3772),
.Y(n_4099)
);

AND2x2_ASAP7_75t_L g4100 ( 
.A(n_3962),
.B(n_3780),
.Y(n_4100)
);

NOR2xp33_ASAP7_75t_SL g4101 ( 
.A(n_3930),
.B(n_3887),
.Y(n_4101)
);

NOR2xp33_ASAP7_75t_L g4102 ( 
.A(n_4031),
.B(n_3870),
.Y(n_4102)
);

INVx1_ASAP7_75t_L g4103 ( 
.A(n_3943),
.Y(n_4103)
);

NAND2xp5_ASAP7_75t_L g4104 ( 
.A(n_3999),
.B(n_3756),
.Y(n_4104)
);

BUFx6f_ASAP7_75t_L g4105 ( 
.A(n_3988),
.Y(n_4105)
);

AND2x4_ASAP7_75t_L g4106 ( 
.A(n_4030),
.B(n_3897),
.Y(n_4106)
);

AND2x2_ASAP7_75t_L g4107 ( 
.A(n_4024),
.B(n_3856),
.Y(n_4107)
);

HB1xp67_ASAP7_75t_L g4108 ( 
.A(n_3980),
.Y(n_4108)
);

OA21x2_ASAP7_75t_L g4109 ( 
.A1(n_3959),
.A2(n_4003),
.B(n_4005),
.Y(n_4109)
);

AND2x2_ASAP7_75t_L g4110 ( 
.A(n_4025),
.B(n_3760),
.Y(n_4110)
);

AND2x2_ASAP7_75t_L g4111 ( 
.A(n_4025),
.B(n_3760),
.Y(n_4111)
);

INVx4_ASAP7_75t_L g4112 ( 
.A(n_3971),
.Y(n_4112)
);

AND2x4_ASAP7_75t_SL g4113 ( 
.A(n_3982),
.B(n_3766),
.Y(n_4113)
);

OR2x2_ASAP7_75t_L g4114 ( 
.A(n_4068),
.B(n_3942),
.Y(n_4114)
);

NAND2xp5_ASAP7_75t_L g4115 ( 
.A(n_4032),
.B(n_3942),
.Y(n_4115)
);

NAND4xp75_ASAP7_75t_L g4116 ( 
.A(n_4054),
.B(n_3930),
.C(n_3953),
.D(n_3994),
.Y(n_4116)
);

INVx1_ASAP7_75t_L g4117 ( 
.A(n_4052),
.Y(n_4117)
);

OR2x2_ASAP7_75t_L g4118 ( 
.A(n_4039),
.B(n_4043),
.Y(n_4118)
);

NAND2xp5_ASAP7_75t_L g4119 ( 
.A(n_4032),
.B(n_4035),
.Y(n_4119)
);

INVx1_ASAP7_75t_L g4120 ( 
.A(n_4037),
.Y(n_4120)
);

AOI22xp5_ASAP7_75t_L g4121 ( 
.A1(n_4033),
.A2(n_3936),
.B1(n_3953),
.B2(n_4102),
.Y(n_4121)
);

OAI22xp5_ASAP7_75t_L g4122 ( 
.A1(n_4050),
.A2(n_3977),
.B1(n_4016),
.B2(n_3994),
.Y(n_4122)
);

OAI22xp5_ASAP7_75t_L g4123 ( 
.A1(n_4089),
.A2(n_3435),
.B1(n_3951),
.B2(n_3937),
.Y(n_4123)
);

OR2x2_ASAP7_75t_L g4124 ( 
.A(n_4092),
.B(n_3948),
.Y(n_4124)
);

AOI21xp33_ASAP7_75t_SL g4125 ( 
.A1(n_4033),
.A2(n_3817),
.B(n_3745),
.Y(n_4125)
);

NAND4xp75_ASAP7_75t_SL g4126 ( 
.A(n_4102),
.B(n_3783),
.C(n_3721),
.D(n_3526),
.Y(n_4126)
);

NAND4xp25_ASAP7_75t_L g4127 ( 
.A(n_4089),
.B(n_3959),
.C(n_3970),
.D(n_3509),
.Y(n_4127)
);

OAI33xp33_ASAP7_75t_L g4128 ( 
.A1(n_4036),
.A2(n_4013),
.A3(n_3957),
.B1(n_3892),
.B2(n_3480),
.B3(n_3475),
.Y(n_4128)
);

INVxp67_ASAP7_75t_SL g4129 ( 
.A(n_4053),
.Y(n_4129)
);

INVx2_ASAP7_75t_L g4130 ( 
.A(n_4098),
.Y(n_4130)
);

NAND2xp5_ASAP7_75t_L g4131 ( 
.A(n_4042),
.B(n_3948),
.Y(n_4131)
);

AND2x2_ASAP7_75t_L g4132 ( 
.A(n_4048),
.B(n_4030),
.Y(n_4132)
);

INVx1_ASAP7_75t_L g4133 ( 
.A(n_4047),
.Y(n_4133)
);

INVx1_ASAP7_75t_L g4134 ( 
.A(n_4053),
.Y(n_4134)
);

NAND2xp5_ASAP7_75t_L g4135 ( 
.A(n_4036),
.B(n_4079),
.Y(n_4135)
);

NAND2xp5_ASAP7_75t_L g4136 ( 
.A(n_4079),
.B(n_3842),
.Y(n_4136)
);

AND2x2_ASAP7_75t_L g4137 ( 
.A(n_4071),
.B(n_3932),
.Y(n_4137)
);

INVx1_ASAP7_75t_L g4138 ( 
.A(n_4104),
.Y(n_4138)
);

AND2x2_ASAP7_75t_L g4139 ( 
.A(n_4099),
.B(n_3997),
.Y(n_4139)
);

INVx1_ASAP7_75t_SL g4140 ( 
.A(n_4097),
.Y(n_4140)
);

INVx1_ASAP7_75t_L g4141 ( 
.A(n_4104),
.Y(n_4141)
);

INVx1_ASAP7_75t_L g4142 ( 
.A(n_4098),
.Y(n_4142)
);

AOI21xp5_ASAP7_75t_L g4143 ( 
.A1(n_4101),
.A2(n_3829),
.B(n_3893),
.Y(n_4143)
);

INVx1_ASAP7_75t_L g4144 ( 
.A(n_4108),
.Y(n_4144)
);

NAND2xp5_ASAP7_75t_L g4145 ( 
.A(n_4080),
.B(n_3865),
.Y(n_4145)
);

INVx1_ASAP7_75t_L g4146 ( 
.A(n_4108),
.Y(n_4146)
);

AOI33xp33_ASAP7_75t_L g4147 ( 
.A1(n_4097),
.A2(n_4045),
.A3(n_4044),
.B1(n_4041),
.B2(n_4085),
.B3(n_4113),
.Y(n_4147)
);

INVx2_ASAP7_75t_L g4148 ( 
.A(n_4086),
.Y(n_4148)
);

NAND2xp33_ASAP7_75t_R g4149 ( 
.A(n_4095),
.B(n_3369),
.Y(n_4149)
);

INVx1_ASAP7_75t_L g4150 ( 
.A(n_4049),
.Y(n_4150)
);

OA222x2_ASAP7_75t_L g4151 ( 
.A1(n_4095),
.A2(n_3893),
.B1(n_3859),
.B2(n_3869),
.C1(n_3883),
.C2(n_3878),
.Y(n_4151)
);

INVx1_ASAP7_75t_L g4152 ( 
.A(n_4060),
.Y(n_4152)
);

OAI211xp5_ASAP7_75t_L g4153 ( 
.A1(n_4082),
.A2(n_3532),
.B(n_3489),
.C(n_3403),
.Y(n_4153)
);

INVx1_ASAP7_75t_L g4154 ( 
.A(n_4064),
.Y(n_4154)
);

NOR2xp33_ASAP7_75t_SL g4155 ( 
.A(n_4112),
.B(n_3834),
.Y(n_4155)
);

AND2x4_ASAP7_75t_L g4156 ( 
.A(n_4112),
.B(n_4088),
.Y(n_4156)
);

INVx1_ASAP7_75t_SL g4157 ( 
.A(n_4087),
.Y(n_4157)
);

INVx2_ASAP7_75t_L g4158 ( 
.A(n_4074),
.Y(n_4158)
);

INVx1_ASAP7_75t_L g4159 ( 
.A(n_4067),
.Y(n_4159)
);

INVx1_ASAP7_75t_L g4160 ( 
.A(n_4069),
.Y(n_4160)
);

INVx1_ASAP7_75t_L g4161 ( 
.A(n_4075),
.Y(n_4161)
);

NOR2x1p5_ASAP7_75t_L g4162 ( 
.A(n_4105),
.B(n_3868),
.Y(n_4162)
);

AND2x2_ASAP7_75t_L g4163 ( 
.A(n_4057),
.B(n_4002),
.Y(n_4163)
);

INVx1_ASAP7_75t_L g4164 ( 
.A(n_4076),
.Y(n_4164)
);

INVx1_ASAP7_75t_L g4165 ( 
.A(n_4080),
.Y(n_4165)
);

INVx2_ASAP7_75t_L g4166 ( 
.A(n_4096),
.Y(n_4166)
);

INVx1_ASAP7_75t_L g4167 ( 
.A(n_4058),
.Y(n_4167)
);

OAI322xp33_ASAP7_75t_L g4168 ( 
.A1(n_4062),
.A2(n_4101),
.A3(n_4083),
.B1(n_4061),
.B2(n_4038),
.C1(n_4058),
.C2(n_3784),
.Y(n_4168)
);

AND2x4_ASAP7_75t_L g4169 ( 
.A(n_4088),
.B(n_3862),
.Y(n_4169)
);

INVx1_ASAP7_75t_L g4170 ( 
.A(n_4078),
.Y(n_4170)
);

INVx1_ASAP7_75t_L g4171 ( 
.A(n_4081),
.Y(n_4171)
);

INVx2_ASAP7_75t_SL g4172 ( 
.A(n_4105),
.Y(n_4172)
);

INVx1_ASAP7_75t_L g4173 ( 
.A(n_4093),
.Y(n_4173)
);

INVx2_ASAP7_75t_SL g4174 ( 
.A(n_4105),
.Y(n_4174)
);

OAI211xp5_ASAP7_75t_L g4175 ( 
.A1(n_4109),
.A2(n_3439),
.B(n_3695),
.C(n_3685),
.Y(n_4175)
);

INVx1_ASAP7_75t_L g4176 ( 
.A(n_4094),
.Y(n_4176)
);

AND2x2_ASAP7_75t_L g4177 ( 
.A(n_4051),
.B(n_4008),
.Y(n_4177)
);

INVx2_ASAP7_75t_SL g4178 ( 
.A(n_4034),
.Y(n_4178)
);

OAI22xp33_ASAP7_75t_L g4179 ( 
.A1(n_4062),
.A2(n_3869),
.B1(n_3878),
.B2(n_3859),
.Y(n_4179)
);

NAND2xp5_ASAP7_75t_L g4180 ( 
.A(n_4083),
.B(n_3945),
.Y(n_4180)
);

INVxp33_ASAP7_75t_L g4181 ( 
.A(n_4046),
.Y(n_4181)
);

OAI22xp5_ASAP7_75t_L g4182 ( 
.A1(n_4040),
.A2(n_3851),
.B1(n_3883),
.B2(n_3799),
.Y(n_4182)
);

AND2x2_ASAP7_75t_L g4183 ( 
.A(n_4070),
.B(n_4020),
.Y(n_4183)
);

INVx1_ASAP7_75t_L g4184 ( 
.A(n_4134),
.Y(n_4184)
);

INVx2_ASAP7_75t_L g4185 ( 
.A(n_4118),
.Y(n_4185)
);

NOR2xp33_ASAP7_75t_L g4186 ( 
.A(n_4155),
.B(n_3560),
.Y(n_4186)
);

OAI22xp33_ASAP7_75t_L g4187 ( 
.A1(n_4125),
.A2(n_4109),
.B1(n_4106),
.B2(n_3864),
.Y(n_4187)
);

OAI22xp5_ASAP7_75t_L g4188 ( 
.A1(n_4125),
.A2(n_4106),
.B1(n_4111),
.B2(n_4110),
.Y(n_4188)
);

INVx1_ASAP7_75t_L g4189 ( 
.A(n_4120),
.Y(n_4189)
);

INVx1_ASAP7_75t_L g4190 ( 
.A(n_4133),
.Y(n_4190)
);

OAI22xp33_ASAP7_75t_L g4191 ( 
.A1(n_4127),
.A2(n_3473),
.B1(n_3630),
.B2(n_3624),
.Y(n_4191)
);

OAI211xp5_ASAP7_75t_L g4192 ( 
.A1(n_4121),
.A2(n_3538),
.B(n_3540),
.C(n_3616),
.Y(n_4192)
);

INVx1_ASAP7_75t_SL g4193 ( 
.A(n_4140),
.Y(n_4193)
);

INVxp33_ASAP7_75t_L g4194 ( 
.A(n_4162),
.Y(n_4194)
);

XOR2xp5_ASAP7_75t_L g4195 ( 
.A(n_4126),
.B(n_3409),
.Y(n_4195)
);

OR2x2_ASAP7_75t_L g4196 ( 
.A(n_4114),
.B(n_4084),
.Y(n_4196)
);

INVx2_ASAP7_75t_L g4197 ( 
.A(n_4130),
.Y(n_4197)
);

OAI221xp5_ASAP7_75t_L g4198 ( 
.A1(n_4121),
.A2(n_3625),
.B1(n_3499),
.B2(n_3495),
.C(n_3401),
.Y(n_4198)
);

INVxp67_ASAP7_75t_L g4199 ( 
.A(n_4149),
.Y(n_4199)
);

AOI22xp5_ASAP7_75t_L g4200 ( 
.A1(n_4123),
.A2(n_3654),
.B1(n_3647),
.B2(n_3906),
.Y(n_4200)
);

AOI21xp33_ASAP7_75t_L g4201 ( 
.A1(n_4175),
.A2(n_3889),
.B(n_3423),
.Y(n_4201)
);

INVx1_ASAP7_75t_L g4202 ( 
.A(n_4119),
.Y(n_4202)
);

AOI221xp5_ASAP7_75t_L g4203 ( 
.A1(n_4168),
.A2(n_4107),
.B1(n_4091),
.B2(n_4100),
.C(n_4090),
.Y(n_4203)
);

INVx1_ASAP7_75t_SL g4204 ( 
.A(n_4157),
.Y(n_4204)
);

INVx1_ASAP7_75t_L g4205 ( 
.A(n_4129),
.Y(n_4205)
);

INVx2_ASAP7_75t_L g4206 ( 
.A(n_4158),
.Y(n_4206)
);

INVx1_ASAP7_75t_L g4207 ( 
.A(n_4180),
.Y(n_4207)
);

NAND2xp5_ASAP7_75t_SL g4208 ( 
.A(n_4147),
.B(n_3586),
.Y(n_4208)
);

INVx1_ASAP7_75t_L g4209 ( 
.A(n_4117),
.Y(n_4209)
);

AOI21xp33_ASAP7_75t_SL g4210 ( 
.A1(n_4122),
.A2(n_3608),
.B(n_3513),
.Y(n_4210)
);

INVxp67_ASAP7_75t_L g4211 ( 
.A(n_4128),
.Y(n_4211)
);

NAND3xp33_ASAP7_75t_SL g4212 ( 
.A(n_4143),
.B(n_3442),
.C(n_3496),
.Y(n_4212)
);

INVx1_ASAP7_75t_L g4213 ( 
.A(n_4138),
.Y(n_4213)
);

NAND2xp5_ASAP7_75t_L g4214 ( 
.A(n_4141),
.B(n_4056),
.Y(n_4214)
);

NAND4xp25_ASAP7_75t_L g4215 ( 
.A(n_4153),
.B(n_3671),
.C(n_3675),
.D(n_3667),
.Y(n_4215)
);

INVx2_ASAP7_75t_SL g4216 ( 
.A(n_4156),
.Y(n_4216)
);

AOI21xp33_ASAP7_75t_L g4217 ( 
.A1(n_4179),
.A2(n_3900),
.B(n_3835),
.Y(n_4217)
);

AOI22xp5_ASAP7_75t_L g4218 ( 
.A1(n_4116),
.A2(n_3854),
.B1(n_3843),
.B2(n_3682),
.Y(n_4218)
);

AOI21xp33_ASAP7_75t_SL g4219 ( 
.A1(n_4182),
.A2(n_3436),
.B(n_3845),
.Y(n_4219)
);

AOI21xp33_ASAP7_75t_SL g4220 ( 
.A1(n_4156),
.A2(n_3389),
.B(n_3636),
.Y(n_4220)
);

OAI21xp5_ASAP7_75t_L g4221 ( 
.A1(n_4181),
.A2(n_3522),
.B(n_3592),
.Y(n_4221)
);

INVx1_ASAP7_75t_L g4222 ( 
.A(n_4167),
.Y(n_4222)
);

NAND2xp5_ASAP7_75t_L g4223 ( 
.A(n_4165),
.B(n_4103),
.Y(n_4223)
);

INVx1_ASAP7_75t_L g4224 ( 
.A(n_4170),
.Y(n_4224)
);

OAI22xp33_ASAP7_75t_L g4225 ( 
.A1(n_4178),
.A2(n_3624),
.B1(n_3907),
.B2(n_3831),
.Y(n_4225)
);

INVx1_ASAP7_75t_L g4226 ( 
.A(n_4171),
.Y(n_4226)
);

INVx2_ASAP7_75t_L g4227 ( 
.A(n_4166),
.Y(n_4227)
);

AOI22xp5_ASAP7_75t_L g4228 ( 
.A1(n_4115),
.A2(n_4059),
.B1(n_4073),
.B2(n_4072),
.Y(n_4228)
);

INVx2_ASAP7_75t_L g4229 ( 
.A(n_4142),
.Y(n_4229)
);

XOR2x2_ASAP7_75t_L g4230 ( 
.A(n_4137),
.B(n_3922),
.Y(n_4230)
);

NAND2xp5_ASAP7_75t_L g4231 ( 
.A(n_4202),
.B(n_4135),
.Y(n_4231)
);

NAND2xp5_ASAP7_75t_L g4232 ( 
.A(n_4207),
.B(n_4131),
.Y(n_4232)
);

AOI21xp33_ASAP7_75t_SL g4233 ( 
.A1(n_4199),
.A2(n_4151),
.B(n_4172),
.Y(n_4233)
);

INVx2_ASAP7_75t_L g4234 ( 
.A(n_4185),
.Y(n_4234)
);

OAI21xp33_ASAP7_75t_SL g4235 ( 
.A1(n_4208),
.A2(n_4151),
.B(n_4132),
.Y(n_4235)
);

OAI21xp5_ASAP7_75t_SL g4236 ( 
.A1(n_4220),
.A2(n_4174),
.B(n_4169),
.Y(n_4236)
);

AND4x1_ASAP7_75t_L g4237 ( 
.A(n_4186),
.B(n_3444),
.C(n_3228),
.D(n_3332),
.Y(n_4237)
);

AND2x2_ASAP7_75t_L g4238 ( 
.A(n_4216),
.B(n_4169),
.Y(n_4238)
);

NOR2xp67_ASAP7_75t_L g4239 ( 
.A(n_4219),
.B(n_4144),
.Y(n_4239)
);

OAI21xp5_ASAP7_75t_L g4240 ( 
.A1(n_4211),
.A2(n_4187),
.B(n_4218),
.Y(n_4240)
);

INVx1_ASAP7_75t_SL g4241 ( 
.A(n_4204),
.Y(n_4241)
);

INVx2_ASAP7_75t_L g4242 ( 
.A(n_4206),
.Y(n_4242)
);

AOI22xp33_ASAP7_75t_L g4243 ( 
.A1(n_4191),
.A2(n_4124),
.B1(n_4065),
.B2(n_4055),
.Y(n_4243)
);

INVx1_ASAP7_75t_L g4244 ( 
.A(n_4223),
.Y(n_4244)
);

NAND2xp5_ASAP7_75t_L g4245 ( 
.A(n_4205),
.B(n_4146),
.Y(n_4245)
);

NAND2xp5_ASAP7_75t_L g4246 ( 
.A(n_4200),
.B(n_4150),
.Y(n_4246)
);

AOI211x1_ASAP7_75t_L g4247 ( 
.A1(n_4192),
.A2(n_4145),
.B(n_4136),
.C(n_4063),
.Y(n_4247)
);

OAI22xp5_ASAP7_75t_L g4248 ( 
.A1(n_4188),
.A2(n_4148),
.B1(n_4163),
.B2(n_4183),
.Y(n_4248)
);

OAI22xp33_ASAP7_75t_L g4249 ( 
.A1(n_4218),
.A2(n_4139),
.B1(n_4177),
.B2(n_4077),
.Y(n_4249)
);

INVx1_ASAP7_75t_L g4250 ( 
.A(n_4189),
.Y(n_4250)
);

AOI22xp5_ASAP7_75t_L g4251 ( 
.A1(n_4200),
.A2(n_4152),
.B1(n_4159),
.B2(n_4154),
.Y(n_4251)
);

NOR3xp33_ASAP7_75t_L g4252 ( 
.A(n_4198),
.B(n_3673),
.C(n_3621),
.Y(n_4252)
);

NAND2xp5_ASAP7_75t_L g4253 ( 
.A(n_4213),
.B(n_4160),
.Y(n_4253)
);

INVx1_ASAP7_75t_L g4254 ( 
.A(n_4190),
.Y(n_4254)
);

INVx1_ASAP7_75t_L g4255 ( 
.A(n_4224),
.Y(n_4255)
);

NAND3xp33_ASAP7_75t_L g4256 ( 
.A(n_4221),
.B(n_4164),
.C(n_4161),
.Y(n_4256)
);

INVx2_ASAP7_75t_L g4257 ( 
.A(n_4227),
.Y(n_4257)
);

OAI32xp33_ASAP7_75t_L g4258 ( 
.A1(n_4194),
.A2(n_4193),
.A3(n_4201),
.B1(n_4196),
.B2(n_4209),
.Y(n_4258)
);

OAI22xp33_ASAP7_75t_SL g4259 ( 
.A1(n_4226),
.A2(n_4173),
.B1(n_4176),
.B2(n_3880),
.Y(n_4259)
);

OAI31xp33_ASAP7_75t_L g4260 ( 
.A1(n_4225),
.A2(n_3593),
.A3(n_4066),
.B(n_3610),
.Y(n_4260)
);

AOI22xp5_ASAP7_75t_L g4261 ( 
.A1(n_4212),
.A2(n_3874),
.B1(n_3909),
.B2(n_3952),
.Y(n_4261)
);

NAND2xp5_ASAP7_75t_L g4262 ( 
.A(n_4222),
.B(n_4203),
.Y(n_4262)
);

INVx1_ASAP7_75t_L g4263 ( 
.A(n_4184),
.Y(n_4263)
);

AOI22xp33_ASAP7_75t_L g4264 ( 
.A1(n_4215),
.A2(n_4217),
.B1(n_4230),
.B2(n_4214),
.Y(n_4264)
);

AOI21xp33_ASAP7_75t_SL g4265 ( 
.A1(n_4195),
.A2(n_3389),
.B(n_3636),
.Y(n_4265)
);

NAND2xp5_ASAP7_75t_L g4266 ( 
.A(n_4228),
.B(n_3955),
.Y(n_4266)
);

OAI21xp33_ASAP7_75t_L g4267 ( 
.A1(n_4210),
.A2(n_4006),
.B(n_4005),
.Y(n_4267)
);

INVx1_ASAP7_75t_L g4268 ( 
.A(n_4229),
.Y(n_4268)
);

OA21x2_ASAP7_75t_L g4269 ( 
.A1(n_4197),
.A2(n_4007),
.B(n_4006),
.Y(n_4269)
);

OAI22xp5_ASAP7_75t_L g4270 ( 
.A1(n_4216),
.A2(n_3177),
.B1(n_3827),
.B2(n_3815),
.Y(n_4270)
);

AOI22xp33_ASAP7_75t_L g4271 ( 
.A1(n_4211),
.A2(n_3852),
.B1(n_3921),
.B2(n_3827),
.Y(n_4271)
);

NAND2xp5_ASAP7_75t_L g4272 ( 
.A(n_4202),
.B(n_3956),
.Y(n_4272)
);

O2A1O1Ixp33_ASAP7_75t_L g4273 ( 
.A1(n_4211),
.A2(n_3659),
.B(n_3311),
.C(n_3559),
.Y(n_4273)
);

AOI22xp5_ASAP7_75t_L g4274 ( 
.A1(n_4211),
.A2(n_3968),
.B1(n_3973),
.B2(n_3965),
.Y(n_4274)
);

NAND2xp5_ASAP7_75t_L g4275 ( 
.A(n_4202),
.B(n_3984),
.Y(n_4275)
);

OAI32xp33_ASAP7_75t_L g4276 ( 
.A1(n_4211),
.A2(n_3802),
.A3(n_3479),
.B1(n_3992),
.B2(n_3991),
.Y(n_4276)
);

OR2x2_ASAP7_75t_L g4277 ( 
.A(n_4202),
.B(n_4007),
.Y(n_4277)
);

AND2x2_ASAP7_75t_L g4278 ( 
.A(n_4216),
.B(n_3825),
.Y(n_4278)
);

NAND2xp5_ASAP7_75t_L g4279 ( 
.A(n_4202),
.B(n_3995),
.Y(n_4279)
);

INVx1_ASAP7_75t_L g4280 ( 
.A(n_4185),
.Y(n_4280)
);

INVx2_ASAP7_75t_L g4281 ( 
.A(n_4185),
.Y(n_4281)
);

OR2x2_ASAP7_75t_L g4282 ( 
.A(n_4277),
.B(n_4023),
.Y(n_4282)
);

AOI21xp5_ASAP7_75t_L g4283 ( 
.A1(n_4235),
.A2(n_3562),
.B(n_3445),
.Y(n_4283)
);

NOR2xp33_ASAP7_75t_L g4284 ( 
.A(n_4241),
.B(n_3719),
.Y(n_4284)
);

OAI21xp33_ASAP7_75t_L g4285 ( 
.A1(n_4240),
.A2(n_4264),
.B(n_4233),
.Y(n_4285)
);

NAND2xp5_ASAP7_75t_SL g4286 ( 
.A(n_4265),
.B(n_3771),
.Y(n_4286)
);

OAI21xp33_ASAP7_75t_L g4287 ( 
.A1(n_4262),
.A2(n_3512),
.B(n_3861),
.Y(n_4287)
);

NOR2xp33_ASAP7_75t_L g4288 ( 
.A(n_4236),
.B(n_3425),
.Y(n_4288)
);

OAI322xp33_ASAP7_75t_L g4289 ( 
.A1(n_4251),
.A2(n_3769),
.A3(n_3770),
.B1(n_3773),
.B2(n_3777),
.C1(n_3823),
.C2(n_3824),
.Y(n_4289)
);

NAND2xp5_ASAP7_75t_L g4290 ( 
.A(n_4244),
.B(n_3855),
.Y(n_4290)
);

NOR2x1_ASAP7_75t_L g4291 ( 
.A(n_4239),
.B(n_3434),
.Y(n_4291)
);

OAI21xp5_ASAP7_75t_SL g4292 ( 
.A1(n_4260),
.A2(n_3568),
.B(n_3323),
.Y(n_4292)
);

AND2x2_ASAP7_75t_L g4293 ( 
.A(n_4239),
.B(n_3815),
.Y(n_4293)
);

NAND3xp33_ASAP7_75t_SL g4294 ( 
.A(n_4273),
.B(n_3355),
.C(n_3545),
.Y(n_4294)
);

INVx2_ASAP7_75t_SL g4295 ( 
.A(n_4238),
.Y(n_4295)
);

NOR2xp33_ASAP7_75t_L g4296 ( 
.A(n_4258),
.B(n_3535),
.Y(n_4296)
);

NAND2xp33_ASAP7_75t_L g4297 ( 
.A(n_4267),
.B(n_3407),
.Y(n_4297)
);

NAND2xp5_ASAP7_75t_SL g4298 ( 
.A(n_4259),
.B(n_3771),
.Y(n_4298)
);

OAI211xp5_ASAP7_75t_SL g4299 ( 
.A1(n_4271),
.A2(n_3082),
.B(n_3125),
.C(n_3601),
.Y(n_4299)
);

INVx2_ASAP7_75t_L g4300 ( 
.A(n_4234),
.Y(n_4300)
);

NOR2xp33_ASAP7_75t_L g4301 ( 
.A(n_4246),
.B(n_3574),
.Y(n_4301)
);

INVx3_ASAP7_75t_L g4302 ( 
.A(n_4269),
.Y(n_4302)
);

AND2x2_ASAP7_75t_L g4303 ( 
.A(n_4281),
.B(n_3832),
.Y(n_4303)
);

INVx2_ASAP7_75t_L g4304 ( 
.A(n_4242),
.Y(n_4304)
);

NAND3xp33_ASAP7_75t_SL g4305 ( 
.A(n_4237),
.B(n_3355),
.C(n_3200),
.Y(n_4305)
);

NAND2xp5_ASAP7_75t_L g4306 ( 
.A(n_4274),
.B(n_3801),
.Y(n_4306)
);

NAND2xp5_ASAP7_75t_L g4307 ( 
.A(n_4247),
.B(n_3828),
.Y(n_4307)
);

INVx1_ASAP7_75t_L g4308 ( 
.A(n_4253),
.Y(n_4308)
);

INVx2_ASAP7_75t_SL g4309 ( 
.A(n_4278),
.Y(n_4309)
);

AOI221xp5_ASAP7_75t_L g4310 ( 
.A1(n_4276),
.A2(n_3789),
.B1(n_3743),
.B2(n_3812),
.C(n_3063),
.Y(n_4310)
);

NOR3x1_ASAP7_75t_L g4311 ( 
.A(n_4256),
.B(n_3454),
.C(n_3078),
.Y(n_4311)
);

INVx1_ASAP7_75t_L g4312 ( 
.A(n_4272),
.Y(n_4312)
);

NOR2x1_ASAP7_75t_SL g4313 ( 
.A(n_4270),
.B(n_3434),
.Y(n_4313)
);

OAI322xp33_ASAP7_75t_L g4314 ( 
.A1(n_4249),
.A2(n_4248),
.A3(n_4245),
.B1(n_4261),
.B2(n_4280),
.C1(n_4266),
.C2(n_4232),
.Y(n_4314)
);

NAND2xp5_ASAP7_75t_L g4315 ( 
.A(n_4231),
.B(n_3840),
.Y(n_4315)
);

NAND3xp33_ASAP7_75t_L g4316 ( 
.A(n_4285),
.B(n_4237),
.C(n_4243),
.Y(n_4316)
);

AOI221xp5_ASAP7_75t_L g4317 ( 
.A1(n_4285),
.A2(n_4254),
.B1(n_4255),
.B2(n_4250),
.C(n_4263),
.Y(n_4317)
);

OR2x2_ASAP7_75t_L g4318 ( 
.A(n_4312),
.B(n_4275),
.Y(n_4318)
);

INVx1_ASAP7_75t_L g4319 ( 
.A(n_4315),
.Y(n_4319)
);

NAND2xp5_ASAP7_75t_L g4320 ( 
.A(n_4287),
.B(n_4268),
.Y(n_4320)
);

NAND2xp5_ASAP7_75t_L g4321 ( 
.A(n_4308),
.B(n_4257),
.Y(n_4321)
);

NOR3x1_ASAP7_75t_L g4322 ( 
.A(n_4305),
.B(n_4279),
.C(n_4252),
.Y(n_4322)
);

AOI21xp5_ASAP7_75t_SL g4323 ( 
.A1(n_4283),
.A2(n_3445),
.B(n_3556),
.Y(n_4323)
);

AND2x2_ASAP7_75t_L g4324 ( 
.A(n_4288),
.B(n_4269),
.Y(n_4324)
);

NAND2xp5_ASAP7_75t_L g4325 ( 
.A(n_4295),
.B(n_3814),
.Y(n_4325)
);

OAI21xp5_ASAP7_75t_L g4326 ( 
.A1(n_4294),
.A2(n_3632),
.B(n_3305),
.Y(n_4326)
);

OA22x2_ASAP7_75t_L g4327 ( 
.A1(n_4309),
.A2(n_3556),
.B1(n_3698),
.B2(n_3832),
.Y(n_4327)
);

OAI21xp33_ASAP7_75t_L g4328 ( 
.A1(n_4296),
.A2(n_3884),
.B(n_3903),
.Y(n_4328)
);

AOI21xp5_ASAP7_75t_L g4329 ( 
.A1(n_4291),
.A2(n_4286),
.B(n_4284),
.Y(n_4329)
);

INVx1_ASAP7_75t_L g4330 ( 
.A(n_4290),
.Y(n_4330)
);

NOR4xp25_ASAP7_75t_L g4331 ( 
.A(n_4314),
.B(n_3275),
.C(n_3111),
.D(n_3169),
.Y(n_4331)
);

AOI211x1_ASAP7_75t_L g4332 ( 
.A1(n_4307),
.A2(n_3268),
.B(n_3282),
.C(n_3588),
.Y(n_4332)
);

AOI211x1_ASAP7_75t_L g4333 ( 
.A1(n_4293),
.A2(n_4298),
.B(n_4306),
.C(n_4303),
.Y(n_4333)
);

NOR3xp33_ASAP7_75t_L g4334 ( 
.A(n_4292),
.B(n_3284),
.C(n_3564),
.Y(n_4334)
);

AOI22xp5_ASAP7_75t_L g4335 ( 
.A1(n_4301),
.A2(n_3844),
.B1(n_3908),
.B2(n_3818),
.Y(n_4335)
);

OAI21xp5_ASAP7_75t_SL g4336 ( 
.A1(n_4310),
.A2(n_3463),
.B(n_3844),
.Y(n_4336)
);

INVx1_ASAP7_75t_L g4337 ( 
.A(n_4300),
.Y(n_4337)
);

HB1xp67_ASAP7_75t_L g4338 ( 
.A(n_4304),
.Y(n_4338)
);

AOI22xp5_ASAP7_75t_L g4339 ( 
.A1(n_4299),
.A2(n_3118),
.B1(n_3690),
.B2(n_2873),
.Y(n_4339)
);

OA22x2_ASAP7_75t_L g4340 ( 
.A1(n_4302),
.A2(n_4313),
.B1(n_4311),
.B2(n_4297),
.Y(n_4340)
);

INVx1_ASAP7_75t_L g4341 ( 
.A(n_4289),
.Y(n_4341)
);

OAI21xp5_ASAP7_75t_SL g4342 ( 
.A1(n_4302),
.A2(n_3124),
.B(n_3041),
.Y(n_4342)
);

INVx1_ASAP7_75t_L g4343 ( 
.A(n_4338),
.Y(n_4343)
);

OAI21xp33_ASAP7_75t_L g4344 ( 
.A1(n_4316),
.A2(n_4282),
.B(n_3800),
.Y(n_4344)
);

AOI211xp5_ASAP7_75t_SL g4345 ( 
.A1(n_4323),
.A2(n_4329),
.B(n_4317),
.C(n_4341),
.Y(n_4345)
);

NOR3xp33_ASAP7_75t_L g4346 ( 
.A(n_4334),
.B(n_2827),
.C(n_2837),
.Y(n_4346)
);

NOR3xp33_ASAP7_75t_SL g4347 ( 
.A(n_4342),
.B(n_649),
.C(n_650),
.Y(n_4347)
);

OAI211xp5_ASAP7_75t_L g4348 ( 
.A1(n_4331),
.A2(n_3582),
.B(n_3542),
.C(n_3424),
.Y(n_4348)
);

NOR2xp33_ASAP7_75t_L g4349 ( 
.A(n_4318),
.B(n_649),
.Y(n_4349)
);

OAI21xp33_ASAP7_75t_SL g4350 ( 
.A1(n_4340),
.A2(n_3620),
.B(n_3333),
.Y(n_4350)
);

AOI22xp5_ASAP7_75t_L g4351 ( 
.A1(n_4336),
.A2(n_3041),
.B1(n_3690),
.B2(n_3007),
.Y(n_4351)
);

AOI221xp5_ASAP7_75t_L g4352 ( 
.A1(n_4333),
.A2(n_3800),
.B1(n_3914),
.B2(n_3923),
.C(n_3702),
.Y(n_4352)
);

NOR3xp33_ASAP7_75t_L g4353 ( 
.A(n_4337),
.B(n_2747),
.C(n_2635),
.Y(n_4353)
);

O2A1O1Ixp33_ASAP7_75t_L g4354 ( 
.A1(n_4320),
.A2(n_2997),
.B(n_3028),
.C(n_2994),
.Y(n_4354)
);

NAND3xp33_ASAP7_75t_SL g4355 ( 
.A(n_4339),
.B(n_2997),
.C(n_2994),
.Y(n_4355)
);

OAI211xp5_ASAP7_75t_L g4356 ( 
.A1(n_4339),
.A2(n_3424),
.B(n_3462),
.C(n_3452),
.Y(n_4356)
);

NAND4xp75_ASAP7_75t_L g4357 ( 
.A(n_4322),
.B(n_4324),
.C(n_4332),
.D(n_4326),
.Y(n_4357)
);

AOI221xp5_ASAP7_75t_L g4358 ( 
.A1(n_4330),
.A2(n_3923),
.B1(n_3914),
.B2(n_3702),
.C(n_3910),
.Y(n_4358)
);

OAI21xp5_ASAP7_75t_SL g4359 ( 
.A1(n_4321),
.A2(n_3173),
.B(n_3133),
.Y(n_4359)
);

OAI322xp33_ASAP7_75t_L g4360 ( 
.A1(n_4319),
.A2(n_3028),
.A3(n_3089),
.B1(n_3904),
.B2(n_3910),
.C1(n_3911),
.C2(n_3805),
.Y(n_4360)
);

XNOR2x1_ASAP7_75t_L g4361 ( 
.A(n_4327),
.B(n_4335),
.Y(n_4361)
);

AOI21xp5_ASAP7_75t_L g4362 ( 
.A1(n_4325),
.A2(n_3579),
.B(n_2846),
.Y(n_4362)
);

XNOR2xp5_ASAP7_75t_L g4363 ( 
.A(n_4328),
.B(n_650),
.Y(n_4363)
);

OAI211xp5_ASAP7_75t_SL g4364 ( 
.A1(n_4317),
.A2(n_653),
.B(n_651),
.C(n_652),
.Y(n_4364)
);

NOR4xp25_ASAP7_75t_L g4365 ( 
.A(n_4316),
.B(n_3911),
.C(n_3904),
.D(n_653),
.Y(n_4365)
);

AOI211xp5_ASAP7_75t_L g4366 ( 
.A1(n_4331),
.A2(n_3462),
.B(n_3483),
.C(n_3452),
.Y(n_4366)
);

OR2x2_ASAP7_75t_L g4367 ( 
.A(n_4343),
.B(n_651),
.Y(n_4367)
);

INVx1_ASAP7_75t_L g4368 ( 
.A(n_4344),
.Y(n_4368)
);

NOR2xp33_ASAP7_75t_SL g4369 ( 
.A(n_4349),
.B(n_3483),
.Y(n_4369)
);

INVxp67_ASAP7_75t_SL g4370 ( 
.A(n_4366),
.Y(n_4370)
);

NOR2x1_ASAP7_75t_SL g4371 ( 
.A(n_4357),
.B(n_3771),
.Y(n_4371)
);

INVx2_ASAP7_75t_L g4372 ( 
.A(n_4363),
.Y(n_4372)
);

INVx1_ASAP7_75t_L g4373 ( 
.A(n_4352),
.Y(n_4373)
);

INVx1_ASAP7_75t_L g4374 ( 
.A(n_4355),
.Y(n_4374)
);

OAI22xp33_ASAP7_75t_L g4375 ( 
.A1(n_4345),
.A2(n_3133),
.B1(n_3173),
.B2(n_3089),
.Y(n_4375)
);

AO22x2_ASAP7_75t_L g4376 ( 
.A1(n_4361),
.A2(n_3007),
.B1(n_3872),
.B2(n_3867),
.Y(n_4376)
);

AO22x1_ASAP7_75t_L g4377 ( 
.A1(n_4365),
.A2(n_3886),
.B1(n_3875),
.B2(n_3340),
.Y(n_4377)
);

NOR2x1_ASAP7_75t_L g4378 ( 
.A(n_4364),
.B(n_4356),
.Y(n_4378)
);

NOR4xp25_ASAP7_75t_L g4379 ( 
.A(n_4350),
.B(n_656),
.C(n_652),
.D(n_655),
.Y(n_4379)
);

NOR2x1_ASAP7_75t_L g4380 ( 
.A(n_4348),
.B(n_2735),
.Y(n_4380)
);

NAND2xp5_ASAP7_75t_L g4381 ( 
.A(n_4347),
.B(n_657),
.Y(n_4381)
);

INVx1_ASAP7_75t_L g4382 ( 
.A(n_4360),
.Y(n_4382)
);

AND2x4_ASAP7_75t_L g4383 ( 
.A(n_4372),
.B(n_4351),
.Y(n_4383)
);

NOR3xp33_ASAP7_75t_SL g4384 ( 
.A(n_4370),
.B(n_4374),
.C(n_4382),
.Y(n_4384)
);

INVx1_ASAP7_75t_L g4385 ( 
.A(n_4367),
.Y(n_4385)
);

INVx4_ASAP7_75t_L g4386 ( 
.A(n_4376),
.Y(n_4386)
);

OR2x2_ASAP7_75t_L g4387 ( 
.A(n_4368),
.B(n_4359),
.Y(n_4387)
);

INVx1_ASAP7_75t_SL g4388 ( 
.A(n_4381),
.Y(n_4388)
);

NAND2xp5_ASAP7_75t_L g4389 ( 
.A(n_4377),
.B(n_4358),
.Y(n_4389)
);

AND2x2_ASAP7_75t_L g4390 ( 
.A(n_4371),
.B(n_4376),
.Y(n_4390)
);

AOI21xp5_ASAP7_75t_L g4391 ( 
.A1(n_4379),
.A2(n_4354),
.B(n_4362),
.Y(n_4391)
);

NAND3xp33_ASAP7_75t_SL g4392 ( 
.A(n_4369),
.B(n_4346),
.C(n_4353),
.Y(n_4392)
);

NOR3x2_ASAP7_75t_L g4393 ( 
.A(n_4378),
.B(n_657),
.C(n_658),
.Y(n_4393)
);

AOI221xp5_ASAP7_75t_L g4394 ( 
.A1(n_4373),
.A2(n_2735),
.B1(n_3763),
.B2(n_3803),
.C(n_3764),
.Y(n_4394)
);

NOR2xp67_ASAP7_75t_L g4395 ( 
.A(n_4380),
.B(n_659),
.Y(n_4395)
);

CKINVDCx5p33_ASAP7_75t_R g4396 ( 
.A(n_4375),
.Y(n_4396)
);

OAI22xp33_ASAP7_75t_L g4397 ( 
.A1(n_4396),
.A2(n_3913),
.B1(n_3768),
.B2(n_3785),
.Y(n_4397)
);

AOI322xp5_ASAP7_75t_L g4398 ( 
.A1(n_4384),
.A2(n_3794),
.A3(n_3791),
.B1(n_3902),
.B2(n_3860),
.C1(n_3245),
.C2(n_3280),
.Y(n_4398)
);

NOR2x1_ASAP7_75t_L g4399 ( 
.A(n_4395),
.B(n_659),
.Y(n_4399)
);

AOI221x1_ASAP7_75t_L g4400 ( 
.A1(n_4385),
.A2(n_660),
.B1(n_662),
.B2(n_663),
.C(n_665),
.Y(n_4400)
);

CKINVDCx5p33_ASAP7_75t_R g4401 ( 
.A(n_4388),
.Y(n_4401)
);

INVx1_ASAP7_75t_L g4402 ( 
.A(n_4393),
.Y(n_4402)
);

INVx2_ASAP7_75t_L g4403 ( 
.A(n_4387),
.Y(n_4403)
);

INVx1_ASAP7_75t_L g4404 ( 
.A(n_4403),
.Y(n_4404)
);

NAND2xp5_ASAP7_75t_L g4405 ( 
.A(n_4400),
.B(n_4386),
.Y(n_4405)
);

XNOR2xp5_ASAP7_75t_L g4406 ( 
.A(n_4401),
.B(n_4383),
.Y(n_4406)
);

INVx2_ASAP7_75t_L g4407 ( 
.A(n_4402),
.Y(n_4407)
);

INVx2_ASAP7_75t_L g4408 ( 
.A(n_4399),
.Y(n_4408)
);

OAI31xp33_ASAP7_75t_L g4409 ( 
.A1(n_4406),
.A2(n_4390),
.A3(n_4397),
.B(n_4391),
.Y(n_4409)
);

OAI22xp33_ASAP7_75t_L g4410 ( 
.A1(n_4404),
.A2(n_4389),
.B1(n_4392),
.B2(n_4394),
.Y(n_4410)
);

INVx2_ASAP7_75t_L g4411 ( 
.A(n_4409),
.Y(n_4411)
);

AOI22x1_ASAP7_75t_SL g4412 ( 
.A1(n_4410),
.A2(n_4407),
.B1(n_4408),
.B2(n_4405),
.Y(n_4412)
);

AOI222xp33_ASAP7_75t_L g4413 ( 
.A1(n_4411),
.A2(n_4398),
.B1(n_2616),
.B2(n_3227),
.C1(n_3340),
.C2(n_2862),
.Y(n_4413)
);

BUFx12f_ASAP7_75t_L g4414 ( 
.A(n_4412),
.Y(n_4414)
);

XNOR2xp5_ASAP7_75t_L g4415 ( 
.A(n_4414),
.B(n_660),
.Y(n_4415)
);

OAI21xp5_ASAP7_75t_L g4416 ( 
.A1(n_4413),
.A2(n_3138),
.B(n_3043),
.Y(n_4416)
);

AOI22xp33_ASAP7_75t_L g4417 ( 
.A1(n_4415),
.A2(n_3256),
.B1(n_3913),
.B2(n_3119),
.Y(n_4417)
);

OR2x6_ASAP7_75t_L g4418 ( 
.A(n_4417),
.B(n_4416),
.Y(n_4418)
);

AOI22xp33_ASAP7_75t_SL g4419 ( 
.A1(n_4418),
.A2(n_3340),
.B1(n_3227),
.B2(n_2865),
.Y(n_4419)
);


endmodule