module fake_aes_8268_n_47 (n_11, n_1, n_2, n_13, n_12, n_6, n_4, n_3, n_9, n_5, n_14, n_7, n_10, n_8, n_0, n_47);
input n_11;
input n_1;
input n_2;
input n_13;
input n_12;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_14;
input n_7;
input n_10;
input n_8;
input n_0;
output n_47;
wire n_45;
wire n_20;
wire n_38;
wire n_44;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_46;
wire n_25;
wire n_30;
wire n_26;
wire n_33;
wire n_16;
wire n_18;
wire n_32;
wire n_41;
wire n_35;
wire n_17;
wire n_15;
wire n_42;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_43;
wire n_40;
wire n_29;
wire n_39;
NOR2xp33_ASAP7_75t_L g15 ( .A(n_5), .B(n_13), .Y(n_15) );
NOR2xp33_ASAP7_75t_R g16 ( .A(n_2), .B(n_4), .Y(n_16) );
XNOR2xp5_ASAP7_75t_L g17 ( .A(n_14), .B(n_11), .Y(n_17) );
AND2x4_ASAP7_75t_L g18 ( .A(n_1), .B(n_7), .Y(n_18) );
AND2x4_ASAP7_75t_L g19 ( .A(n_8), .B(n_10), .Y(n_19) );
AND2x2_ASAP7_75t_SL g20 ( .A(n_6), .B(n_9), .Y(n_20) );
NAND2xp5_ASAP7_75t_SL g21 ( .A(n_4), .B(n_5), .Y(n_21) );
BUFx2_ASAP7_75t_L g22 ( .A(n_0), .Y(n_22) );
NOR2xp33_ASAP7_75t_L g23 ( .A(n_22), .B(n_0), .Y(n_23) );
BUFx3_ASAP7_75t_L g24 ( .A(n_19), .Y(n_24) );
INVx2_ASAP7_75t_SL g25 ( .A(n_18), .Y(n_25) );
AOI22xp5_ASAP7_75t_L g26 ( .A1(n_18), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_26) );
O2A1O1Ixp33_ASAP7_75t_L g27 ( .A1(n_23), .A2(n_21), .B(n_15), .C(n_19), .Y(n_27) );
BUFx12f_ASAP7_75t_L g28 ( .A(n_25), .Y(n_28) );
INVx2_ASAP7_75t_L g29 ( .A(n_24), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_29), .B(n_23), .Y(n_30) );
INVxp67_ASAP7_75t_SL g31 ( .A(n_28), .Y(n_31) );
NAND2xp5_ASAP7_75t_L g32 ( .A(n_30), .B(n_27), .Y(n_32) );
AND2x2_ASAP7_75t_L g33 ( .A(n_30), .B(n_26), .Y(n_33) );
AND2x4_ASAP7_75t_L g34 ( .A(n_32), .B(n_31), .Y(n_34) );
AND2x2_ASAP7_75t_L g35 ( .A(n_33), .B(n_31), .Y(n_35) );
INVx1_ASAP7_75t_L g36 ( .A(n_32), .Y(n_36) );
BUFx3_ASAP7_75t_L g37 ( .A(n_34), .Y(n_37) );
AOI31xp33_ASAP7_75t_SL g38 ( .A1(n_35), .A2(n_17), .A3(n_15), .B(n_16), .Y(n_38) );
AOI21xp33_ASAP7_75t_L g39 ( .A1(n_36), .A2(n_27), .B(n_20), .Y(n_39) );
NOR3xp33_ASAP7_75t_L g40 ( .A(n_39), .B(n_35), .C(n_34), .Y(n_40) );
AND2x4_ASAP7_75t_L g41 ( .A(n_37), .B(n_34), .Y(n_41) );
NAND3xp33_ASAP7_75t_L g42 ( .A(n_37), .B(n_20), .C(n_34), .Y(n_42) );
NOR2xp33_ASAP7_75t_L g43 ( .A(n_42), .B(n_36), .Y(n_43) );
INVx1_ASAP7_75t_L g44 ( .A(n_41), .Y(n_44) );
AOI22xp5_ASAP7_75t_L g45 ( .A1(n_40), .A2(n_38), .B1(n_16), .B2(n_3), .Y(n_45) );
INVx1_ASAP7_75t_L g46 ( .A(n_44), .Y(n_46) );
OAI22xp33_ASAP7_75t_L g47 ( .A1(n_46), .A2(n_45), .B1(n_43), .B2(n_12), .Y(n_47) );
endmodule