module fake_jpeg_22652_n_340 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_340);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_340;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_7),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

CKINVDCx11_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_5),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_5),
.Y(n_28)
);

CKINVDCx20_ASAP7_75t_R g29 ( 
.A(n_16),
.Y(n_29)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

BUFx3_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_15),
.Y(n_33)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_3),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_13),
.Y(n_36)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_28),
.Y(n_37)
);

INVx5_ASAP7_75t_L g57 ( 
.A(n_37),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_31),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_38),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

BUFx4f_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g42 ( 
.A(n_21),
.Y(n_42)
);

BUFx3_ASAP7_75t_L g58 ( 
.A(n_42),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_24),
.B(n_0),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_43),
.B(n_48),
.Y(n_59)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

INVx2_ASAP7_75t_L g65 ( 
.A(n_45),
.Y(n_65)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_SL g49 ( 
.A1(n_46),
.A2(n_28),
.B1(n_47),
.B2(n_30),
.Y(n_49)
);

BUFx5_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_29),
.B(n_19),
.Y(n_48)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_49),
.A2(n_27),
.B1(n_24),
.B2(n_25),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g50 ( 
.A1(n_46),
.A2(n_37),
.B1(n_44),
.B2(n_42),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g66 ( 
.A1(n_50),
.A2(n_42),
.B1(n_30),
.B2(n_40),
.Y(n_66)
);

AND2x2_ASAP7_75t_L g53 ( 
.A(n_40),
.B(n_0),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_53),
.B(n_21),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_43),
.B(n_33),
.Y(n_61)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_61),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_33),
.Y(n_63)
);

OR2x2_ASAP7_75t_L g77 ( 
.A(n_63),
.B(n_29),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_47),
.A2(n_28),
.B1(n_30),
.B2(n_17),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g70 ( 
.A1(n_64),
.A2(n_17),
.B1(n_27),
.B2(n_24),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_66),
.A2(n_70),
.B1(n_76),
.B2(n_81),
.Y(n_124)
);

OAI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_57),
.A2(n_40),
.B1(n_17),
.B2(n_19),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g110 ( 
.A1(n_67),
.A2(n_72),
.B1(n_89),
.B2(n_92),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_63),
.Y(n_68)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_68),
.Y(n_121)
);

OAI22xp33_ASAP7_75t_L g69 ( 
.A1(n_51),
.A2(n_40),
.B1(n_41),
.B2(n_45),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_69),
.A2(n_84),
.B1(n_65),
.B2(n_55),
.Y(n_113)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_71),
.B(n_59),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_58),
.Y(n_73)
);

CKINVDCx16_ASAP7_75t_R g104 ( 
.A(n_73),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_39),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_74),
.B(n_97),
.Y(n_117)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_58),
.Y(n_75)
);

BUFx4f_ASAP7_75t_L g99 ( 
.A(n_75),
.Y(n_99)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_64),
.A2(n_25),
.B1(n_27),
.B2(n_29),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g126 ( 
.A(n_77),
.B(n_86),
.Y(n_126)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_78),
.Y(n_102)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_54),
.Y(n_79)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_79),
.Y(n_106)
);

INVx3_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

BUFx2_ASAP7_75t_L g120 ( 
.A(n_80),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_SL g81 ( 
.A1(n_49),
.A2(n_41),
.B1(n_45),
.B2(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_SL g82 ( 
.A(n_54),
.Y(n_82)
);

NAND4xp25_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_95),
.C(n_56),
.D(n_65),
.Y(n_100)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_54),
.Y(n_83)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_83),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_L g84 ( 
.A1(n_51),
.A2(n_60),
.B1(n_45),
.B2(n_50),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_54),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g115 ( 
.A(n_85),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g86 ( 
.A(n_62),
.B(n_18),
.Y(n_86)
);

INVx3_ASAP7_75t_L g87 ( 
.A(n_52),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_SL g103 ( 
.A1(n_87),
.A2(n_88),
.B1(n_91),
.B2(n_56),
.Y(n_103)
);

INVx6_ASAP7_75t_L g88 ( 
.A(n_56),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_L g89 ( 
.A1(n_53),
.A2(n_18),
.B1(n_36),
.B2(n_26),
.Y(n_89)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_57),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_53),
.A2(n_36),
.B1(n_26),
.B2(n_35),
.Y(n_92)
);

OAI22xp5_ASAP7_75t_L g93 ( 
.A1(n_59),
.A2(n_35),
.B1(n_21),
.B2(n_32),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_93),
.A2(n_23),
.B1(n_32),
.B2(n_22),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_52),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g116 ( 
.A(n_96),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_61),
.B(n_39),
.Y(n_97)
);

INVx2_ASAP7_75t_L g98 ( 
.A(n_75),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_98),
.B(n_107),
.Y(n_130)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_100),
.Y(n_136)
);

OAI22xp33_ASAP7_75t_L g101 ( 
.A1(n_95),
.A2(n_51),
.B1(n_60),
.B2(n_55),
.Y(n_101)
);

OAI22xp5_ASAP7_75t_L g143 ( 
.A1(n_101),
.A2(n_114),
.B1(n_127),
.B2(n_128),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_103),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g105 ( 
.A(n_80),
.Y(n_105)
);

BUFx3_ASAP7_75t_L g132 ( 
.A(n_105),
.Y(n_132)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_78),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g108 ( 
.A1(n_90),
.A2(n_60),
.B1(n_57),
.B2(n_65),
.Y(n_108)
);

INVxp67_ASAP7_75t_L g147 ( 
.A(n_108),
.Y(n_147)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g134 ( 
.A(n_109),
.B(n_123),
.Y(n_134)
);

MAJIxp5_ASAP7_75t_L g141 ( 
.A(n_111),
.B(n_23),
.C(n_39),
.Y(n_141)
);

OR2x2_ASAP7_75t_L g112 ( 
.A(n_77),
.B(n_90),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g129 ( 
.A(n_112),
.B(n_94),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_113),
.A2(n_81),
.B1(n_88),
.B2(n_87),
.Y(n_140)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_66),
.A2(n_32),
.B1(n_22),
.B2(n_21),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g153 ( 
.A(n_119),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g122 ( 
.A(n_85),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g154 ( 
.A(n_122),
.Y(n_154)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_91),
.Y(n_123)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_97),
.B(n_52),
.Y(n_125)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_71),
.Y(n_133)
);

AOI22xp33_ASAP7_75t_L g127 ( 
.A1(n_84),
.A2(n_32),
.B1(n_22),
.B2(n_38),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_SL g187 ( 
.A(n_129),
.B(n_131),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_SL g131 ( 
.A(n_112),
.B(n_94),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_133),
.B(n_135),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_L g135 ( 
.A(n_117),
.B(n_111),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g137 ( 
.A(n_117),
.B(n_74),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_149),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_120),
.Y(n_139)
);

CKINVDCx20_ASAP7_75t_R g158 ( 
.A(n_139),
.Y(n_158)
);

OAI22xp5_ASAP7_75t_L g157 ( 
.A1(n_140),
.A2(n_124),
.B1(n_128),
.B2(n_101),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_141),
.B(n_150),
.C(n_119),
.Y(n_168)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_102),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_142),
.B(n_145),
.Y(n_173)
);

AND2x2_ASAP7_75t_SL g144 ( 
.A(n_125),
.B(n_69),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g184 ( 
.A1(n_144),
.A2(n_34),
.B(n_96),
.Y(n_184)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_102),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_146),
.B(n_148),
.Y(n_181)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_102),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_121),
.B(n_83),
.Y(n_149)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_124),
.B(n_79),
.C(n_38),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g151 ( 
.A(n_126),
.B(n_1),
.Y(n_151)
);

INVxp33_ASAP7_75t_L g174 ( 
.A(n_151),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_120),
.B(n_1),
.Y(n_152)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_152),
.Y(n_162)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_99),
.Y(n_155)
);

INVxp67_ASAP7_75t_SL g179 ( 
.A(n_155),
.Y(n_179)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_99),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_156),
.A2(n_107),
.B1(n_98),
.B2(n_119),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_161),
.B1(n_175),
.B2(n_143),
.Y(n_190)
);

INVxp67_ASAP7_75t_L g159 ( 
.A(n_134),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_159),
.B(n_167),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g160 ( 
.A(n_144),
.B(n_99),
.Y(n_160)
);

MAJIxp5_ASAP7_75t_SL g204 ( 
.A(n_160),
.B(n_168),
.C(n_185),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_140),
.A2(n_110),
.B1(n_113),
.B2(n_123),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_130),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_163),
.B(n_166),
.Y(n_191)
);

XNOR2xp5_ASAP7_75t_L g164 ( 
.A(n_135),
.B(n_119),
.Y(n_164)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_164),
.B(n_153),
.Y(n_198)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_130),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_134),
.Y(n_167)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_170),
.B(n_172),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g195 ( 
.A(n_171),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_139),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_SL g175 ( 
.A1(n_150),
.A2(n_116),
.B1(n_52),
.B2(n_109),
.Y(n_175)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_143),
.A2(n_116),
.B1(n_118),
.B2(n_106),
.Y(n_176)
);

OAI22xp5_ASAP7_75t_SL g194 ( 
.A1(n_176),
.A2(n_145),
.B1(n_136),
.B2(n_147),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_137),
.B(n_38),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_178),
.Y(n_188)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_133),
.Y(n_178)
);

AO21x1_ASAP7_75t_L g180 ( 
.A1(n_136),
.A2(n_34),
.B(n_22),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g206 ( 
.A1(n_180),
.A2(n_155),
.B(n_146),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g182 ( 
.A(n_153),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g220 ( 
.A1(n_182),
.A2(n_183),
.B(n_4),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_132),
.Y(n_183)
);

OAI21xp5_ASAP7_75t_L g196 ( 
.A1(n_184),
.A2(n_138),
.B(n_152),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g185 ( 
.A(n_141),
.B(n_2),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_144),
.B(n_34),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_186),
.B(n_144),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g189 ( 
.A(n_181),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_189),
.B(n_193),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_L g233 ( 
.A1(n_190),
.A2(n_208),
.B1(n_215),
.B2(n_217),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_192),
.B(n_207),
.Y(n_228)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_179),
.Y(n_193)
);

AOI22xp5_ASAP7_75t_L g229 ( 
.A1(n_194),
.A2(n_203),
.B1(n_166),
.B2(n_162),
.Y(n_229)
);

OAI21xp5_ASAP7_75t_L g244 ( 
.A1(n_196),
.A2(n_200),
.B(n_209),
.Y(n_244)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_169),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_197),
.B(n_202),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_198),
.B(n_201),
.Y(n_227)
);

OAI21xp5_ASAP7_75t_L g200 ( 
.A1(n_186),
.A2(n_129),
.B(n_131),
.Y(n_200)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_164),
.B(n_165),
.Y(n_201)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_169),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_176),
.A2(n_148),
.B1(n_156),
.B2(n_151),
.Y(n_203)
);

AOI32xp33_ASAP7_75t_L g205 ( 
.A1(n_184),
.A2(n_153),
.A3(n_132),
.B1(n_105),
.B2(n_154),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_205),
.B(n_210),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_206),
.A2(n_218),
.B(n_220),
.Y(n_222)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_173),
.Y(n_207)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_180),
.A2(n_160),
.B1(n_170),
.B2(n_167),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_L g209 ( 
.A1(n_165),
.A2(n_132),
.B(n_105),
.Y(n_209)
);

XNOR2xp5_ASAP7_75t_SL g210 ( 
.A(n_178),
.B(n_105),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_211),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_168),
.B(n_104),
.C(n_115),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_213),
.B(n_219),
.C(n_6),
.Y(n_246)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_177),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_214),
.B(n_216),
.Y(n_230)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_175),
.A2(n_142),
.B1(n_122),
.B2(n_34),
.Y(n_215)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_187),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_160),
.A2(n_2),
.B1(n_3),
.B2(n_4),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_159),
.A2(n_2),
.B(n_3),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_163),
.B(n_3),
.C(n_4),
.Y(n_219)
);

AOI21xp5_ASAP7_75t_L g224 ( 
.A1(n_220),
.A2(n_158),
.B(n_172),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_SL g248 ( 
.A1(n_224),
.A2(n_218),
.B1(n_217),
.B2(n_195),
.Y(n_248)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_199),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_225),
.B(n_229),
.Y(n_263)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_212),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g256 ( 
.A(n_226),
.B(n_231),
.Y(n_256)
);

INVx1_ASAP7_75t_SL g231 ( 
.A(n_206),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g235 ( 
.A(n_198),
.B(n_158),
.C(n_183),
.Y(n_235)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_235),
.B(n_245),
.C(n_246),
.Y(n_250)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_191),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_SL g247 ( 
.A(n_236),
.B(n_239),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g237 ( 
.A(n_201),
.B(n_210),
.Y(n_237)
);

XOR2xp5_ASAP7_75t_L g258 ( 
.A(n_237),
.B(n_204),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_188),
.B(n_162),
.Y(n_238)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_238),
.Y(n_251)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_188),
.Y(n_239)
);

FAx1_ASAP7_75t_SL g240 ( 
.A(n_192),
.B(n_185),
.CI(n_187),
.CON(n_240),
.SN(n_240)
);

OAI21xp33_ASAP7_75t_L g260 ( 
.A1(n_240),
.A2(n_194),
.B(n_219),
.Y(n_260)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_241),
.Y(n_252)
);

CKINVDCx16_ASAP7_75t_R g242 ( 
.A(n_215),
.Y(n_242)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_242),
.B(n_203),
.Y(n_253)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_190),
.A2(n_180),
.B1(n_174),
.B2(n_185),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_243),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_213),
.B(n_5),
.C(n_16),
.Y(n_245)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g249 ( 
.A(n_234),
.Y(n_249)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_249),
.Y(n_268)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_253),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_226),
.B(n_200),
.Y(n_254)
);

CKINVDCx14_ASAP7_75t_R g281 ( 
.A(n_254),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_227),
.B(n_204),
.C(n_196),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_255),
.B(n_264),
.C(n_221),
.Y(n_270)
);

CKINVDCx20_ASAP7_75t_R g257 ( 
.A(n_228),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g275 ( 
.A(n_257),
.Y(n_275)
);

XOR2xp5_ASAP7_75t_L g271 ( 
.A(n_258),
.B(n_261),
.Y(n_271)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_228),
.Y(n_259)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_259),
.Y(n_276)
);

MAJx2_ASAP7_75t_L g284 ( 
.A(n_260),
.B(n_240),
.C(n_245),
.Y(n_284)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_227),
.B(n_211),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_266),
.B1(n_224),
.B2(n_222),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_235),
.B(n_6),
.C(n_7),
.Y(n_264)
);

XNOR2xp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_8),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g285 ( 
.A(n_265),
.B(n_264),
.Y(n_285)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_238),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_241),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_267)
);

AOI22xp5_ASAP7_75t_L g273 ( 
.A1(n_267),
.A2(n_233),
.B1(n_225),
.B2(n_230),
.Y(n_273)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_282),
.C(n_285),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_255),
.B(n_236),
.C(n_221),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_272),
.B(n_274),
.C(n_278),
.Y(n_299)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_273),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g274 ( 
.A(n_250),
.B(n_244),
.C(n_223),
.Y(n_274)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_277),
.Y(n_292)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_250),
.B(n_244),
.C(n_230),
.Y(n_278)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_252),
.A2(n_231),
.B1(n_232),
.B2(n_222),
.Y(n_279)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_279),
.Y(n_293)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_258),
.B(n_246),
.C(n_229),
.Y(n_282)
);

CKINVDCx16_ASAP7_75t_R g283 ( 
.A(n_263),
.Y(n_283)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_283),
.Y(n_295)
);

XOR2x1_ASAP7_75t_SL g287 ( 
.A(n_284),
.B(n_265),
.Y(n_287)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_273),
.B(n_267),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_286),
.B(n_279),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g307 ( 
.A(n_287),
.B(n_288),
.Y(n_307)
);

XOR2xp5_ASAP7_75t_L g288 ( 
.A(n_271),
.B(n_261),
.Y(n_288)
);

XOR2xp5_ASAP7_75t_L g290 ( 
.A(n_271),
.B(n_256),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_290),
.B(n_281),
.C(n_280),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_L g294 ( 
.A(n_272),
.B(n_247),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g306 ( 
.A(n_294),
.B(n_298),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_256),
.C(n_252),
.Y(n_296)
);

MAJIxp5_ASAP7_75t_L g309 ( 
.A(n_296),
.B(n_300),
.C(n_290),
.Y(n_309)
);

AOI22xp33_ASAP7_75t_SL g297 ( 
.A1(n_275),
.A2(n_251),
.B1(n_248),
.B2(n_262),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_L g310 ( 
.A1(n_297),
.A2(n_269),
.B1(n_293),
.B2(n_291),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_270),
.B(n_249),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_282),
.B(n_251),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g301 ( 
.A(n_299),
.B(n_274),
.C(n_268),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_301),
.B(n_303),
.C(n_304),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g316 ( 
.A(n_302),
.Y(n_316)
);

INVx1_ASAP7_75t_SL g303 ( 
.A(n_295),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_299),
.B(n_268),
.C(n_276),
.Y(n_304)
);

NOR2xp67_ASAP7_75t_SL g305 ( 
.A(n_287),
.B(n_284),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_SL g313 ( 
.A(n_305),
.B(n_308),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_289),
.B(n_285),
.Y(n_308)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_309),
.B(n_9),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g318 ( 
.A(n_310),
.B(n_311),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g311 ( 
.A(n_288),
.B(n_300),
.Y(n_311)
);

XOR2xp5_ASAP7_75t_L g317 ( 
.A(n_312),
.B(n_10),
.Y(n_317)
);

OAI22xp5_ASAP7_75t_SL g314 ( 
.A1(n_304),
.A2(n_292),
.B1(n_297),
.B2(n_240),
.Y(n_314)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_314),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_SL g324 ( 
.A(n_315),
.B(n_317),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g319 ( 
.A1(n_301),
.A2(n_16),
.B1(n_12),
.B2(n_14),
.Y(n_319)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_319),
.Y(n_325)
);

AO21x1_ASAP7_75t_L g320 ( 
.A1(n_307),
.A2(n_303),
.B(n_306),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g326 ( 
.A(n_320),
.B(n_11),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_SL g323 ( 
.A1(n_313),
.A2(n_307),
.B(n_12),
.Y(n_323)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_323),
.B(n_326),
.C(n_314),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_316),
.B(n_11),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g332 ( 
.A(n_327),
.B(n_328),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_321),
.B(n_315),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g333 ( 
.A1(n_329),
.A2(n_330),
.B(n_331),
.Y(n_333)
);

AO21x1_ASAP7_75t_L g330 ( 
.A1(n_322),
.A2(n_320),
.B(n_321),
.Y(n_330)
);

XNOR2x1_ASAP7_75t_SL g331 ( 
.A(n_328),
.B(n_317),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_333),
.B(n_332),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g335 ( 
.A(n_334),
.B(n_324),
.Y(n_335)
);

HB1xp67_ASAP7_75t_L g336 ( 
.A(n_335),
.Y(n_336)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_336),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g338 ( 
.A1(n_337),
.A2(n_325),
.B(n_318),
.Y(n_338)
);

AOI21xp5_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_12),
.B(n_14),
.Y(n_339)
);

MAJIxp5_ASAP7_75t_L g340 ( 
.A(n_339),
.B(n_15),
.C(n_329),
.Y(n_340)
);


endmodule