module fake_netlist_1_7962_n_895 (n_117, n_44, n_133, n_149, n_81, n_69, n_204, n_185, n_22, n_203, n_57, n_88, n_52, n_26, n_50, n_33, n_102, n_73, n_49, n_119, n_141, n_115, n_97, n_80, n_167, n_107, n_158, n_60, n_114, n_121, n_41, n_35, n_94, n_65, n_171, n_196, n_125, n_192, n_9, n_161, n_10, n_177, n_130, n_189, n_103, n_19, n_87, n_137, n_180, n_104, n_160, n_98, n_74, n_206, n_154, n_7, n_29, n_195, n_165, n_146, n_45, n_85, n_181, n_101, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_91, n_108, n_116, n_155, n_209, n_139, n_16, n_13, n_198, n_169, n_193, n_152, n_113, n_95, n_124, n_156, n_128, n_120, n_129, n_70, n_17, n_63, n_14, n_71, n_90, n_56, n_135, n_42, n_188, n_24, n_78, n_197, n_201, n_6, n_4, n_127, n_170, n_40, n_111, n_157, n_79, n_202, n_38, n_64, n_142, n_184, n_191, n_200, n_46, n_31, n_208, n_58, n_122, n_187, n_138, n_126, n_178, n_118, n_32, n_0, n_179, n_84, n_131, n_112, n_55, n_205, n_12, n_86, n_143, n_182, n_166, n_162, n_186, n_75, n_163, n_105, n_159, n_174, n_72, n_136, n_43, n_76, n_89, n_176, n_68, n_144, n_27, n_53, n_183, n_67, n_77, n_20, n_2, n_147, n_199, n_54, n_148, n_123, n_83, n_172, n_28, n_48, n_100, n_92, n_11, n_25, n_30, n_59, n_150, n_168, n_194, n_3, n_18, n_110, n_66, n_134, n_1, n_164, n_82, n_106, n_175, n_15, n_173, n_190, n_145, n_153, n_61, n_21, n_99, n_109, n_93, n_132, n_151, n_51, n_140, n_207, n_96, n_39, n_895);
input n_117;
input n_44;
input n_133;
input n_149;
input n_81;
input n_69;
input n_204;
input n_185;
input n_22;
input n_203;
input n_57;
input n_88;
input n_52;
input n_26;
input n_50;
input n_33;
input n_102;
input n_73;
input n_49;
input n_119;
input n_141;
input n_115;
input n_97;
input n_80;
input n_167;
input n_107;
input n_158;
input n_60;
input n_114;
input n_121;
input n_41;
input n_35;
input n_94;
input n_65;
input n_171;
input n_196;
input n_125;
input n_192;
input n_9;
input n_161;
input n_10;
input n_177;
input n_130;
input n_189;
input n_103;
input n_19;
input n_87;
input n_137;
input n_180;
input n_104;
input n_160;
input n_98;
input n_74;
input n_206;
input n_154;
input n_7;
input n_29;
input n_195;
input n_165;
input n_146;
input n_45;
input n_85;
input n_181;
input n_101;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_91;
input n_108;
input n_116;
input n_155;
input n_209;
input n_139;
input n_16;
input n_13;
input n_198;
input n_169;
input n_193;
input n_152;
input n_113;
input n_95;
input n_124;
input n_156;
input n_128;
input n_120;
input n_129;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_90;
input n_56;
input n_135;
input n_42;
input n_188;
input n_24;
input n_78;
input n_197;
input n_201;
input n_6;
input n_4;
input n_127;
input n_170;
input n_40;
input n_111;
input n_157;
input n_79;
input n_202;
input n_38;
input n_64;
input n_142;
input n_184;
input n_191;
input n_200;
input n_46;
input n_31;
input n_208;
input n_58;
input n_122;
input n_187;
input n_138;
input n_126;
input n_178;
input n_118;
input n_32;
input n_0;
input n_179;
input n_84;
input n_131;
input n_112;
input n_55;
input n_205;
input n_12;
input n_86;
input n_143;
input n_182;
input n_166;
input n_162;
input n_186;
input n_75;
input n_163;
input n_105;
input n_159;
input n_174;
input n_72;
input n_136;
input n_43;
input n_76;
input n_89;
input n_176;
input n_68;
input n_144;
input n_27;
input n_53;
input n_183;
input n_67;
input n_77;
input n_20;
input n_2;
input n_147;
input n_199;
input n_54;
input n_148;
input n_123;
input n_83;
input n_172;
input n_28;
input n_48;
input n_100;
input n_92;
input n_11;
input n_25;
input n_30;
input n_59;
input n_150;
input n_168;
input n_194;
input n_3;
input n_18;
input n_110;
input n_66;
input n_134;
input n_1;
input n_164;
input n_82;
input n_106;
input n_175;
input n_15;
input n_173;
input n_190;
input n_145;
input n_153;
input n_61;
input n_21;
input n_99;
input n_109;
input n_93;
input n_132;
input n_151;
input n_51;
input n_140;
input n_207;
input n_96;
input n_39;
output n_895;
wire n_663;
wire n_707;
wire n_791;
wire n_361;
wire n_513;
wire n_838;
wire n_705;
wire n_603;
wire n_604;
wire n_858;
wire n_590;
wire n_407;
wire n_885;
wire n_755;
wire n_646;
wire n_792;
wire n_284;
wire n_278;
wire n_500;
wire n_848;
wire n_607;
wire n_808;
wire n_829;
wire n_431;
wire n_484;
wire n_852;
wire n_862;
wire n_496;
wire n_667;
wire n_311;
wire n_801;
wire n_292;
wire n_309;
wire n_701;
wire n_612;
wire n_328;
wire n_655;
wire n_468;
wire n_743;
wire n_523;
wire n_229;
wire n_757;
wire n_750;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_770;
wire n_252;
wire n_878;
wire n_814;
wire n_637;
wire n_817;
wire n_802;
wire n_856;
wire n_353;
wire n_564;
wire n_779;
wire n_528;
wire n_288;
wire n_383;
wire n_661;
wire n_850;
wire n_762;
wire n_672;
wire n_532;
wire n_627;
wire n_758;
wire n_544;
wire n_890;
wire n_400;
wire n_787;
wire n_853;
wire n_296;
wire n_765;
wire n_386;
wire n_432;
wire n_659;
wire n_807;
wire n_877;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_783;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_789;
wire n_330;
wire n_587;
wire n_662;
wire n_678;
wire n_387;
wire n_434;
wire n_384;
wire n_227;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_812;
wire n_598;
wire n_489;
wire n_777;
wire n_732;
wire n_752;
wire n_351;
wire n_860;
wire n_401;
wire n_461;
wire n_305;
wire n_599;
wire n_228;
wire n_724;
wire n_786;
wire n_857;
wire n_345;
wire n_360;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_796;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_773;
wire n_847;
wire n_840;
wire n_392;
wire n_668;
wire n_846;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_563;
wire n_638;
wire n_830;
wire n_560;
wire n_517;
wire n_479;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_726;
wire n_780;
wire n_712;
wire n_447;
wire n_872;
wire n_608;
wire n_567;
wire n_809;
wire n_888;
wire n_580;
wire n_502;
wire n_543;
wire n_854;
wire n_312;
wire n_455;
wire n_529;
wire n_880;
wire n_630;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_865;
wire n_647;
wire n_367;
wire n_644;
wire n_250;
wire n_764;
wire n_314;
wire n_237;
wire n_255;
wire n_426;
wire n_624;
wire n_725;
wire n_769;
wire n_818;
wire n_844;
wire n_230;
wire n_274;
wire n_738;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_798;
wire n_241;
wire n_575;
wire n_238;
wire n_711;
wire n_318;
wire n_884;
wire n_887;
wire n_471;
wire n_632;
wire n_767;
wire n_828;
wire n_293;
wire n_506;
wire n_533;
wire n_393;
wire n_490;
wire n_247;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_826;
wire n_304;
wire n_399;
wire n_892;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_863;
wire n_322;
wire n_310;
wire n_708;
wire n_307;
wire n_634;
wire n_610;
wire n_730;
wire n_735;
wire n_696;
wire n_771;
wire n_784;
wire n_474;
wire n_354;
wire n_402;
wire n_893;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_415;
wire n_243;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_813;
wire n_352;
wire n_746;
wire n_619;
wire n_882;
wire n_268;
wire n_501;
wire n_248;
wire n_871;
wire n_803;
wire n_299;
wire n_338;
wire n_519;
wire n_699;
wire n_729;
wire n_805;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_849;
wire n_864;
wire n_810;
wire n_329;
wire n_251;
wire n_747;
wire n_635;
wire n_889;
wire n_731;
wire n_689;
wire n_525;
wire n_218;
wire n_876;
wire n_886;
wire n_507;
wire n_605;
wire n_719;
wire n_611;
wire n_704;
wire n_633;
wire n_873;
wire n_271;
wire n_760;
wire n_751;
wire n_800;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_259;
wire n_308;
wire n_546;
wire n_412;
wire n_664;
wire n_827;
wire n_565;
wire n_224;
wire n_788;
wire n_219;
wire n_475;
wire n_578;
wire n_542;
wire n_537;
wire n_214;
wire n_660;
wire n_430;
wire n_839;
wire n_450;
wire n_579;
wire n_776;
wire n_879;
wire n_403;
wire n_557;
wire n_516;
wire n_842;
wire n_254;
wire n_549;
wire n_622;
wire n_832;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_526;
wire n_276;
wire n_649;
wire n_320;
wire n_768;
wire n_869;
wire n_797;
wire n_285;
wire n_420;
wire n_446;
wire n_423;
wire n_342;
wire n_666;
wire n_621;
wire n_799;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_874;
wire n_217;
wire n_388;
wire n_454;
wire n_687;
wire n_273;
wire n_505;
wire n_706;
wire n_823;
wire n_822;
wire n_390;
wire n_682;
wire n_514;
wire n_486;
wire n_720;
wire n_568;
wire n_245;
wire n_357;
wire n_653;
wire n_716;
wire n_881;
wire n_260;
wire n_806;
wire n_539;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_718;
wire n_536;
wire n_816;
wire n_265;
wire n_264;
wire n_522;
wire n_883;
wire n_573;
wire n_673;
wire n_669;
wire n_754;
wire n_775;
wire n_616;
wire n_365;
wire n_717;
wire n_541;
wire n_363;
wire n_315;
wire n_409;
wire n_733;
wire n_861;
wire n_295;
wire n_654;
wire n_263;
wire n_894;
wire n_495;
wire n_364;
wire n_428;
wire n_566;
wire n_794;
wire n_376;
wire n_639;
wire n_552;
wire n_744;
wire n_677;
wire n_344;
wire n_503;
wire n_283;
wire n_756;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_870;
wire n_790;
wire n_761;
wire n_615;
wire n_212;
wire n_472;
wire n_419;
wire n_851;
wire n_825;
wire n_396;
wire n_804;
wire n_477;
wire n_815;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_721;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_821;
wire n_745;
wire n_684;
wire n_440;
wire n_553;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_723;
wire n_811;
wire n_749;
wire n_835;
wire n_225;
wire n_535;
wire n_530;
wire n_737;
wire n_778;
wire n_220;
wire n_358;
wire n_795;
wire n_267;
wire n_221;
wire n_456;
wire n_782;
wire n_449;
wire n_300;
wire n_734;
wire n_524;
wire n_584;
wire n_875;
wire n_497;
wire n_728;
wire n_339;
wire n_657;
wire n_583;
wire n_763;
wire n_620;
wire n_240;
wire n_841;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_441;
wire n_836;
wire n_561;
wire n_335;
wire n_272;
wire n_741;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_766;
wire n_602;
wire n_831;
wire n_859;
wire n_424;
wire n_714;
wire n_629;
wire n_569;
wire n_297;
wire n_837;
wire n_410;
wire n_774;
wire n_867;
wire n_377;
wire n_510;
wire n_343;
wire n_675;
wire n_291;
wire n_504;
wire n_581;
wire n_458;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_855;
wire n_722;
wire n_618;
wire n_834;
wire n_727;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_785;
wire n_375;
wire n_451;
wire n_487;
wire n_748;
wire n_371;
wire n_688;
wire n_868;
wire n_323;
wire n_473;
wire n_347;
wire n_820;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_843;
wire n_266;
wire n_683;
wire n_213;
wire n_824;
wire n_538;
wire n_793;
wire n_492;
wire n_592;
wire n_753;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_521;
wire n_625;
wire n_650;
wire n_695;
wire n_469;
wire n_742;
wire n_585;
wire n_845;
wire n_713;
wire n_891;
wire n_457;
wire n_595;
wire n_759;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_833;
wire n_866;
wire n_736;
wire n_287;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_781;
wire n_421;
wire n_709;
wire n_739;
wire n_740;
wire n_483;
wire n_408;
wire n_772;
wire n_290;
wire n_405;
wire n_819;
wire n_280;
wire n_395;
wire n_406;
wire n_491;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g210 ( .A(n_14), .Y(n_210) );
INVx1_ASAP7_75t_L g211 ( .A(n_125), .Y(n_211) );
INVx1_ASAP7_75t_L g212 ( .A(n_136), .Y(n_212) );
INVxp33_ASAP7_75t_SL g213 ( .A(n_129), .Y(n_213) );
INVx1_ASAP7_75t_L g214 ( .A(n_33), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g215 ( .A(n_95), .Y(n_215) );
BUFx6f_ASAP7_75t_L g216 ( .A(n_2), .Y(n_216) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_102), .Y(n_217) );
CKINVDCx20_ASAP7_75t_R g218 ( .A(n_137), .Y(n_218) );
INVx2_ASAP7_75t_L g219 ( .A(n_74), .Y(n_219) );
INVx1_ASAP7_75t_L g220 ( .A(n_201), .Y(n_220) );
INVx1_ASAP7_75t_L g221 ( .A(n_121), .Y(n_221) );
INVx1_ASAP7_75t_L g222 ( .A(n_17), .Y(n_222) );
BUFx2_ASAP7_75t_L g223 ( .A(n_118), .Y(n_223) );
CKINVDCx5p33_ASAP7_75t_R g224 ( .A(n_194), .Y(n_224) );
INVx1_ASAP7_75t_L g225 ( .A(n_204), .Y(n_225) );
CKINVDCx14_ASAP7_75t_R g226 ( .A(n_0), .Y(n_226) );
BUFx3_ASAP7_75t_L g227 ( .A(n_206), .Y(n_227) );
BUFx6f_ASAP7_75t_L g228 ( .A(n_177), .Y(n_228) );
INVx2_ASAP7_75t_L g229 ( .A(n_110), .Y(n_229) );
INVx1_ASAP7_75t_L g230 ( .A(n_107), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_18), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_109), .Y(n_232) );
BUFx2_ASAP7_75t_L g233 ( .A(n_113), .Y(n_233) );
INVxp67_ASAP7_75t_SL g234 ( .A(n_87), .Y(n_234) );
INVx1_ASAP7_75t_L g235 ( .A(n_209), .Y(n_235) );
CKINVDCx5p33_ASAP7_75t_R g236 ( .A(n_191), .Y(n_236) );
INVx1_ASAP7_75t_L g237 ( .A(n_190), .Y(n_237) );
INVxp67_ASAP7_75t_SL g238 ( .A(n_178), .Y(n_238) );
BUFx6f_ASAP7_75t_L g239 ( .A(n_154), .Y(n_239) );
CKINVDCx5p33_ASAP7_75t_R g240 ( .A(n_122), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_161), .Y(n_241) );
INVx1_ASAP7_75t_L g242 ( .A(n_172), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_112), .Y(n_243) );
CKINVDCx20_ASAP7_75t_R g244 ( .A(n_205), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_49), .Y(n_245) );
INVx1_ASAP7_75t_L g246 ( .A(n_3), .Y(n_246) );
CKINVDCx20_ASAP7_75t_R g247 ( .A(n_9), .Y(n_247) );
INVx1_ASAP7_75t_L g248 ( .A(n_119), .Y(n_248) );
CKINVDCx20_ASAP7_75t_R g249 ( .A(n_207), .Y(n_249) );
CKINVDCx20_ASAP7_75t_R g250 ( .A(n_189), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_141), .Y(n_251) );
INVx1_ASAP7_75t_L g252 ( .A(n_203), .Y(n_252) );
INVx2_ASAP7_75t_L g253 ( .A(n_159), .Y(n_253) );
INVx1_ASAP7_75t_L g254 ( .A(n_86), .Y(n_254) );
INVx1_ASAP7_75t_L g255 ( .A(n_155), .Y(n_255) );
INVx1_ASAP7_75t_L g256 ( .A(n_81), .Y(n_256) );
CKINVDCx20_ASAP7_75t_R g257 ( .A(n_39), .Y(n_257) );
BUFx6f_ASAP7_75t_L g258 ( .A(n_111), .Y(n_258) );
CKINVDCx5p33_ASAP7_75t_R g259 ( .A(n_164), .Y(n_259) );
INVx2_ASAP7_75t_SL g260 ( .A(n_24), .Y(n_260) );
INVx1_ASAP7_75t_L g261 ( .A(n_208), .Y(n_261) );
CKINVDCx5p33_ASAP7_75t_R g262 ( .A(n_188), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_187), .Y(n_263) );
INVx1_ASAP7_75t_L g264 ( .A(n_138), .Y(n_264) );
OR2x2_ASAP7_75t_L g265 ( .A(n_3), .B(n_160), .Y(n_265) );
INVx2_ASAP7_75t_SL g266 ( .A(n_199), .Y(n_266) );
CKINVDCx5p33_ASAP7_75t_R g267 ( .A(n_57), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_40), .Y(n_268) );
BUFx3_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
INVx1_ASAP7_75t_L g270 ( .A(n_64), .Y(n_270) );
INVx1_ASAP7_75t_L g271 ( .A(n_179), .Y(n_271) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_12), .Y(n_272) );
INVx1_ASAP7_75t_L g273 ( .A(n_1), .Y(n_273) );
CKINVDCx16_ASAP7_75t_R g274 ( .A(n_139), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_38), .Y(n_275) );
INVx1_ASAP7_75t_L g276 ( .A(n_7), .Y(n_276) );
INVxp67_ASAP7_75t_SL g277 ( .A(n_17), .Y(n_277) );
INVx1_ASAP7_75t_L g278 ( .A(n_148), .Y(n_278) );
INVx1_ASAP7_75t_L g279 ( .A(n_92), .Y(n_279) );
INVx1_ASAP7_75t_L g280 ( .A(n_75), .Y(n_280) );
INVx1_ASAP7_75t_L g281 ( .A(n_69), .Y(n_281) );
INVx1_ASAP7_75t_L g282 ( .A(n_7), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_6), .Y(n_283) );
INVx1_ASAP7_75t_L g284 ( .A(n_165), .Y(n_284) );
INVx1_ASAP7_75t_L g285 ( .A(n_183), .Y(n_285) );
INVx1_ASAP7_75t_L g286 ( .A(n_140), .Y(n_286) );
BUFx2_ASAP7_75t_L g287 ( .A(n_26), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_126), .Y(n_288) );
INVx1_ASAP7_75t_L g289 ( .A(n_175), .Y(n_289) );
INVxp67_ASAP7_75t_SL g290 ( .A(n_128), .Y(n_290) );
INVx2_ASAP7_75t_L g291 ( .A(n_94), .Y(n_291) );
CKINVDCx20_ASAP7_75t_R g292 ( .A(n_51), .Y(n_292) );
INVx2_ASAP7_75t_L g293 ( .A(n_98), .Y(n_293) );
INVx2_ASAP7_75t_L g294 ( .A(n_198), .Y(n_294) );
INVx1_ASAP7_75t_L g295 ( .A(n_18), .Y(n_295) );
CKINVDCx5p33_ASAP7_75t_R g296 ( .A(n_58), .Y(n_296) );
INVxp67_ASAP7_75t_L g297 ( .A(n_91), .Y(n_297) );
INVx1_ASAP7_75t_L g298 ( .A(n_36), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_197), .Y(n_299) );
INVx1_ASAP7_75t_L g300 ( .A(n_57), .Y(n_300) );
CKINVDCx20_ASAP7_75t_R g301 ( .A(n_93), .Y(n_301) );
CKINVDCx5p33_ASAP7_75t_R g302 ( .A(n_186), .Y(n_302) );
CKINVDCx5p33_ASAP7_75t_R g303 ( .A(n_108), .Y(n_303) );
INVx1_ASAP7_75t_L g304 ( .A(n_34), .Y(n_304) );
INVx1_ASAP7_75t_L g305 ( .A(n_149), .Y(n_305) );
INVxp67_ASAP7_75t_SL g306 ( .A(n_67), .Y(n_306) );
INVx1_ASAP7_75t_L g307 ( .A(n_5), .Y(n_307) );
INVx1_ASAP7_75t_L g308 ( .A(n_116), .Y(n_308) );
BUFx3_ASAP7_75t_L g309 ( .A(n_152), .Y(n_309) );
NOR2xp67_ASAP7_75t_L g310 ( .A(n_176), .B(n_185), .Y(n_310) );
HB1xp67_ASAP7_75t_L g311 ( .A(n_28), .Y(n_311) );
INVx1_ASAP7_75t_L g312 ( .A(n_78), .Y(n_312) );
XOR2xp5_ASAP7_75t_L g313 ( .A(n_120), .B(n_90), .Y(n_313) );
INVx2_ASAP7_75t_L g314 ( .A(n_163), .Y(n_314) );
CKINVDCx20_ASAP7_75t_R g315 ( .A(n_162), .Y(n_315) );
CKINVDCx16_ASAP7_75t_R g316 ( .A(n_33), .Y(n_316) );
CKINVDCx5p33_ASAP7_75t_R g317 ( .A(n_5), .Y(n_317) );
INVx1_ASAP7_75t_L g318 ( .A(n_167), .Y(n_318) );
CKINVDCx20_ASAP7_75t_R g319 ( .A(n_19), .Y(n_319) );
BUFx6f_ASAP7_75t_L g320 ( .A(n_158), .Y(n_320) );
CKINVDCx5p33_ASAP7_75t_R g321 ( .A(n_24), .Y(n_321) );
INVx1_ASAP7_75t_L g322 ( .A(n_173), .Y(n_322) );
INVx2_ASAP7_75t_L g323 ( .A(n_37), .Y(n_323) );
INVxp33_ASAP7_75t_L g324 ( .A(n_142), .Y(n_324) );
CKINVDCx20_ASAP7_75t_R g325 ( .A(n_49), .Y(n_325) );
CKINVDCx5p33_ASAP7_75t_R g326 ( .A(n_130), .Y(n_326) );
CKINVDCx14_ASAP7_75t_R g327 ( .A(n_65), .Y(n_327) );
BUFx6f_ASAP7_75t_L g328 ( .A(n_73), .Y(n_328) );
XNOR2x1_ASAP7_75t_L g329 ( .A(n_202), .B(n_115), .Y(n_329) );
INVx1_ASAP7_75t_L g330 ( .A(n_200), .Y(n_330) );
BUFx5_ASAP7_75t_L g331 ( .A(n_184), .Y(n_331) );
INVx1_ASAP7_75t_L g332 ( .A(n_39), .Y(n_332) );
INVxp67_ASAP7_75t_L g333 ( .A(n_169), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_323), .Y(n_334) );
INVx2_ASAP7_75t_L g335 ( .A(n_331), .Y(n_335) );
AND2x2_ASAP7_75t_L g336 ( .A(n_324), .B(n_0), .Y(n_336) );
NOR2xp33_ASAP7_75t_L g337 ( .A(n_266), .B(n_1), .Y(n_337) );
INVx2_ASAP7_75t_L g338 ( .A(n_331), .Y(n_338) );
CKINVDCx5p33_ASAP7_75t_R g339 ( .A(n_274), .Y(n_339) );
OA21x2_ASAP7_75t_L g340 ( .A1(n_219), .A2(n_77), .B(n_76), .Y(n_340) );
AND2x4_ASAP7_75t_L g341 ( .A(n_223), .B(n_2), .Y(n_341) );
INVx2_ASAP7_75t_L g342 ( .A(n_331), .Y(n_342) );
NOR2xp33_ASAP7_75t_L g343 ( .A(n_233), .B(n_4), .Y(n_343) );
INVx1_ASAP7_75t_L g344 ( .A(n_211), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_227), .B(n_4), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_226), .A2(n_8), .B1(n_10), .B2(n_11), .Y(n_346) );
INVx5_ASAP7_75t_L g347 ( .A(n_228), .Y(n_347) );
AND2x2_ASAP7_75t_L g348 ( .A(n_324), .B(n_8), .Y(n_348) );
BUFx6f_ASAP7_75t_L g349 ( .A(n_228), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_212), .Y(n_350) );
BUFx2_ASAP7_75t_L g351 ( .A(n_226), .Y(n_351) );
BUFx6f_ASAP7_75t_L g352 ( .A(n_228), .Y(n_352) );
OAI22xp5_ASAP7_75t_L g353 ( .A1(n_327), .A2(n_10), .B1(n_11), .B2(n_12), .Y(n_353) );
AND2x4_ASAP7_75t_L g354 ( .A(n_227), .B(n_13), .Y(n_354) );
BUFx12f_ASAP7_75t_L g355 ( .A(n_236), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g356 ( .A(n_260), .B(n_13), .Y(n_356) );
INVx2_ASAP7_75t_L g357 ( .A(n_331), .Y(n_357) );
AND2x4_ASAP7_75t_L g358 ( .A(n_269), .B(n_14), .Y(n_358) );
INVx1_ASAP7_75t_L g359 ( .A(n_220), .Y(n_359) );
NOR2xp33_ASAP7_75t_L g360 ( .A(n_221), .B(n_15), .Y(n_360) );
AOI22xp33_ASAP7_75t_SL g361 ( .A1(n_247), .A2(n_15), .B1(n_16), .B2(n_19), .Y(n_361) );
INVx2_ASAP7_75t_L g362 ( .A(n_331), .Y(n_362) );
INVx2_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
INVx1_ASAP7_75t_L g364 ( .A(n_225), .Y(n_364) );
INVx2_ASAP7_75t_L g365 ( .A(n_331), .Y(n_365) );
AND2x4_ASAP7_75t_L g366 ( .A(n_269), .B(n_16), .Y(n_366) );
OAI22xp5_ASAP7_75t_SL g367 ( .A1(n_247), .A2(n_20), .B1(n_21), .B2(n_22), .Y(n_367) );
BUFx8_ASAP7_75t_SL g368 ( .A(n_257), .Y(n_368) );
INVx1_ASAP7_75t_L g369 ( .A(n_230), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_349), .Y(n_370) );
INVxp67_ASAP7_75t_L g371 ( .A(n_351), .Y(n_371) );
AND2x6_ASAP7_75t_L g372 ( .A(n_345), .B(n_288), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g373 ( .A(n_344), .B(n_219), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_335), .Y(n_374) );
BUFx6f_ASAP7_75t_L g375 ( .A(n_349), .Y(n_375) );
INVx1_ASAP7_75t_L g376 ( .A(n_335), .Y(n_376) );
INVx1_ASAP7_75t_L g377 ( .A(n_335), .Y(n_377) );
AND2x2_ASAP7_75t_L g378 ( .A(n_351), .B(n_287), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_338), .Y(n_379) );
INVx4_ASAP7_75t_L g380 ( .A(n_345), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_344), .B(n_229), .Y(n_381) );
AND2x2_ASAP7_75t_L g382 ( .A(n_336), .B(n_327), .Y(n_382) );
AND2x2_ASAP7_75t_L g383 ( .A(n_336), .B(n_311), .Y(n_383) );
INVx2_ASAP7_75t_L g384 ( .A(n_349), .Y(n_384) );
INVx2_ASAP7_75t_L g385 ( .A(n_349), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g386 ( .A1(n_350), .A2(n_214), .B1(n_222), .B2(n_210), .Y(n_386) );
NOR2xp33_ASAP7_75t_L g387 ( .A(n_350), .B(n_297), .Y(n_387) );
AND2x6_ASAP7_75t_L g388 ( .A(n_345), .B(n_354), .Y(n_388) );
INVx3_ASAP7_75t_L g389 ( .A(n_345), .Y(n_389) );
AND2x2_ASAP7_75t_L g390 ( .A(n_336), .B(n_316), .Y(n_390) );
NAND2xp5_ASAP7_75t_SL g391 ( .A(n_341), .B(n_236), .Y(n_391) );
INVx2_ASAP7_75t_L g392 ( .A(n_349), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_338), .Y(n_393) );
AND2x2_ASAP7_75t_L g394 ( .A(n_348), .B(n_240), .Y(n_394) );
BUFx6f_ASAP7_75t_L g395 ( .A(n_349), .Y(n_395) );
INVx3_ASAP7_75t_L g396 ( .A(n_354), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_359), .B(n_229), .Y(n_397) );
INVx2_ASAP7_75t_L g398 ( .A(n_349), .Y(n_398) );
NOR2xp33_ASAP7_75t_L g399 ( .A(n_359), .B(n_333), .Y(n_399) );
NOR2xp33_ASAP7_75t_L g400 ( .A(n_364), .B(n_241), .Y(n_400) );
BUFx2_ASAP7_75t_L g401 ( .A(n_355), .Y(n_401) );
INVx1_ASAP7_75t_SL g402 ( .A(n_348), .Y(n_402) );
INVx3_ASAP7_75t_L g403 ( .A(n_354), .Y(n_403) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_355), .Y(n_404) );
BUFx2_ASAP7_75t_L g405 ( .A(n_355), .Y(n_405) );
INVx1_ASAP7_75t_L g406 ( .A(n_342), .Y(n_406) );
OR2x2_ASAP7_75t_L g407 ( .A(n_341), .B(n_364), .Y(n_407) );
INVx1_ASAP7_75t_SL g408 ( .A(n_339), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_342), .Y(n_409) );
BUFx3_ASAP7_75t_L g410 ( .A(n_354), .Y(n_410) );
AOI22xp33_ASAP7_75t_L g411 ( .A1(n_369), .A2(n_231), .B1(n_246), .B2(n_245), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_369), .B(n_241), .Y(n_412) );
INVx2_ASAP7_75t_L g413 ( .A(n_352), .Y(n_413) );
INVx1_ASAP7_75t_L g414 ( .A(n_342), .Y(n_414) );
INVx1_ASAP7_75t_L g415 ( .A(n_357), .Y(n_415) );
INVx2_ASAP7_75t_L g416 ( .A(n_352), .Y(n_416) );
AOI22xp5_ASAP7_75t_L g417 ( .A1(n_341), .A2(n_329), .B1(n_218), .B2(n_249), .Y(n_417) );
CKINVDCx20_ASAP7_75t_R g418 ( .A(n_401), .Y(n_418) );
INVx1_ASAP7_75t_L g419 ( .A(n_382), .Y(n_419) );
CKINVDCx20_ASAP7_75t_R g420 ( .A(n_401), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_382), .B(n_358), .Y(n_421) );
INVx2_ASAP7_75t_L g422 ( .A(n_374), .Y(n_422) );
AND2x4_ASAP7_75t_SL g423 ( .A(n_390), .B(n_218), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_376), .Y(n_424) );
NAND2x1p5_ASAP7_75t_L g425 ( .A(n_405), .B(n_329), .Y(n_425) );
HB1xp67_ASAP7_75t_L g426 ( .A(n_394), .Y(n_426) );
AOI22xp5_ASAP7_75t_L g427 ( .A1(n_390), .A2(n_366), .B1(n_358), .B2(n_343), .Y(n_427) );
AND2x4_ASAP7_75t_L g428 ( .A(n_394), .B(n_358), .Y(n_428) );
INVx2_ASAP7_75t_L g429 ( .A(n_376), .Y(n_429) );
OAI22xp5_ASAP7_75t_L g430 ( .A1(n_417), .A2(n_249), .B1(n_250), .B2(n_244), .Y(n_430) );
INVx1_ASAP7_75t_L g431 ( .A(n_407), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_377), .Y(n_432) );
BUFx2_ASAP7_75t_L g433 ( .A(n_371), .Y(n_433) );
OAI22xp33_ASAP7_75t_L g434 ( .A1(n_417), .A2(n_353), .B1(n_346), .B2(n_244), .Y(n_434) );
INVx4_ASAP7_75t_L g435 ( .A(n_380), .Y(n_435) );
AOI22xp5_ASAP7_75t_L g436 ( .A1(n_390), .A2(n_366), .B1(n_356), .B2(n_337), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_407), .Y(n_437) );
NOR2xp33_ASAP7_75t_L g438 ( .A(n_407), .B(n_356), .Y(n_438) );
NOR2xp33_ASAP7_75t_L g439 ( .A(n_391), .B(n_360), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_410), .Y(n_440) );
AOI22xp5_ASAP7_75t_L g441 ( .A1(n_383), .A2(n_353), .B1(n_346), .B2(n_250), .Y(n_441) );
INVx8_ASAP7_75t_L g442 ( .A(n_388), .Y(n_442) );
INVx2_ASAP7_75t_L g443 ( .A(n_380), .Y(n_443) );
INVx2_ASAP7_75t_SL g444 ( .A(n_378), .Y(n_444) );
AO22x1_ASAP7_75t_L g445 ( .A1(n_408), .A2(n_213), .B1(n_296), .B2(n_302), .Y(n_445) );
HB1xp67_ASAP7_75t_L g446 ( .A(n_371), .Y(n_446) );
NAND2xp5_ASAP7_75t_L g447 ( .A(n_387), .B(n_302), .Y(n_447) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_387), .B(n_303), .Y(n_448) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_380), .B(n_357), .Y(n_449) );
BUFx4f_ASAP7_75t_L g450 ( .A(n_405), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_399), .B(n_303), .Y(n_451) );
INVx2_ASAP7_75t_SL g452 ( .A(n_378), .Y(n_452) );
NAND2xp5_ASAP7_75t_SL g453 ( .A(n_380), .B(n_357), .Y(n_453) );
O2A1O1Ixp5_ASAP7_75t_L g454 ( .A1(n_389), .A2(n_234), .B(n_238), .C(n_217), .Y(n_454) );
INVx2_ASAP7_75t_L g455 ( .A(n_377), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g456 ( .A(n_388), .B(n_334), .Y(n_456) );
INVx1_ASAP7_75t_L g457 ( .A(n_373), .Y(n_457) );
BUFx6f_ASAP7_75t_L g458 ( .A(n_388), .Y(n_458) );
AOI22xp33_ASAP7_75t_L g459 ( .A1(n_388), .A2(n_363), .B1(n_365), .B2(n_362), .Y(n_459) );
CKINVDCx5p33_ASAP7_75t_R g460 ( .A(n_404), .Y(n_460) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_388), .B(n_215), .Y(n_461) );
INVx3_ASAP7_75t_L g462 ( .A(n_389), .Y(n_462) );
INVx1_ASAP7_75t_L g463 ( .A(n_373), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g464 ( .A1(n_388), .A2(n_363), .B1(n_365), .B2(n_362), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g465 ( .A(n_389), .B(n_362), .Y(n_465) );
INVx1_ASAP7_75t_L g466 ( .A(n_381), .Y(n_466) );
INVx2_ASAP7_75t_L g467 ( .A(n_379), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_408), .B(n_296), .Y(n_468) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_372), .A2(n_315), .B1(n_301), .B2(n_367), .Y(n_469) );
NAND2xp5_ASAP7_75t_L g470 ( .A(n_372), .B(n_224), .Y(n_470) );
INVx1_ASAP7_75t_L g471 ( .A(n_381), .Y(n_471) );
AOI22xp33_ASAP7_75t_SL g472 ( .A1(n_389), .A2(n_367), .B1(n_257), .B2(n_292), .Y(n_472) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_396), .B(n_259), .Y(n_473) );
AOI21xp5_ASAP7_75t_L g474 ( .A1(n_396), .A2(n_340), .B(n_291), .Y(n_474) );
INVx2_ASAP7_75t_L g475 ( .A(n_379), .Y(n_475) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_396), .B(n_232), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_403), .B(n_262), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_397), .Y(n_478) );
AOI22xp5_ASAP7_75t_L g479 ( .A1(n_403), .A2(n_315), .B1(n_317), .B2(n_267), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_412), .Y(n_480) );
NOR2xp33_ASAP7_75t_L g481 ( .A(n_403), .B(n_235), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_412), .B(n_326), .Y(n_482) );
NOR2xp33_ASAP7_75t_L g483 ( .A(n_400), .B(n_237), .Y(n_483) );
INVx1_ASAP7_75t_L g484 ( .A(n_400), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_386), .B(n_321), .Y(n_485) );
AND2x6_ASAP7_75t_SL g486 ( .A(n_386), .B(n_368), .Y(n_486) );
NAND2xp5_ASAP7_75t_L g487 ( .A(n_393), .B(n_290), .Y(n_487) );
NAND2x1_ASAP7_75t_L g488 ( .A(n_393), .B(n_340), .Y(n_488) );
INVx4_ASAP7_75t_L g489 ( .A(n_406), .Y(n_489) );
AOI21xp5_ASAP7_75t_L g490 ( .A1(n_406), .A2(n_340), .B(n_291), .Y(n_490) );
INVx1_ASAP7_75t_L g491 ( .A(n_463), .Y(n_491) );
OAI22xp5_ASAP7_75t_L g492 ( .A1(n_427), .A2(n_411), .B1(n_313), .B2(n_361), .Y(n_492) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_474), .A2(n_414), .B(n_409), .Y(n_493) );
NOR2xp33_ASAP7_75t_R g494 ( .A(n_418), .B(n_272), .Y(n_494) );
NOR3xp33_ASAP7_75t_SL g495 ( .A(n_434), .B(n_306), .C(n_277), .Y(n_495) );
CKINVDCx14_ASAP7_75t_R g496 ( .A(n_420), .Y(n_496) );
OAI21xp5_ASAP7_75t_L g497 ( .A1(n_490), .A2(n_415), .B(n_414), .Y(n_497) );
AOI21xp5_ASAP7_75t_L g498 ( .A1(n_465), .A2(n_415), .B(n_340), .Y(n_498) );
A2O1A1Ixp33_ASAP7_75t_L g499 ( .A1(n_438), .A2(n_270), .B(n_273), .C(n_268), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_466), .B(n_275), .Y(n_500) );
INVx1_ASAP7_75t_L g501 ( .A(n_471), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g502 ( .A(n_478), .B(n_276), .Y(n_502) );
NOR2x1p5_ASAP7_75t_L g503 ( .A(n_460), .B(n_468), .Y(n_503) );
NAND2xp5_ASAP7_75t_L g504 ( .A(n_480), .B(n_428), .Y(n_504) );
INVx3_ASAP7_75t_L g505 ( .A(n_435), .Y(n_505) );
CKINVDCx11_ASAP7_75t_R g506 ( .A(n_486), .Y(n_506) );
A2O1A1Ixp33_ASAP7_75t_L g507 ( .A1(n_438), .A2(n_282), .B(n_283), .C(n_281), .Y(n_507) );
INVx1_ASAP7_75t_L g508 ( .A(n_431), .Y(n_508) );
INVx1_ASAP7_75t_L g509 ( .A(n_437), .Y(n_509) );
BUFx3_ASAP7_75t_L g510 ( .A(n_450), .Y(n_510) );
OAI22xp5_ASAP7_75t_L g511 ( .A1(n_426), .A2(n_361), .B1(n_292), .B2(n_325), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g512 ( .A1(n_426), .A2(n_319), .B1(n_325), .B2(n_265), .Y(n_512) );
O2A1O1Ixp33_ASAP7_75t_L g513 ( .A1(n_444), .A2(n_295), .B(n_300), .C(n_298), .Y(n_513) );
AND2x4_ASAP7_75t_L g514 ( .A(n_419), .B(n_304), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g515 ( .A1(n_449), .A2(n_384), .B(n_370), .Y(n_515) );
OAI21xp33_ASAP7_75t_SL g516 ( .A1(n_481), .A2(n_332), .B(n_307), .Y(n_516) );
NAND2xp5_ASAP7_75t_L g517 ( .A(n_436), .B(n_216), .Y(n_517) );
AND2x6_ASAP7_75t_L g518 ( .A(n_458), .B(n_288), .Y(n_518) );
A2O1A1Ixp33_ASAP7_75t_L g519 ( .A1(n_481), .A2(n_243), .B(n_248), .C(n_242), .Y(n_519) );
OAI22xp5_ASAP7_75t_L g520 ( .A1(n_442), .A2(n_216), .B1(n_252), .B2(n_251), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_462), .Y(n_521) );
INVx5_ASAP7_75t_L g522 ( .A(n_442), .Y(n_522) );
AOI22xp5_ASAP7_75t_L g523 ( .A1(n_434), .A2(n_255), .B1(n_256), .B2(n_254), .Y(n_523) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_450), .B(n_261), .Y(n_524) );
BUFx8_ASAP7_75t_L g525 ( .A(n_452), .Y(n_525) );
INVx4_ASAP7_75t_L g526 ( .A(n_442), .Y(n_526) );
INVx2_ASAP7_75t_L g527 ( .A(n_443), .Y(n_527) );
O2A1O1Ixp5_ASAP7_75t_L g528 ( .A1(n_488), .A2(n_253), .B(n_294), .C(n_293), .Y(n_528) );
AOI21xp5_ASAP7_75t_L g529 ( .A1(n_449), .A2(n_384), .B(n_370), .Y(n_529) );
AOI22xp5_ASAP7_75t_L g530 ( .A1(n_485), .A2(n_263), .B1(n_271), .B2(n_264), .Y(n_530) );
AOI21xp5_ASAP7_75t_L g531 ( .A1(n_453), .A2(n_392), .B(n_385), .Y(n_531) );
AOI21xp5_ASAP7_75t_L g532 ( .A1(n_453), .A2(n_392), .B(n_385), .Y(n_532) );
BUFx6f_ASAP7_75t_SL g533 ( .A(n_484), .Y(n_533) );
A2O1A1Ixp33_ASAP7_75t_L g534 ( .A1(n_454), .A2(n_278), .B(n_280), .C(n_279), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g535 ( .A(n_439), .B(n_482), .Y(n_535) );
O2A1O1Ixp5_ASAP7_75t_SL g536 ( .A1(n_476), .A2(n_285), .B(n_286), .C(n_284), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_439), .B(n_289), .Y(n_537) );
A2O1A1Ixp33_ASAP7_75t_L g538 ( .A1(n_421), .A2(n_305), .B(n_308), .C(n_299), .Y(n_538) );
OAI22xp5_ASAP7_75t_L g539 ( .A1(n_425), .A2(n_318), .B1(n_322), .B2(n_312), .Y(n_539) );
BUFx2_ASAP7_75t_L g540 ( .A(n_479), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_422), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g542 ( .A(n_447), .B(n_330), .Y(n_542) );
NAND2x1p5_ASAP7_75t_L g543 ( .A(n_469), .B(n_309), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g544 ( .A(n_448), .B(n_309), .Y(n_544) );
BUFx3_ASAP7_75t_L g545 ( .A(n_423), .Y(n_545) );
AOI21xp5_ASAP7_75t_L g546 ( .A1(n_473), .A2(n_413), .B(n_398), .Y(n_546) );
AND2x2_ASAP7_75t_L g547 ( .A(n_441), .B(n_21), .Y(n_547) );
OR2x6_ASAP7_75t_L g548 ( .A(n_445), .B(n_310), .Y(n_548) );
NOR2xp67_ASAP7_75t_L g549 ( .A(n_424), .B(n_79), .Y(n_549) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_477), .A2(n_413), .B(n_398), .Y(n_550) );
AND2x2_ASAP7_75t_SL g551 ( .A(n_472), .B(n_314), .Y(n_551) );
INVx4_ASAP7_75t_L g552 ( .A(n_424), .Y(n_552) );
AOI21x1_ASAP7_75t_L g553 ( .A1(n_456), .A2(n_416), .B(n_347), .Y(n_553) );
NOR2xp33_ASAP7_75t_L g554 ( .A(n_451), .B(n_22), .Y(n_554) );
AND2x4_ASAP7_75t_L g555 ( .A(n_440), .B(n_23), .Y(n_555) );
NOR2xp33_ASAP7_75t_R g556 ( .A(n_470), .B(n_23), .Y(n_556) );
NOR2xp67_ASAP7_75t_SL g557 ( .A(n_461), .B(n_239), .Y(n_557) );
A2O1A1Ixp33_ASAP7_75t_L g558 ( .A1(n_483), .A2(n_239), .B(n_258), .C(n_320), .Y(n_558) );
OAI22xp5_ASAP7_75t_L g559 ( .A1(n_429), .A2(n_328), .B1(n_320), .B2(n_258), .Y(n_559) );
NAND2xp5_ASAP7_75t_L g560 ( .A(n_432), .B(n_25), .Y(n_560) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_455), .B(n_27), .Y(n_561) );
CKINVDCx5p33_ASAP7_75t_R g562 ( .A(n_487), .Y(n_562) );
OAI21x1_ASAP7_75t_L g563 ( .A1(n_459), .A2(n_395), .B(n_375), .Y(n_563) );
INVx4_ASAP7_75t_L g564 ( .A(n_467), .Y(n_564) );
BUFx3_ASAP7_75t_L g565 ( .A(n_475), .Y(n_565) );
INVx2_ASAP7_75t_L g566 ( .A(n_464), .Y(n_566) );
AND2x6_ASAP7_75t_L g567 ( .A(n_464), .B(n_239), .Y(n_567) );
NOR3xp33_ASAP7_75t_L g568 ( .A(n_430), .B(n_29), .C(n_30), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_457), .B(n_31), .Y(n_569) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_446), .A2(n_328), .B1(n_258), .B2(n_352), .Y(n_570) );
AOI21xp5_ASAP7_75t_L g571 ( .A1(n_474), .A2(n_395), .B(n_375), .Y(n_571) );
NAND2xp5_ASAP7_75t_L g572 ( .A(n_457), .B(n_31), .Y(n_572) );
INVx3_ASAP7_75t_L g573 ( .A(n_489), .Y(n_573) );
AOI21xp5_ASAP7_75t_L g574 ( .A1(n_474), .A2(n_395), .B(n_375), .Y(n_574) );
AND2x2_ASAP7_75t_L g575 ( .A(n_433), .B(n_32), .Y(n_575) );
BUFx3_ASAP7_75t_L g576 ( .A(n_418), .Y(n_576) );
A2O1A1Ixp33_ASAP7_75t_L g577 ( .A1(n_438), .A2(n_328), .B(n_352), .C(n_375), .Y(n_577) );
BUFx6f_ASAP7_75t_L g578 ( .A(n_458), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g579 ( .A1(n_474), .A2(n_395), .B(n_352), .Y(n_579) );
AND2x4_ASAP7_75t_L g580 ( .A(n_419), .B(n_32), .Y(n_580) );
A2O1A1Ixp33_ASAP7_75t_L g581 ( .A1(n_438), .A2(n_352), .B(n_395), .C(n_35), .Y(n_581) );
BUFx6f_ASAP7_75t_L g582 ( .A(n_458), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_535), .A2(n_395), .B(n_82), .Y(n_583) );
BUFx8_ASAP7_75t_SL g584 ( .A(n_576), .Y(n_584) );
NOR2xp33_ASAP7_75t_SL g585 ( .A(n_567), .B(n_526), .Y(n_585) );
AND2x2_ASAP7_75t_L g586 ( .A(n_495), .B(n_38), .Y(n_586) );
NOR2xp33_ASAP7_75t_R g587 ( .A(n_496), .B(n_506), .Y(n_587) );
NAND3xp33_ASAP7_75t_L g588 ( .A(n_581), .B(n_41), .C(n_42), .Y(n_588) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_580), .A2(n_42), .B1(n_43), .B2(n_44), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_552), .Y(n_590) );
INVx2_ASAP7_75t_L g591 ( .A(n_552), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_491), .B(n_43), .Y(n_592) );
INVx5_ASAP7_75t_L g593 ( .A(n_518), .Y(n_593) );
INVx1_ASAP7_75t_L g594 ( .A(n_501), .Y(n_594) );
AOI21xp5_ASAP7_75t_L g595 ( .A1(n_498), .A2(n_83), .B(n_80), .Y(n_595) );
AOI21xp5_ASAP7_75t_L g596 ( .A1(n_493), .A2(n_497), .B(n_571), .Y(n_596) );
BUFx6f_ASAP7_75t_L g597 ( .A(n_578), .Y(n_597) );
AOI21xp5_ASAP7_75t_L g598 ( .A1(n_574), .A2(n_85), .B(n_84), .Y(n_598) );
AO31x2_ASAP7_75t_L g599 ( .A1(n_577), .A2(n_44), .A3(n_45), .B(n_46), .Y(n_599) );
O2A1O1Ixp33_ASAP7_75t_L g600 ( .A1(n_516), .A2(n_45), .B(n_46), .C(n_47), .Y(n_600) );
NOR2xp33_ASAP7_75t_L g601 ( .A(n_540), .B(n_47), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g602 ( .A1(n_492), .A2(n_48), .B1(n_50), .B2(n_51), .Y(n_602) );
INVx3_ASAP7_75t_L g603 ( .A(n_564), .Y(n_603) );
NAND2xp5_ASAP7_75t_SL g604 ( .A(n_562), .B(n_48), .Y(n_604) );
O2A1O1Ixp33_ASAP7_75t_L g605 ( .A1(n_516), .A2(n_50), .B(n_52), .C(n_53), .Y(n_605) );
NAND2x1p5_ASAP7_75t_L g606 ( .A(n_510), .B(n_52), .Y(n_606) );
AO21x1_ASAP7_75t_L g607 ( .A1(n_560), .A2(n_89), .B(n_88), .Y(n_607) );
OAI211xp5_ASAP7_75t_SL g608 ( .A1(n_523), .A2(n_54), .B(n_55), .C(n_56), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g609 ( .A(n_504), .B(n_508), .Y(n_609) );
BUFx3_ASAP7_75t_L g610 ( .A(n_525), .Y(n_610) );
NAND2x1p5_ASAP7_75t_L g611 ( .A(n_522), .B(n_545), .Y(n_611) );
INVx3_ASAP7_75t_L g612 ( .A(n_573), .Y(n_612) );
OAI21xp5_ASAP7_75t_L g613 ( .A1(n_528), .A2(n_59), .B(n_60), .Y(n_613) );
INVx2_ASAP7_75t_SL g614 ( .A(n_525), .Y(n_614) );
NOR2x1_ASAP7_75t_R g615 ( .A(n_522), .B(n_60), .Y(n_615) );
AO31x2_ASAP7_75t_L g616 ( .A1(n_558), .A2(n_519), .A3(n_534), .B(n_517), .Y(n_616) );
AOI22xp5_ASAP7_75t_L g617 ( .A1(n_551), .A2(n_61), .B1(n_62), .B2(n_63), .Y(n_617) );
INVx2_ASAP7_75t_L g618 ( .A(n_565), .Y(n_618) );
A2O1A1Ixp33_ASAP7_75t_L g619 ( .A1(n_569), .A2(n_66), .B(n_67), .C(n_68), .Y(n_619) );
NAND2xp5_ASAP7_75t_L g620 ( .A(n_509), .B(n_530), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_572), .Y(n_621) );
BUFx12f_ASAP7_75t_L g622 ( .A(n_503), .Y(n_622) );
AOI21xp5_ASAP7_75t_L g623 ( .A1(n_546), .A2(n_143), .B(n_196), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_580), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_522), .B(n_69), .Y(n_625) );
O2A1O1Ixp33_ASAP7_75t_L g626 ( .A1(n_513), .A2(n_70), .B(n_71), .C(n_72), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g627 ( .A1(n_550), .A2(n_144), .B(n_195), .Y(n_627) );
BUFx2_ASAP7_75t_SL g628 ( .A(n_533), .Y(n_628) );
BUFx10_ASAP7_75t_L g629 ( .A(n_533), .Y(n_629) );
CKINVDCx8_ASAP7_75t_R g630 ( .A(n_555), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_514), .B(n_72), .Y(n_631) );
INVx1_ASAP7_75t_SL g632 ( .A(n_555), .Y(n_632) );
HB1xp67_ASAP7_75t_L g633 ( .A(n_512), .Y(n_633) );
OAI21xp5_ASAP7_75t_L g634 ( .A1(n_566), .A2(n_96), .B(n_97), .Y(n_634) );
INVx2_ASAP7_75t_L g635 ( .A(n_541), .Y(n_635) );
BUFx12f_ASAP7_75t_L g636 ( .A(n_548), .Y(n_636) );
AO31x2_ASAP7_75t_L g637 ( .A1(n_561), .A2(n_99), .A3(n_100), .B(n_101), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_536), .B(n_103), .C(n_104), .Y(n_638) );
AOI21xp5_ASAP7_75t_L g639 ( .A1(n_515), .A2(n_105), .B(n_106), .Y(n_639) );
AND2x4_ASAP7_75t_L g640 ( .A(n_526), .B(n_114), .Y(n_640) );
AOI31xp67_ASAP7_75t_L g641 ( .A1(n_570), .A2(n_544), .A3(n_537), .B(n_542), .Y(n_641) );
BUFx3_ASAP7_75t_L g642 ( .A(n_573), .Y(n_642) );
INVx2_ASAP7_75t_L g643 ( .A(n_527), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_500), .Y(n_644) );
NAND2xp5_ASAP7_75t_L g645 ( .A(n_514), .B(n_117), .Y(n_645) );
BUFx10_ASAP7_75t_L g646 ( .A(n_518), .Y(n_646) );
BUFx3_ASAP7_75t_L g647 ( .A(n_547), .Y(n_647) );
OAI21xp5_ASAP7_75t_L g648 ( .A1(n_529), .A2(n_123), .B(n_124), .Y(n_648) );
HB1xp67_ASAP7_75t_L g649 ( .A(n_575), .Y(n_649) );
AOI22xp33_ASAP7_75t_L g650 ( .A1(n_511), .A2(n_127), .B1(n_131), .B2(n_132), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g651 ( .A1(n_568), .A2(n_133), .B1(n_134), .B2(n_135), .Y(n_651) );
OAI21xp5_ASAP7_75t_L g652 ( .A1(n_531), .A2(n_145), .B(n_146), .Y(n_652) );
AOI21xp5_ASAP7_75t_L g653 ( .A1(n_532), .A2(n_147), .B(n_150), .Y(n_653) );
AO32x2_ASAP7_75t_L g654 ( .A1(n_539), .A2(n_151), .A3(n_153), .B1(n_156), .B2(n_157), .Y(n_654) );
OR2x6_ASAP7_75t_L g655 ( .A(n_543), .B(n_166), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_502), .B(n_168), .Y(n_656) );
BUFx12f_ASAP7_75t_L g657 ( .A(n_518), .Y(n_657) );
OAI21xp5_ASAP7_75t_L g658 ( .A1(n_549), .A2(n_170), .B(n_171), .Y(n_658) );
AND2x2_ASAP7_75t_L g659 ( .A(n_524), .B(n_174), .Y(n_659) );
INVx2_ASAP7_75t_L g660 ( .A(n_505), .Y(n_660) );
OAI21x1_ASAP7_75t_L g661 ( .A1(n_553), .A2(n_180), .B(n_181), .Y(n_661) );
OA21x2_ASAP7_75t_L g662 ( .A1(n_549), .A2(n_192), .B(n_193), .Y(n_662) );
INVx2_ASAP7_75t_L g663 ( .A(n_521), .Y(n_663) );
AO31x2_ASAP7_75t_L g664 ( .A1(n_559), .A2(n_520), .A3(n_567), .B(n_557), .Y(n_664) );
O2A1O1Ixp33_ASAP7_75t_L g665 ( .A1(n_556), .A2(n_567), .B(n_578), .C(n_582), .Y(n_665) );
AOI22xp5_ASAP7_75t_L g666 ( .A1(n_578), .A2(n_551), .B1(n_492), .B2(n_568), .Y(n_666) );
NAND2xp5_ASAP7_75t_L g667 ( .A(n_491), .B(n_402), .Y(n_667) );
OAI21xp5_ASAP7_75t_L g668 ( .A1(n_493), .A2(n_498), .B(n_474), .Y(n_668) );
OAI21x1_ASAP7_75t_L g669 ( .A1(n_579), .A2(n_563), .B(n_571), .Y(n_669) );
INVx2_ASAP7_75t_L g670 ( .A(n_552), .Y(n_670) );
CKINVDCx5p33_ASAP7_75t_R g671 ( .A(n_494), .Y(n_671) );
A2O1A1Ixp33_ASAP7_75t_L g672 ( .A1(n_535), .A2(n_554), .B(n_516), .C(n_438), .Y(n_672) );
O2A1O1Ixp33_ASAP7_75t_L g673 ( .A1(n_499), .A2(n_507), .B(n_516), .C(n_538), .Y(n_673) );
AND2x2_ASAP7_75t_L g674 ( .A(n_495), .B(n_390), .Y(n_674) );
INVx1_ASAP7_75t_L g675 ( .A(n_491), .Y(n_675) );
OA21x2_ASAP7_75t_L g676 ( .A1(n_669), .A2(n_668), .B(n_596), .Y(n_676) );
A2O1A1Ixp33_ASAP7_75t_L g677 ( .A1(n_672), .A2(n_673), .B(n_666), .C(n_617), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g678 ( .A1(n_630), .A2(n_617), .B1(n_632), .B2(n_666), .Y(n_678) );
AND2x4_ASAP7_75t_L g679 ( .A(n_644), .B(n_640), .Y(n_679) );
INVx3_ASAP7_75t_L g680 ( .A(n_603), .Y(n_680) );
CKINVDCx5p33_ASAP7_75t_R g681 ( .A(n_587), .Y(n_681) );
AND2x4_ASAP7_75t_L g682 ( .A(n_640), .B(n_603), .Y(n_682) );
AOI211xp5_ASAP7_75t_L g683 ( .A1(n_589), .A2(n_615), .B(n_601), .C(n_633), .Y(n_683) );
NAND2xp5_ASAP7_75t_L g684 ( .A(n_675), .B(n_609), .Y(n_684) );
INVx1_ASAP7_75t_L g685 ( .A(n_592), .Y(n_685) );
BUFx3_ASAP7_75t_L g686 ( .A(n_584), .Y(n_686) );
OR2x6_ASAP7_75t_L g687 ( .A(n_628), .B(n_614), .Y(n_687) );
AOI21xp33_ASAP7_75t_SL g688 ( .A1(n_606), .A2(n_604), .B(n_611), .Y(n_688) );
NAND2x1p5_ASAP7_75t_L g689 ( .A(n_625), .B(n_593), .Y(n_689) );
NAND2xp5_ASAP7_75t_L g690 ( .A(n_620), .B(n_667), .Y(n_690) );
BUFx12f_ASAP7_75t_L g691 ( .A(n_629), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_631), .Y(n_692) );
INVx2_ASAP7_75t_L g693 ( .A(n_643), .Y(n_693) );
CKINVDCx20_ASAP7_75t_R g694 ( .A(n_671), .Y(n_694) );
NAND2xp5_ASAP7_75t_L g695 ( .A(n_649), .B(n_624), .Y(n_695) );
AOI22xp33_ASAP7_75t_L g696 ( .A1(n_621), .A2(n_622), .B1(n_608), .B2(n_586), .Y(n_696) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_600), .A2(n_605), .B(n_626), .Y(n_697) );
INVx1_ASAP7_75t_L g698 ( .A(n_625), .Y(n_698) );
OAI21xp5_ASAP7_75t_L g699 ( .A1(n_613), .A2(n_588), .B(n_641), .Y(n_699) );
AOI21xp5_ASAP7_75t_L g700 ( .A1(n_656), .A2(n_583), .B(n_595), .Y(n_700) );
INVx4_ASAP7_75t_L g701 ( .A(n_629), .Y(n_701) );
INVx2_ASAP7_75t_L g702 ( .A(n_590), .Y(n_702) );
BUFx6f_ASAP7_75t_L g703 ( .A(n_597), .Y(n_703) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_585), .A2(n_665), .B(n_638), .Y(n_704) );
INVx3_ASAP7_75t_L g705 ( .A(n_657), .Y(n_705) );
OAI21x1_ASAP7_75t_L g706 ( .A1(n_661), .A2(n_658), .B(n_598), .Y(n_706) );
AND2x4_ASAP7_75t_L g707 ( .A(n_655), .B(n_642), .Y(n_707) );
HB1xp67_ASAP7_75t_L g708 ( .A(n_618), .Y(n_708) );
INVx8_ASAP7_75t_L g709 ( .A(n_655), .Y(n_709) );
INVx3_ASAP7_75t_L g710 ( .A(n_646), .Y(n_710) );
INVx2_ASAP7_75t_L g711 ( .A(n_670), .Y(n_711) );
BUFx3_ASAP7_75t_L g712 ( .A(n_636), .Y(n_712) );
AND2x2_ASAP7_75t_L g713 ( .A(n_591), .B(n_663), .Y(n_713) );
AOI21xp5_ASAP7_75t_L g714 ( .A1(n_623), .A2(n_627), .B(n_607), .Y(n_714) );
BUFx5_ASAP7_75t_L g715 ( .A(n_646), .Y(n_715) );
INVx1_ASAP7_75t_L g716 ( .A(n_599), .Y(n_716) );
NAND2xp5_ASAP7_75t_L g717 ( .A(n_616), .B(n_612), .Y(n_717) );
NAND2xp5_ASAP7_75t_L g718 ( .A(n_616), .B(n_659), .Y(n_718) );
OA21x2_ASAP7_75t_L g719 ( .A1(n_634), .A2(n_658), .B(n_652), .Y(n_719) );
OAI22xp5_ASAP7_75t_L g720 ( .A1(n_651), .A2(n_650), .B1(n_593), .B2(n_645), .Y(n_720) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_639), .A2(n_653), .B(n_648), .Y(n_721) );
INVx1_ASAP7_75t_L g722 ( .A(n_619), .Y(n_722) );
INVx2_ASAP7_75t_L g723 ( .A(n_660), .Y(n_723) );
OAI21xp5_ASAP7_75t_L g724 ( .A1(n_662), .A2(n_664), .B(n_654), .Y(n_724) );
OR2x6_ASAP7_75t_L g725 ( .A(n_654), .B(n_664), .Y(n_725) );
AOI21xp5_ASAP7_75t_L g726 ( .A1(n_637), .A2(n_579), .B(n_596), .Y(n_726) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_637), .A2(n_579), .B(n_596), .Y(n_727) );
INVx4_ASAP7_75t_SL g728 ( .A(n_610), .Y(n_728) );
NOR2x1_ASAP7_75t_L g729 ( .A(n_610), .B(n_628), .Y(n_729) );
INVx2_ASAP7_75t_L g730 ( .A(n_635), .Y(n_730) );
A2O1A1Ixp33_ASAP7_75t_L g731 ( .A1(n_672), .A2(n_673), .B(n_666), .C(n_617), .Y(n_731) );
INVx3_ASAP7_75t_L g732 ( .A(n_603), .Y(n_732) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_647), .A2(n_551), .B1(n_674), .B2(n_492), .Y(n_733) );
BUFx8_ASAP7_75t_L g734 ( .A(n_610), .Y(n_734) );
INVx2_ASAP7_75t_L g735 ( .A(n_635), .Y(n_735) );
AOI22xp5_ASAP7_75t_L g736 ( .A1(n_674), .A2(n_434), .B1(n_551), .B2(n_492), .Y(n_736) );
AOI22xp33_ASAP7_75t_L g737 ( .A1(n_647), .A2(n_551), .B1(n_674), .B2(n_492), .Y(n_737) );
AOI22xp33_ASAP7_75t_L g738 ( .A1(n_647), .A2(n_551), .B1(n_674), .B2(n_492), .Y(n_738) );
OR2x6_ASAP7_75t_L g739 ( .A(n_628), .B(n_610), .Y(n_739) );
BUFx6f_ASAP7_75t_L g740 ( .A(n_597), .Y(n_740) );
AND2x4_ASAP7_75t_L g741 ( .A(n_644), .B(n_491), .Y(n_741) );
INVx2_ASAP7_75t_L g742 ( .A(n_635), .Y(n_742) );
INVx1_ASAP7_75t_L g743 ( .A(n_594), .Y(n_743) );
OAI21xp33_ASAP7_75t_L g744 ( .A1(n_672), .A2(n_617), .B(n_602), .Y(n_744) );
NOR2x1_ASAP7_75t_SL g745 ( .A(n_655), .B(n_657), .Y(n_745) );
INVx1_ASAP7_75t_L g746 ( .A(n_594), .Y(n_746) );
INVx2_ASAP7_75t_L g747 ( .A(n_635), .Y(n_747) );
INVx2_ASAP7_75t_L g748 ( .A(n_676), .Y(n_748) );
AND2x2_ASAP7_75t_L g749 ( .A(n_730), .B(n_735), .Y(n_749) );
INVx1_ASAP7_75t_L g750 ( .A(n_717), .Y(n_750) );
BUFx3_ASAP7_75t_L g751 ( .A(n_734), .Y(n_751) );
AO21x2_ASAP7_75t_L g752 ( .A1(n_724), .A2(n_699), .B(n_726), .Y(n_752) );
AO21x2_ASAP7_75t_L g753 ( .A1(n_724), .A2(n_699), .B(n_727), .Y(n_753) );
AND2x2_ASAP7_75t_L g754 ( .A(n_742), .B(n_747), .Y(n_754) );
OR2x2_ASAP7_75t_L g755 ( .A(n_684), .B(n_690), .Y(n_755) );
OAI22xp5_ASAP7_75t_L g756 ( .A1(n_683), .A2(n_709), .B1(n_736), .B2(n_738), .Y(n_756) );
INVx3_ASAP7_75t_L g757 ( .A(n_703), .Y(n_757) );
AND2x2_ASAP7_75t_L g758 ( .A(n_684), .B(n_693), .Y(n_758) );
INVx2_ASAP7_75t_SL g759 ( .A(n_709), .Y(n_759) );
INVx3_ASAP7_75t_L g760 ( .A(n_703), .Y(n_760) );
INVx1_ASAP7_75t_L g761 ( .A(n_717), .Y(n_761) );
INVx1_ASAP7_75t_L g762 ( .A(n_716), .Y(n_762) );
AND2x2_ASAP7_75t_L g763 ( .A(n_679), .B(n_741), .Y(n_763) );
AND2x4_ASAP7_75t_L g764 ( .A(n_682), .B(n_745), .Y(n_764) );
OAI211xp5_ASAP7_75t_L g765 ( .A1(n_733), .A2(n_737), .B(n_696), .C(n_688), .Y(n_765) );
AND2x2_ASAP7_75t_L g766 ( .A(n_743), .B(n_746), .Y(n_766) );
AND2x4_ASAP7_75t_L g767 ( .A(n_707), .B(n_680), .Y(n_767) );
OR2x2_ASAP7_75t_L g768 ( .A(n_678), .B(n_718), .Y(n_768) );
OR2x2_ASAP7_75t_L g769 ( .A(n_678), .B(n_677), .Y(n_769) );
AND2x4_ASAP7_75t_L g770 ( .A(n_680), .B(n_732), .Y(n_770) );
OR2x6_ASAP7_75t_L g771 ( .A(n_689), .B(n_687), .Y(n_771) );
OA21x2_ASAP7_75t_L g772 ( .A1(n_731), .A2(n_706), .B(n_704), .Y(n_772) );
OR2x2_ASAP7_75t_L g773 ( .A(n_695), .B(n_698), .Y(n_773) );
AOI221xp5_ASAP7_75t_L g774 ( .A1(n_744), .A2(n_697), .B1(n_692), .B2(n_685), .C(n_722), .Y(n_774) );
OR2x2_ASAP7_75t_L g775 ( .A(n_725), .B(n_708), .Y(n_775) );
AND2x2_ASAP7_75t_L g776 ( .A(n_713), .B(n_711), .Y(n_776) );
AOI21xp5_ASAP7_75t_SL g777 ( .A1(n_719), .A2(n_720), .B(n_725), .Y(n_777) );
OA21x2_ASAP7_75t_L g778 ( .A1(n_721), .A2(n_700), .B(n_714), .Y(n_778) );
INVx1_ASAP7_75t_L g779 ( .A(n_723), .Y(n_779) );
INVx1_ASAP7_75t_L g780 ( .A(n_702), .Y(n_780) );
OR2x6_ASAP7_75t_L g781 ( .A(n_687), .B(n_739), .Y(n_781) );
BUFx2_ASAP7_75t_L g782 ( .A(n_740), .Y(n_782) );
AND2x4_ASAP7_75t_L g783 ( .A(n_710), .B(n_705), .Y(n_783) );
OR2x6_ASAP7_75t_L g784 ( .A(n_739), .B(n_701), .Y(n_784) );
AND2x2_ASAP7_75t_L g785 ( .A(n_715), .B(n_739), .Y(n_785) );
AOI21xp5_ASAP7_75t_SL g786 ( .A1(n_715), .A2(n_686), .B(n_712), .Y(n_786) );
INVx2_ASAP7_75t_L g787 ( .A(n_715), .Y(n_787) );
AND2x2_ASAP7_75t_L g788 ( .A(n_715), .B(n_729), .Y(n_788) );
INVx1_ASAP7_75t_L g789 ( .A(n_728), .Y(n_789) );
OAI21x1_ASAP7_75t_L g790 ( .A1(n_691), .A2(n_681), .B(n_694), .Y(n_790) );
AND2x2_ASAP7_75t_L g791 ( .A(n_730), .B(n_735), .Y(n_791) );
AO21x2_ASAP7_75t_L g792 ( .A1(n_724), .A2(n_699), .B(n_726), .Y(n_792) );
AND2x2_ASAP7_75t_L g793 ( .A(n_750), .B(n_761), .Y(n_793) );
AND2x2_ASAP7_75t_L g794 ( .A(n_750), .B(n_761), .Y(n_794) );
OAI22xp33_ASAP7_75t_L g795 ( .A1(n_781), .A2(n_756), .B1(n_771), .B2(n_784), .Y(n_795) );
INVx1_ASAP7_75t_L g796 ( .A(n_762), .Y(n_796) );
INVx1_ASAP7_75t_L g797 ( .A(n_762), .Y(n_797) );
CKINVDCx5p33_ASAP7_75t_R g798 ( .A(n_751), .Y(n_798) );
INVx2_ASAP7_75t_L g799 ( .A(n_748), .Y(n_799) );
AND2x2_ASAP7_75t_SL g800 ( .A(n_768), .B(n_769), .Y(n_800) );
NAND2xp5_ASAP7_75t_L g801 ( .A(n_769), .B(n_774), .Y(n_801) );
BUFx2_ASAP7_75t_L g802 ( .A(n_782), .Y(n_802) );
NAND2xp5_ASAP7_75t_L g803 ( .A(n_755), .B(n_758), .Y(n_803) );
NAND2xp5_ASAP7_75t_L g804 ( .A(n_755), .B(n_758), .Y(n_804) );
INVx4_ASAP7_75t_L g805 ( .A(n_781), .Y(n_805) );
INVx4_ASAP7_75t_L g806 ( .A(n_781), .Y(n_806) );
INVx4_ASAP7_75t_L g807 ( .A(n_781), .Y(n_807) );
AND2x2_ASAP7_75t_L g808 ( .A(n_766), .B(n_776), .Y(n_808) );
NOR2x1p5_ASAP7_75t_L g809 ( .A(n_751), .B(n_787), .Y(n_809) );
INVx1_ASAP7_75t_L g810 ( .A(n_775), .Y(n_810) );
AND2x2_ASAP7_75t_SL g811 ( .A(n_777), .B(n_764), .Y(n_811) );
AND2x2_ASAP7_75t_L g812 ( .A(n_752), .B(n_753), .Y(n_812) );
AND2x2_ASAP7_75t_L g813 ( .A(n_753), .B(n_792), .Y(n_813) );
INVx1_ASAP7_75t_L g814 ( .A(n_796), .Y(n_814) );
INVx1_ASAP7_75t_SL g815 ( .A(n_798), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g816 ( .A(n_809), .Y(n_816) );
CKINVDCx14_ASAP7_75t_R g817 ( .A(n_808), .Y(n_817) );
INVx1_ASAP7_75t_L g818 ( .A(n_796), .Y(n_818) );
INVx1_ASAP7_75t_L g819 ( .A(n_797), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_797), .Y(n_820) );
AND2x2_ASAP7_75t_L g821 ( .A(n_793), .B(n_772), .Y(n_821) );
INVx2_ASAP7_75t_SL g822 ( .A(n_809), .Y(n_822) );
OAI21xp5_ASAP7_75t_L g823 ( .A1(n_801), .A2(n_765), .B(n_786), .Y(n_823) );
AND2x2_ASAP7_75t_SL g824 ( .A(n_811), .B(n_764), .Y(n_824) );
INVx2_ASAP7_75t_L g825 ( .A(n_799), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g826 ( .A(n_803), .B(n_791), .Y(n_826) );
INVxp67_ASAP7_75t_L g827 ( .A(n_802), .Y(n_827) );
OR2x2_ASAP7_75t_L g828 ( .A(n_810), .B(n_773), .Y(n_828) );
AND2x4_ASAP7_75t_L g829 ( .A(n_805), .B(n_767), .Y(n_829) );
NAND2xp5_ASAP7_75t_L g830 ( .A(n_803), .B(n_749), .Y(n_830) );
INVx3_ASAP7_75t_L g831 ( .A(n_811), .Y(n_831) );
NAND2xp5_ASAP7_75t_L g832 ( .A(n_804), .B(n_749), .Y(n_832) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_804), .B(n_791), .Y(n_833) );
AND2x2_ASAP7_75t_L g834 ( .A(n_794), .B(n_778), .Y(n_834) );
INVx3_ASAP7_75t_L g835 ( .A(n_831), .Y(n_835) );
INVx1_ASAP7_75t_L g836 ( .A(n_814), .Y(n_836) );
INVx1_ASAP7_75t_L g837 ( .A(n_814), .Y(n_837) );
OR2x6_ASAP7_75t_L g838 ( .A(n_831), .B(n_805), .Y(n_838) );
NOR2xp33_ASAP7_75t_SL g839 ( .A(n_815), .B(n_784), .Y(n_839) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_817), .A2(n_800), .B1(n_795), .B2(n_805), .Y(n_840) );
NAND2x1_ASAP7_75t_L g841 ( .A(n_831), .B(n_806), .Y(n_841) );
AND2x4_ASAP7_75t_SL g842 ( .A(n_829), .B(n_806), .Y(n_842) );
INVx1_ASAP7_75t_L g843 ( .A(n_818), .Y(n_843) );
AND3x2_ASAP7_75t_L g844 ( .A(n_823), .B(n_785), .C(n_789), .Y(n_844) );
AND2x2_ASAP7_75t_L g845 ( .A(n_834), .B(n_812), .Y(n_845) );
INVx1_ASAP7_75t_L g846 ( .A(n_818), .Y(n_846) );
INVx2_ASAP7_75t_L g847 ( .A(n_825), .Y(n_847) );
INVx1_ASAP7_75t_L g848 ( .A(n_819), .Y(n_848) );
INVx1_ASAP7_75t_L g849 ( .A(n_819), .Y(n_849) );
CKINVDCx5p33_ASAP7_75t_R g850 ( .A(n_816), .Y(n_850) );
INVx1_ASAP7_75t_L g851 ( .A(n_820), .Y(n_851) );
AND2x2_ASAP7_75t_L g852 ( .A(n_821), .B(n_813), .Y(n_852) );
INVx1_ASAP7_75t_L g853 ( .A(n_836), .Y(n_853) );
AOI22x1_ASAP7_75t_SL g854 ( .A1(n_850), .A2(n_816), .B1(n_807), .B2(n_806), .Y(n_854) );
CKINVDCx14_ASAP7_75t_R g855 ( .A(n_850), .Y(n_855) );
INVx2_ASAP7_75t_L g856 ( .A(n_847), .Y(n_856) );
INVx2_ASAP7_75t_L g857 ( .A(n_847), .Y(n_857) );
AOI21xp33_ASAP7_75t_SL g858 ( .A1(n_840), .A2(n_824), .B(n_822), .Y(n_858) );
AND2x2_ASAP7_75t_L g859 ( .A(n_852), .B(n_845), .Y(n_859) );
AOI22xp5_ASAP7_75t_L g860 ( .A1(n_839), .A2(n_824), .B1(n_807), .B2(n_806), .Y(n_860) );
INVx1_ASAP7_75t_L g861 ( .A(n_837), .Y(n_861) );
XNOR2x1_ASAP7_75t_L g862 ( .A(n_859), .B(n_790), .Y(n_862) );
INVx1_ASAP7_75t_L g863 ( .A(n_853), .Y(n_863) );
A2O1A1Ixp33_ASAP7_75t_L g864 ( .A1(n_858), .A2(n_842), .B(n_841), .C(n_759), .Y(n_864) );
INVx1_ASAP7_75t_L g865 ( .A(n_853), .Y(n_865) );
INVx1_ASAP7_75t_L g866 ( .A(n_861), .Y(n_866) );
HB1xp67_ASAP7_75t_L g867 ( .A(n_856), .Y(n_867) );
NAND2xp33_ASAP7_75t_L g868 ( .A(n_860), .B(n_835), .Y(n_868) );
INVx1_ASAP7_75t_L g869 ( .A(n_861), .Y(n_869) );
AOI22xp33_ASAP7_75t_SL g870 ( .A1(n_862), .A2(n_854), .B1(n_855), .B2(n_842), .Y(n_870) );
OAI21xp5_ASAP7_75t_SL g871 ( .A1(n_864), .A2(n_844), .B(n_854), .Y(n_871) );
O2A1O1Ixp5_ASAP7_75t_L g872 ( .A1(n_864), .A2(n_807), .B(n_835), .C(n_783), .Y(n_872) );
NOR3xp33_ASAP7_75t_L g873 ( .A(n_868), .B(n_783), .C(n_788), .Y(n_873) );
A2O1A1Ixp33_ASAP7_75t_SL g874 ( .A1(n_868), .A2(n_827), .B(n_757), .C(n_760), .Y(n_874) );
INVx1_ASAP7_75t_L g875 ( .A(n_863), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g876 ( .A1(n_870), .A2(n_869), .B1(n_865), .B2(n_866), .Y(n_876) );
INVx1_ASAP7_75t_L g877 ( .A(n_875), .Y(n_877) );
AOI211xp5_ASAP7_75t_L g878 ( .A1(n_871), .A2(n_785), .B(n_829), .C(n_867), .Y(n_878) );
INVx1_ASAP7_75t_L g879 ( .A(n_877), .Y(n_879) );
NAND4xp25_ASAP7_75t_L g880 ( .A(n_878), .B(n_872), .C(n_874), .D(n_873), .Y(n_880) );
NAND3xp33_ASAP7_75t_L g881 ( .A(n_876), .B(n_783), .C(n_856), .Y(n_881) );
INVx2_ASAP7_75t_L g882 ( .A(n_879), .Y(n_882) );
NAND4xp25_ASAP7_75t_SL g883 ( .A(n_881), .B(n_763), .C(n_828), .D(n_826), .Y(n_883) );
NOR2x1_ASAP7_75t_L g884 ( .A(n_880), .B(n_838), .Y(n_884) );
BUFx2_ASAP7_75t_L g885 ( .A(n_884), .Y(n_885) );
INVx2_ASAP7_75t_L g886 ( .A(n_882), .Y(n_886) );
INVx2_ASAP7_75t_L g887 ( .A(n_886), .Y(n_887) );
OAI22xp5_ASAP7_75t_L g888 ( .A1(n_885), .A2(n_883), .B1(n_857), .B2(n_833), .Y(n_888) );
INVx1_ASAP7_75t_L g889 ( .A(n_887), .Y(n_889) );
INVx1_ASAP7_75t_L g890 ( .A(n_888), .Y(n_890) );
AOI222xp33_ASAP7_75t_L g891 ( .A1(n_889), .A2(n_767), .B1(n_779), .B2(n_780), .C1(n_770), .C2(n_846), .Y(n_891) );
AOI222xp33_ASAP7_75t_L g892 ( .A1(n_890), .A2(n_780), .B1(n_770), .B2(n_849), .C1(n_851), .C2(n_848), .Y(n_892) );
OAI21xp5_ASAP7_75t_L g893 ( .A1(n_891), .A2(n_770), .B(n_754), .Y(n_893) );
OA21x2_ASAP7_75t_L g894 ( .A1(n_893), .A2(n_892), .B(n_843), .Y(n_894) );
AOI21xp33_ASAP7_75t_SL g895 ( .A1(n_894), .A2(n_830), .B(n_832), .Y(n_895) );
endmodule