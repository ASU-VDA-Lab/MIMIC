module fake_netlist_1_10283_n_40 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_40);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_40;
wire n_20;
wire n_38;
wire n_36;
wire n_37;
wire n_34;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_33;
wire n_18;
wire n_32;
wire n_35;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_27;
wire n_21;
wire n_29;
wire n_39;
INVx2_ASAP7_75t_L g12 ( .A(n_4), .Y(n_12) );
NAND2xp5_ASAP7_75t_L g13 ( .A(n_2), .B(n_6), .Y(n_13) );
NAND2xp5_ASAP7_75t_L g14 ( .A(n_6), .B(n_7), .Y(n_14) );
INVx1_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
NAND2xp5_ASAP7_75t_L g16 ( .A(n_4), .B(n_11), .Y(n_16) );
AND2x2_ASAP7_75t_L g17 ( .A(n_3), .B(n_10), .Y(n_17) );
AO21x1_ASAP7_75t_L g18 ( .A1(n_13), .A2(n_0), .B(n_1), .Y(n_18) );
CKINVDCx5p33_ASAP7_75t_R g19 ( .A(n_17), .Y(n_19) );
OAI22xp5_ASAP7_75t_L g20 ( .A1(n_15), .A2(n_0), .B1(n_1), .B2(n_2), .Y(n_20) );
OAI21xp5_ASAP7_75t_L g21 ( .A1(n_15), .A2(n_0), .B(n_3), .Y(n_21) );
INVx1_ASAP7_75t_L g22 ( .A(n_18), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_18), .Y(n_23) );
INVx1_ASAP7_75t_SL g24 ( .A(n_19), .Y(n_24) );
HB1xp67_ASAP7_75t_L g25 ( .A(n_24), .Y(n_25) );
AND2x2_ASAP7_75t_L g26 ( .A(n_22), .B(n_21), .Y(n_26) );
NAND2xp5_ASAP7_75t_L g27 ( .A(n_26), .B(n_23), .Y(n_27) );
AND2x2_ASAP7_75t_L g28 ( .A(n_26), .B(n_23), .Y(n_28) );
INVxp67_ASAP7_75t_L g29 ( .A(n_28), .Y(n_29) );
AND2x2_ASAP7_75t_L g30 ( .A(n_28), .B(n_25), .Y(n_30) );
AOI21xp5_ASAP7_75t_L g31 ( .A1(n_29), .A2(n_27), .B(n_22), .Y(n_31) );
OAI322xp33_ASAP7_75t_L g32 ( .A1(n_29), .A2(n_20), .A3(n_16), .B1(n_14), .B2(n_12), .C1(n_17), .C2(n_21), .Y(n_32) );
O2A1O1Ixp5_ASAP7_75t_L g33 ( .A1(n_30), .A2(n_12), .B(n_7), .C(n_8), .Y(n_33) );
NAND3xp33_ASAP7_75t_L g34 ( .A(n_33), .B(n_30), .C(n_8), .Y(n_34) );
INVx1_ASAP7_75t_L g35 ( .A(n_32), .Y(n_35) );
AND2x2_ASAP7_75t_L g36 ( .A(n_31), .B(n_5), .Y(n_36) );
INVx1_ASAP7_75t_L g37 ( .A(n_36), .Y(n_37) );
OAI21x1_ASAP7_75t_SL g38 ( .A1(n_34), .A2(n_10), .B(n_5), .Y(n_38) );
OAI22xp5_ASAP7_75t_SL g39 ( .A1(n_37), .A2(n_35), .B1(n_36), .B2(n_9), .Y(n_39) );
AOI22xp5_ASAP7_75t_L g40 ( .A1(n_39), .A2(n_9), .B1(n_38), .B2(n_35), .Y(n_40) );
endmodule