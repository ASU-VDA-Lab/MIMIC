module fake_jpeg_18510_n_345 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_345);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_345;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_260;
wire n_199;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

INVx2_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx5_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_0),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_12),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_1),
.Y(n_22)
);

INVx6_ASAP7_75t_L g23 ( 
.A(n_5),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_1),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_4),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_8),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

BUFx8_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_6),
.Y(n_31)
);

CKINVDCx16_ASAP7_75t_R g32 ( 
.A(n_12),
.Y(n_32)
);

INVx2_ASAP7_75t_L g33 ( 
.A(n_8),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

BUFx5_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_11),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_7),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_30),
.Y(n_38)
);

INVx5_ASAP7_75t_SL g57 ( 
.A(n_38),
.Y(n_57)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_20),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_44),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_18),
.Y(n_40)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_18),
.Y(n_41)
);

INVx4_ASAP7_75t_L g55 ( 
.A(n_41),
.Y(n_55)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_19),
.Y(n_42)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_42),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_18),
.Y(n_43)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_43),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_31),
.B(n_36),
.Y(n_44)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_30),
.Y(n_45)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_45),
.Y(n_62)
);

INVx3_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g50 ( 
.A(n_46),
.Y(n_50)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_18),
.Y(n_47)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_47),
.Y(n_51)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_17),
.B(n_1),
.C(n_2),
.Y(n_48)
);

MAJIxp5_ASAP7_75t_L g59 ( 
.A(n_48),
.B(n_32),
.C(n_28),
.Y(n_59)
);

BUFx12_ASAP7_75t_L g49 ( 
.A(n_30),
.Y(n_49)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_49),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_42),
.A2(n_33),
.B1(n_19),
.B2(n_16),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_52),
.A2(n_61),
.B1(n_46),
.B2(n_25),
.Y(n_69)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_45),
.Y(n_53)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_53),
.Y(n_66)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g85 ( 
.A(n_59),
.B(n_38),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_48),
.B(n_33),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g80 ( 
.A(n_60),
.B(n_38),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g61 ( 
.A1(n_42),
.A2(n_33),
.B1(n_16),
.B2(n_25),
.Y(n_61)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_53),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_67),
.Y(n_113)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_62),
.Y(n_68)
);

INVx2_ASAP7_75t_SL g122 ( 
.A(n_68),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_69),
.A2(n_84),
.B1(n_85),
.B2(n_41),
.Y(n_136)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_56),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_71),
.B(n_74),
.Y(n_124)
);

INVx6_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_72),
.A2(n_97),
.B1(n_104),
.B2(n_105),
.Y(n_137)
);

INVx3_ASAP7_75t_L g73 ( 
.A(n_62),
.Y(n_73)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_73),
.Y(n_120)
);

CKINVDCx20_ASAP7_75t_R g74 ( 
.A(n_51),
.Y(n_74)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

INVx6_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

INVx3_ASAP7_75t_L g109 ( 
.A(n_76),
.Y(n_109)
);

INVx3_ASAP7_75t_L g77 ( 
.A(n_63),
.Y(n_77)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_77),
.Y(n_134)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_55),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g111 ( 
.A(n_78),
.Y(n_111)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_63),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_79),
.B(n_89),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_80),
.B(n_103),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g81 ( 
.A(n_51),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_81),
.B(n_87),
.Y(n_130)
);

INVx4_ASAP7_75t_L g82 ( 
.A(n_58),
.Y(n_82)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_82),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_44),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_SL g114 ( 
.A(n_83),
.B(n_99),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_64),
.A2(n_46),
.B1(n_25),
.B2(n_23),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g133 ( 
.A(n_86),
.Y(n_133)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g88 ( 
.A(n_64),
.Y(n_88)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_88),
.Y(n_115)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_65),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_90),
.B(n_91),
.Y(n_119)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_50),
.Y(n_91)
);

HAxp5_ASAP7_75t_SL g92 ( 
.A(n_59),
.B(n_49),
.CON(n_92),
.SN(n_92)
);

OR2x2_ASAP7_75t_SL g121 ( 
.A(n_92),
.B(n_103),
.Y(n_121)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_93),
.B(n_94),
.Y(n_128)
);

INVx3_ASAP7_75t_L g94 ( 
.A(n_57),
.Y(n_94)
);

INVx4_ASAP7_75t_L g95 ( 
.A(n_57),
.Y(n_95)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_95),
.Y(n_116)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_57),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_96),
.B(n_98),
.Y(n_131)
);

INVx11_ASAP7_75t_L g97 ( 
.A(n_52),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_60),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_54),
.B(n_31),
.Y(n_99)
);

BUFx16f_ASAP7_75t_L g100 ( 
.A(n_65),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_100),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_58),
.Y(n_101)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_101),
.Y(n_129)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_53),
.Y(n_102)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_102),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g103 ( 
.A(n_54),
.B(n_38),
.Y(n_103)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_62),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_53),
.Y(n_105)
);

OAI21xp5_ASAP7_75t_L g106 ( 
.A1(n_60),
.A2(n_36),
.B(n_29),
.Y(n_106)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_106),
.B(n_22),
.Y(n_110)
);

OA22x2_ASAP7_75t_L g107 ( 
.A1(n_97),
.A2(n_23),
.B1(n_49),
.B2(n_43),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_107),
.A2(n_136),
.B1(n_24),
.B2(n_35),
.Y(n_162)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_110),
.B(n_26),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_92),
.A2(n_23),
.B1(n_40),
.B2(n_43),
.Y(n_117)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_117),
.A2(n_127),
.B1(n_32),
.B2(n_30),
.Y(n_157)
);

MAJIxp5_ASAP7_75t_L g118 ( 
.A(n_85),
.B(n_38),
.C(n_40),
.Y(n_118)
);

XNOR2xp5_ASAP7_75t_L g145 ( 
.A(n_118),
.B(n_30),
.Y(n_145)
);

OR2x2_ASAP7_75t_L g123 ( 
.A(n_84),
.B(n_49),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g141 ( 
.A1(n_123),
.A2(n_47),
.B(n_82),
.Y(n_141)
);

AOI22xp33_ASAP7_75t_L g125 ( 
.A1(n_70),
.A2(n_17),
.B1(n_37),
.B2(n_34),
.Y(n_125)
);

AOI22xp33_ASAP7_75t_L g156 ( 
.A1(n_125),
.A2(n_27),
.B1(n_37),
.B2(n_20),
.Y(n_156)
);

OAI22xp5_ASAP7_75t_L g127 ( 
.A1(n_72),
.A2(n_17),
.B1(n_47),
.B2(n_41),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_138),
.B(n_95),
.Y(n_140)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_116),
.Y(n_139)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_139),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_140),
.B(n_144),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g186 ( 
.A1(n_141),
.A2(n_151),
.B(n_155),
.Y(n_186)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_116),
.Y(n_142)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_142),
.Y(n_184)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_124),
.Y(n_143)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_143),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_124),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_145),
.B(n_127),
.Y(n_167)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_146),
.Y(n_194)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_112),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_147),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g175 ( 
.A(n_148),
.B(n_114),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_121),
.A2(n_78),
.B1(n_76),
.B2(n_75),
.Y(n_149)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_149),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_135),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g190 ( 
.A(n_150),
.B(n_108),
.Y(n_190)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_121),
.A2(n_22),
.B(n_26),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_131),
.B(n_101),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_160),
.Y(n_174)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_133),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_156),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_136),
.A2(n_66),
.B1(n_73),
.B2(n_88),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_154),
.A2(n_158),
.B1(n_162),
.B2(n_165),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_117),
.A2(n_138),
.B(n_123),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g172 ( 
.A1(n_157),
.A2(n_159),
.B1(n_110),
.B2(n_115),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_137),
.A2(n_27),
.B1(n_21),
.B2(n_29),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g159 ( 
.A1(n_107),
.A2(n_21),
.B1(n_34),
.B2(n_24),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_130),
.B(n_28),
.Y(n_160)
);

INVx8_ASAP7_75t_L g161 ( 
.A(n_109),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_161),
.B(n_111),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_130),
.B(n_100),
.Y(n_163)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_163),
.B(n_164),
.Y(n_187)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_118),
.B(n_28),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_123),
.A2(n_28),
.B1(n_35),
.B2(n_3),
.Y(n_165)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_162),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g168 ( 
.A(n_143),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_168),
.B(n_169),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g169 ( 
.A(n_139),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_172),
.A2(n_188),
.B1(n_189),
.B2(n_196),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_175),
.B(n_147),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_142),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_177),
.B(n_178),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g178 ( 
.A(n_152),
.Y(n_178)
);

BUFx24_ASAP7_75t_SL g179 ( 
.A(n_148),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_179),
.B(n_193),
.Y(n_212)
);

CKINVDCx14_ASAP7_75t_R g181 ( 
.A(n_163),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_181),
.B(n_195),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_151),
.A2(n_107),
.B1(n_132),
.B2(n_110),
.Y(n_182)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_182),
.A2(n_159),
.B(n_158),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_145),
.B(n_114),
.C(n_119),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_183),
.B(n_165),
.C(n_157),
.Y(n_204)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_185),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g188 ( 
.A1(n_155),
.A2(n_107),
.B1(n_115),
.B2(n_129),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g189 ( 
.A1(n_164),
.A2(n_129),
.B1(n_108),
.B2(n_135),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_190),
.B(n_197),
.Y(n_206)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_144),
.A2(n_126),
.B(n_133),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g213 ( 
.A1(n_192),
.A2(n_134),
.B(n_120),
.Y(n_213)
);

INVxp33_ASAP7_75t_L g193 ( 
.A(n_160),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_146),
.B(n_109),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_141),
.A2(n_134),
.B1(n_122),
.B2(n_120),
.Y(n_196)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_140),
.B(n_113),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_197),
.Y(n_198)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

XOR2xp5_ASAP7_75t_L g238 ( 
.A(n_200),
.B(n_225),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_201),
.B(n_207),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_186),
.A2(n_150),
.B1(n_154),
.B2(n_132),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g249 ( 
.A1(n_203),
.A2(n_227),
.B1(n_216),
.B2(n_213),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_204),
.B(n_223),
.C(n_167),
.Y(n_229)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_171),
.Y(n_205)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_205),
.Y(n_251)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_171),
.Y(n_207)
);

OAI21xp5_ASAP7_75t_L g237 ( 
.A1(n_208),
.A2(n_209),
.B(n_213),
.Y(n_237)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_170),
.A2(n_153),
.B(n_126),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_173),
.B(n_156),
.Y(n_210)
);

CKINVDCx16_ASAP7_75t_R g248 ( 
.A(n_210),
.Y(n_248)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_184),
.Y(n_214)
);

INVx1_ASAP7_75t_SL g253 ( 
.A(n_214),
.Y(n_253)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_184),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g230 ( 
.A(n_215),
.Y(n_230)
);

AOI21xp5_ASAP7_75t_L g216 ( 
.A1(n_170),
.A2(n_153),
.B(n_161),
.Y(n_216)
);

OAI21xp5_ASAP7_75t_L g252 ( 
.A1(n_216),
.A2(n_86),
.B(n_175),
.Y(n_252)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_191),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g235 ( 
.A(n_217),
.Y(n_235)
);

BUFx2_ASAP7_75t_L g218 ( 
.A(n_196),
.Y(n_218)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_218),
.Y(n_242)
);

OA21x2_ASAP7_75t_L g219 ( 
.A1(n_180),
.A2(n_161),
.B(n_122),
.Y(n_219)
);

OA21x2_ASAP7_75t_L g233 ( 
.A1(n_219),
.A2(n_192),
.B(n_174),
.Y(n_233)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_191),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_220),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g221 ( 
.A(n_194),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g244 ( 
.A(n_221),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_183),
.B(n_113),
.C(n_111),
.Y(n_223)
);

CKINVDCx20_ASAP7_75t_R g224 ( 
.A(n_194),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_224),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g225 ( 
.A(n_186),
.B(n_122),
.Y(n_225)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_188),
.B(n_113),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_L g246 ( 
.A1(n_226),
.A2(n_177),
.B(n_169),
.Y(n_246)
);

NAND2xp33_ASAP7_75t_R g227 ( 
.A(n_182),
.B(n_35),
.Y(n_227)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_229),
.B(n_240),
.Y(n_255)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_223),
.B(n_187),
.C(n_189),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_231),
.B(n_247),
.Y(n_270)
);

XNOR2x2_ASAP7_75t_L g232 ( 
.A(n_225),
.B(n_178),
.Y(n_232)
);

OAI21xp33_ASAP7_75t_L g267 ( 
.A1(n_232),
.A2(n_209),
.B(n_219),
.Y(n_267)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_233),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g239 ( 
.A1(n_226),
.A2(n_172),
.B1(n_187),
.B2(n_176),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g265 ( 
.A1(n_239),
.A2(n_252),
.B1(n_206),
.B2(n_220),
.Y(n_265)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_200),
.B(n_174),
.Y(n_240)
);

HB1xp67_ASAP7_75t_L g241 ( 
.A(n_203),
.Y(n_241)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_241),
.Y(n_259)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_204),
.B(n_176),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g261 ( 
.A(n_245),
.B(n_249),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_246),
.Y(n_262)
);

MAJIxp5_ASAP7_75t_L g247 ( 
.A(n_222),
.B(n_168),
.C(n_166),
.Y(n_247)
);

XOR2xp5_ASAP7_75t_L g250 ( 
.A(n_222),
.B(n_166),
.Y(n_250)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_250),
.B(n_228),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_242),
.A2(n_226),
.B1(n_198),
.B2(n_218),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_257),
.A2(n_264),
.B1(n_253),
.B2(n_9),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g258 ( 
.A(n_254),
.B(n_210),
.Y(n_258)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_258),
.Y(n_281)
);

OA21x2_ASAP7_75t_SL g260 ( 
.A1(n_232),
.A2(n_211),
.B(n_212),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_SL g277 ( 
.A(n_260),
.B(n_273),
.Y(n_277)
);

INVxp67_ASAP7_75t_SL g263 ( 
.A(n_244),
.Y(n_263)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_263),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_242),
.A2(n_202),
.B1(n_206),
.B2(n_208),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_265),
.A2(n_266),
.B1(n_233),
.B2(n_250),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_239),
.A2(n_217),
.B1(n_199),
.B2(n_228),
.Y(n_266)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_267),
.B(n_268),
.Y(n_278)
);

OAI21xp33_ASAP7_75t_L g269 ( 
.A1(n_234),
.A2(n_215),
.B(n_214),
.Y(n_269)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_269),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_243),
.B(n_205),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_271),
.B(n_272),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_243),
.B(n_219),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g273 ( 
.A(n_230),
.B(n_7),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_251),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_274),
.B(n_275),
.Y(n_286)
);

CKINVDCx5p33_ASAP7_75t_R g275 ( 
.A(n_235),
.Y(n_275)
);

BUFx24_ASAP7_75t_SL g276 ( 
.A(n_255),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_276),
.B(n_266),
.Y(n_300)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_259),
.A2(n_247),
.B1(n_248),
.B2(n_233),
.Y(n_280)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_280),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_282),
.A2(n_267),
.B1(n_265),
.B2(n_269),
.Y(n_301)
);

AOI21xp5_ASAP7_75t_L g283 ( 
.A1(n_256),
.A2(n_237),
.B(n_246),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_SL g303 ( 
.A(n_283),
.B(n_291),
.Y(n_303)
);

OAI22xp5_ASAP7_75t_L g285 ( 
.A1(n_264),
.A2(n_237),
.B1(n_236),
.B2(n_252),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_9),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_255),
.B(n_229),
.C(n_231),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_288),
.B(n_289),
.C(n_292),
.Y(n_295)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_270),
.B(n_245),
.C(n_238),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_SL g290 ( 
.A(n_268),
.B(n_238),
.Y(n_290)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_290),
.B(n_289),
.Y(n_298)
);

INVx4_ASAP7_75t_L g291 ( 
.A(n_275),
.Y(n_291)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_291),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g292 ( 
.A(n_261),
.B(n_240),
.C(n_253),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g305 ( 
.A(n_293),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g294 ( 
.A(n_286),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_294),
.A2(n_296),
.B1(n_281),
.B2(n_279),
.Y(n_311)
);

CKINVDCx20_ASAP7_75t_R g296 ( 
.A(n_286),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_L g297 ( 
.A(n_288),
.B(n_261),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g309 ( 
.A(n_297),
.B(n_300),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g310 ( 
.A(n_298),
.B(n_301),
.Y(n_310)
);

AOI21xp5_ASAP7_75t_L g299 ( 
.A1(n_287),
.A2(n_262),
.B(n_257),
.Y(n_299)
);

CKINVDCx16_ASAP7_75t_R g314 ( 
.A(n_299),
.Y(n_314)
);

FAx1_ASAP7_75t_SL g302 ( 
.A(n_278),
.B(n_9),
.CI(n_14),
.CON(n_302),
.SN(n_302)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_302),
.B(n_306),
.Y(n_318)
);

XOR2xp5_ASAP7_75t_L g315 ( 
.A(n_303),
.B(n_304),
.Y(n_315)
);

FAx1_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_1),
.CI(n_2),
.CON(n_304),
.SN(n_304)
);

OAI321xp33_ASAP7_75t_L g317 ( 
.A1(n_306),
.A2(n_283),
.A3(n_277),
.B1(n_12),
.B2(n_15),
.C(n_6),
.Y(n_317)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_311),
.Y(n_322)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_292),
.C(n_290),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g325 ( 
.A(n_312),
.B(n_313),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_295),
.B(n_297),
.C(n_298),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_307),
.B(n_293),
.C(n_278),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g328 ( 
.A(n_316),
.B(n_318),
.Y(n_328)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_317),
.Y(n_324)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_301),
.C(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_319),
.B(n_304),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_310),
.B(n_308),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g332 ( 
.A(n_320),
.B(n_314),
.Y(n_332)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_310),
.B(n_316),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_321),
.B(n_327),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_323),
.B(n_315),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g326 ( 
.A(n_315),
.B(n_284),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g329 ( 
.A(n_326),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_SL g327 ( 
.A1(n_319),
.A2(n_305),
.B1(n_304),
.B2(n_302),
.Y(n_327)
);

CKINVDCx14_ASAP7_75t_R g330 ( 
.A(n_328),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g335 ( 
.A(n_330),
.B(n_332),
.Y(n_335)
);

AOI21xp5_ASAP7_75t_L g336 ( 
.A1(n_331),
.A2(n_334),
.B(n_321),
.Y(n_336)
);

NOR2xp33_ASAP7_75t_L g334 ( 
.A(n_324),
.B(n_309),
.Y(n_334)
);

NAND4xp25_ASAP7_75t_L g338 ( 
.A(n_336),
.B(n_337),
.C(n_329),
.D(n_325),
.Y(n_338)
);

XOR2xp5_ASAP7_75t_L g337 ( 
.A(n_333),
.B(n_320),
.Y(n_337)
);

OAI321xp33_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_331),
.A3(n_335),
.B1(n_322),
.B2(n_302),
.C(n_10),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g340 ( 
.A1(n_339),
.A2(n_10),
.B1(n_14),
.B2(n_13),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

A2O1A1Ixp33_ASAP7_75t_SL g342 ( 
.A1(n_341),
.A2(n_10),
.B(n_14),
.C(n_13),
.Y(n_342)
);

BUFx24_ASAP7_75t_SL g343 ( 
.A(n_342),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g344 ( 
.A(n_343),
.B(n_15),
.C(n_3),
.Y(n_344)
);

AOI21xp5_ASAP7_75t_L g345 ( 
.A1(n_344),
.A2(n_15),
.B(n_3),
.Y(n_345)
);


endmodule