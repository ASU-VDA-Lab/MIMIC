module fake_jpeg_830_n_54 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_7, n_54);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;
input n_7;

output n_54;

wire n_13;
wire n_21;
wire n_53;
wire n_33;
wire n_45;
wire n_10;
wire n_23;
wire n_27;
wire n_22;
wire n_47;
wire n_51;
wire n_14;
wire n_40;
wire n_19;
wire n_18;
wire n_20;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_37;
wire n_50;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;

BUFx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

NAND2xp5_ASAP7_75t_SL g9 ( 
.A(n_3),
.B(n_5),
.Y(n_9)
);

INVx4_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_4),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g12 ( 
.A(n_0),
.B(n_2),
.Y(n_12)
);

BUFx16f_ASAP7_75t_L g13 ( 
.A(n_3),
.Y(n_13)
);

NOR2xp33_ASAP7_75t_L g14 ( 
.A(n_1),
.B(n_0),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_6),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_15),
.Y(n_18)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_18),
.Y(n_35)
);

INVx5_ASAP7_75t_L g19 ( 
.A(n_10),
.Y(n_19)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_19),
.Y(n_30)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_15),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_20),
.B(n_22),
.Y(n_32)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_21),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_12),
.B(n_4),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_14),
.B(n_1),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_23),
.A2(n_24),
.B(n_27),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g24 ( 
.A(n_16),
.B(n_1),
.Y(n_24)
);

AOI22xp33_ASAP7_75t_L g25 ( 
.A1(n_16),
.A2(n_17),
.B1(n_10),
.B2(n_11),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_25),
.A2(n_8),
.B1(n_9),
.B2(n_7),
.Y(n_29)
);

OAI22xp5_ASAP7_75t_SL g26 ( 
.A1(n_17),
.A2(n_6),
.B1(n_7),
.B2(n_11),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g34 ( 
.A1(n_26),
.A2(n_28),
.B1(n_19),
.B2(n_24),
.Y(n_34)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_13),
.Y(n_28)
);

NAND2xp33_ASAP7_75t_R g37 ( 
.A(n_29),
.B(n_34),
.Y(n_37)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_22),
.B(n_8),
.Y(n_31)
);

AND2x6_ASAP7_75t_L g39 ( 
.A(n_31),
.B(n_26),
.Y(n_39)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_35),
.Y(n_38)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_38),
.B(n_39),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_32),
.B(n_23),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_40),
.B(n_36),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g47 ( 
.A(n_41),
.B(n_33),
.Y(n_47)
);

XOR2x2_ASAP7_75t_L g42 ( 
.A(n_39),
.B(n_36),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_42),
.B(n_44),
.C(n_31),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_34),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_45),
.B(n_46),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g46 ( 
.A1(n_44),
.A2(n_20),
.B1(n_35),
.B2(n_18),
.Y(n_46)
);

NOR5xp2_ASAP7_75t_L g49 ( 
.A(n_47),
.B(n_42),
.C(n_28),
.D(n_30),
.E(n_21),
.Y(n_49)
);

CKINVDCx5p33_ASAP7_75t_R g51 ( 
.A(n_49),
.Y(n_51)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_48),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g52 ( 
.A1(n_50),
.A2(n_43),
.B1(n_45),
.B2(n_30),
.Y(n_52)
);

HB1xp67_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

XNOR2xp5_ASAP7_75t_L g54 ( 
.A(n_53),
.B(n_51),
.Y(n_54)
);


endmodule