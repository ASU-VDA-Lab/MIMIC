module fake_jpeg_133_n_408 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_408);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_408;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_370;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_3),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_1),
.Y(n_20)
);

BUFx12_ASAP7_75t_L g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_15),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_6),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_2),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_12),
.Y(n_26)
);

INVx6_ASAP7_75t_SL g27 ( 
.A(n_0),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx8_ASAP7_75t_L g29 ( 
.A(n_7),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_11),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx5_ASAP7_75t_L g34 ( 
.A(n_7),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_9),
.B(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_2),
.Y(n_39)
);

INVx4_ASAP7_75t_L g40 ( 
.A(n_0),
.Y(n_40)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx10_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_9),
.Y(n_43)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_7),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_13),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_2),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_5),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_4),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_11),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_0),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_4),
.Y(n_51)
);

INVx4_ASAP7_75t_L g52 ( 
.A(n_5),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_17),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_53),
.Y(n_121)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_17),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_54),
.Y(n_140)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_27),
.Y(n_55)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_55),
.Y(n_116)
);

INVx8_ASAP7_75t_L g56 ( 
.A(n_27),
.Y(n_56)
);

INVx5_ASAP7_75t_L g138 ( 
.A(n_56),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g57 ( 
.A1(n_37),
.A2(n_16),
.B1(n_15),
.B2(n_14),
.Y(n_57)
);

OAI22xp5_ASAP7_75t_SL g139 ( 
.A1(n_57),
.A2(n_47),
.B1(n_48),
.B2(n_30),
.Y(n_139)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_40),
.Y(n_58)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_58),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_37),
.B(n_15),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_59),
.B(n_66),
.Y(n_115)
);

INVx5_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g141 ( 
.A(n_60),
.Y(n_141)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_23),
.Y(n_61)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_40),
.Y(n_62)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_62),
.Y(n_135)
);

INVx4_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

INVx2_ASAP7_75t_SL g161 ( 
.A(n_63),
.Y(n_161)
);

INVx5_ASAP7_75t_L g64 ( 
.A(n_23),
.Y(n_64)
);

INVx4_ASAP7_75t_L g153 ( 
.A(n_64),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g65 ( 
.A(n_29),
.Y(n_65)
);

INVx4_ASAP7_75t_SL g136 ( 
.A(n_65),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g66 ( 
.A(n_22),
.B(n_16),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g169 ( 
.A(n_67),
.Y(n_169)
);

HB1xp67_ASAP7_75t_L g68 ( 
.A(n_52),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_29),
.Y(n_69)
);

INVx3_ASAP7_75t_L g134 ( 
.A(n_69),
.Y(n_134)
);

BUFx5_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

INVx5_ASAP7_75t_SL g126 ( 
.A(n_70),
.Y(n_126)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_23),
.Y(n_71)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_71),
.Y(n_177)
);

INVx11_ASAP7_75t_L g72 ( 
.A(n_29),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g152 ( 
.A(n_72),
.Y(n_152)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_17),
.Y(n_73)
);

INVx6_ASAP7_75t_L g147 ( 
.A(n_73),
.Y(n_147)
);

BUFx3_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

HB1xp67_ASAP7_75t_L g178 ( 
.A(n_74),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_22),
.B(n_38),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_75),
.B(n_76),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_25),
.B(n_14),
.Y(n_76)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_32),
.Y(n_77)
);

INVx8_ASAP7_75t_L g155 ( 
.A(n_77),
.Y(n_155)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_32),
.Y(n_78)
);

INVx8_ASAP7_75t_L g170 ( 
.A(n_78),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_19),
.B(n_1),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_79),
.B(n_80),
.Y(n_124)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_19),
.Y(n_80)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_52),
.Y(n_81)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_81),
.Y(n_137)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_29),
.Y(n_82)
);

CKINVDCx14_ASAP7_75t_R g131 ( 
.A(n_82),
.Y(n_131)
);

INVx8_ASAP7_75t_L g83 ( 
.A(n_32),
.Y(n_83)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_83),
.Y(n_145)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_19),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_84),
.B(n_85),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_3),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_52),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_86)
);

OR2x2_ASAP7_75t_L g122 ( 
.A(n_86),
.B(n_88),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_26),
.B(n_4),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_87),
.B(n_97),
.Y(n_142)
);

INVx13_ASAP7_75t_L g88 ( 
.A(n_42),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g89 ( 
.A1(n_44),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_107),
.B1(n_33),
.B2(n_31),
.Y(n_111)
);

AOI21xp5_ASAP7_75t_L g90 ( 
.A1(n_26),
.A2(n_8),
.B(n_9),
.Y(n_90)
);

OAI21xp5_ASAP7_75t_L g130 ( 
.A1(n_90),
.A2(n_50),
.B(n_39),
.Y(n_130)
);

BUFx3_ASAP7_75t_L g91 ( 
.A(n_44),
.Y(n_91)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_91),
.Y(n_180)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_92),
.Y(n_128)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_51),
.Y(n_93)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_93),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_51),
.Y(n_94)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_94),
.Y(n_168)
);

INVx8_ASAP7_75t_L g95 ( 
.A(n_51),
.Y(n_95)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_95),
.Y(n_175)
);

BUFx4f_ASAP7_75t_L g96 ( 
.A(n_42),
.Y(n_96)
);

AND2x2_ASAP7_75t_L g148 ( 
.A(n_96),
.B(n_98),
.Y(n_148)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_18),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_51),
.Y(n_98)
);

INVx11_ASAP7_75t_L g99 ( 
.A(n_42),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g171 ( 
.A(n_99),
.B(n_103),
.Y(n_171)
);

INVx6_ASAP7_75t_L g100 ( 
.A(n_46),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_100),
.B(n_101),
.Y(n_172)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_46),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_35),
.B(n_8),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_102),
.B(n_104),
.Y(n_144)
);

INVx4_ASAP7_75t_L g103 ( 
.A(n_34),
.Y(n_103)
);

INVx8_ASAP7_75t_L g104 ( 
.A(n_42),
.Y(n_104)
);

INVx2_ASAP7_75t_L g105 ( 
.A(n_46),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g157 ( 
.A(n_105),
.B(n_110),
.Y(n_157)
);

INVx5_ASAP7_75t_L g106 ( 
.A(n_42),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_106),
.B(n_108),
.Y(n_146)
);

INVx11_ASAP7_75t_L g107 ( 
.A(n_42),
.Y(n_107)
);

BUFx12_ASAP7_75t_L g108 ( 
.A(n_21),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_35),
.B(n_8),
.Y(n_109)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_109),
.B(n_9),
.Y(n_150)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_18),
.Y(n_110)
);

OAI21xp33_ASAP7_75t_L g182 ( 
.A1(n_111),
.A2(n_150),
.B(n_108),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_65),
.B(n_50),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_SL g201 ( 
.A(n_112),
.B(n_158),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_89),
.A2(n_33),
.B1(n_31),
.B2(n_28),
.Y(n_113)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_113),
.A2(n_119),
.B1(n_123),
.B2(n_129),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_72),
.A2(n_28),
.B1(n_33),
.B2(n_31),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g191 ( 
.A1(n_117),
.A2(n_132),
.B1(n_143),
.B2(n_149),
.Y(n_191)
);

AOI22xp33_ASAP7_75t_L g119 ( 
.A1(n_53),
.A2(n_39),
.B1(n_38),
.B2(n_47),
.Y(n_119)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_63),
.B(n_45),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_120),
.B(n_159),
.Y(n_186)
);

AOI22xp5_ASAP7_75t_L g123 ( 
.A1(n_54),
.A2(n_24),
.B1(n_49),
.B2(n_48),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_24),
.B1(n_49),
.B2(n_48),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g216 ( 
.A1(n_130),
.A2(n_125),
.B(n_122),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_82),
.A2(n_28),
.B1(n_49),
.B2(n_30),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_139),
.A2(n_166),
.B1(n_113),
.B2(n_133),
.Y(n_198)
);

AOI22xp33_ASAP7_75t_SL g143 ( 
.A1(n_82),
.A2(n_24),
.B1(n_43),
.B2(n_41),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_69),
.A2(n_45),
.B1(n_43),
.B2(n_41),
.Y(n_149)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_103),
.A2(n_20),
.B1(n_41),
.B2(n_45),
.Y(n_151)
);

AOI22xp33_ASAP7_75t_SL g199 ( 
.A1(n_151),
.A2(n_154),
.B1(n_162),
.B2(n_174),
.Y(n_199)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_96),
.A2(n_43),
.B1(n_36),
.B2(n_18),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_60),
.B(n_36),
.Y(n_156)
);

INVxp67_ASAP7_75t_L g230 ( 
.A(n_156),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_SL g158 ( 
.A(n_61),
.B(n_36),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_73),
.B(n_20),
.Y(n_159)
);

NOR2xp33_ASAP7_75t_SL g160 ( 
.A(n_74),
.B(n_20),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_SL g210 ( 
.A(n_160),
.B(n_142),
.Y(n_210)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_64),
.A2(n_30),
.B1(n_34),
.B2(n_21),
.Y(n_162)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_77),
.A2(n_34),
.B1(n_21),
.B2(n_13),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_163),
.A2(n_165),
.B1(n_166),
.B2(n_173),
.Y(n_214)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_56),
.B(n_10),
.Y(n_164)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_164),
.B(n_176),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g165 ( 
.A1(n_78),
.A2(n_10),
.B1(n_11),
.B2(n_13),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_92),
.A2(n_21),
.B1(n_10),
.B2(n_13),
.Y(n_166)
);

AOI22xp5_ASAP7_75t_L g173 ( 
.A1(n_93),
.A2(n_10),
.B1(n_21),
.B2(n_98),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g174 ( 
.A1(n_91),
.A2(n_99),
.B1(n_107),
.B2(n_106),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_100),
.B(n_104),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g179 ( 
.A1(n_83),
.A2(n_95),
.B1(n_94),
.B2(n_88),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_SL g204 ( 
.A1(n_179),
.A2(n_148),
.B1(n_134),
.B2(n_172),
.Y(n_204)
);

CKINVDCx14_ASAP7_75t_R g261 ( 
.A(n_182),
.Y(n_261)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_161),
.Y(n_183)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_183),
.Y(n_252)
);

INVx3_ASAP7_75t_L g184 ( 
.A(n_153),
.Y(n_184)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_122),
.A2(n_108),
.B1(n_159),
.B2(n_157),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_185),
.A2(n_196),
.B1(n_198),
.B2(n_209),
.Y(n_240)
);

CKINVDCx20_ASAP7_75t_R g187 ( 
.A(n_118),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g264 ( 
.A(n_187),
.B(n_190),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g188 ( 
.A(n_136),
.Y(n_188)
);

HB1xp67_ASAP7_75t_L g263 ( 
.A(n_188),
.Y(n_263)
);

NAND2xp5_ASAP7_75t_SL g189 ( 
.A(n_120),
.B(n_124),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_189),
.B(n_215),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_112),
.Y(n_190)
);

INVx4_ASAP7_75t_L g192 ( 
.A(n_161),
.Y(n_192)
);

BUFx6f_ASAP7_75t_L g244 ( 
.A(n_192),
.Y(n_244)
);

CKINVDCx16_ASAP7_75t_R g193 ( 
.A(n_171),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g270 ( 
.A(n_193),
.B(n_208),
.Y(n_270)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_136),
.Y(n_194)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_194),
.Y(n_243)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_136),
.Y(n_195)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_195),
.Y(n_253)
);

OAI22xp33_ASAP7_75t_L g196 ( 
.A1(n_123),
.A2(n_129),
.B1(n_165),
.B2(n_173),
.Y(n_196)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_153),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g275 ( 
.A(n_200),
.Y(n_275)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_161),
.Y(n_202)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_202),
.Y(n_256)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_138),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_210),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_204),
.A2(n_206),
.B1(n_211),
.B2(n_221),
.Y(n_246)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_130),
.A2(n_157),
.B1(n_168),
.B2(n_167),
.Y(n_205)
);

OAI22xp5_ASAP7_75t_L g254 ( 
.A1(n_205),
.A2(n_222),
.B1(n_228),
.B2(n_233),
.Y(n_254)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_144),
.A2(n_134),
.B1(n_139),
.B2(n_177),
.Y(n_206)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_115),
.B(n_172),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_207),
.B(n_189),
.C(n_230),
.Y(n_250)
);

AO22x1_ASAP7_75t_L g208 ( 
.A1(n_172),
.A2(n_122),
.B1(n_148),
.B2(n_135),
.Y(n_208)
);

OAI22xp33_ASAP7_75t_L g209 ( 
.A1(n_128),
.A2(n_168),
.B1(n_167),
.B2(n_137),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g211 ( 
.A1(n_177),
.A2(n_178),
.B1(n_116),
.B2(n_137),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g212 ( 
.A(n_138),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g248 ( 
.A(n_212),
.B(n_227),
.Y(n_248)
);

INVx6_ASAP7_75t_L g213 ( 
.A(n_121),
.Y(n_213)
);

BUFx6f_ASAP7_75t_L g257 ( 
.A(n_213),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_158),
.B(n_160),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g268 ( 
.A(n_216),
.B(n_217),
.Y(n_268)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_148),
.Y(n_217)
);

OR2x2_ASAP7_75t_L g218 ( 
.A(n_126),
.B(n_116),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_218),
.B(n_219),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_171),
.B(n_114),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_171),
.A2(n_128),
.B1(n_147),
.B2(n_114),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_220),
.A2(n_223),
.B1(n_224),
.B2(n_226),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g221 ( 
.A1(n_127),
.A2(n_180),
.B1(n_145),
.B2(n_141),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_147),
.A2(n_121),
.B1(n_169),
.B2(n_140),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_135),
.A2(n_121),
.B1(n_169),
.B2(n_140),
.Y(n_223)
);

AOI22xp33_ASAP7_75t_SL g224 ( 
.A1(n_127),
.A2(n_180),
.B1(n_145),
.B2(n_141),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_146),
.B(n_175),
.Y(n_225)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_225),
.B(n_234),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g226 ( 
.A1(n_140),
.A2(n_169),
.B1(n_155),
.B2(n_170),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g227 ( 
.A(n_131),
.Y(n_227)
);

OAI22xp5_ASAP7_75t_L g228 ( 
.A1(n_155),
.A2(n_170),
.B1(n_175),
.B2(n_152),
.Y(n_228)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_152),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_229),
.B(n_231),
.Y(n_260)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_126),
.Y(n_231)
);

INVx2_ASAP7_75t_L g232 ( 
.A(n_161),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_232),
.B(n_236),
.Y(n_272)
);

AOI22xp33_ASAP7_75t_L g233 ( 
.A1(n_113),
.A2(n_120),
.B1(n_130),
.B2(n_159),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_157),
.B(n_120),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_122),
.A2(n_159),
.B1(n_157),
.B2(n_165),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_L g258 ( 
.A1(n_235),
.A2(n_238),
.B1(n_199),
.B2(n_218),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_133),
.B(n_142),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_121),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g245 ( 
.A(n_237),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_113),
.A2(n_65),
.B1(n_72),
.B2(n_82),
.Y(n_238)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_136),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_239),
.B(n_195),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_198),
.A2(n_186),
.B1(n_234),
.B2(n_193),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_247),
.A2(n_258),
.B1(n_266),
.B2(n_267),
.Y(n_291)
);

OAI32xp33_ASAP7_75t_L g249 ( 
.A1(n_186),
.A2(n_219),
.A3(n_215),
.B1(n_185),
.B2(n_235),
.Y(n_249)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_249),
.B(n_241),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_250),
.B(n_255),
.C(n_184),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g251 ( 
.A(n_218),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_251),
.B(n_265),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g255 ( 
.A(n_207),
.B(n_225),
.C(n_217),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g265 ( 
.A(n_228),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_191),
.A2(n_190),
.B1(n_197),
.B2(n_181),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g267 ( 
.A1(n_197),
.A2(n_181),
.B1(n_214),
.B2(n_208),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_213),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g285 ( 
.A(n_269),
.B(n_274),
.Y(n_285)
);

AO21x2_ASAP7_75t_SL g271 ( 
.A1(n_208),
.A2(n_220),
.B(n_214),
.Y(n_271)
);

OA21x2_ASAP7_75t_L g294 ( 
.A1(n_271),
.A2(n_273),
.B(n_270),
.Y(n_294)
);

NOR2x1p5_ASAP7_75t_L g273 ( 
.A(n_194),
.B(n_239),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_213),
.Y(n_274)
);

CKINVDCx20_ASAP7_75t_R g276 ( 
.A(n_237),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_276),
.B(n_279),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_201),
.A2(n_212),
.B1(n_203),
.B2(n_210),
.Y(n_277)
);

AO22x2_ASAP7_75t_L g297 ( 
.A1(n_277),
.A2(n_271),
.B1(n_267),
.B2(n_266),
.Y(n_297)
);

HAxp5_ASAP7_75t_SL g311 ( 
.A(n_278),
.B(n_260),
.CON(n_311),
.SN(n_311)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_201),
.B(n_236),
.Y(n_279)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_243),
.Y(n_281)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_281),
.Y(n_313)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_270),
.A2(n_227),
.B(n_192),
.Y(n_282)
);

OAI21xp5_ASAP7_75t_SL g318 ( 
.A1(n_282),
.A2(n_295),
.B(n_273),
.Y(n_318)
);

OAI22xp33_ASAP7_75t_L g283 ( 
.A1(n_271),
.A2(n_237),
.B1(n_226),
.B2(n_200),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_283),
.A2(n_254),
.B1(n_273),
.B2(n_271),
.Y(n_317)
);

INVxp67_ASAP7_75t_L g315 ( 
.A(n_284),
.Y(n_315)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_255),
.B(n_188),
.C(n_223),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g314 ( 
.A(n_286),
.B(n_292),
.Y(n_314)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_243),
.Y(n_287)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_287),
.Y(n_316)
);

BUFx6f_ASAP7_75t_L g288 ( 
.A(n_257),
.Y(n_288)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_288),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_241),
.B(n_247),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_289),
.B(n_297),
.Y(n_329)
);

NOR2x1_ASAP7_75t_L g290 ( 
.A(n_270),
.B(n_268),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_290),
.B(n_308),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_248),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

NOR2xp33_ASAP7_75t_L g327 ( 
.A(n_293),
.B(n_299),
.Y(n_327)
);

OR2x2_ASAP7_75t_L g328 ( 
.A(n_294),
.B(n_280),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_251),
.A2(n_258),
.B(n_246),
.Y(n_295)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_253),
.Y(n_298)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_298),
.Y(n_325)
);

INVx2_ASAP7_75t_L g299 ( 
.A(n_244),
.Y(n_299)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_256),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_256),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_301),
.B(n_305),
.Y(n_332)
);

INVx3_ASAP7_75t_L g303 ( 
.A(n_244),
.Y(n_303)
);

AOI22xp33_ASAP7_75t_SL g322 ( 
.A1(n_303),
.A2(n_304),
.B1(n_245),
.B2(n_276),
.Y(n_322)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_265),
.A2(n_254),
.B1(n_271),
.B2(n_245),
.Y(n_304)
);

INVx2_ASAP7_75t_L g305 ( 
.A(n_244),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_252),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_306),
.B(n_307),
.Y(n_333)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_252),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_242),
.B(n_272),
.Y(n_308)
);

INVxp67_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_309),
.Y(n_330)
);

CKINVDCx14_ASAP7_75t_R g326 ( 
.A(n_311),
.Y(n_326)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_312),
.B(n_250),
.Y(n_334)
);

OAI22xp5_ASAP7_75t_L g343 ( 
.A1(n_317),
.A2(n_319),
.B1(n_322),
.B2(n_323),
.Y(n_343)
);

AOI21xp5_ASAP7_75t_L g353 ( 
.A1(n_318),
.A2(n_297),
.B(n_309),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_283),
.A2(n_240),
.B1(n_277),
.B2(n_261),
.Y(n_319)
);

OAI22xp33_ASAP7_75t_SL g321 ( 
.A1(n_295),
.A2(n_240),
.B1(n_259),
.B2(n_264),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_249),
.B1(n_280),
.B2(n_264),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g338 ( 
.A1(n_328),
.A2(n_294),
.B(n_291),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_291),
.A2(n_259),
.B1(n_262),
.B2(n_268),
.Y(n_331)
);

INVx2_ASAP7_75t_L g344 ( 
.A(n_331),
.Y(n_344)
);

AOI221xp5_ASAP7_75t_L g341 ( 
.A1(n_334),
.A2(n_292),
.B1(n_310),
.B2(n_286),
.C(n_262),
.Y(n_341)
);

NOR2x1_ASAP7_75t_L g336 ( 
.A(n_323),
.B(n_290),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g356 ( 
.A(n_336),
.B(n_338),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_315),
.B(n_284),
.C(n_289),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_337),
.B(n_345),
.C(n_346),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g339 ( 
.A(n_334),
.B(n_312),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_339),
.B(n_340),
.Y(n_365)
);

XNOR2x1_ASAP7_75t_L g340 ( 
.A(n_331),
.B(n_312),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_341),
.A2(n_326),
.B1(n_319),
.B2(n_317),
.Y(n_363)
);

OAI21xp5_ASAP7_75t_L g342 ( 
.A1(n_328),
.A2(n_282),
.B(n_302),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_342),
.B(n_349),
.Y(n_358)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_314),
.B(n_296),
.C(n_287),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_298),
.C(n_281),
.Y(n_346)
);

HB1xp67_ASAP7_75t_L g347 ( 
.A(n_327),
.Y(n_347)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_347),
.Y(n_361)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_333),
.Y(n_348)
);

INVx1_ASAP7_75t_L g354 ( 
.A(n_348),
.Y(n_354)
);

FAx1_ASAP7_75t_SL g349 ( 
.A(n_328),
.B(n_323),
.CI(n_320),
.CON(n_349),
.SN(n_349)
);

XNOR2xp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_297),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g359 ( 
.A(n_350),
.B(n_351),
.C(n_352),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g351 ( 
.A(n_329),
.B(n_293),
.C(n_297),
.Y(n_351)
);

OAI322xp33_ASAP7_75t_L g352 ( 
.A1(n_326),
.A2(n_285),
.A3(n_297),
.B1(n_301),
.B2(n_300),
.C1(n_269),
.C2(n_274),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_353),
.B(n_318),
.Y(n_364)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_348),
.Y(n_355)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_355),
.Y(n_368)
);

AOI22xp5_ASAP7_75t_L g360 ( 
.A1(n_343),
.A2(n_321),
.B1(n_317),
.B2(n_329),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g371 ( 
.A1(n_360),
.A2(n_344),
.B1(n_335),
.B2(n_342),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_337),
.B(n_328),
.C(n_318),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g375 ( 
.A(n_362),
.B(n_367),
.C(n_340),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g370 ( 
.A(n_363),
.B(n_350),
.Y(n_370)
);

OAI21xp5_ASAP7_75t_SL g369 ( 
.A1(n_364),
.A2(n_353),
.B(n_338),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g366 ( 
.A(n_345),
.B(n_327),
.Y(n_366)
);

NAND2xp5_ASAP7_75t_SL g377 ( 
.A(n_366),
.B(n_330),
.Y(n_377)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_346),
.B(n_330),
.C(n_319),
.Y(n_367)
);

AOI21xp5_ASAP7_75t_SL g387 ( 
.A1(n_369),
.A2(n_377),
.B(n_362),
.Y(n_387)
);

XOR2xp5_ASAP7_75t_L g379 ( 
.A(n_370),
.B(n_377),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_371),
.B(n_372),
.Y(n_382)
);

INVxp33_ASAP7_75t_SL g372 ( 
.A(n_366),
.Y(n_372)
);

OAI22xp5_ASAP7_75t_SL g373 ( 
.A1(n_360),
.A2(n_344),
.B1(n_335),
.B2(n_322),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g383 ( 
.A(n_373),
.B(n_376),
.Y(n_383)
);

AOI21xp5_ASAP7_75t_L g374 ( 
.A1(n_364),
.A2(n_343),
.B(n_351),
.Y(n_374)
);

OAI21xp5_ASAP7_75t_SL g380 ( 
.A1(n_374),
.A2(n_378),
.B(n_356),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_375),
.B(n_357),
.C(n_365),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g376 ( 
.A1(n_358),
.A2(n_349),
.B1(n_339),
.B2(n_336),
.Y(n_376)
);

AOI321xp33_ASAP7_75t_L g378 ( 
.A1(n_354),
.A2(n_349),
.A3(n_336),
.B1(n_313),
.B2(n_316),
.C(n_325),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_380),
.B(n_385),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_381),
.B(n_384),
.Y(n_391)
);

OAI21xp5_ASAP7_75t_SL g384 ( 
.A1(n_374),
.A2(n_356),
.B(n_359),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_375),
.B(n_357),
.C(n_359),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_370),
.B(n_367),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_386),
.B(n_376),
.Y(n_389)
);

AOI31xp33_ASAP7_75t_SL g393 ( 
.A1(n_387),
.A2(n_378),
.A3(n_371),
.B(n_369),
.Y(n_393)
);

OAI21xp5_ASAP7_75t_L g399 ( 
.A1(n_389),
.A2(n_393),
.B(n_394),
.Y(n_399)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_382),
.B(n_361),
.Y(n_390)
);

AOI21xp5_ASAP7_75t_L g396 ( 
.A1(n_390),
.A2(n_392),
.B(n_388),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_355),
.Y(n_392)
);

NOR2x1_ASAP7_75t_L g394 ( 
.A(n_379),
.B(n_354),
.Y(n_394)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_391),
.B(n_387),
.C(n_386),
.Y(n_395)
);

NAND2xp5_ASAP7_75t_L g402 ( 
.A(n_395),
.B(n_332),
.Y(n_402)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_396),
.B(n_333),
.Y(n_401)
);

XOR2xp5_ASAP7_75t_L g397 ( 
.A(n_394),
.B(n_383),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_397),
.B(n_398),
.C(n_368),
.Y(n_400)
);

AOI22xp5_ASAP7_75t_SL g398 ( 
.A1(n_393),
.A2(n_373),
.B1(n_368),
.B2(n_365),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_400),
.B(n_401),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_402),
.B(n_399),
.Y(n_403)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_403),
.B(n_397),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_405),
.B(n_406),
.C(n_313),
.Y(n_407)
);

OAI21xp5_ASAP7_75t_SL g406 ( 
.A1(n_404),
.A2(n_324),
.B(n_332),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_407),
.B(n_325),
.Y(n_408)
);


endmodule