module real_aes_15703_n_344 (n_76, n_113, n_187, n_90, n_257, n_65, n_74, n_185, n_285, n_30, n_222, n_61, n_20, n_287, n_64, n_254, n_207, n_10, n_83, n_181, n_124, n_191, n_209, n_299, n_322, n_328, n_19, n_40, n_318, n_239, n_100, n_54, n_112, n_319, n_35, n_42, n_329, n_132, n_131, n_144, n_169, n_242, n_308, n_172, n_341, n_232, n_6, n_69, n_317, n_321, n_73, n_320, n_77, n_260, n_37, n_97, n_186, n_138, n_26, n_235, n_245, n_161, n_189, n_271, n_2, n_145, n_227, n_92, n_330, n_332, n_292, n_116, n_94, n_289, n_280, n_333, n_213, n_184, n_28, n_202, n_56, n_34, n_98, n_121, n_125, n_216, n_82, n_327, n_47, n_106, n_32, n_263, n_230, n_51, n_248, n_301, n_27, n_343, n_174, n_18, n_104, n_211, n_281, n_173, n_234, n_284, n_153, n_316, n_75, n_178, n_298, n_49, n_43, n_297, n_9, n_119, n_310, n_164, n_231, n_44, n_102, n_122, n_141, n_128, n_111, n_167, n_80, n_179, n_12, n_68, n_129, n_304, n_311, n_324, n_25, n_278, n_236, n_267, n_218, n_48, n_204, n_339, n_89, n_277, n_331, n_93, n_182, n_323, n_199, n_142, n_223, n_67, n_250, n_85, n_45, n_5, n_244, n_118, n_139, n_87, n_171, n_78, n_146, n_17, n_226, n_255, n_286, n_120, n_261, n_238, n_58, n_165, n_246, n_176, n_163, n_29, n_52, n_251, n_220, n_197, n_296, n_3, n_41, n_256, n_71, n_302, n_126, n_200, n_115, n_96, n_110, n_150, n_147, n_288, n_23, n_334, n_274, n_160, n_303, n_95, n_188, n_269, n_201, n_306, n_158, n_4, n_193, n_293, n_162, n_275, n_214, n_46, n_109, n_59, n_203, n_81, n_133, n_273, n_114, n_276, n_295, n_265, n_154, n_127, n_326, n_24, n_217, n_55, n_1748, n_62, n_291, n_148, n_88, n_159, n_11, n_108, n_60, n_233, n_290, n_155, n_243, n_268, n_136, n_157, n_282, n_101, n_309, n_229, n_107, n_33, n_53, n_36, n_149, n_190, n_262, n_134, n_336, n_195, n_300, n_252, n_283, n_314, n_249, n_221, n_156, n_57, n_66, n_21, n_31, n_8, n_312, n_183, n_266, n_205, n_335, n_177, n_313, n_22, n_140, n_219, n_180, n_212, n_210, n_325, n_338, n_103, n_166, n_224, n_151, n_130, n_253, n_99, n_15, n_72, n_152, n_198, n_7, n_228, n_272, n_196, n_315, n_123, n_279, n_79, n_270, n_305, n_117, n_208, n_215, n_135, n_70, n_50, n_170, n_86, n_340, n_13, n_168, n_175, n_241, n_105, n_84, n_294, n_258, n_206, n_307, n_342, n_14, n_194, n_137, n_225, n_16, n_39, n_337, n_247, n_240, n_38, n_259, n_143, n_192, n_0, n_264, n_63, n_1, n_237, n_91, n_344);
input n_76;
input n_113;
input n_187;
input n_90;
input n_257;
input n_65;
input n_74;
input n_185;
input n_285;
input n_30;
input n_222;
input n_61;
input n_20;
input n_287;
input n_64;
input n_254;
input n_207;
input n_10;
input n_83;
input n_181;
input n_124;
input n_191;
input n_209;
input n_299;
input n_322;
input n_328;
input n_19;
input n_40;
input n_318;
input n_239;
input n_100;
input n_54;
input n_112;
input n_319;
input n_35;
input n_42;
input n_329;
input n_132;
input n_131;
input n_144;
input n_169;
input n_242;
input n_308;
input n_172;
input n_341;
input n_232;
input n_6;
input n_69;
input n_317;
input n_321;
input n_73;
input n_320;
input n_77;
input n_260;
input n_37;
input n_97;
input n_186;
input n_138;
input n_26;
input n_235;
input n_245;
input n_161;
input n_189;
input n_271;
input n_2;
input n_145;
input n_227;
input n_92;
input n_330;
input n_332;
input n_292;
input n_116;
input n_94;
input n_289;
input n_280;
input n_333;
input n_213;
input n_184;
input n_28;
input n_202;
input n_56;
input n_34;
input n_98;
input n_121;
input n_125;
input n_216;
input n_82;
input n_327;
input n_47;
input n_106;
input n_32;
input n_263;
input n_230;
input n_51;
input n_248;
input n_301;
input n_27;
input n_343;
input n_174;
input n_18;
input n_104;
input n_211;
input n_281;
input n_173;
input n_234;
input n_284;
input n_153;
input n_316;
input n_75;
input n_178;
input n_298;
input n_49;
input n_43;
input n_297;
input n_9;
input n_119;
input n_310;
input n_164;
input n_231;
input n_44;
input n_102;
input n_122;
input n_141;
input n_128;
input n_111;
input n_167;
input n_80;
input n_179;
input n_12;
input n_68;
input n_129;
input n_304;
input n_311;
input n_324;
input n_25;
input n_278;
input n_236;
input n_267;
input n_218;
input n_48;
input n_204;
input n_339;
input n_89;
input n_277;
input n_331;
input n_93;
input n_182;
input n_323;
input n_199;
input n_142;
input n_223;
input n_67;
input n_250;
input n_85;
input n_45;
input n_5;
input n_244;
input n_118;
input n_139;
input n_87;
input n_171;
input n_78;
input n_146;
input n_17;
input n_226;
input n_255;
input n_286;
input n_120;
input n_261;
input n_238;
input n_58;
input n_165;
input n_246;
input n_176;
input n_163;
input n_29;
input n_52;
input n_251;
input n_220;
input n_197;
input n_296;
input n_3;
input n_41;
input n_256;
input n_71;
input n_302;
input n_126;
input n_200;
input n_115;
input n_96;
input n_110;
input n_150;
input n_147;
input n_288;
input n_23;
input n_334;
input n_274;
input n_160;
input n_303;
input n_95;
input n_188;
input n_269;
input n_201;
input n_306;
input n_158;
input n_4;
input n_193;
input n_293;
input n_162;
input n_275;
input n_214;
input n_46;
input n_109;
input n_59;
input n_203;
input n_81;
input n_133;
input n_273;
input n_114;
input n_276;
input n_295;
input n_265;
input n_154;
input n_127;
input n_326;
input n_24;
input n_217;
input n_55;
input n_1748;
input n_62;
input n_291;
input n_148;
input n_88;
input n_159;
input n_11;
input n_108;
input n_60;
input n_233;
input n_290;
input n_155;
input n_243;
input n_268;
input n_136;
input n_157;
input n_282;
input n_101;
input n_309;
input n_229;
input n_107;
input n_33;
input n_53;
input n_36;
input n_149;
input n_190;
input n_262;
input n_134;
input n_336;
input n_195;
input n_300;
input n_252;
input n_283;
input n_314;
input n_249;
input n_221;
input n_156;
input n_57;
input n_66;
input n_21;
input n_31;
input n_8;
input n_312;
input n_183;
input n_266;
input n_205;
input n_335;
input n_177;
input n_313;
input n_22;
input n_140;
input n_219;
input n_180;
input n_212;
input n_210;
input n_325;
input n_338;
input n_103;
input n_166;
input n_224;
input n_151;
input n_130;
input n_253;
input n_99;
input n_15;
input n_72;
input n_152;
input n_198;
input n_7;
input n_228;
input n_272;
input n_196;
input n_315;
input n_123;
input n_279;
input n_79;
input n_270;
input n_305;
input n_117;
input n_208;
input n_215;
input n_135;
input n_70;
input n_50;
input n_170;
input n_86;
input n_340;
input n_13;
input n_168;
input n_175;
input n_241;
input n_105;
input n_84;
input n_294;
input n_258;
input n_206;
input n_307;
input n_342;
input n_14;
input n_194;
input n_137;
input n_225;
input n_16;
input n_39;
input n_337;
input n_247;
input n_240;
input n_38;
input n_259;
input n_143;
input n_192;
input n_0;
input n_264;
input n_63;
input n_1;
input n_237;
input n_91;
output n_344;
wire n_476;
wire n_599;
wire n_887;
wire n_1314;
wire n_1279;
wire n_830;
wire n_1371;
wire n_624;
wire n_618;
wire n_933;
wire n_485;
wire n_822;
wire n_750;
wire n_1641;
wire n_503;
wire n_1591;
wire n_469;
wire n_1310;
wire n_1376;
wire n_592;
wire n_1621;
wire n_1729;
wire n_1737;
wire n_761;
wire n_421;
wire n_919;
wire n_1217;
wire n_1423;
wire n_1034;
wire n_549;
wire n_571;
wire n_1328;
wire n_1219;
wire n_952;
wire n_1166;
wire n_752;
wire n_448;
wire n_556;
wire n_593;
wire n_989;
wire n_431;
wire n_1044;
wire n_1730;
wire n_1744;
wire n_963;
wire n_551;
wire n_884;
wire n_814;
wire n_944;
wire n_1283;
wire n_983;
wire n_955;
wire n_975;
wire n_941;
wire n_1313;
wire n_1468;
wire n_1713;
wire n_870;
wire n_1248;
wire n_1602;
wire n_548;
wire n_572;
wire n_815;
wire n_1140;
wire n_1453;
wire n_1520;
wire n_786;
wire n_512;
wire n_395;
wire n_795;
wire n_1379;
wire n_400;
wire n_1597;
wire n_1415;
wire n_1160;
wire n_1287;
wire n_883;
wire n_478;
wire n_1575;
wire n_1687;
wire n_553;
wire n_1367;
wire n_744;
wire n_1325;
wire n_1225;
wire n_1382;
wire n_875;
wire n_951;
wire n_1199;
wire n_1441;
wire n_1543;
wire n_791;
wire n_976;
wire n_636;
wire n_906;
wire n_477;
wire n_1477;
wire n_595;
wire n_1282;
wire n_683;
wire n_840;
wire n_570;
wire n_675;
wire n_835;
wire n_732;
wire n_784;
wire n_962;
wire n_1599;
wire n_755;
wire n_409;
wire n_781;
wire n_576;
wire n_1688;
wire n_956;
wire n_1242;
wire n_1537;
wire n_796;
wire n_874;
wire n_1126;
wire n_383;
wire n_1607;
wire n_455;
wire n_682;
wire n_1745;
wire n_812;
wire n_782;
wire n_817;
wire n_760;
wire n_608;
wire n_534;
wire n_1454;
wire n_708;
wire n_1020;
wire n_885;
wire n_950;
wire n_381;
wire n_1196;
wire n_1013;
wire n_808;
wire n_1639;
wire n_1224;
wire n_1694;
wire n_688;
wire n_1042;
wire n_1588;
wire n_363;
wire n_1317;
wire n_417;
wire n_690;
wire n_1419;
wire n_499;
wire n_1142;
wire n_1731;
wire n_1589;
wire n_947;
wire n_970;
wire n_1677;
wire n_1149;
wire n_368;
wire n_527;
wire n_1676;
wire n_1342;
wire n_1440;
wire n_552;
wire n_1383;
wire n_1346;
wire n_1675;
wire n_590;
wire n_1293;
wire n_432;
wire n_1131;
wire n_1008;
wire n_1491;
wire n_805;
wire n_1600;
wire n_619;
wire n_1095;
wire n_1250;
wire n_1284;
wire n_360;
wire n_1583;
wire n_1465;
wire n_859;
wire n_1486;
wire n_1304;
wire n_685;
wire n_1080;
wire n_917;
wire n_1247;
wire n_501;
wire n_1380;
wire n_488;
wire n_1658;
wire n_954;
wire n_702;
wire n_1007;
wire n_351;
wire n_898;
wire n_562;
wire n_1022;
wire n_1502;
wire n_404;
wire n_1073;
wire n_728;
wire n_1301;
wire n_1632;
wire n_1201;
wire n_997;
wire n_1105;
wire n_1243;
wire n_1003;
wire n_346;
wire n_749;
wire n_914;
wire n_1286;
wire n_494;
wire n_1661;
wire n_927;
wire n_723;
wire n_972;
wire n_1351;
wire n_1628;
wire n_1587;
wire n_1570;
wire n_1209;
wire n_411;
wire n_498;
wire n_765;
wire n_1397;
wire n_1554;
wire n_648;
wire n_1487;
wire n_939;
wire n_1615;
wire n_928;
wire n_1384;
wire n_789;
wire n_1515;
wire n_738;
wire n_1387;
wire n_922;
wire n_1048;
wire n_1422;
wire n_787;
wire n_1214;
wire n_806;
wire n_715;
wire n_1714;
wire n_420;
wire n_1666;
wire n_1490;
wire n_1258;
wire n_873;
wire n_438;
wire n_446;
wire n_1281;
wire n_1559;
wire n_1510;
wire n_1495;
wire n_1727;
wire n_712;
wire n_422;
wire n_861;
wire n_1574;
wire n_479;
wire n_825;
wire n_541;
wire n_839;
wire n_811;
wire n_558;
wire n_1742;
wire n_724;
wire n_1648;
wire n_440;
wire n_1231;
wire n_1305;
wire n_1161;
wire n_686;
wire n_1299;
wire n_949;
wire n_586;
wire n_1508;
wire n_1421;
wire n_788;
wire n_441;
wire n_1045;
wire n_1339;
wire n_837;
wire n_1349;
wire n_1708;
wire n_1445;
wire n_1631;
wire n_829;
wire n_1030;
wire n_1348;
wire n_375;
wire n_1391;
wire n_597;
wire n_1036;
wire n_687;
wire n_652;
wire n_1538;
wire n_500;
wire n_804;
wire n_1173;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_1488;
wire n_1572;
wire n_1514;
wire n_480;
wire n_1652;
wire n_684;
wire n_1178;
wire n_1531;
wire n_821;
wire n_1657;
wire n_1616;
wire n_1563;
wire n_1018;
wire n_980;
wire n_1233;
wire n_1106;
wire n_1205;
wire n_838;
wire n_1561;
wire n_635;
wire n_792;
wire n_1392;
wire n_1542;
wire n_665;
wire n_991;
wire n_667;
wire n_1712;
wire n_1556;
wire n_580;
wire n_1004;
wire n_1417;
wire n_1370;
wire n_1703;
wire n_1717;
wire n_1723;
wire n_979;
wire n_445;
wire n_596;
wire n_1740;
wire n_1197;
wire n_657;
wire n_1260;
wire n_355;
wire n_1606;
wire n_1129;
wire n_1285;
wire n_742;
wire n_1014;
wire n_1385;
wire n_1629;
wire n_1618;
wire n_461;
wire n_1047;
wire n_1016;
wire n_1545;
wire n_694;
wire n_1350;
wire n_894;
wire n_545;
wire n_1459;
wire n_1530;
wire n_401;
wire n_538;
wire n_1594;
wire n_537;
wire n_1651;
wire n_560;
wire n_1094;
wire n_1719;
wire n_1220;
wire n_696;
wire n_1147;
wire n_1425;
wire n_1613;
wire n_1504;
wire n_704;
wire n_453;
wire n_647;
wire n_399;
wire n_948;
wire n_700;
wire n_1499;
wire n_677;
wire n_1269;
wire n_378;
wire n_591;
wire n_1635;
wire n_1518;
wire n_1702;
wire n_1366;
wire n_678;
wire n_415;
wire n_1400;
wire n_564;
wire n_638;
wire n_510;
wire n_1361;
wire n_1358;
wire n_1577;
wire n_1642;
wire n_1406;
wire n_550;
wire n_966;
wire n_1568;
wire n_1368;
wire n_994;
wire n_384;
wire n_1612;
wire n_1479;
wire n_1128;
wire n_1098;
wire n_824;
wire n_1238;
wire n_1611;
wire n_992;
wire n_813;
wire n_981;
wire n_1338;
wire n_1182;
wire n_872;
wire n_1401;
wire n_1086;
wire n_1189;
wire n_1070;
wire n_1665;
wire n_535;
wire n_882;
wire n_1741;
wire n_1210;
wire n_1456;
wire n_746;
wire n_656;
wire n_1614;
wire n_1148;
wire n_748;
wire n_860;
wire n_1261;
wire n_1062;
wire n_1439;
wire n_651;
wire n_1585;
wire n_1500;
wire n_801;
wire n_1271;
wire n_1653;
wire n_529;
wire n_504;
wire n_973;
wire n_1364;
wire n_659;
wire n_634;
wire n_903;
wire n_1668;
wire n_565;
wire n_925;
wire n_1389;
wire n_1393;
wire n_457;
wire n_1121;
wire n_1059;
wire n_493;
wire n_1362;
wire n_610;
wire n_1035;
wire n_620;
wire n_722;
wire n_1174;
wire n_1193;
wire n_1553;
wire n_754;
wire n_508;
wire n_1141;
wire n_1112;
wire n_1485;
wire n_1408;
wire n_1680;
wire n_428;
wire n_783;
wire n_1107;
wire n_1564;
wire n_505;
wire n_600;
wire n_731;
wire n_964;
wire n_605;
wire n_1516;
wire n_1386;
wire n_406;
wire n_1493;
wire n_1579;
wire n_617;
wire n_733;
wire n_402;
wire n_602;
wire n_1404;
wire n_658;
wire n_676;
wire n_531;
wire n_1031;
wire n_1394;
wire n_807;
wire n_1011;
wire n_416;
wire n_1567;
wire n_895;
wire n_1569;
wire n_799;
wire n_490;
wire n_391;
wire n_695;
wire n_1181;
wire n_881;
wire n_1626;
wire n_1145;
wire n_645;
wire n_1529;
wire n_557;
wire n_1681;
wire n_1620;
wire n_777;
wire n_985;
wire n_1659;
wire n_910;
wire n_642;
wire n_613;
wire n_1125;
wire n_1347;
wire n_1655;
wire n_1522;
wire n_1163;
wire n_1278;
wire n_734;
wire n_1623;
wire n_735;
wire n_1179;
wire n_569;
wire n_1171;
wire n_785;
wire n_1203;
wire n_1716;
wire n_1232;
wire n_471;
wire n_853;
wire n_810;
wire n_1136;
wire n_699;
wire n_1187;
wire n_1000;
wire n_1580;
wire n_649;
wire n_358;
wire n_1234;
wire n_622;
wire n_1634;
wire n_1002;
wire n_1353;
wire n_1165;
wire n_1551;
wire n_1667;
wire n_1058;
wire n_1216;
wire n_662;
wire n_850;
wire n_354;
wire n_720;
wire n_1026;
wire n_492;
wire n_407;
wire n_419;
wire n_1023;
wire n_730;
wire n_1699;
wire n_643;
wire n_1403;
wire n_486;
wire n_779;
wire n_481;
wire n_691;
wire n_589;
wire n_365;
wire n_526;
wire n_1513;
wire n_1194;
wire n_389;
wire n_1609;
wire n_1462;
wire n_701;
wire n_809;
wire n_1532;
wire n_520;
wire n_679;
wire n_926;
wire n_1643;
wire n_942;
wire n_1374;
wire n_1120;
wire n_1497;
wire n_1548;
wire n_1526;
wire n_689;
wire n_1483;
wire n_946;
wire n_753;
wire n_1409;
wire n_1188;
wire n_623;
wire n_1032;
wire n_1474;
wire n_721;
wire n_1431;
wire n_1133;
wire n_1593;
wire n_739;
wire n_1322;
wire n_1525;
wire n_1732;
wire n_1162;
wire n_1463;
wire n_762;
wire n_1524;
wire n_1298;
wire n_1633;
wire n_442;
wire n_740;
wire n_1686;
wire n_1357;
wire n_639;
wire n_1186;
wire n_1365;
wire n_459;
wire n_1172;
wire n_1689;
wire n_998;
wire n_1625;
wire n_1395;
wire n_1276;
wire n_836;
wire n_1733;
wire n_1184;
wire n_583;
wire n_347;
wire n_414;
wire n_1336;
wire n_776;
wire n_1138;
wire n_890;
wire n_1306;
wire n_1413;
wire n_1266;
wire n_497;
wire n_911;
wire n_450;
wire n_1578;
wire n_473;
wire n_967;
wire n_1709;
wire n_1159;
wire n_474;
wire n_1315;
wire n_1055;
wire n_611;
wire n_380;
wire n_1576;
wire n_844;
wire n_968;
wire n_710;
wire n_1040;
wire n_1102;
wire n_661;
wire n_1185;
wire n_447;
wire n_403;
wire n_1039;
wire n_1119;
wire n_574;
wire n_1069;
wire n_1451;
wire n_842;
wire n_798;
wire n_1700;
wire n_668;
wire n_862;
wire n_869;
wire n_1066;
wire n_1377;
wire n_800;
wire n_778;
wire n_1170;
wire n_1175;
wire n_522;
wire n_1475;
wire n_977;
wire n_943;
wire n_357;
wire n_905;
wire n_386;
wire n_878;
wire n_1734;
wire n_1333;
wire n_577;
wire n_1610;
wire n_759;
wire n_1235;
wire n_900;
wire n_841;
wire n_1724;
wire n_1218;
wire n_736;
wire n_1706;
wire n_766;
wire n_1113;
wire n_1268;
wire n_852;
wire n_1695;
wire n_1089;
wire n_1122;
wire n_908;
wire n_1123;
wire n_923;
wire n_1302;
wire n_1289;
wire n_937;
wire n_1442;
wire n_773;
wire n_353;
wire n_1446;
wire n_865;
wire n_1644;
wire n_1736;
wire n_1707;
wire n_856;
wire n_594;
wire n_1146;
wire n_1685;
wire n_1435;
wire n_374;
wire n_932;
wire n_958;
wire n_775;
wire n_763;
wire n_1093;
wire n_427;
wire n_1540;
wire n_519;
wire n_1116;
wire n_709;
wire n_388;
wire n_1470;
wire n_816;
wire n_625;
wire n_953;
wire n_1565;
wire n_1373;
wire n_1558;
wire n_716;
wire n_1683;
wire n_356;
wire n_584;
wire n_896;
wire n_1722;
wire n_528;
wire n_1078;
wire n_495;
wire n_1072;
wire n_1638;
wire n_370;
wire n_1663;
wire n_352;
wire n_935;
wire n_1505;
wire n_467;
wire n_1213;
wire n_1053;
wire n_515;
wire n_1019;
wire n_680;
wire n_1180;
wire n_904;
wire n_920;
wire n_1117;
wire n_1168;
wire n_1598;
wire n_1309;
wire n_909;
wire n_523;
wire n_996;
wire n_439;
wire n_506;
wire n_606;
wire n_513;
wire n_1332;
wire n_1411;
wire n_1263;
wire n_1115;
wire n_725;
wire n_960;
wire n_671;
wire n_1084;
wire n_1726;
wire n_1656;
wire n_454;
wire n_1303;
wire n_1471;
wire n_443;
wire n_1029;
wire n_345;
wire n_1207;
wire n_1555;
wire n_664;
wire n_367;
wire n_1017;
wire n_581;
wire n_936;
wire n_1215;
wire n_582;
wire n_641;
wire n_1738;
wire n_940;
wire n_745;
wire n_1608;
wire n_1167;
wire n_1327;
wire n_609;
wire n_1743;
wire n_1006;
wire n_1259;
wire n_350;
wire n_561;
wire n_437;
wire n_1560;
wire n_405;
wire n_1223;
wire n_621;
wire n_1012;
wire n_1241;
wire n_1414;
wire n_1671;
wire n_502;
wire n_434;
wire n_769;
wire n_1212;
wire n_1455;
wire n_1054;
wire n_1669;
wire n_1308;
wire n_1050;
wire n_426;
wire n_1550;
wire n_1134;
wire n_1670;
wire n_1319;
wire n_1363;
wire n_616;
wire n_880;
wire n_1103;
wire n_1274;
wire n_832;
wire n_1321;
wire n_1429;
wire n_1660;
wire n_1060;
wire n_1154;
wire n_361;
wire n_632;
wire n_1344;
wire n_1450;
wire n_1603;
wire n_1720;
wire n_1331;
wire n_714;
wire n_1222;
wire n_1041;
wire n_1512;
wire n_957;
wire n_1255;
wire n_995;
wire n_1124;
wire n_1335;
wire n_1405;
wire n_912;
wire n_464;
wire n_1227;
wire n_1509;
wire n_945;
wire n_392;
wire n_563;
wire n_891;
wire n_568;
wire n_1586;
wire n_413;
wire n_1157;
wire n_902;
wire n_1158;
wire n_1079;
wire n_1330;
wire n_1033;
wire n_1464;
wire n_1028;
wire n_366;
wire n_727;
wire n_1083;
wire n_397;
wire n_1056;
wire n_1592;
wire n_1605;
wire n_663;
wire n_588;
wire n_1682;
wire n_1698;
wire n_1448;
wire n_707;
wire n_915;
wire n_1001;
wire n_1418;
wire n_711;
wire n_864;
wire n_1169;
wire n_377;
wire n_1139;
wire n_1482;
wire n_1038;
wire n_1085;
wire n_845;
wire n_1673;
wire n_1619;
wire n_1127;
wire n_1718;
wire n_484;
wire n_893;
wire n_1068;
wire n_747;
wire n_1672;
wire n_1244;
wire n_1581;
wire n_697;
wire n_978;
wire n_847;
wire n_1452;
wire n_826;
wire n_373;
wire n_628;
wire n_487;
wire n_831;
wire n_653;
wire n_1725;
wire n_692;
wire n_1433;
wire n_1051;
wire n_1696;
wire n_1355;
wire n_1494;
wire n_1517;
wire n_827;
wire n_472;
wire n_866;
wire n_452;
wire n_630;
wire n_820;
wire n_1208;
wire n_612;
wire n_1426;
wire n_858;
wire n_764;
wire n_741;
wire n_1090;
wire n_456;
wire n_359;
wire n_1469;
wire n_1164;
wire n_433;
wire n_627;
wire n_1693;
wire n_418;
wire n_771;
wire n_1378;
wire n_524;
wire n_1496;
wire n_1191;
wire n_705;
wire n_1206;
wire n_1270;
wire n_1566;
wire n_1399;
wire n_546;
wire n_1010;
wire n_1375;
wire n_1015;
wire n_863;
wire n_525;
wire n_1226;
wire n_1617;
wire n_644;
wire n_1150;
wire n_1341;
wire n_833;
wire n_1229;
wire n_1690;
wire n_929;
wire n_1143;
wire n_1190;
wire n_1728;
wire n_543;
wire n_1710;
wire n_585;
wire n_1343;
wire n_465;
wire n_719;
wire n_1457;
wire n_1604;
wire n_1156;
wire n_988;
wire n_1466;
wire n_921;
wire n_1396;
wire n_640;
wire n_1176;
wire n_1721;
wire n_1691;
wire n_1511;
wire n_1151;
wire n_1501;
wire n_1254;
wire n_1458;
wire n_646;
wire n_1211;
wire n_650;
wire n_743;
wire n_823;
wire n_393;
wire n_1480;
wire n_1101;
wire n_1251;
wire n_1076;
wire n_1434;
wire n_1461;
wire n_1449;
wire n_1715;
wire n_1407;
wire n_1104;
wire n_849;
wire n_1061;
wire n_554;
wire n_1153;
wire n_1337;
wire n_797;
wire n_1704;
wire n_1177;
wire n_758;
wire n_436;
wire n_390;
wire n_1096;
wire n_1316;
wire n_1590;
wire n_1420;
wire n_1552;
wire n_1544;
wire n_1571;
wire n_1092;
wire n_846;
wire n_631;
wire n_673;
wire n_1410;
wire n_1067;
wire n_518;
wire n_1292;
wire n_1192;
wire n_1478;
wire n_1507;
wire n_1240;
wire n_987;
wire n_1596;
wire n_362;
wire n_1065;
wire n_540;
wire n_1064;
wire n_1075;
wire n_718;
wire n_669;
wire n_1091;
wire n_423;
wire n_1221;
wire n_458;
wire n_1200;
wire n_444;
wire n_364;
wire n_555;
wire n_1295;
wire n_974;
wire n_1329;
wire n_857;
wire n_1424;
wire n_1674;
wire n_376;
wire n_491;
wire n_1294;
wire n_1110;
wire n_1137;
wire n_1533;
wire n_460;
wire n_1679;
wire n_1595;
wire n_1735;
wire n_666;
wire n_660;
wire n_1359;
wire n_886;
wire n_767;
wire n_889;
wire n_1398;
wire n_379;
wire n_1432;
wire n_1021;
wire n_1297;
wire n_1046;
wire n_1109;
wire n_961;
wire n_1447;
wire n_489;
wire n_1622;
wire n_1381;
wire n_1582;
wire n_573;
wire n_1099;
wire n_1654;
wire n_626;
wire n_539;
wire n_462;
wire n_615;
wire n_1118;
wire n_990;
wire n_1108;
wire n_670;
wire n_818;
wire n_918;
wire n_1272;
wire n_1541;
wire n_408;
wire n_892;
wire n_578;
wire n_372;
wire n_938;
wire n_774;
wire n_466;
wire n_559;
wire n_1049;
wire n_1277;
wire n_1584;
wire n_984;
wire n_726;
wire n_369;
wire n_517;
wire n_931;
wire n_780;
wire n_530;
wire n_834;
wire n_693;
wire n_496;
wire n_1360;
wire n_1082;
wire n_1257;
wire n_468;
wire n_532;
wire n_1025;
wire n_924;
wire n_1264;
wire n_1527;
wire n_1245;
wire n_1152;
wire n_1539;
wire n_1081;
wire n_547;
wire n_1324;
wire n_1198;
wire n_1678;
wire n_1307;
wire n_993;
wire n_819;
wire n_737;
wire n_1489;
wire n_1637;
wire n_1318;
wire n_1290;
wire n_1135;
wire n_1063;
wire n_828;
wire n_770;
wire n_867;
wire n_1100;
wire n_398;
wire n_1519;
wire n_425;
wire n_1650;
wire n_879;
wire n_1640;
wire n_449;
wire n_1340;
wire n_1562;
wire n_607;
wire n_629;
wire n_706;
wire n_901;
wire n_876;
wire n_1443;
wire n_655;
wire n_654;
wire n_1521;
wire n_672;
wire n_567;
wire n_916;
wire n_1354;
wire n_1547;
wire n_1334;
wire n_1291;
wire n_1437;
wire n_1473;
wire n_986;
wire n_451;
wire n_1037;
wire n_1267;
wire n_790;
wire n_1262;
wire n_410;
wire n_1684;
wire n_1444;
wire n_751;
wire n_999;
wire n_913;
wire n_1237;
wire n_1506;
wire n_1356;
wire n_1646;
wire n_768;
wire n_412;
wire n_542;
wire n_1256;
wire n_1427;
wire n_1077;
wire n_1111;
wire n_1503;
wire n_1249;
wire n_1416;
wire n_387;
wire n_1239;
wire n_1662;
wire n_969;
wire n_1535;
wire n_1009;
wire n_1202;
wire n_1498;
wire n_1549;
wire n_604;
wire n_848;
wire n_756;
wire n_713;
wire n_598;
wire n_430;
wire n_1252;
wire n_1647;
wire n_1132;
wire n_1649;
wire n_1275;
wire n_843;
wire n_579;
wire n_533;
wire n_1472;
wire n_385;
wire n_536;
wire n_470;
wire n_851;
wire n_1155;
wire n_934;
wire n_1636;
wire n_1027;
wire n_965;
wire n_1296;
wire n_382;
wire n_1484;
wire n_1043;
wire n_435;
wire n_511;
wire n_1492;
wire n_1467;
wire n_509;
wire n_1204;
wire n_930;
wire n_1265;
wire n_1057;
wire n_907;
wire n_1430;
wire n_1481;
wire n_1005;
wire n_1312;
wire n_1697;
wire n_899;
wire n_637;
wire n_544;
wire n_1476;
wire n_1087;
wire n_1536;
wire n_1746;
wire n_1711;
wire n_482;
wire n_633;
wire n_971;
wire n_1052;
wire n_1071;
wire n_1311;
wire n_1601;
wire n_1438;
wire n_1273;
wire n_959;
wire n_349;
wire n_1573;
wire n_1130;
wire n_794;
wire n_1228;
wire n_681;
wire n_982;
wire n_717;
wire n_1624;
wire n_1253;
wire n_1183;
wire n_516;
wire n_1460;
wire n_521;
wire n_1195;
wire n_575;
wire n_1300;
wire n_1372;
wire n_698;
wire n_371;
wire n_1345;
wire n_587;
wire n_1701;
wire n_1664;
wire n_1428;
wire n_1246;
wire n_1074;
wire n_674;
wire n_888;
wire n_1546;
wire n_1436;
wire n_793;
wire n_1390;
wire n_1412;
wire n_757;
wire n_1534;
wire n_803;
wire n_514;
wire n_507;
wire n_1557;
wire n_614;
wire n_772;
wire n_1114;
wire n_566;
wire n_871;
wire n_1739;
wire n_1088;
wire n_1230;
wire n_1326;
wire n_1402;
wire n_1388;
wire n_483;
wire n_1630;
wire n_1352;
wire n_729;
wire n_394;
wire n_1280;
wire n_1323;
wire n_703;
wire n_1097;
wire n_1369;
wire n_601;
wire n_463;
wire n_396;
wire n_1236;
wire n_1523;
wire n_348;
wire n_1528;
wire n_603;
wire n_1692;
wire n_1288;
wire n_868;
wire n_1705;
wire n_1024;
wire n_1144;
wire n_1627;
wire n_475;
wire n_897;
wire n_1320;
wire n_855;
wire n_1645;
wire n_429;
INVx1_ASAP7_75t_L g1645 ( .A(n_0), .Y(n_1645) );
AO22x1_ASAP7_75t_L g1669 ( .A1(n_0), .A2(n_231), .B1(n_385), .B2(n_572), .Y(n_1669) );
AND2x2_ASAP7_75t_L g363 ( .A(n_1), .B(n_364), .Y(n_363) );
INVx1_ASAP7_75t_L g383 ( .A(n_1), .Y(n_383) );
AND2x2_ASAP7_75t_L g410 ( .A(n_1), .B(n_248), .Y(n_410) );
NOR2xp33_ASAP7_75t_L g912 ( .A(n_1), .B(n_382), .Y(n_912) );
INVx1_ASAP7_75t_L g1653 ( .A(n_2), .Y(n_1653) );
AOI22xp33_ASAP7_75t_L g1668 ( .A1(n_2), .A2(n_128), .B1(n_373), .B2(n_375), .Y(n_1668) );
AOI22xp33_ASAP7_75t_SL g529 ( .A1(n_3), .A2(n_47), .B1(n_440), .B2(n_530), .Y(n_529) );
INVxp67_ASAP7_75t_SL g606 ( .A(n_3), .Y(n_606) );
INVx1_ASAP7_75t_L g1704 ( .A(n_4), .Y(n_1704) );
INVx1_ASAP7_75t_L g1350 ( .A(n_5), .Y(n_1350) );
OAI22xp5_ASAP7_75t_L g1367 ( .A1(n_5), .A2(n_331), .B1(n_562), .B2(n_567), .Y(n_1367) );
AOI22xp33_ASAP7_75t_L g1702 ( .A1(n_6), .A2(n_73), .B1(n_544), .B2(n_644), .Y(n_1702) );
AOI221xp5_ASAP7_75t_L g1720 ( .A1(n_6), .A2(n_14), .B1(n_656), .B2(n_657), .C(n_1721), .Y(n_1720) );
INVx1_ASAP7_75t_L g843 ( .A(n_7), .Y(n_843) );
AOI22xp33_ASAP7_75t_SL g1186 ( .A1(n_8), .A2(n_223), .B1(n_638), .B2(n_1187), .Y(n_1186) );
INVxp67_ASAP7_75t_SL g1212 ( .A(n_8), .Y(n_1212) );
AOI221xp5_ASAP7_75t_L g857 ( .A1(n_9), .A2(n_295), .B1(n_379), .B2(n_729), .C(n_858), .Y(n_857) );
AOI22xp33_ASAP7_75t_SL g877 ( .A1(n_9), .A2(n_315), .B1(n_451), .B2(n_534), .Y(n_877) );
AOI22xp33_ASAP7_75t_L g646 ( .A1(n_10), .A2(n_280), .B1(n_644), .B2(n_647), .Y(n_646) );
AOI221xp5_ASAP7_75t_L g652 ( .A1(n_10), .A2(n_87), .B1(n_375), .B2(n_614), .C(n_653), .Y(n_652) );
AOI22xp33_ASAP7_75t_L g757 ( .A1(n_11), .A2(n_317), .B1(n_371), .B2(n_758), .Y(n_757) );
INVx1_ASAP7_75t_L g777 ( .A(n_11), .Y(n_777) );
INVxp67_ASAP7_75t_SL g1123 ( .A(n_12), .Y(n_1123) );
AND4x1_ASAP7_75t_L g1164 ( .A(n_12), .B(n_1125), .C(n_1128), .D(n_1147), .Y(n_1164) );
OAI22xp5_ASAP7_75t_L g1632 ( .A1(n_13), .A2(n_1633), .B1(n_1634), .B2(n_1635), .Y(n_1632) );
CKINVDCx5p33_ASAP7_75t_R g1633 ( .A(n_13), .Y(n_1633) );
AOI22xp33_ASAP7_75t_SL g1712 ( .A1(n_14), .A2(n_242), .B1(n_440), .B2(n_1088), .Y(n_1712) );
INVx2_ASAP7_75t_L g428 ( .A(n_15), .Y(n_428) );
OAI22xp5_ASAP7_75t_SL g1286 ( .A1(n_16), .A2(n_276), .B1(n_724), .B2(n_1287), .Y(n_1286) );
OAI221xp5_ASAP7_75t_L g1297 ( .A1(n_16), .A2(n_276), .B1(n_598), .B2(n_600), .C(n_1298), .Y(n_1297) );
XNOR2x1_ASAP7_75t_L g1267 ( .A(n_17), .B(n_1268), .Y(n_1267) );
AOI22xp5_ASAP7_75t_L g1461 ( .A1(n_17), .A2(n_19), .B1(n_1407), .B2(n_1415), .Y(n_1461) );
INVx1_ASAP7_75t_L g797 ( .A(n_18), .Y(n_797) );
OAI222xp33_ASAP7_75t_L g826 ( .A1(n_18), .A2(n_166), .B1(n_664), .B2(n_682), .C1(n_827), .C2(n_832), .Y(n_826) );
AOI22xp33_ASAP7_75t_L g645 ( .A1(n_20), .A2(n_228), .B1(n_451), .B2(n_640), .Y(n_645) );
AOI22xp33_ASAP7_75t_L g654 ( .A1(n_20), .A2(n_142), .B1(n_655), .B2(n_657), .Y(n_654) );
INVx1_ASAP7_75t_L g1069 ( .A(n_21), .Y(n_1069) );
AOI22xp33_ASAP7_75t_L g861 ( .A1(n_22), .A2(n_261), .B1(n_583), .B2(n_585), .Y(n_861) );
AOI22xp33_ASAP7_75t_L g879 ( .A1(n_22), .A2(n_255), .B1(n_440), .B2(n_458), .Y(n_879) );
INVx1_ASAP7_75t_L g1708 ( .A(n_23), .Y(n_1708) );
OAI22xp5_ASAP7_75t_L g1127 ( .A1(n_24), .A2(n_160), .B1(n_562), .B2(n_567), .Y(n_1127) );
OAI211xp5_ASAP7_75t_L g1129 ( .A1(n_24), .A2(n_1097), .B(n_1130), .C(n_1133), .Y(n_1129) );
OAI22xp5_ASAP7_75t_L g1094 ( .A1(n_25), .A2(n_296), .B1(n_562), .B2(n_567), .Y(n_1094) );
AOI22xp33_ASAP7_75t_L g1137 ( .A1(n_26), .A2(n_95), .B1(n_385), .B2(n_742), .Y(n_1137) );
AOI22xp33_ASAP7_75t_L g1157 ( .A1(n_26), .A2(n_37), .B1(n_535), .B2(n_1155), .Y(n_1157) );
CKINVDCx5p33_ASAP7_75t_R g688 ( .A(n_27), .Y(n_688) );
INVx1_ASAP7_75t_L g1296 ( .A(n_28), .Y(n_1296) );
HB1xp67_ASAP7_75t_L g1391 ( .A(n_29), .Y(n_1391) );
AND2x2_ASAP7_75t_L g1408 ( .A(n_29), .B(n_1389), .Y(n_1408) );
AOI22xp33_ASAP7_75t_L g1541 ( .A1(n_30), .A2(n_193), .B1(n_1415), .B2(n_1436), .Y(n_1541) );
OAI22xp5_ASAP7_75t_SL g1038 ( .A1(n_31), .A2(n_281), .B1(n_1039), .B2(n_1040), .Y(n_1038) );
INVxp67_ASAP7_75t_SL g1072 ( .A(n_31), .Y(n_1072) );
AOI22xp33_ASAP7_75t_L g1086 ( .A1(n_32), .A2(n_221), .B1(n_451), .B2(n_1084), .Y(n_1086) );
AOI221xp5_ASAP7_75t_L g1114 ( .A1(n_32), .A2(n_306), .B1(n_617), .B2(n_1115), .C(n_1117), .Y(n_1114) );
CKINVDCx5p33_ASAP7_75t_R g1168 ( .A(n_33), .Y(n_1168) );
INVx1_ASAP7_75t_L g1225 ( .A(n_34), .Y(n_1225) );
OAI211xp5_ASAP7_75t_L g1233 ( .A1(n_34), .A2(n_825), .B(n_1206), .C(n_1234), .Y(n_1233) );
CKINVDCx5p33_ASAP7_75t_R g1126 ( .A(n_35), .Y(n_1126) );
AOI22xp5_ASAP7_75t_L g865 ( .A1(n_36), .A2(n_315), .B1(n_371), .B2(n_583), .Y(n_865) );
AOI22xp5_ASAP7_75t_L g878 ( .A1(n_36), .A2(n_295), .B1(n_451), .B2(n_804), .Y(n_878) );
AOI221xp5_ASAP7_75t_L g1144 ( .A1(n_37), .A2(n_324), .B1(n_375), .B2(n_617), .C(n_1145), .Y(n_1144) );
AOI22xp33_ASAP7_75t_L g1000 ( .A1(n_38), .A2(n_57), .B1(n_452), .B2(n_942), .Y(n_1000) );
INVx1_ASAP7_75t_L g1010 ( .A(n_38), .Y(n_1010) );
INVx1_ASAP7_75t_L g1080 ( .A(n_39), .Y(n_1080) );
OAI221xp5_ASAP7_75t_L g1108 ( .A1(n_39), .A2(n_244), .B1(n_596), .B2(n_600), .C(n_1109), .Y(n_1108) );
INVx1_ASAP7_75t_L g921 ( .A(n_40), .Y(n_921) );
INVx1_ASAP7_75t_L g823 ( .A(n_41), .Y(n_823) );
AOI22xp5_ASAP7_75t_L g887 ( .A1(n_42), .A2(n_53), .B1(n_888), .B2(n_889), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g940 ( .A1(n_42), .A2(n_159), .B1(n_451), .B2(n_941), .Y(n_940) );
AOI221xp5_ASAP7_75t_L g1244 ( .A1(n_43), .A2(n_297), .B1(n_375), .B2(n_379), .C(n_614), .Y(n_1244) );
INVxp67_ASAP7_75t_SL g1252 ( .A(n_43), .Y(n_1252) );
INVxp67_ASAP7_75t_SL g1707 ( .A(n_44), .Y(n_1707) );
OAI22xp5_ASAP7_75t_L g1729 ( .A1(n_44), .A2(n_163), .B1(n_678), .B2(n_1730), .Y(n_1729) );
INVx1_ASAP7_75t_L g1230 ( .A(n_45), .Y(n_1230) );
OAI22xp5_ASAP7_75t_L g1245 ( .A1(n_45), .A2(n_212), .B1(n_1097), .B2(n_1246), .Y(n_1245) );
AOI221xp5_ASAP7_75t_L g989 ( .A1(n_46), .A2(n_334), .B1(n_443), .B2(n_990), .C(n_991), .Y(n_989) );
AOI221xp5_ASAP7_75t_L g1008 ( .A1(n_46), .A2(n_122), .B1(n_729), .B2(n_754), .C(n_1009), .Y(n_1008) );
AOI221xp5_ASAP7_75t_L g574 ( .A1(n_47), .A2(n_106), .B1(n_575), .B2(n_577), .C(n_580), .Y(n_574) );
INVx1_ASAP7_75t_L g761 ( .A(n_48), .Y(n_761) );
AOI22xp33_ASAP7_75t_L g1183 ( .A1(n_49), .A2(n_275), .B1(n_447), .B2(n_1184), .Y(n_1183) );
INVx1_ASAP7_75t_L g1208 ( .A(n_49), .Y(n_1208) );
OAI21xp5_ASAP7_75t_L g869 ( .A1(n_50), .A2(n_699), .B(n_870), .Y(n_869) );
INVx1_ASAP7_75t_L g1716 ( .A(n_51), .Y(n_1716) );
NAND5xp2_ASAP7_75t_L g352 ( .A(n_52), .B(n_353), .C(n_435), .D(n_479), .E(n_495), .Y(n_352) );
INVx1_ASAP7_75t_L g514 ( .A(n_52), .Y(n_514) );
AOI22xp33_ASAP7_75t_SL g932 ( .A1(n_53), .A2(n_170), .B1(n_933), .B2(n_934), .Y(n_932) );
INVx1_ASAP7_75t_L g760 ( .A(n_54), .Y(n_760) );
INVx1_ASAP7_75t_L g822 ( .A(n_55), .Y(n_822) );
AOI22xp33_ASAP7_75t_L g1355 ( .A1(n_56), .A2(n_184), .B1(n_731), .B2(n_1101), .Y(n_1355) );
AOI22xp33_ASAP7_75t_SL g1374 ( .A1(n_56), .A2(n_309), .B1(n_440), .B2(n_1153), .Y(n_1374) );
INVx1_ASAP7_75t_L g1005 ( .A(n_57), .Y(n_1005) );
INVxp67_ASAP7_75t_SL g1243 ( .A(n_58), .Y(n_1243) );
AOI22xp33_ASAP7_75t_L g1263 ( .A1(n_58), .A2(n_140), .B1(n_644), .B2(n_1264), .Y(n_1263) );
AOI22xp5_ASAP7_75t_L g1434 ( .A1(n_59), .A2(n_213), .B1(n_1407), .B2(n_1412), .Y(n_1434) );
CKINVDCx5p33_ASAP7_75t_R g1706 ( .A(n_60), .Y(n_1706) );
AOI22xp5_ASAP7_75t_L g1422 ( .A1(n_61), .A2(n_321), .B1(n_1415), .B2(n_1423), .Y(n_1422) );
AOI22xp33_ASAP7_75t_L g1694 ( .A1(n_61), .A2(n_1695), .B1(n_1739), .B2(n_1741), .Y(n_1694) );
INVx1_ASAP7_75t_L g1738 ( .A(n_61), .Y(n_1738) );
BUFx6f_ASAP7_75t_L g360 ( .A(n_62), .Y(n_360) );
INVx1_ASAP7_75t_L g1131 ( .A(n_63), .Y(n_1131) );
OAI22xp33_ASAP7_75t_L g1149 ( .A1(n_63), .A2(n_108), .B1(n_546), .B2(n_1150), .Y(n_1149) );
XOR2x2_ASAP7_75t_L g1342 ( .A(n_64), .B(n_1343), .Y(n_1342) );
AOI22xp5_ASAP7_75t_L g1435 ( .A1(n_65), .A2(n_302), .B1(n_1415), .B2(n_1436), .Y(n_1435) );
INVx1_ASAP7_75t_L g1177 ( .A(n_66), .Y(n_1177) );
AOI22xp5_ASAP7_75t_L g1441 ( .A1(n_67), .A2(n_130), .B1(n_1407), .B2(n_1412), .Y(n_1441) );
INVx1_ASAP7_75t_L g630 ( .A(n_68), .Y(n_630) );
OAI222xp33_ASAP7_75t_L g663 ( .A1(n_68), .A2(n_342), .B1(n_664), .B2(n_665), .C1(n_675), .C2(n_681), .Y(n_663) );
INVx1_ASAP7_75t_L g1295 ( .A(n_69), .Y(n_1295) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_70), .A2(n_257), .B1(n_532), .B2(n_535), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g582 ( .A1(n_70), .A2(n_144), .B1(n_583), .B2(n_584), .Y(n_582) );
CKINVDCx5p33_ASAP7_75t_R g662 ( .A(n_71), .Y(n_662) );
AOI221xp5_ASAP7_75t_L g372 ( .A1(n_72), .A2(n_167), .B1(n_373), .B2(n_375), .C(n_379), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g455 ( .A1(n_72), .A2(n_237), .B1(n_451), .B2(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g1737 ( .A(n_73), .Y(n_1737) );
AOI22xp33_ASAP7_75t_L g384 ( .A1(n_74), .A2(n_237), .B1(n_371), .B2(n_385), .Y(n_384) );
AOI22xp33_ASAP7_75t_L g446 ( .A1(n_74), .A2(n_167), .B1(n_447), .B2(n_451), .Y(n_446) );
AOI221xp5_ASAP7_75t_L g1134 ( .A1(n_75), .A2(n_323), .B1(n_653), .B2(n_1115), .C(n_1135), .Y(n_1134) );
AOI22xp33_ASAP7_75t_SL g1159 ( .A1(n_75), .A2(n_289), .B1(n_802), .B2(n_941), .Y(n_1159) );
AOI22xp5_ASAP7_75t_L g844 ( .A1(n_76), .A2(n_845), .B1(n_846), .B2(n_881), .Y(n_844) );
INVxp67_ASAP7_75t_SL g881 ( .A(n_76), .Y(n_881) );
AOI221xp5_ASAP7_75t_L g890 ( .A1(n_77), .A2(n_320), .B1(n_891), .B2(n_892), .C(n_894), .Y(n_890) );
AOI221xp5_ASAP7_75t_L g936 ( .A1(n_77), .A2(n_283), .B1(n_783), .B2(n_937), .C(n_939), .Y(n_936) );
AOI22xp33_ASAP7_75t_SL g1179 ( .A1(n_78), .A2(n_173), .B1(n_783), .B2(n_1180), .Y(n_1179) );
INVxp67_ASAP7_75t_SL g1211 ( .A(n_78), .Y(n_1211) );
OAI211xp5_ASAP7_75t_SL g980 ( .A1(n_79), .A2(n_951), .B(n_958), .C(n_981), .Y(n_980) );
INVx1_ASAP7_75t_L g1015 ( .A(n_79), .Y(n_1015) );
INVx1_ASAP7_75t_L g854 ( .A(n_80), .Y(n_854) );
CKINVDCx5p33_ASAP7_75t_R g404 ( .A(n_81), .Y(n_404) );
INVxp67_ASAP7_75t_SL g926 ( .A(n_82), .Y(n_926) );
OAI22xp5_ASAP7_75t_L g943 ( .A1(n_82), .A2(n_328), .B1(n_944), .B2(n_947), .Y(n_943) );
AOI22xp33_ASAP7_75t_SL g1087 ( .A1(n_83), .A2(n_336), .B1(n_440), .B2(n_1088), .Y(n_1087) );
AOI221xp5_ASAP7_75t_L g1102 ( .A1(n_83), .A2(n_146), .B1(n_389), .B2(n_1045), .C(n_1103), .Y(n_1102) );
AOI22xp33_ASAP7_75t_L g541 ( .A1(n_84), .A2(n_106), .B1(n_530), .B2(n_542), .Y(n_541) );
INVxp67_ASAP7_75t_SL g612 ( .A(n_84), .Y(n_612) );
INVx1_ASAP7_75t_L g856 ( .A(n_85), .Y(n_856) );
OR2x2_ASAP7_75t_L g1228 ( .A(n_86), .B(n_557), .Y(n_1228) );
AOI22xp33_ASAP7_75t_L g639 ( .A1(n_87), .A2(n_134), .B1(n_640), .B2(n_644), .Y(n_639) );
OAI221xp5_ASAP7_75t_L g1239 ( .A1(n_88), .A2(n_209), .B1(n_600), .B2(n_1240), .C(n_1241), .Y(n_1239) );
OAI322xp33_ASAP7_75t_L g1250 ( .A1(n_88), .A2(n_551), .A3(n_1056), .B1(n_1251), .B2(n_1253), .C1(n_1259), .C2(n_1260), .Y(n_1250) );
AOI22xp33_ASAP7_75t_SL g1323 ( .A1(n_89), .A2(n_204), .B1(n_447), .B2(n_451), .Y(n_1323) );
AOI22xp33_ASAP7_75t_L g1334 ( .A1(n_89), .A2(n_99), .B1(n_585), .B2(n_758), .Y(n_1334) );
AOI22xp33_ASAP7_75t_SL g1043 ( .A1(n_90), .A2(n_158), .B1(n_572), .B2(n_820), .Y(n_1043) );
INVxp67_ASAP7_75t_SL g1065 ( .A(n_90), .Y(n_1065) );
INVx1_ASAP7_75t_L g1271 ( .A(n_91), .Y(n_1271) );
AOI22xp33_ASAP7_75t_SL g1279 ( .A1(n_92), .A2(n_277), .B1(n_442), .B2(n_1067), .Y(n_1279) );
AOI221xp5_ASAP7_75t_L g1291 ( .A1(n_92), .A2(n_101), .B1(n_389), .B2(n_818), .C(n_1045), .Y(n_1291) );
INVx1_ASAP7_75t_L g1215 ( .A(n_93), .Y(n_1215) );
AOI22xp5_ASAP7_75t_L g1426 ( .A1(n_94), .A2(n_335), .B1(n_1407), .B2(n_1412), .Y(n_1426) );
AOI22xp33_ASAP7_75t_L g1154 ( .A1(n_95), .A2(n_324), .B1(n_535), .B2(n_1155), .Y(n_1154) );
AOI22xp33_ASAP7_75t_L g722 ( .A1(n_96), .A2(n_267), .B1(n_440), .B2(n_442), .Y(n_722) );
AOI221xp5_ASAP7_75t_L g728 ( .A1(n_96), .A2(n_262), .B1(n_576), .B2(n_581), .C(n_729), .Y(n_728) );
OAI21xp33_ASAP7_75t_L g683 ( .A1(n_97), .A2(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g1273 ( .A(n_98), .Y(n_1273) );
AOI22xp33_ASAP7_75t_SL g1326 ( .A1(n_99), .A2(n_279), .B1(n_447), .B2(n_451), .Y(n_1326) );
INVx1_ASAP7_75t_L g712 ( .A(n_100), .Y(n_712) );
AOI22xp33_ASAP7_75t_L g730 ( .A1(n_100), .A2(n_287), .B1(n_585), .B2(n_731), .Y(n_730) );
AOI22xp33_ASAP7_75t_L g1285 ( .A1(n_101), .A2(n_191), .B1(n_783), .B2(n_1264), .Y(n_1285) );
CKINVDCx5p33_ASAP7_75t_R g1715 ( .A(n_102), .Y(n_1715) );
AOI22xp33_ASAP7_75t_L g1710 ( .A1(n_103), .A2(n_311), .B1(n_808), .B2(n_1711), .Y(n_1710) );
AOI221xp5_ASAP7_75t_L g1734 ( .A1(n_103), .A2(n_210), .B1(n_367), .B2(n_371), .C(n_1735), .Y(n_1734) );
AOI22xp33_ASAP7_75t_SL g809 ( .A1(n_104), .A2(n_313), .B1(n_440), .B2(n_442), .Y(n_809) );
INVxp67_ASAP7_75t_SL g815 ( .A(n_104), .Y(n_815) );
CKINVDCx5p33_ASAP7_75t_R g1319 ( .A(n_105), .Y(n_1319) );
XNOR2xp5_ASAP7_75t_L g748 ( .A(n_107), .B(n_749), .Y(n_748) );
AOI22xp5_ASAP7_75t_SL g1427 ( .A1(n_107), .A2(n_225), .B1(n_1415), .B2(n_1423), .Y(n_1427) );
INVx1_ASAP7_75t_L g1132 ( .A(n_108), .Y(n_1132) );
OAI211xp5_ASAP7_75t_L g392 ( .A1(n_109), .A2(n_393), .B(n_397), .C(n_401), .Y(n_392) );
INVx1_ASAP7_75t_L g510 ( .A(n_109), .Y(n_510) );
INVx1_ASAP7_75t_L g1242 ( .A(n_110), .Y(n_1242) );
AOI22xp33_ASAP7_75t_L g1049 ( .A1(n_111), .A2(n_236), .B1(n_367), .B2(n_572), .Y(n_1049) );
AOI22xp33_ASAP7_75t_L g1062 ( .A1(n_111), .A2(n_251), .B1(n_530), .B2(n_544), .Y(n_1062) );
AOI21xp33_ASAP7_75t_L g767 ( .A1(n_112), .A2(n_729), .B(n_768), .Y(n_767) );
INVx1_ASAP7_75t_L g776 ( .A(n_112), .Y(n_776) );
INVx1_ASAP7_75t_L g697 ( .A(n_113), .Y(n_697) );
INVx1_ASAP7_75t_L g1031 ( .A(n_114), .Y(n_1031) );
OAI221xp5_ASAP7_75t_L g1138 ( .A1(n_115), .A2(n_264), .B1(n_596), .B2(n_681), .C(n_1139), .Y(n_1138) );
INVx1_ASAP7_75t_L g1163 ( .A(n_115), .Y(n_1163) );
INVx1_ASAP7_75t_L g1389 ( .A(n_116), .Y(n_1389) );
AOI221xp5_ASAP7_75t_L g753 ( .A1(n_117), .A2(n_249), .B1(n_581), .B2(n_754), .C(n_755), .Y(n_753) );
AOI22xp33_ASAP7_75t_L g778 ( .A1(n_117), .A2(n_176), .B1(n_440), .B2(n_478), .Y(n_778) );
INVx1_ASAP7_75t_L g1315 ( .A(n_118), .Y(n_1315) );
INVx1_ASAP7_75t_L g1314 ( .A(n_119), .Y(n_1314) );
AOI221xp5_ASAP7_75t_L g1321 ( .A1(n_120), .A2(n_278), .B1(n_1189), .B2(n_1264), .C(n_1322), .Y(n_1321) );
AOI221xp5_ASAP7_75t_L g1333 ( .A1(n_120), .A2(n_232), .B1(n_389), .B2(n_576), .C(n_578), .Y(n_1333) );
AOI22xp33_ASAP7_75t_L g1182 ( .A1(n_121), .A2(n_182), .B1(n_447), .B2(n_808), .Y(n_1182) );
INVx1_ASAP7_75t_L g1209 ( .A(n_121), .Y(n_1209) );
INVx1_ASAP7_75t_L g996 ( .A(n_122), .Y(n_996) );
AOI22xp5_ASAP7_75t_L g1429 ( .A1(n_123), .A2(n_312), .B1(n_1412), .B2(n_1423), .Y(n_1429) );
OAI222xp33_ASAP7_75t_L g1659 ( .A1(n_124), .A2(n_319), .B1(n_954), .B2(n_956), .C1(n_1660), .C2(n_1662), .Y(n_1659) );
INVx1_ASAP7_75t_L g1672 ( .A(n_124), .Y(n_1672) );
INVx1_ASAP7_75t_L g526 ( .A(n_125), .Y(n_526) );
OAI221xp5_ASAP7_75t_L g595 ( .A1(n_125), .A2(n_126), .B1(n_596), .B2(n_600), .C(n_603), .Y(n_595) );
INVx1_ASAP7_75t_L g523 ( .A(n_126), .Y(n_523) );
OAI211xp5_ASAP7_75t_L g1033 ( .A1(n_127), .A2(n_828), .B(n_1034), .C(n_1035), .Y(n_1033) );
INVxp33_ASAP7_75t_SL g1053 ( .A(n_127), .Y(n_1053) );
INVx1_ASAP7_75t_L g1650 ( .A(n_128), .Y(n_1650) );
CKINVDCx5p33_ASAP7_75t_R g718 ( .A(n_129), .Y(n_718) );
OAI22xp33_ASAP7_75t_L g961 ( .A1(n_131), .A2(n_164), .B1(n_962), .B2(n_965), .Y(n_961) );
INVxp67_ASAP7_75t_SL g969 ( .A(n_131), .Y(n_969) );
INVxp67_ASAP7_75t_SL g1359 ( .A(n_132), .Y(n_1359) );
AOI22xp33_ASAP7_75t_L g1375 ( .A1(n_132), .A2(n_253), .B1(n_805), .B2(n_1376), .Y(n_1375) );
INVx1_ASAP7_75t_L g863 ( .A(n_133), .Y(n_863) );
INVx1_ASAP7_75t_L g673 ( .A(n_134), .Y(n_673) );
INVx1_ASAP7_75t_L g707 ( .A(n_135), .Y(n_707) );
AOI21xp33_ASAP7_75t_L g740 ( .A1(n_135), .A2(n_617), .B(n_729), .Y(n_740) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_136), .A2(n_162), .B1(n_567), .B2(n_699), .Y(n_698) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_136), .A2(n_570), .B(n_727), .C(n_733), .Y(n_726) );
INVx1_ASAP7_75t_L g1172 ( .A(n_137), .Y(n_1172) );
OAI222xp33_ASAP7_75t_L g1205 ( .A1(n_137), .A2(n_206), .B1(n_681), .B2(n_1206), .C1(n_1207), .C2(n_1210), .Y(n_1205) );
INVx1_ASAP7_75t_L g1349 ( .A(n_138), .Y(n_1349) );
OAI22xp33_ASAP7_75t_L g1381 ( .A1(n_138), .A2(n_175), .B1(n_1090), .B2(n_1150), .Y(n_1381) );
INVxp67_ASAP7_75t_SL g1353 ( .A(n_139), .Y(n_1353) );
AOI22xp33_ASAP7_75t_SL g1377 ( .A1(n_139), .A2(n_197), .B1(n_535), .B2(n_1378), .Y(n_1377) );
AOI221xp5_ASAP7_75t_L g1238 ( .A1(n_140), .A2(n_220), .B1(n_375), .B2(n_581), .C(n_1045), .Y(n_1238) );
AOI221xp5_ASAP7_75t_L g864 ( .A1(n_141), .A2(n_255), .B1(n_389), .B2(n_578), .C(n_754), .Y(n_864) );
AOI22xp33_ASAP7_75t_L g876 ( .A1(n_141), .A2(n_261), .B1(n_440), .B2(n_478), .Y(n_876) );
AOI22xp33_ASAP7_75t_SL g637 ( .A1(n_142), .A2(n_230), .B1(n_451), .B2(n_638), .Y(n_637) );
OAI22xp33_ASAP7_75t_L g979 ( .A1(n_143), .A2(n_341), .B1(n_962), .B2(n_965), .Y(n_979) );
INVxp33_ASAP7_75t_SL g1019 ( .A(n_143), .Y(n_1019) );
AOI22xp33_ASAP7_75t_L g536 ( .A1(n_144), .A2(n_172), .B1(n_532), .B2(n_535), .Y(n_536) );
CKINVDCx5p33_ASAP7_75t_R g982 ( .A(n_145), .Y(n_982) );
AOI22xp33_ASAP7_75t_SL g1082 ( .A1(n_146), .A2(n_192), .B1(n_440), .B2(n_530), .Y(n_1082) );
OA21x2_ASAP7_75t_L g1269 ( .A1(n_147), .A2(n_557), .B(n_1270), .Y(n_1269) );
INVx1_ASAP7_75t_L g986 ( .A(n_148), .Y(n_986) );
AOI221xp5_ASAP7_75t_L g1003 ( .A1(n_148), .A2(n_245), .B1(n_729), .B2(n_754), .C(n_1004), .Y(n_1003) );
AOI221xp5_ASAP7_75t_L g905 ( .A1(n_149), .A2(n_159), .B1(n_889), .B2(n_906), .C(n_908), .Y(n_905) );
AOI221xp5_ASAP7_75t_L g935 ( .A1(n_149), .A2(n_320), .B1(n_440), .B2(n_463), .C(n_530), .Y(n_935) );
AOI22xp33_ASAP7_75t_L g1083 ( .A1(n_150), .A2(n_306), .B1(n_805), .B2(n_1084), .Y(n_1083) );
AOI22xp33_ASAP7_75t_L g1099 ( .A1(n_150), .A2(n_221), .B1(n_1100), .B2(n_1101), .Y(n_1099) );
OAI22xp33_ASAP7_75t_L g545 ( .A1(n_151), .A2(n_274), .B1(n_546), .B2(n_551), .Y(n_545) );
INVx1_ASAP7_75t_L g592 ( .A(n_151), .Y(n_592) );
INVx1_ASAP7_75t_L g848 ( .A(n_152), .Y(n_848) );
INVx1_ASAP7_75t_L g1193 ( .A(n_153), .Y(n_1193) );
CKINVDCx5p33_ASAP7_75t_R g1093 ( .A(n_154), .Y(n_1093) );
OAI221xp5_ASAP7_75t_L g762 ( .A1(n_155), .A2(n_329), .B1(n_664), .B2(n_682), .C(n_763), .Y(n_762) );
OAI22xp33_ASAP7_75t_L g784 ( .A1(n_155), .A2(n_329), .B1(n_525), .B2(n_724), .Y(n_784) );
INVx1_ASAP7_75t_L g689 ( .A(n_156), .Y(n_689) );
INVx1_ASAP7_75t_L g494 ( .A(n_157), .Y(n_494) );
INVx1_ASAP7_75t_L g1061 ( .A(n_158), .Y(n_1061) );
CKINVDCx5p33_ASAP7_75t_R g1037 ( .A(n_161), .Y(n_1037) );
INVxp67_ASAP7_75t_SL g1718 ( .A(n_163), .Y(n_1718) );
INVxp67_ASAP7_75t_SL g917 ( .A(n_164), .Y(n_917) );
OAI22xp5_ASAP7_75t_L g561 ( .A1(n_165), .A2(n_188), .B1(n_562), .B2(n_567), .Y(n_561) );
OAI211xp5_ASAP7_75t_L g569 ( .A1(n_165), .A2(n_570), .B(n_573), .C(n_587), .Y(n_569) );
INVx1_ASAP7_75t_L g796 ( .A(n_166), .Y(n_796) );
INVx1_ASAP7_75t_L g1647 ( .A(n_168), .Y(n_1647) );
AOI22xp33_ASAP7_75t_L g1680 ( .A1(n_168), .A2(n_258), .B1(n_371), .B2(n_385), .Y(n_1680) );
INVx1_ASAP7_75t_L g1538 ( .A(n_169), .Y(n_1538) );
INVx1_ASAP7_75t_L g909 ( .A(n_170), .Y(n_909) );
AOI22xp5_ASAP7_75t_SL g1440 ( .A1(n_171), .A2(n_181), .B1(n_1415), .B2(n_1423), .Y(n_1440) );
AOI221xp5_ASAP7_75t_L g613 ( .A1(n_172), .A2(n_257), .B1(n_614), .B2(n_615), .C(n_617), .Y(n_613) );
AOI221xp5_ASAP7_75t_L g1198 ( .A1(n_173), .A2(n_223), .B1(n_653), .B2(n_1199), .C(n_1200), .Y(n_1198) );
CKINVDCx5p33_ASAP7_75t_R g1036 ( .A(n_174), .Y(n_1036) );
INVx1_ASAP7_75t_L g1347 ( .A(n_175), .Y(n_1347) );
AOI22xp33_ASAP7_75t_SL g769 ( .A1(n_176), .A2(n_301), .B1(n_572), .B2(n_583), .Y(n_769) );
OAI211xp5_ASAP7_75t_L g751 ( .A1(n_177), .A2(n_570), .B(n_752), .C(n_759), .Y(n_751) );
OAI22xp5_ASAP7_75t_L g787 ( .A1(n_177), .A2(n_322), .B1(n_567), .B2(n_699), .Y(n_787) );
INVx1_ASAP7_75t_L g1047 ( .A(n_178), .Y(n_1047) );
INVx1_ASAP7_75t_L g1278 ( .A(n_179), .Y(n_1278) );
AOI221xp5_ASAP7_75t_L g1304 ( .A1(n_179), .A2(n_226), .B1(n_578), .B2(n_1305), .C(n_1308), .Y(n_1304) );
OAI211xp5_ASAP7_75t_L g354 ( .A1(n_180), .A2(n_355), .B(n_365), .C(n_391), .Y(n_354) );
NOR2xp33_ASAP7_75t_L g417 ( .A(n_180), .B(n_418), .Y(n_417) );
XNOR2x2_ASAP7_75t_L g1074 ( .A(n_181), .B(n_1075), .Y(n_1074) );
AOI22xp33_ASAP7_75t_L g1201 ( .A1(n_182), .A2(n_275), .B1(n_1100), .B2(n_1202), .Y(n_1201) );
AOI221xp5_ASAP7_75t_L g1324 ( .A1(n_183), .A2(n_232), .B1(n_783), .B2(n_1264), .C(n_1325), .Y(n_1324) );
AOI22xp33_ASAP7_75t_L g1336 ( .A1(n_183), .A2(n_278), .B1(n_585), .B2(n_820), .Y(n_1336) );
AOI22xp33_ASAP7_75t_SL g1380 ( .A1(n_184), .A2(n_338), .B1(n_440), .B2(n_802), .Y(n_1380) );
INVx2_ASAP7_75t_L g1410 ( .A(n_185), .Y(n_1410) );
AND2x2_ASAP7_75t_L g1413 ( .A(n_185), .B(n_1411), .Y(n_1413) );
AND2x2_ASAP7_75t_L g1418 ( .A(n_185), .B(n_288), .Y(n_1418) );
AOI22xp33_ASAP7_75t_L g803 ( .A1(n_186), .A2(n_333), .B1(n_804), .B2(n_805), .Y(n_803) );
INVx1_ASAP7_75t_L g831 ( .A(n_186), .Y(n_831) );
CKINVDCx5p33_ASAP7_75t_R g1249 ( .A(n_187), .Y(n_1249) );
INVx1_ASAP7_75t_L g736 ( .A(n_189), .Y(n_736) );
AOI22xp5_ASAP7_75t_SL g1460 ( .A1(n_190), .A2(n_252), .B1(n_1412), .B2(n_1417), .Y(n_1460) );
INVx1_ASAP7_75t_L g1303 ( .A(n_191), .Y(n_1303) );
INVxp67_ASAP7_75t_SL g1110 ( .A(n_192), .Y(n_1110) );
XOR2x2_ASAP7_75t_L g518 ( .A(n_194), .B(n_519), .Y(n_518) );
AOI22xp5_ASAP7_75t_L g1414 ( .A1(n_194), .A2(n_310), .B1(n_1415), .B2(n_1417), .Y(n_1414) );
OAI22xp33_ASAP7_75t_L g1089 ( .A1(n_195), .A2(n_260), .B1(n_551), .B2(n_1090), .Y(n_1089) );
INVx1_ASAP7_75t_L g1106 ( .A(n_195), .Y(n_1106) );
AOI22xp5_ASAP7_75t_L g1421 ( .A1(n_196), .A2(n_256), .B1(n_1407), .B2(n_1412), .Y(n_1421) );
INVxp67_ASAP7_75t_SL g1360 ( .A(n_197), .Y(n_1360) );
INVx1_ASAP7_75t_L g1687 ( .A(n_198), .Y(n_1687) );
NOR2xp33_ASAP7_75t_L g1362 ( .A(n_199), .B(n_664), .Y(n_1362) );
INVx1_ASAP7_75t_L g1372 ( .A(n_199), .Y(n_1372) );
INVx1_ASAP7_75t_L g1192 ( .A(n_200), .Y(n_1192) );
AOI22xp33_ASAP7_75t_L g366 ( .A1(n_201), .A2(n_272), .B1(n_367), .B2(n_371), .Y(n_366) );
AOI22xp33_ASAP7_75t_SL g457 ( .A1(n_201), .A2(n_286), .B1(n_440), .B2(n_458), .Y(n_457) );
AOI22xp33_ASAP7_75t_SL g713 ( .A1(n_202), .A2(n_262), .B1(n_440), .B2(n_442), .Y(n_713) );
AOI22xp33_ASAP7_75t_SL g741 ( .A1(n_202), .A2(n_267), .B1(n_583), .B2(n_742), .Y(n_741) );
INVx1_ASAP7_75t_L g842 ( .A(n_203), .Y(n_842) );
AOI221xp5_ASAP7_75t_L g1337 ( .A1(n_204), .A2(n_279), .B1(n_578), .B2(n_617), .C(n_754), .Y(n_1337) );
INVx1_ASAP7_75t_L g1284 ( .A(n_205), .Y(n_1284) );
AOI22xp33_ASAP7_75t_L g1292 ( .A1(n_205), .A2(n_266), .B1(n_371), .B2(n_1293), .Y(n_1292) );
INVx1_ASAP7_75t_L g1174 ( .A(n_206), .Y(n_1174) );
INVx1_ASAP7_75t_L g633 ( .A(n_207), .Y(n_633) );
OAI211xp5_ASAP7_75t_L g650 ( .A1(n_207), .A2(n_570), .B(n_651), .C(n_659), .Y(n_650) );
AOI22xp5_ASAP7_75t_L g1430 ( .A1(n_208), .A2(n_271), .B1(n_1407), .B2(n_1415), .Y(n_1430) );
INVx1_ASAP7_75t_L g1224 ( .A(n_209), .Y(n_1224) );
AOI22xp33_ASAP7_75t_L g1700 ( .A1(n_210), .A2(n_293), .B1(n_535), .B2(n_1701), .Y(n_1700) );
CKINVDCx5p33_ASAP7_75t_R g1649 ( .A(n_211), .Y(n_1649) );
INVx1_ASAP7_75t_L g1227 ( .A(n_212), .Y(n_1227) );
CKINVDCx5p33_ASAP7_75t_R g764 ( .A(n_214), .Y(n_764) );
INVx1_ASAP7_75t_L g1265 ( .A(n_215), .Y(n_1265) );
CKINVDCx5p33_ASAP7_75t_R g407 ( .A(n_216), .Y(n_407) );
INVx2_ASAP7_75t_L g430 ( .A(n_217), .Y(n_430) );
INVx1_ASAP7_75t_L g464 ( .A(n_217), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_217), .B(n_428), .Y(n_488) );
CKINVDCx5p33_ASAP7_75t_R g660 ( .A(n_218), .Y(n_660) );
INVx1_ASAP7_75t_L g1657 ( .A(n_219), .Y(n_1657) );
NAND2xp33_ASAP7_75t_SL g1681 ( .A(n_219), .B(n_373), .Y(n_1681) );
INVx1_ASAP7_75t_L g1257 ( .A(n_220), .Y(n_1257) );
AOI22xp33_ASAP7_75t_L g807 ( .A1(n_222), .A2(n_303), .B1(n_448), .B2(n_808), .Y(n_807) );
INVx1_ASAP7_75t_L g829 ( .A(n_222), .Y(n_829) );
AOI22xp33_ASAP7_75t_SL g801 ( .A1(n_224), .A2(n_247), .B1(n_440), .B2(n_802), .Y(n_801) );
INVxp67_ASAP7_75t_SL g833 ( .A(n_224), .Y(n_833) );
INVx1_ASAP7_75t_L g1283 ( .A(n_226), .Y(n_1283) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_227), .A2(n_292), .B1(n_393), .B2(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g504 ( .A(n_227), .Y(n_504) );
INVx1_ASAP7_75t_L g668 ( .A(n_228), .Y(n_668) );
INVx1_ASAP7_75t_L g1237 ( .A(n_229), .Y(n_1237) );
INVx1_ASAP7_75t_L g676 ( .A(n_230), .Y(n_676) );
AOI21xp5_ASAP7_75t_L g1658 ( .A1(n_231), .A2(n_463), .B(n_942), .Y(n_1658) );
OAI21xp5_ASAP7_75t_L g839 ( .A1(n_233), .A2(n_699), .B(n_840), .Y(n_839) );
INVx1_ASAP7_75t_L g1683 ( .A(n_234), .Y(n_1683) );
BUFx3_ASAP7_75t_L g422 ( .A(n_235), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g1066 ( .A1(n_236), .A2(n_268), .B1(n_530), .B2(n_1067), .Y(n_1066) );
INVx1_ASAP7_75t_L g1331 ( .A(n_238), .Y(n_1331) );
CKINVDCx5p33_ASAP7_75t_R g983 ( .A(n_239), .Y(n_983) );
AOI22xp5_ASAP7_75t_L g1406 ( .A1(n_240), .A2(n_269), .B1(n_1407), .B2(n_1412), .Y(n_1406) );
INVx1_ASAP7_75t_L g1640 ( .A(n_241), .Y(n_1640) );
NOR2xp33_ASAP7_75t_L g1642 ( .A(n_241), .B(n_962), .Y(n_1642) );
INVx1_ASAP7_75t_L g1736 ( .A(n_242), .Y(n_1736) );
AOI21xp33_ASAP7_75t_L g1048 ( .A1(n_243), .A2(n_379), .B(n_729), .Y(n_1048) );
INVx1_ASAP7_75t_L g1059 ( .A(n_243), .Y(n_1059) );
INVx1_ASAP7_75t_L g1079 ( .A(n_244), .Y(n_1079) );
AOI21xp33_ASAP7_75t_L g999 ( .A1(n_245), .A2(n_643), .B(n_939), .Y(n_999) );
XOR2x2_ASAP7_75t_L g1026 ( .A(n_246), .B(n_1027), .Y(n_1026) );
AOI21xp33_ASAP7_75t_L g817 ( .A1(n_247), .A2(n_389), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g364 ( .A(n_248), .Y(n_364) );
BUFx3_ASAP7_75t_L g382 ( .A(n_248), .Y(n_382) );
AOI22xp33_ASAP7_75t_L g782 ( .A1(n_249), .A2(n_301), .B1(n_440), .B2(n_783), .Y(n_782) );
XNOR2x1_ASAP7_75t_L g1311 ( .A(n_250), .B(n_1312), .Y(n_1311) );
NAND2xp5_ASAP7_75t_SL g1042 ( .A(n_251), .B(n_729), .Y(n_1042) );
AOI21xp5_ASAP7_75t_L g1356 ( .A1(n_253), .A2(n_379), .B(n_1357), .Y(n_1356) );
CKINVDCx5p33_ASAP7_75t_R g988 ( .A(n_254), .Y(n_988) );
INVx1_ASAP7_75t_L g1655 ( .A(n_258), .Y(n_1655) );
INVx1_ASAP7_75t_L g1330 ( .A(n_259), .Y(n_1330) );
INVx1_ASAP7_75t_L g1107 ( .A(n_260), .Y(n_1107) );
INVx1_ASAP7_75t_L g1235 ( .A(n_263), .Y(n_1235) );
INVx1_ASAP7_75t_L g1161 ( .A(n_264), .Y(n_1161) );
INVx1_ASAP7_75t_L g734 ( .A(n_265), .Y(n_734) );
NAND2xp33_ASAP7_75t_SL g1280 ( .A(n_266), .B(n_808), .Y(n_1280) );
NAND2xp5_ASAP7_75t_SL g1044 ( .A(n_268), .B(n_1045), .Y(n_1044) );
INVx1_ASAP7_75t_L g970 ( .A(n_270), .Y(n_970) );
AOI22xp33_ASAP7_75t_SL g439 ( .A1(n_272), .A2(n_343), .B1(n_440), .B2(n_442), .Y(n_439) );
INVx1_ASAP7_75t_L g425 ( .A(n_273), .Y(n_425) );
INVx1_ASAP7_75t_L g445 ( .A(n_273), .Y(n_445) );
INVx1_ASAP7_75t_L g588 ( .A(n_274), .Y(n_588) );
INVx1_ASAP7_75t_L g1300 ( .A(n_277), .Y(n_1300) );
INVx1_ASAP7_75t_L g680 ( .A(n_280), .Y(n_680) );
OAI21xp33_ASAP7_75t_L g1051 ( .A1(n_281), .A2(n_481), .B(n_1052), .Y(n_1051) );
INVx1_ASAP7_75t_L g799 ( .A(n_282), .Y(n_799) );
INVx1_ASAP7_75t_L g910 ( .A(n_283), .Y(n_910) );
CKINVDCx5p33_ASAP7_75t_R g1639 ( .A(n_284), .Y(n_1639) );
CKINVDCx5p33_ASAP7_75t_R g1318 ( .A(n_285), .Y(n_1318) );
AOI221xp5_ASAP7_75t_SL g387 ( .A1(n_286), .A2(n_343), .B1(n_373), .B2(n_388), .C(n_389), .Y(n_387) );
INVx1_ASAP7_75t_L g721 ( .A(n_287), .Y(n_721) );
INVx1_ASAP7_75t_L g1411 ( .A(n_288), .Y(n_1411) );
AND2x2_ASAP7_75t_L g1416 ( .A(n_288), .B(n_1410), .Y(n_1416) );
INVxp67_ASAP7_75t_SL g1143 ( .A(n_289), .Y(n_1143) );
OAI211xp5_ASAP7_75t_SL g1351 ( .A1(n_290), .A2(n_600), .B(n_1352), .C(n_1358), .Y(n_1351) );
INVx1_ASAP7_75t_L g1371 ( .A(n_290), .Y(n_1371) );
INVx1_ASAP7_75t_L g868 ( .A(n_291), .Y(n_868) );
INVx1_ASAP7_75t_L g476 ( .A(n_292), .Y(n_476) );
INVx1_ASAP7_75t_L g1723 ( .A(n_293), .Y(n_1723) );
XNOR2xp5_ASAP7_75t_L g971 ( .A(n_294), .B(n_972), .Y(n_971) );
OAI211xp5_ASAP7_75t_L g1096 ( .A1(n_296), .A2(n_1097), .B(n_1098), .C(n_1105), .Y(n_1096) );
INVxp67_ASAP7_75t_SL g1261 ( .A(n_297), .Y(n_1261) );
INVx1_ASAP7_75t_L g867 ( .A(n_298), .Y(n_867) );
INVx1_ASAP7_75t_L g1540 ( .A(n_299), .Y(n_1540) );
CKINVDCx16_ASAP7_75t_R g1661 ( .A(n_300), .Y(n_1661) );
AOI22xp5_ASAP7_75t_L g819 ( .A1(n_303), .A2(n_333), .B1(n_585), .B2(n_820), .Y(n_819) );
OAI21xp33_ASAP7_75t_L g1190 ( .A1(n_304), .A2(n_562), .B(n_1191), .Y(n_1190) );
INVx1_ASAP7_75t_L g974 ( .A(n_305), .Y(n_974) );
OAI21xp5_ASAP7_75t_SL g1338 ( .A1(n_307), .A2(n_699), .B(n_1339), .Y(n_1338) );
INVx1_ASAP7_75t_L g994 ( .A(n_308), .Y(n_994) );
AOI221xp5_ASAP7_75t_L g1361 ( .A1(n_309), .A2(n_338), .B1(n_581), .B2(n_1115), .C(n_1117), .Y(n_1361) );
INVx1_ASAP7_75t_L g1722 ( .A(n_311), .Y(n_1722) );
INVxp67_ASAP7_75t_SL g837 ( .A(n_313), .Y(n_837) );
INVxp67_ASAP7_75t_SL g1142 ( .A(n_314), .Y(n_1142) );
AOI22xp33_ASAP7_75t_SL g1152 ( .A1(n_314), .A2(n_323), .B1(n_544), .B2(n_1153), .Y(n_1152) );
BUFx6f_ASAP7_75t_L g362 ( .A(n_316), .Y(n_362) );
INVx1_ASAP7_75t_L g781 ( .A(n_317), .Y(n_781) );
INVx1_ASAP7_75t_L g1366 ( .A(n_318), .Y(n_1366) );
NOR2xp33_ASAP7_75t_R g1674 ( .A(n_319), .B(n_1675), .Y(n_1674) );
INVxp67_ASAP7_75t_SL g924 ( .A(n_325), .Y(n_924) );
OAI221xp5_ASAP7_75t_L g953 ( .A1(n_325), .A2(n_327), .B1(n_954), .B2(n_956), .C(n_958), .Y(n_953) );
INVx1_ASAP7_75t_L g786 ( .A(n_326), .Y(n_786) );
OAI221xp5_ASAP7_75t_L g896 ( .A1(n_327), .A2(n_328), .B1(n_897), .B2(n_902), .C(n_903), .Y(n_896) );
INVx2_ASAP7_75t_L g416 ( .A(n_330), .Y(n_416) );
INVx1_ASAP7_75t_L g434 ( .A(n_330), .Y(n_434) );
INVx1_ASAP7_75t_L g469 ( .A(n_330), .Y(n_469) );
CKINVDCx5p33_ASAP7_75t_R g560 ( .A(n_332), .Y(n_560) );
INVx1_ASAP7_75t_L g1006 ( .A(n_334), .Y(n_1006) );
INVxp67_ASAP7_75t_SL g1113 ( .A(n_336), .Y(n_1113) );
OAI22xp33_ASAP7_75t_SL g723 ( .A1(n_337), .A2(n_340), .B1(n_525), .B2(n_724), .Y(n_723) );
OAI221xp5_ASAP7_75t_L g737 ( .A1(n_337), .A2(n_340), .B1(n_596), .B2(n_682), .C(n_738), .Y(n_737) );
XNOR2xp5_ASAP7_75t_L g694 ( .A(n_339), .B(n_695), .Y(n_694) );
INVxp67_ASAP7_75t_SL g977 ( .A(n_341), .Y(n_977) );
INVx1_ASAP7_75t_L g629 ( .A(n_342), .Y(n_629) );
AOI21xp5_ASAP7_75t_L g344 ( .A1(n_345), .A2(n_1384), .B(n_1399), .Y(n_344) );
XNOR2xp5_ASAP7_75t_L g345 ( .A(n_346), .B(n_619), .Y(n_345) );
HB1xp67_ASAP7_75t_L g346 ( .A(n_347), .Y(n_346) );
XNOR2xp5_ASAP7_75t_L g347 ( .A(n_348), .B(n_518), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
NAND3xp33_ASAP7_75t_L g351 ( .A(n_352), .B(n_511), .C(n_515), .Y(n_351) );
INVx1_ASAP7_75t_L g512 ( .A(n_353), .Y(n_512) );
AOI21x1_ASAP7_75t_L g353 ( .A1(n_354), .A2(n_414), .B(n_417), .Y(n_353) );
INVx2_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
AOI221xp5_ASAP7_75t_L g862 ( .A1(n_356), .A2(n_586), .B1(n_863), .B2(n_864), .C(n_865), .Y(n_862) );
AOI221xp5_ASAP7_75t_L g1290 ( .A1(n_356), .A2(n_586), .B1(n_1273), .B2(n_1291), .C(n_1292), .Y(n_1290) );
AOI221xp5_ASAP7_75t_L g1332 ( .A1(n_356), .A2(n_586), .B1(n_1314), .B2(n_1333), .C(n_1334), .Y(n_1332) );
AND2x2_ASAP7_75t_L g356 ( .A(n_357), .B(n_363), .Y(n_356) );
AND2x4_ASAP7_75t_L g918 ( .A(n_357), .B(n_919), .Y(n_918) );
INVx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g742 ( .A(n_358), .Y(n_742) );
INVx2_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
BUFx3_ASAP7_75t_L g371 ( .A(n_359), .Y(n_371) );
BUFx6f_ASAP7_75t_L g572 ( .A(n_359), .Y(n_572) );
BUFx3_ASAP7_75t_L g585 ( .A(n_359), .Y(n_585) );
AND2x2_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g370 ( .A(n_360), .Y(n_370) );
AND2x2_ASAP7_75t_L g374 ( .A(n_360), .B(n_362), .Y(n_374) );
INVx2_ASAP7_75t_L g378 ( .A(n_360), .Y(n_378) );
OR2x2_ASAP7_75t_L g396 ( .A(n_360), .B(n_362), .Y(n_396) );
NAND2x1_ASAP7_75t_L g400 ( .A(n_360), .B(n_362), .Y(n_400) );
BUFx2_ASAP7_75t_L g403 ( .A(n_360), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_360), .B(n_361), .Y(n_611) );
OR2x2_ASAP7_75t_L g672 ( .A(n_360), .B(n_369), .Y(n_672) );
INVx2_ASAP7_75t_L g361 ( .A(n_362), .Y(n_361) );
INVx2_ASAP7_75t_L g369 ( .A(n_362), .Y(n_369) );
AND2x2_ASAP7_75t_L g377 ( .A(n_362), .B(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g566 ( .A(n_362), .Y(n_566) );
BUFx2_ASAP7_75t_L g411 ( .A(n_363), .Y(n_411) );
AND2x2_ASAP7_75t_L g492 ( .A(n_363), .B(n_493), .Y(n_492) );
AND2x4_ASAP7_75t_L g571 ( .A(n_363), .B(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g591 ( .A(n_363), .B(n_368), .Y(n_591) );
AND2x4_ASAP7_75t_L g594 ( .A(n_363), .B(n_493), .Y(n_594) );
AND2x4_ASAP7_75t_SL g599 ( .A(n_363), .B(n_373), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g920 ( .A(n_363), .B(n_469), .Y(n_920) );
AOI22xp5_ASAP7_75t_L g365 ( .A1(n_366), .A2(n_372), .B1(n_384), .B2(n_387), .Y(n_365) );
BUFx6f_ASAP7_75t_L g656 ( .A(n_367), .Y(n_656) );
INVx3_ASAP7_75t_L g732 ( .A(n_367), .Y(n_732) );
A2O1A1Ixp33_ASAP7_75t_L g1731 ( .A1(n_367), .A2(n_408), .B(n_1708), .C(n_1732), .Y(n_1731) );
BUFx6f_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
INVx3_ASAP7_75t_L g386 ( .A(n_368), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g559 ( .A(n_368), .B(n_410), .Y(n_559) );
AND2x2_ASAP7_75t_L g368 ( .A(n_369), .B(n_370), .Y(n_368) );
HB1xp67_ASAP7_75t_L g406 ( .A(n_369), .Y(n_406) );
BUFx6f_ASAP7_75t_L g576 ( .A(n_373), .Y(n_576) );
AND2x6_ASAP7_75t_L g586 ( .A(n_373), .B(n_410), .Y(n_586) );
BUFx3_ASAP7_75t_L g614 ( .A(n_373), .Y(n_614) );
BUFx3_ASAP7_75t_L g754 ( .A(n_373), .Y(n_754) );
BUFx3_ASAP7_75t_L g1045 ( .A(n_373), .Y(n_1045) );
BUFx3_ASAP7_75t_L g1117 ( .A(n_373), .Y(n_1117) );
INVx1_ASAP7_75t_L g1136 ( .A(n_373), .Y(n_1136) );
BUFx6f_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g860 ( .A(n_374), .Y(n_860) );
INVx2_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
INVx2_ASAP7_75t_L g388 ( .A(n_376), .Y(n_388) );
INVx2_ASAP7_75t_L g376 ( .A(n_377), .Y(n_376) );
BUFx6f_ASAP7_75t_L g493 ( .A(n_377), .Y(n_493) );
BUFx3_ASAP7_75t_L g729 ( .A(n_377), .Y(n_729) );
INVx3_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
INVx2_ASAP7_75t_L g617 ( .A(n_380), .Y(n_617) );
INVx1_ASAP7_75t_L g768 ( .A(n_380), .Y(n_768) );
OAI221xp5_ASAP7_75t_L g1207 ( .A1(n_380), .A2(n_669), .B1(n_893), .B2(n_1208), .C(n_1209), .Y(n_1207) );
INVx2_ASAP7_75t_L g1308 ( .A(n_380), .Y(n_1308) );
OAI221xp5_ASAP7_75t_L g1721 ( .A1(n_380), .A2(n_397), .B1(n_1722), .B2(n_1723), .C(n_1724), .Y(n_1721) );
AND2x4_ASAP7_75t_L g380 ( .A(n_381), .B(n_383), .Y(n_380) );
INVxp67_ASAP7_75t_L g1398 ( .A(n_381), .Y(n_1398) );
INVx2_ASAP7_75t_L g381 ( .A(n_382), .Y(n_381) );
AND2x4_ASAP7_75t_L g390 ( .A(n_382), .B(n_383), .Y(n_390) );
INVx1_ASAP7_75t_L g1395 ( .A(n_383), .Y(n_1395) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
INVx2_ASAP7_75t_SL g583 ( .A(n_386), .Y(n_583) );
INVx2_ASAP7_75t_L g758 ( .A(n_386), .Y(n_758) );
INVx1_ASAP7_75t_L g820 ( .A(n_386), .Y(n_820) );
INVx2_ASAP7_75t_L g1100 ( .A(n_386), .Y(n_1100) );
INVx2_ASAP7_75t_L g616 ( .A(n_388), .Y(n_616) );
INVx1_ASAP7_75t_L g1116 ( .A(n_388), .Y(n_1116) );
INVx4_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx4_ASAP7_75t_L g581 ( .A(n_390), .Y(n_581) );
INVx1_ASAP7_75t_SL g653 ( .A(n_390), .Y(n_653) );
AND2x2_ASAP7_75t_SL g895 ( .A(n_390), .B(n_487), .Y(n_895) );
AND2x4_ASAP7_75t_L g1011 ( .A(n_390), .B(n_1012), .Y(n_1011) );
NAND4xp25_ASAP7_75t_L g1041 ( .A(n_390), .B(n_1042), .C(n_1043), .D(n_1044), .Y(n_1041) );
OAI221xp5_ASAP7_75t_L g1735 ( .A1(n_390), .A2(n_399), .B1(n_830), .B2(n_1736), .C(n_1737), .Y(n_1735) );
AOI22xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_408), .B1(n_411), .B2(n_412), .Y(n_391) );
INVx3_ASAP7_75t_L g393 ( .A(n_394), .Y(n_393) );
BUFx6f_ASAP7_75t_L g605 ( .A(n_394), .Y(n_605) );
INVx4_ASAP7_75t_L g1034 ( .A(n_394), .Y(n_1034) );
BUFx4f_ASAP7_75t_L g394 ( .A(n_395), .Y(n_394) );
INVx3_ASAP7_75t_L g678 ( .A(n_395), .Y(n_678) );
INVx2_ASAP7_75t_L g836 ( .A(n_395), .Y(n_836) );
INVx3_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
INVx2_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g739 ( .A(n_398), .Y(n_739) );
INVx2_ASAP7_75t_L g828 ( .A(n_398), .Y(n_828) );
INVx4_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
BUFx4f_ASAP7_75t_L g413 ( .A(n_399), .Y(n_413) );
BUFx4f_ASAP7_75t_L g816 ( .A(n_399), .Y(n_816) );
BUFx4f_ASAP7_75t_L g893 ( .A(n_399), .Y(n_893) );
OR2x6_ASAP7_75t_L g903 ( .A(n_399), .B(n_904), .Y(n_903) );
BUFx4f_ASAP7_75t_L g1354 ( .A(n_399), .Y(n_1354) );
BUFx6f_ASAP7_75t_L g399 ( .A(n_400), .Y(n_399) );
BUFx3_ASAP7_75t_L g667 ( .A(n_400), .Y(n_667) );
AOI22xp5_ASAP7_75t_L g401 ( .A1(n_402), .A2(n_404), .B1(n_405), .B2(n_407), .Y(n_401) );
AND2x2_ASAP7_75t_L g853 ( .A(n_402), .B(n_410), .Y(n_853) );
AOI22xp33_ASAP7_75t_L g1035 ( .A1(n_402), .A2(n_405), .B1(n_1036), .B2(n_1037), .Y(n_1035) );
AOI22xp5_ASAP7_75t_L g1733 ( .A1(n_402), .A2(n_405), .B1(n_1706), .B2(n_1715), .Y(n_1733) );
BUFx2_ASAP7_75t_L g402 ( .A(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g602 ( .A(n_403), .Y(n_602) );
INVx1_ASAP7_75t_L g901 ( .A(n_403), .Y(n_901) );
AOI221xp5_ASAP7_75t_L g465 ( .A1(n_404), .A2(n_466), .B1(n_472), .B2(n_476), .C(n_477), .Y(n_465) );
INVx1_ASAP7_75t_L g405 ( .A(n_406), .Y(n_405) );
AOI222xp33_ASAP7_75t_L g495 ( .A1(n_407), .A2(n_496), .B1(n_501), .B2(n_504), .C1(n_505), .C2(n_510), .Y(n_495) );
AOI22xp5_ASAP7_75t_L g1032 ( .A1(n_408), .A2(n_411), .B1(n_1033), .B2(n_1038), .Y(n_1032) );
INVx1_ASAP7_75t_L g408 ( .A(n_409), .Y(n_408) );
NOR2x1_ASAP7_75t_L g601 ( .A(n_409), .B(n_602), .Y(n_601) );
INVx1_ASAP7_75t_L g409 ( .A(n_410), .Y(n_409) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_410), .B(n_565), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g899 ( .A(n_410), .B(n_416), .Y(n_899) );
INVxp67_ASAP7_75t_L g1727 ( .A(n_411), .Y(n_1727) );
BUFx2_ASAP7_75t_L g770 ( .A(n_414), .Y(n_770) );
BUFx2_ASAP7_75t_L g967 ( .A(n_414), .Y(n_967) );
OAI31xp33_ASAP7_75t_L g1719 ( .A1(n_414), .A2(n_1720), .A3(n_1726), .B(n_1734), .Y(n_1719) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
AND3x4_ASAP7_75t_L g437 ( .A(n_415), .B(n_430), .C(n_438), .Y(n_437) );
INVx2_ASAP7_75t_SL g618 ( .A(n_415), .Y(n_618) );
OAI31xp33_ASAP7_75t_SL g978 ( .A1(n_415), .A2(n_979), .A3(n_980), .B(n_984), .Y(n_978) );
OAI31xp33_ASAP7_75t_L g1641 ( .A1(n_415), .A2(n_1642), .A3(n_1643), .B(n_1659), .Y(n_1641) );
INVx2_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
BUFx2_ASAP7_75t_L g462 ( .A(n_416), .Y(n_462) );
INVx5_ASAP7_75t_L g634 ( .A(n_418), .Y(n_634) );
INVx3_ASAP7_75t_L g872 ( .A(n_418), .Y(n_872) );
OR2x6_ASAP7_75t_L g418 ( .A(n_419), .B(n_431), .Y(n_418) );
OR2x2_ASAP7_75t_L g567 ( .A(n_419), .B(n_431), .Y(n_567) );
INVx2_ASAP7_75t_L g952 ( .A(n_419), .Y(n_952) );
NAND2x1p5_ASAP7_75t_L g419 ( .A(n_420), .B(n_426), .Y(n_419) );
INVx8_ASAP7_75t_L g441 ( .A(n_420), .Y(n_441) );
BUFx3_ASAP7_75t_L g544 ( .A(n_420), .Y(n_544) );
BUFx3_ASAP7_75t_L g942 ( .A(n_420), .Y(n_942) );
AND2x2_ASAP7_75t_L g945 ( .A(n_420), .B(n_946), .Y(n_945) );
HB1xp67_ASAP7_75t_L g1067 ( .A(n_420), .Y(n_1067) );
AND2x4_ASAP7_75t_L g420 ( .A(n_421), .B(n_423), .Y(n_420) );
AND2x4_ASAP7_75t_L g449 ( .A(n_421), .B(n_450), .Y(n_449) );
INVx2_ASAP7_75t_L g421 ( .A(n_422), .Y(n_421) );
AND2x4_ASAP7_75t_L g443 ( .A(n_422), .B(n_444), .Y(n_443) );
BUFx6f_ASAP7_75t_L g453 ( .A(n_422), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g509 ( .A(n_422), .B(n_445), .Y(n_509) );
OR2x2_ASAP7_75t_L g549 ( .A(n_422), .B(n_424), .Y(n_549) );
INVx1_ASAP7_75t_L g423 ( .A(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g424 ( .A(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_L g450 ( .A(n_425), .Y(n_450) );
AND2x4_ASAP7_75t_L g467 ( .A(n_426), .B(n_468), .Y(n_467) );
AND2x6_ASAP7_75t_L g955 ( .A(n_426), .B(n_470), .Y(n_955) );
AND2x2_ASAP7_75t_L g957 ( .A(n_426), .B(n_475), .Y(n_957) );
INVx1_ASAP7_75t_L g960 ( .A(n_426), .Y(n_960) );
AND2x4_ASAP7_75t_L g426 ( .A(n_427), .B(n_429), .Y(n_426) );
NAND2x1p5_ASAP7_75t_L g463 ( .A(n_427), .B(n_464), .Y(n_463) );
NAND3x1_ASAP7_75t_L g539 ( .A(n_427), .B(n_464), .C(n_540), .Y(n_539) );
INVx3_ASAP7_75t_L g427 ( .A(n_428), .Y(n_427) );
BUFx3_ASAP7_75t_L g438 ( .A(n_428), .Y(n_438) );
NAND2xp33_ASAP7_75t_SL g705 ( .A(n_428), .B(n_430), .Y(n_705) );
INVx1_ASAP7_75t_L g429 ( .A(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g1651 ( .A(n_430), .B(n_438), .Y(n_1651) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g491 ( .A(n_432), .Y(n_491) );
OR2x2_ASAP7_75t_L g563 ( .A(n_432), .B(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g902 ( .A(n_432), .B(n_564), .Y(n_902) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
INVx2_ASAP7_75t_L g487 ( .A(n_433), .Y(n_487) );
INVx1_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
INVx1_ASAP7_75t_L g513 ( .A(n_435), .Y(n_513) );
AND2x2_ASAP7_75t_L g435 ( .A(n_436), .B(n_465), .Y(n_435) );
AOI33xp33_ASAP7_75t_L g436 ( .A1(n_437), .A2(n_439), .A3(n_446), .B1(n_455), .B2(n_457), .B3(n_460), .Y(n_436) );
AOI33xp33_ASAP7_75t_L g528 ( .A1(n_437), .A2(n_529), .A3(n_531), .B1(n_536), .B2(n_537), .B3(n_541), .Y(n_528) );
BUFx3_ASAP7_75t_L g636 ( .A(n_437), .Y(n_636) );
AOI33xp33_ASAP7_75t_L g800 ( .A1(n_437), .A2(n_801), .A3(n_803), .B1(n_807), .B2(n_809), .B3(n_810), .Y(n_800) );
AOI33xp33_ASAP7_75t_L g875 ( .A1(n_437), .A2(n_876), .A3(n_877), .B1(n_878), .B2(n_879), .B3(n_880), .Y(n_875) );
AOI33xp33_ASAP7_75t_L g1081 ( .A1(n_437), .A2(n_537), .A3(n_1082), .B1(n_1083), .B2(n_1086), .B3(n_1087), .Y(n_1081) );
AOI33xp33_ASAP7_75t_L g1151 ( .A1(n_437), .A2(n_1152), .A3(n_1154), .B1(n_1157), .B2(n_1158), .B3(n_1159), .Y(n_1151) );
INVx1_ASAP7_75t_L g1325 ( .A(n_437), .Y(n_1325) );
AOI33xp33_ASAP7_75t_L g1373 ( .A1(n_437), .A2(n_537), .A3(n_1374), .B1(n_1375), .B2(n_1377), .B3(n_1380), .Y(n_1373) );
NAND3xp33_ASAP7_75t_L g1699 ( .A(n_437), .B(n_1700), .C(n_1702), .Y(n_1699) );
BUFx2_ASAP7_75t_L g647 ( .A(n_440), .Y(n_647) );
INVx8_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx2_ASAP7_75t_L g502 ( .A(n_441), .Y(n_502) );
INVx3_ASAP7_75t_L g638 ( .A(n_441), .Y(n_638) );
CKINVDCx5p33_ASAP7_75t_R g990 ( .A(n_441), .Y(n_990) );
INVx2_ASAP7_75t_L g1264 ( .A(n_441), .Y(n_1264) );
BUFx2_ASAP7_75t_L g442 ( .A(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g459 ( .A(n_443), .Y(n_459) );
BUFx2_ASAP7_75t_L g478 ( .A(n_443), .Y(n_478) );
BUFx3_ASAP7_75t_L g530 ( .A(n_443), .Y(n_530) );
AND2x2_ASAP7_75t_L g948 ( .A(n_443), .B(n_946), .Y(n_948) );
BUFx2_ASAP7_75t_L g1088 ( .A(n_443), .Y(n_1088) );
BUFx2_ASAP7_75t_L g1153 ( .A(n_443), .Y(n_1153) );
BUFx2_ASAP7_75t_L g1189 ( .A(n_443), .Y(n_1189) );
INVx1_ASAP7_75t_L g454 ( .A(n_444), .Y(n_454) );
INVx2_ASAP7_75t_L g444 ( .A(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g500 ( .A(n_445), .Y(n_500) );
BUFx6f_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g456 ( .A(n_448), .Y(n_456) );
INVx2_ASAP7_75t_L g717 ( .A(n_448), .Y(n_717) );
INVx2_ASAP7_75t_L g1085 ( .A(n_448), .Y(n_1085) );
INVx2_ASAP7_75t_L g1156 ( .A(n_448), .Y(n_1156) );
BUFx6f_ASAP7_75t_L g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_L g484 ( .A(n_449), .Y(n_484) );
BUFx8_ASAP7_75t_L g534 ( .A(n_449), .Y(n_534) );
BUFx6f_ASAP7_75t_L g643 ( .A(n_449), .Y(n_643) );
BUFx2_ASAP7_75t_L g1184 ( .A(n_451), .Y(n_1184) );
BUFx12f_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
BUFx3_ASAP7_75t_L g535 ( .A(n_452), .Y(n_535) );
INVx5_ASAP7_75t_L g806 ( .A(n_452), .Y(n_806) );
BUFx2_ASAP7_75t_L g934 ( .A(n_452), .Y(n_934) );
AND2x4_ASAP7_75t_L g966 ( .A(n_452), .B(n_964), .Y(n_966) );
AND2x4_ASAP7_75t_L g452 ( .A(n_453), .B(n_454), .Y(n_452) );
INVx2_ASAP7_75t_L g471 ( .A(n_453), .Y(n_471) );
NAND2x1p5_ASAP7_75t_L g499 ( .A(n_453), .B(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g475 ( .A(n_454), .Y(n_475) );
AOI22xp5_ASAP7_75t_L g1660 ( .A1(n_458), .A2(n_502), .B1(n_1639), .B2(n_1661), .Y(n_1660) );
INVx2_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g644 ( .A(n_459), .Y(n_644) );
INVx2_ASAP7_75t_L g783 ( .A(n_459), .Y(n_783) );
INVx1_ASAP7_75t_L g802 ( .A(n_459), .Y(n_802) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx1_ASAP7_75t_L g810 ( .A(n_461), .Y(n_810) );
INVx1_ASAP7_75t_SL g880 ( .A(n_461), .Y(n_880) );
OR2x6_ASAP7_75t_L g461 ( .A(n_462), .B(n_463), .Y(n_461) );
INVx1_ASAP7_75t_L g745 ( .A(n_462), .Y(n_745) );
AND2x4_ASAP7_75t_L g911 ( .A(n_462), .B(n_912), .Y(n_911) );
OR2x2_ASAP7_75t_L g1322 ( .A(n_462), .B(n_463), .Y(n_1322) );
INVx3_ASAP7_75t_L g992 ( .A(n_463), .Y(n_992) );
AOI22xp5_ASAP7_75t_L g795 ( .A1(n_466), .A2(n_472), .B1(n_796), .B2(n_797), .Y(n_795) );
AOI22xp33_ASAP7_75t_L g874 ( .A1(n_466), .A2(n_472), .B1(n_854), .B2(n_856), .Y(n_874) );
AOI22xp5_ASAP7_75t_L g1317 ( .A1(n_466), .A2(n_472), .B1(n_1318), .B2(n_1319), .Y(n_1317) );
AOI221xp5_ASAP7_75t_L g1714 ( .A1(n_466), .A2(n_472), .B1(n_477), .B2(n_1715), .C(n_1716), .Y(n_1714) );
AND2x4_ASAP7_75t_SL g466 ( .A(n_467), .B(n_470), .Y(n_466) );
AND2x4_ASAP7_75t_SL g472 ( .A(n_467), .B(n_473), .Y(n_472) );
AND2x4_ASAP7_75t_L g477 ( .A(n_467), .B(n_478), .Y(n_477) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_467), .B(n_470), .Y(n_525) );
AND2x4_ASAP7_75t_L g527 ( .A(n_467), .B(n_473), .Y(n_527) );
AND2x2_ASAP7_75t_L g1162 ( .A(n_467), .B(n_470), .Y(n_1162) );
AND2x2_ASAP7_75t_L g1173 ( .A(n_467), .B(n_470), .Y(n_1173) );
OR2x2_ASAP7_75t_L g558 ( .A(n_468), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g915 ( .A(n_468), .Y(n_915) );
INVx1_ASAP7_75t_L g468 ( .A(n_469), .Y(n_468) );
INVx1_ASAP7_75t_L g540 ( .A(n_469), .Y(n_540) );
INVx3_ASAP7_75t_L g470 ( .A(n_471), .Y(n_470) );
INVx1_ASAP7_75t_L g724 ( .A(n_472), .Y(n_724) );
INVx2_ASAP7_75t_L g473 ( .A(n_474), .Y(n_473) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx3_ASAP7_75t_L g554 ( .A(n_477), .Y(n_554) );
HB1xp67_ASAP7_75t_L g701 ( .A(n_477), .Y(n_701) );
NOR3xp33_ASAP7_75t_L g771 ( .A(n_477), .B(n_772), .C(n_784), .Y(n_771) );
INVx3_ASAP7_75t_L g811 ( .A(n_477), .Y(n_811) );
AOI211xp5_ASAP7_75t_L g871 ( .A1(n_477), .A2(n_863), .B(n_872), .C(n_873), .Y(n_871) );
NOR3xp33_ASAP7_75t_SL g1274 ( .A(n_477), .B(n_1275), .C(n_1286), .Y(n_1274) );
INVx1_ASAP7_75t_L g517 ( .A(n_479), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_494), .Y(n_479) );
NAND2x1_ASAP7_75t_L g480 ( .A(n_481), .B(n_489), .Y(n_480) );
INVx2_ASAP7_75t_SL g481 ( .A(n_482), .Y(n_481) );
AOI22xp33_ASAP7_75t_L g840 ( .A1(n_482), .A2(n_501), .B1(n_822), .B2(n_823), .Y(n_840) );
AOI22xp33_ASAP7_75t_L g870 ( .A1(n_482), .A2(n_686), .B1(n_867), .B2(n_868), .Y(n_870) );
AOI22xp33_ASAP7_75t_L g1339 ( .A1(n_482), .A2(n_501), .B1(n_1330), .B2(n_1331), .Y(n_1339) );
AND2x2_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx2_ASAP7_75t_L g1282 ( .A(n_483), .Y(n_1282) );
INVx3_ASAP7_75t_L g483 ( .A(n_484), .Y(n_483) );
OAI221xp5_ASAP7_75t_L g706 ( .A1(n_484), .A2(n_707), .B1(n_708), .B2(n_712), .C(n_713), .Y(n_706) );
INVx1_ASAP7_75t_L g933 ( .A(n_484), .Y(n_933) );
OR2x6_ASAP7_75t_SL g962 ( .A(n_484), .B(n_963), .Y(n_962) );
INVxp67_ASAP7_75t_L g550 ( .A(n_485), .Y(n_550) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
OR2x2_ASAP7_75t_L g497 ( .A(n_486), .B(n_498), .Y(n_497) );
INVx1_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
OR2x2_ASAP7_75t_L g506 ( .A(n_486), .B(n_507), .Y(n_506) );
OR2x2_ASAP7_75t_L g486 ( .A(n_487), .B(n_488), .Y(n_486) );
OR2x2_ASAP7_75t_L g704 ( .A(n_487), .B(n_705), .Y(n_704) );
INVx1_ASAP7_75t_L g1013 ( .A(n_487), .Y(n_1013) );
INVx1_ASAP7_75t_L g946 ( .A(n_488), .Y(n_946) );
INVx1_ASAP7_75t_L g964 ( .A(n_488), .Y(n_964) );
INVx2_ASAP7_75t_L g489 ( .A(n_490), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g968 ( .A(n_490), .B(n_969), .Y(n_968) );
NAND2xp5_ASAP7_75t_L g976 ( .A(n_490), .B(n_977), .Y(n_976) );
AOI22xp33_ASAP7_75t_L g1638 ( .A1(n_490), .A2(n_929), .B1(n_1639), .B2(n_1640), .Y(n_1638) );
AND2x4_ASAP7_75t_L g490 ( .A(n_491), .B(n_492), .Y(n_490) );
AND2x4_ASAP7_75t_L g929 ( .A(n_491), .B(n_591), .Y(n_929) );
INVx2_ASAP7_75t_L g579 ( .A(n_493), .Y(n_579) );
INVx1_ASAP7_75t_L g756 ( .A(n_493), .Y(n_756) );
BUFx6f_ASAP7_75t_L g818 ( .A(n_493), .Y(n_818) );
INVx1_ASAP7_75t_L g516 ( .A(n_495), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g1052 ( .A1(n_496), .A2(n_505), .B1(n_1037), .B2(n_1053), .Y(n_1052) );
AOI222xp33_ASAP7_75t_L g1705 ( .A1(n_496), .A2(n_501), .B1(n_505), .B2(n_1706), .C1(n_1707), .C2(n_1708), .Y(n_1705) );
INVx2_ASAP7_75t_L g496 ( .A(n_497), .Y(n_496) );
AND2x4_ASAP7_75t_L g562 ( .A(n_497), .B(n_563), .Y(n_562) );
AND2x4_ASAP7_75t_L g699 ( .A(n_497), .B(n_563), .Y(n_699) );
INVx3_ASAP7_75t_L g998 ( .A(n_498), .Y(n_998) );
BUFx6f_ASAP7_75t_L g498 ( .A(n_499), .Y(n_498) );
BUFx2_ASAP7_75t_L g959 ( .A(n_499), .Y(n_959) );
AND2x4_ASAP7_75t_L g501 ( .A(n_502), .B(n_503), .Y(n_501) );
AND2x4_ASAP7_75t_L g686 ( .A(n_502), .B(n_503), .Y(n_686) );
AND2x4_ASAP7_75t_L g552 ( .A(n_503), .B(n_534), .Y(n_552) );
INVx1_ASAP7_75t_L g505 ( .A(n_506), .Y(n_505) );
AND2x4_ASAP7_75t_L g557 ( .A(n_506), .B(n_558), .Y(n_557) );
BUFx3_ASAP7_75t_L g987 ( .A(n_507), .Y(n_987) );
INVx1_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
BUFx6f_ASAP7_75t_L g720 ( .A(n_508), .Y(n_720) );
INVx1_ASAP7_75t_L g508 ( .A(n_509), .Y(n_508) );
BUFx2_ASAP7_75t_L g711 ( .A(n_509), .Y(n_711) );
OAI21xp5_ASAP7_75t_L g511 ( .A1(n_512), .A2(n_513), .B(n_514), .Y(n_511) );
OAI21xp33_ASAP7_75t_L g515 ( .A1(n_514), .A2(n_516), .B(n_517), .Y(n_515) );
NAND3xp33_ASAP7_75t_L g519 ( .A(n_520), .B(n_555), .C(n_568), .Y(n_519) );
NOR3xp33_ASAP7_75t_L g520 ( .A(n_521), .B(n_545), .C(n_553), .Y(n_520) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_528), .Y(n_521) );
AOI22xp33_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B1(n_526), .B2(n_527), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g628 ( .A1(n_524), .A2(n_629), .B1(n_630), .B2(n_631), .Y(n_628) );
AOI221x1_ASAP7_75t_L g1054 ( .A1(n_524), .A2(n_527), .B1(n_1031), .B2(n_1036), .C(n_1055), .Y(n_1054) );
AOI22xp33_ASAP7_75t_L g1078 ( .A1(n_524), .A2(n_527), .B1(n_1079), .B2(n_1080), .Y(n_1078) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
HB1xp67_ASAP7_75t_L g631 ( .A(n_527), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g1160 ( .A1(n_527), .A2(n_1161), .B1(n_1162), .B2(n_1163), .Y(n_1160) );
AO22x1_ASAP7_75t_L g1171 ( .A1(n_527), .A2(n_1172), .B1(n_1173), .B2(n_1174), .Y(n_1171) );
AOI22xp33_ASAP7_75t_L g1223 ( .A1(n_527), .A2(n_1173), .B1(n_1224), .B2(n_1225), .Y(n_1223) );
AOI22xp33_ASAP7_75t_L g1370 ( .A1(n_527), .A2(n_1162), .B1(n_1371), .B2(n_1372), .Y(n_1370) );
INVx1_ASAP7_75t_L g532 ( .A(n_533), .Y(n_532) );
INVx3_ASAP7_75t_L g533 ( .A(n_534), .Y(n_533) );
INVx2_ASAP7_75t_SL g775 ( .A(n_534), .Y(n_775) );
BUFx2_ASAP7_75t_L g537 ( .A(n_538), .Y(n_537) );
BUFx2_ASAP7_75t_L g648 ( .A(n_538), .Y(n_648) );
BUFx2_ASAP7_75t_L g1158 ( .A(n_538), .Y(n_1158) );
BUFx2_ASAP7_75t_L g1185 ( .A(n_538), .Y(n_1185) );
INVx3_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
INVx3_ASAP7_75t_L g715 ( .A(n_539), .Y(n_715) );
INVx1_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
INVx2_ASAP7_75t_SL g1181 ( .A(n_544), .Y(n_1181) );
NAND2xp5_ASAP7_75t_L g1070 ( .A(n_546), .B(n_928), .Y(n_1070) );
OR2x6_ASAP7_75t_L g546 ( .A(n_547), .B(n_550), .Y(n_546) );
OR2x2_ASAP7_75t_L g1090 ( .A(n_547), .B(n_550), .Y(n_1090) );
INVx2_ASAP7_75t_SL g547 ( .A(n_548), .Y(n_547) );
INVx2_ASAP7_75t_L g548 ( .A(n_549), .Y(n_548) );
BUFx4f_ASAP7_75t_L g1256 ( .A(n_549), .Y(n_1256) );
INVxp67_ASAP7_75t_L g1310 ( .A(n_551), .Y(n_1310) );
INVx2_ASAP7_75t_L g551 ( .A(n_552), .Y(n_551) );
AOI22xp33_ASAP7_75t_L g685 ( .A1(n_552), .A2(n_660), .B1(n_662), .B2(n_686), .Y(n_685) );
AOI22xp33_ASAP7_75t_L g746 ( .A1(n_552), .A2(n_686), .B1(n_734), .B2(n_736), .Y(n_746) );
AOI22xp33_ASAP7_75t_L g788 ( .A1(n_552), .A2(n_686), .B1(n_760), .B2(n_761), .Y(n_788) );
INVx2_ASAP7_75t_L g1150 ( .A(n_552), .Y(n_1150) );
AOI22xp33_ASAP7_75t_L g1191 ( .A1(n_552), .A2(n_686), .B1(n_1192), .B2(n_1193), .Y(n_1191) );
NAND2xp5_ASAP7_75t_L g1703 ( .A(n_552), .B(n_1704), .Y(n_1703) );
INVx2_ASAP7_75t_SL g553 ( .A(n_554), .Y(n_553) );
AND4x1_ASAP7_75t_L g627 ( .A(n_554), .B(n_628), .C(n_632), .D(n_635), .Y(n_627) );
AND5x1_ASAP7_75t_L g1027 ( .A(n_554), .B(n_1028), .C(n_1054), .D(n_1068), .E(n_1071), .Y(n_1027) );
AND4x1_ASAP7_75t_L g1147 ( .A(n_554), .B(n_1148), .C(n_1151), .D(n_1160), .Y(n_1147) );
NAND5xp2_ASAP7_75t_L g1222 ( .A(n_554), .B(n_1223), .C(n_1226), .D(n_1228), .E(n_1229), .Y(n_1222) );
NAND3xp33_ASAP7_75t_SL g1316 ( .A(n_554), .B(n_1317), .C(n_1320), .Y(n_1316) );
AOI21xp33_ASAP7_75t_SL g555 ( .A1(n_556), .A2(n_560), .B(n_561), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_556), .B(n_688), .Y(n_687) );
AOI21xp5_ASAP7_75t_L g696 ( .A1(n_556), .A2(n_697), .B(n_698), .Y(n_696) );
AOI21xp5_ASAP7_75t_L g785 ( .A1(n_556), .A2(n_786), .B(n_787), .Y(n_785) );
NAND2xp5_ASAP7_75t_L g841 ( .A(n_556), .B(n_842), .Y(n_841) );
NAND2xp5_ASAP7_75t_L g847 ( .A(n_556), .B(n_848), .Y(n_847) );
AOI21xp33_ASAP7_75t_SL g1092 ( .A1(n_556), .A2(n_1093), .B(n_1094), .Y(n_1092) );
AOI21xp33_ASAP7_75t_L g1125 ( .A1(n_556), .A2(n_1126), .B(n_1127), .Y(n_1125) );
AOI211x1_ASAP7_75t_L g1167 ( .A1(n_556), .A2(n_1168), .B(n_1169), .C(n_1190), .Y(n_1167) );
AOI221xp5_ASAP7_75t_L g1313 ( .A1(n_556), .A2(n_872), .B1(n_1314), .B2(n_1315), .C(n_1316), .Y(n_1313) );
AOI21xp33_ASAP7_75t_SL g1365 ( .A1(n_556), .A2(n_1366), .B(n_1367), .Y(n_1365) );
INVx8_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g1688 ( .A(n_558), .B(n_1689), .Y(n_1688) );
INVx1_ASAP7_75t_L g916 ( .A(n_559), .Y(n_916) );
HB1xp67_ASAP7_75t_L g684 ( .A(n_562), .Y(n_684) );
INVx2_ASAP7_75t_L g1248 ( .A(n_562), .Y(n_1248) );
INVx2_ASAP7_75t_SL g1017 ( .A(n_563), .Y(n_1017) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g1684 ( .A(n_567), .B(n_1685), .Y(n_1684) );
OAI21xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_595), .B(n_618), .Y(n_568) );
INVx2_ASAP7_75t_SL g570 ( .A(n_571), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g824 ( .A(n_571), .B(n_799), .Y(n_824) );
INVx3_ASAP7_75t_L g1097 ( .A(n_571), .Y(n_1097) );
NAND2xp5_ASAP7_75t_R g1204 ( .A(n_571), .B(n_1177), .Y(n_1204) );
AOI22xp33_ASAP7_75t_L g1348 ( .A1(n_571), .A2(n_735), .B1(n_1349), .B2(n_1350), .Y(n_1348) );
INVx1_ASAP7_75t_L g658 ( .A(n_572), .Y(n_658) );
BUFx2_ASAP7_75t_L g1101 ( .A(n_572), .Y(n_1101) );
AOI21xp5_ASAP7_75t_SL g573 ( .A1(n_574), .A2(n_582), .B(n_586), .Y(n_573) );
BUFx2_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AOI221xp5_ASAP7_75t_L g1728 ( .A1(n_576), .A2(n_1104), .B1(n_1704), .B2(n_1716), .C(n_1729), .Y(n_1728) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
INVx2_ASAP7_75t_L g578 ( .A(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g1104 ( .A(n_579), .Y(n_1104) );
HB1xp67_ASAP7_75t_SL g580 ( .A(n_581), .Y(n_580) );
BUFx3_ASAP7_75t_L g584 ( .A(n_585), .Y(n_584) );
INVx1_ASAP7_75t_SL g1203 ( .A(n_585), .Y(n_1203) );
AOI21xp5_ASAP7_75t_L g651 ( .A1(n_586), .A2(n_652), .B(n_654), .Y(n_651) );
AOI21xp5_ASAP7_75t_L g727 ( .A1(n_586), .A2(n_728), .B(n_730), .Y(n_727) );
AOI21xp5_ASAP7_75t_L g752 ( .A1(n_586), .A2(n_753), .B(n_757), .Y(n_752) );
INVx1_ASAP7_75t_L g825 ( .A(n_586), .Y(n_825) );
AOI21xp5_ASAP7_75t_L g1098 ( .A1(n_586), .A2(n_1099), .B(n_1102), .Y(n_1098) );
AOI21xp5_ASAP7_75t_L g1133 ( .A1(n_586), .A2(n_1134), .B(n_1137), .Y(n_1133) );
AOI21xp5_ASAP7_75t_L g1197 ( .A1(n_586), .A2(n_1198), .B(n_1201), .Y(n_1197) );
AOI21xp5_ASAP7_75t_L g1346 ( .A1(n_586), .A2(n_593), .B(n_1347), .Y(n_1346) );
AOI22xp33_ASAP7_75t_L g587 ( .A1(n_588), .A2(n_589), .B1(n_592), .B2(n_593), .Y(n_587) );
AOI22xp33_ASAP7_75t_L g659 ( .A1(n_589), .A2(n_660), .B1(n_661), .B2(n_662), .Y(n_659) );
AOI22xp5_ASAP7_75t_L g1105 ( .A1(n_589), .A2(n_593), .B1(n_1106), .B2(n_1107), .Y(n_1105) );
AOI22xp33_ASAP7_75t_L g1196 ( .A1(n_589), .A2(n_594), .B1(n_1192), .B2(n_1193), .Y(n_1196) );
INVx2_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g590 ( .A(n_591), .Y(n_590) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_591), .Y(n_735) );
AOI22xp33_ASAP7_75t_L g759 ( .A1(n_591), .A2(n_594), .B1(n_760), .B2(n_761), .Y(n_759) );
AOI22xp33_ASAP7_75t_L g1130 ( .A1(n_593), .A2(n_735), .B1(n_1131), .B2(n_1132), .Y(n_1130) );
INVxp67_ASAP7_75t_SL g1240 ( .A(n_593), .Y(n_1240) );
BUFx6f_ASAP7_75t_L g593 ( .A(n_594), .Y(n_593) );
HB1xp67_ASAP7_75t_L g661 ( .A(n_594), .Y(n_661) );
AOI22xp33_ASAP7_75t_L g733 ( .A1(n_594), .A2(n_734), .B1(n_735), .B2(n_736), .Y(n_733) );
AOI22xp5_ASAP7_75t_L g821 ( .A1(n_594), .A2(n_735), .B1(n_822), .B2(n_823), .Y(n_821) );
AOI22xp33_ASAP7_75t_L g866 ( .A1(n_594), .A2(n_735), .B1(n_867), .B2(n_868), .Y(n_866) );
AOI22xp5_ASAP7_75t_L g1294 ( .A1(n_594), .A2(n_735), .B1(n_1295), .B2(n_1296), .Y(n_1294) );
AOI22xp5_ASAP7_75t_L g1329 ( .A1(n_594), .A2(n_735), .B1(n_1330), .B2(n_1331), .Y(n_1329) );
INVx2_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
INVx2_ASAP7_75t_L g664 ( .A(n_597), .Y(n_664) );
INVx1_ASAP7_75t_L g1206 ( .A(n_597), .Y(n_1206) );
INVx4_ASAP7_75t_L g597 ( .A(n_598), .Y(n_597) );
INVx2_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
BUFx3_ASAP7_75t_L g855 ( .A(n_599), .Y(n_855) );
INVx2_ASAP7_75t_L g600 ( .A(n_601), .Y(n_600) );
INVx2_ASAP7_75t_L g682 ( .A(n_601), .Y(n_682) );
OAI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_606), .B1(n_607), .B2(n_612), .C(n_613), .Y(n_603) );
OAI22xp5_ASAP7_75t_L g1210 ( .A1(n_604), .A2(n_1211), .B1(n_1212), .B2(n_1213), .Y(n_1210) );
INVx2_ASAP7_75t_L g604 ( .A(n_605), .Y(n_604) );
BUFx2_ASAP7_75t_L g679 ( .A(n_607), .Y(n_679) );
INVx1_ASAP7_75t_L g888 ( .A(n_607), .Y(n_888) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_608), .Y(n_607) );
INVx2_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
INVx2_ASAP7_75t_L g838 ( .A(n_609), .Y(n_838) );
INVx4_ASAP7_75t_L g1040 ( .A(n_609), .Y(n_1040) );
INVx2_ASAP7_75t_SL g1112 ( .A(n_609), .Y(n_1112) );
BUFx6f_ASAP7_75t_L g1214 ( .A(n_609), .Y(n_1214) );
INVx1_ASAP7_75t_L g1302 ( .A(n_609), .Y(n_1302) );
INVx2_ASAP7_75t_L g1730 ( .A(n_609), .Y(n_1730) );
INVx8_ASAP7_75t_L g609 ( .A(n_610), .Y(n_609) );
BUFx2_ASAP7_75t_L g907 ( .A(n_610), .Y(n_907) );
BUFx6f_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx2_ASAP7_75t_L g615 ( .A(n_616), .Y(n_615) );
INVx2_ASAP7_75t_L g1357 ( .A(n_616), .Y(n_1357) );
INVx1_ASAP7_75t_L g674 ( .A(n_617), .Y(n_674) );
O2A1O1Ixp5_ASAP7_75t_L g649 ( .A1(n_618), .A2(n_650), .B(n_663), .C(n_683), .Y(n_649) );
OAI21xp5_ASAP7_75t_L g1095 ( .A1(n_618), .A2(n_1096), .B(n_1108), .Y(n_1095) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_620), .B(n_1382), .C(n_1383), .Y(n_619) );
NAND3xp33_ASAP7_75t_L g620 ( .A(n_621), .B(n_1021), .C(n_1341), .Y(n_620) );
INVx1_ASAP7_75t_L g621 ( .A(n_622), .Y(n_621) );
NAND3xp33_ASAP7_75t_L g1382 ( .A(n_622), .B(n_1021), .C(n_1342), .Y(n_1382) );
AOI33xp33_ASAP7_75t_L g1383 ( .A1(n_622), .A2(n_623), .A3(n_1022), .B1(n_1341), .B2(n_1342), .B3(n_1748), .Y(n_1383) );
INVx2_ASAP7_75t_L g622 ( .A(n_623), .Y(n_622) );
OA22x2_ASAP7_75t_L g623 ( .A1(n_624), .A2(n_625), .B1(n_690), .B2(n_691), .Y(n_623) );
INVx1_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
XOR2x2_ASAP7_75t_L g625 ( .A(n_626), .B(n_689), .Y(n_625) );
NAND3x1_ASAP7_75t_SL g626 ( .A(n_627), .B(n_649), .C(n_687), .Y(n_626) );
NAND2xp5_ASAP7_75t_L g632 ( .A(n_633), .B(n_634), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g798 ( .A(n_634), .B(n_799), .Y(n_798) );
NAND2xp5_ASAP7_75t_L g1071 ( .A(n_634), .B(n_1072), .Y(n_1071) );
NAND2xp5_ASAP7_75t_L g1176 ( .A(n_634), .B(n_1177), .Y(n_1176) );
NAND2xp5_ASAP7_75t_L g1717 ( .A(n_634), .B(n_1718), .Y(n_1717) );
AOI33xp33_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_637), .A3(n_639), .B1(n_645), .B2(n_646), .B3(n_648), .Y(n_635) );
AOI33xp33_ASAP7_75t_L g1178 ( .A1(n_636), .A2(n_1179), .A3(n_1182), .B1(n_1183), .B2(n_1185), .B3(n_1186), .Y(n_1178) );
INVx1_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
OAI221xp5_ASAP7_75t_L g1260 ( .A1(n_641), .A2(n_1237), .B1(n_1261), .B2(n_1262), .C(n_1263), .Y(n_1260) );
BUFx3_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
OAI221xp5_ASAP7_75t_L g1064 ( .A1(n_642), .A2(n_987), .B1(n_1047), .B2(n_1065), .C(n_1066), .Y(n_1064) );
INVx8_ASAP7_75t_L g1701 ( .A(n_642), .Y(n_1701) );
INVx5_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx3_ASAP7_75t_L g938 ( .A(n_643), .Y(n_938) );
INVx2_ASAP7_75t_SL g1058 ( .A(n_643), .Y(n_1058) );
HB1xp67_ASAP7_75t_L g1376 ( .A(n_643), .Y(n_1376) );
INVx2_ASAP7_75t_SL g1379 ( .A(n_643), .Y(n_1379) );
HB1xp67_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx1_ASAP7_75t_L g657 ( .A(n_658), .Y(n_657) );
OAI221xp5_ASAP7_75t_L g665 ( .A1(n_666), .A2(n_668), .B1(n_669), .B2(n_673), .C(n_674), .Y(n_665) );
BUFx2_ASAP7_75t_SL g666 ( .A(n_667), .Y(n_666) );
INVx2_ASAP7_75t_SL g766 ( .A(n_667), .Y(n_766) );
OR2x2_ASAP7_75t_L g923 ( .A(n_667), .B(n_920), .Y(n_923) );
OR2x2_ASAP7_75t_L g1675 ( .A(n_667), .B(n_920), .Y(n_1675) );
NAND2xp5_ASAP7_75t_L g1732 ( .A(n_667), .B(n_1733), .Y(n_1732) );
INVx2_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx4_ASAP7_75t_L g670 ( .A(n_671), .Y(n_670) );
BUFx2_ASAP7_75t_L g671 ( .A(n_672), .Y(n_671) );
BUFx3_ASAP7_75t_L g830 ( .A(n_672), .Y(n_830) );
BUFx2_ASAP7_75t_L g1039 ( .A(n_672), .Y(n_1039) );
INVx1_ASAP7_75t_L g1679 ( .A(n_672), .Y(n_1679) );
INVx2_ASAP7_75t_L g1725 ( .A(n_672), .Y(n_1725) );
OAI221xp5_ASAP7_75t_L g827 ( .A1(n_674), .A2(n_828), .B1(n_829), .B2(n_830), .C(n_831), .Y(n_827) );
OAI22xp5_ASAP7_75t_L g675 ( .A1(n_676), .A2(n_677), .B1(n_679), .B2(n_680), .Y(n_675) );
INVx1_ASAP7_75t_L g889 ( .A(n_677), .Y(n_889) );
OAI221xp5_ASAP7_75t_L g1109 ( .A1(n_677), .A2(n_1110), .B1(n_1111), .B2(n_1113), .C(n_1114), .Y(n_1109) );
OAI221xp5_ASAP7_75t_L g1234 ( .A1(n_677), .A2(n_1235), .B1(n_1236), .B2(n_1237), .C(n_1238), .Y(n_1234) );
OAI221xp5_ASAP7_75t_L g1241 ( .A1(n_677), .A2(n_907), .B1(n_1242), .B2(n_1243), .C(n_1244), .Y(n_1241) );
OAI221xp5_ASAP7_75t_L g1358 ( .A1(n_677), .A2(n_1111), .B1(n_1359), .B2(n_1360), .C(n_1361), .Y(n_1358) );
BUFx6f_ASAP7_75t_L g677 ( .A(n_678), .Y(n_677) );
OAI22xp5_ASAP7_75t_L g1004 ( .A1(n_678), .A2(n_838), .B1(n_1005), .B2(n_1006), .Y(n_1004) );
OAI22x1_ASAP7_75t_SL g1009 ( .A1(n_678), .A2(n_838), .B1(n_988), .B2(n_1010), .Y(n_1009) );
INVx2_ASAP7_75t_SL g1141 ( .A(n_678), .Y(n_1141) );
BUFx3_ASAP7_75t_L g1299 ( .A(n_678), .Y(n_1299) );
OAI221xp5_ASAP7_75t_L g1139 ( .A1(n_679), .A2(n_1140), .B1(n_1142), .B2(n_1143), .C(n_1144), .Y(n_1139) );
BUFx2_ASAP7_75t_L g681 ( .A(n_682), .Y(n_681) );
NAND2xp5_ASAP7_75t_L g1229 ( .A(n_686), .B(n_1230), .Y(n_1229) );
AOI22xp5_ASAP7_75t_L g1309 ( .A1(n_686), .A2(n_1295), .B1(n_1296), .B2(n_1310), .Y(n_1309) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
XNOR2x1_ASAP7_75t_L g691 ( .A(n_692), .B(n_790), .Y(n_691) );
INVx1_ASAP7_75t_L g692 ( .A(n_693), .Y(n_692) );
AO22x2_ASAP7_75t_L g693 ( .A1(n_694), .A2(n_747), .B1(n_748), .B2(n_789), .Y(n_693) );
INVx1_ASAP7_75t_L g789 ( .A(n_694), .Y(n_789) );
AND4x1_ASAP7_75t_L g695 ( .A(n_696), .B(n_700), .C(n_725), .D(n_746), .Y(n_695) );
INVx1_ASAP7_75t_SL g1272 ( .A(n_699), .Y(n_1272) );
NOR3xp33_ASAP7_75t_L g700 ( .A(n_701), .B(n_702), .C(n_723), .Y(n_700) );
OAI22xp5_ASAP7_75t_SL g702 ( .A1(n_703), .A2(n_706), .B1(n_714), .B2(n_716), .Y(n_702) );
BUFx4f_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
BUFx8_ASAP7_75t_L g773 ( .A(n_704), .Y(n_773) );
BUFx2_ASAP7_75t_L g1056 ( .A(n_704), .Y(n_1056) );
BUFx4f_ASAP7_75t_L g1276 ( .A(n_704), .Y(n_1276) );
BUFx2_ASAP7_75t_L g939 ( .A(n_705), .Y(n_939) );
OAI221xp5_ASAP7_75t_L g774 ( .A1(n_708), .A2(n_775), .B1(n_776), .B2(n_777), .C(n_778), .Y(n_774) );
INVx3_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
BUFx2_ASAP7_75t_L g709 ( .A(n_710), .Y(n_709) );
INVx1_ASAP7_75t_L g710 ( .A(n_711), .Y(n_710) );
BUFx3_ASAP7_75t_L g1262 ( .A(n_711), .Y(n_1262) );
INVx2_ASAP7_75t_L g714 ( .A(n_715), .Y(n_714) );
CKINVDCx5p33_ASAP7_75t_R g779 ( .A(n_715), .Y(n_779) );
INVx2_ASAP7_75t_L g1063 ( .A(n_715), .Y(n_1063) );
OAI221xp5_ASAP7_75t_L g716 ( .A1(n_717), .A2(n_718), .B1(n_719), .B2(n_721), .C(n_722), .Y(n_716) );
INVx1_ASAP7_75t_L g804 ( .A(n_717), .Y(n_804) );
OAI211xp5_ASAP7_75t_L g738 ( .A1(n_718), .A2(n_739), .B(n_740), .C(n_741), .Y(n_738) );
OAI221xp5_ASAP7_75t_L g780 ( .A1(n_719), .A2(n_764), .B1(n_775), .B2(n_781), .C(n_782), .Y(n_780) );
CKINVDCx8_ASAP7_75t_R g719 ( .A(n_720), .Y(n_719) );
INVx3_ASAP7_75t_L g1060 ( .A(n_720), .Y(n_1060) );
INVx3_ASAP7_75t_L g1646 ( .A(n_720), .Y(n_1646) );
INVx3_ASAP7_75t_L g1654 ( .A(n_720), .Y(n_1654) );
OAI21xp5_ASAP7_75t_L g725 ( .A1(n_726), .A2(n_737), .B(n_743), .Y(n_725) );
INVx2_ASAP7_75t_SL g731 ( .A(n_732), .Y(n_731) );
INVx1_ASAP7_75t_L g1293 ( .A(n_732), .Y(n_1293) );
INVx1_ASAP7_75t_L g1246 ( .A(n_735), .Y(n_1246) );
OAI21xp5_ASAP7_75t_L g1194 ( .A1(n_743), .A2(n_1195), .B(n_1205), .Y(n_1194) );
AOI21xp5_ASAP7_75t_L g1327 ( .A1(n_743), .A2(n_1328), .B(n_1338), .Y(n_1327) );
INVx2_ASAP7_75t_L g743 ( .A(n_744), .Y(n_743) );
INVx1_ASAP7_75t_L g850 ( .A(n_744), .Y(n_850) );
BUFx2_ASAP7_75t_L g744 ( .A(n_745), .Y(n_744) );
INVx1_ASAP7_75t_L g1146 ( .A(n_745), .Y(n_1146) );
NAND2xp5_ASAP7_75t_L g1689 ( .A(n_745), .B(n_966), .Y(n_1689) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
AND4x1_ASAP7_75t_L g749 ( .A(n_750), .B(n_771), .C(n_785), .D(n_788), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g750 ( .A1(n_751), .A2(n_762), .B(n_770), .Y(n_750) );
INVx2_ASAP7_75t_SL g755 ( .A(n_756), .Y(n_755) );
OAI211xp5_ASAP7_75t_L g763 ( .A1(n_764), .A2(n_765), .B(n_767), .C(n_769), .Y(n_763) );
OAI211xp5_ASAP7_75t_L g1046 ( .A1(n_765), .A2(n_1047), .B(n_1048), .C(n_1049), .Y(n_1046) );
INVx5_ASAP7_75t_L g765 ( .A(n_766), .Y(n_765) );
O2A1O1Ixp5_ASAP7_75t_SL g812 ( .A1(n_770), .A2(n_813), .B(n_826), .C(n_839), .Y(n_812) );
OAI22xp5_ASAP7_75t_SL g772 ( .A1(n_773), .A2(n_774), .B1(n_779), .B2(n_780), .Y(n_772) );
XOR2xp5_ASAP7_75t_L g790 ( .A(n_791), .B(n_882), .Y(n_790) );
XNOR2xp5_ASAP7_75t_L g791 ( .A(n_792), .B(n_844), .Y(n_791) );
XOR2xp5_ASAP7_75t_L g792 ( .A(n_793), .B(n_843), .Y(n_792) );
NAND3xp33_ASAP7_75t_L g793 ( .A(n_794), .B(n_812), .C(n_841), .Y(n_793) );
AND4x1_ASAP7_75t_L g794 ( .A(n_795), .B(n_798), .C(n_800), .D(n_811), .Y(n_794) );
INVx2_ASAP7_75t_R g805 ( .A(n_806), .Y(n_805) );
INVx2_ASAP7_75t_L g808 ( .A(n_806), .Y(n_808) );
NAND3xp33_ASAP7_75t_L g1709 ( .A(n_810), .B(n_1710), .C(n_1712), .Y(n_1709) );
INVx1_ASAP7_75t_L g1091 ( .A(n_811), .Y(n_1091) );
NAND2xp5_ASAP7_75t_SL g1175 ( .A(n_811), .B(n_1176), .Y(n_1175) );
NAND4xp25_ASAP7_75t_L g813 ( .A(n_814), .B(n_821), .C(n_824), .D(n_825), .Y(n_813) );
OAI211xp5_ASAP7_75t_L g814 ( .A1(n_815), .A2(n_816), .B(n_817), .C(n_819), .Y(n_814) );
BUFx3_ASAP7_75t_L g1200 ( .A(n_818), .Y(n_1200) );
INVx2_ASAP7_75t_L g891 ( .A(n_830), .Y(n_891) );
OAI221xp5_ASAP7_75t_L g908 ( .A1(n_830), .A2(n_893), .B1(n_909), .B2(n_910), .C(n_911), .Y(n_908) );
OAI22xp5_ASAP7_75t_L g832 ( .A1(n_833), .A2(n_834), .B1(n_837), .B2(n_838), .Y(n_832) );
INVx1_ASAP7_75t_L g834 ( .A(n_835), .Y(n_834) );
INVxp67_ASAP7_75t_L g835 ( .A(n_836), .Y(n_835) );
OR2x6_ASAP7_75t_L g1397 ( .A(n_836), .B(n_1398), .Y(n_1397) );
INVx1_ASAP7_75t_L g845 ( .A(n_846), .Y(n_845) );
NAND3xp33_ASAP7_75t_L g846 ( .A(n_847), .B(n_849), .C(n_871), .Y(n_846) );
AOI21xp5_ASAP7_75t_L g849 ( .A1(n_850), .A2(n_851), .B(n_869), .Y(n_849) );
OAI21xp5_ASAP7_75t_L g1288 ( .A1(n_850), .A2(n_1289), .B(n_1297), .Y(n_1288) );
NAND3xp33_ASAP7_75t_L g851 ( .A(n_852), .B(n_862), .C(n_866), .Y(n_851) );
AOI222xp33_ASAP7_75t_L g852 ( .A1(n_853), .A2(n_854), .B1(n_855), .B2(n_856), .C1(n_857), .C2(n_861), .Y(n_852) );
AOI222xp33_ASAP7_75t_L g1335 ( .A1(n_853), .A2(n_855), .B1(n_1318), .B2(n_1319), .C1(n_1336), .C2(n_1337), .Y(n_1335) );
NAND2xp5_ASAP7_75t_L g1030 ( .A(n_855), .B(n_1031), .Y(n_1030) );
INVx1_ASAP7_75t_L g858 ( .A(n_859), .Y(n_858) );
INVx1_ASAP7_75t_L g1199 ( .A(n_859), .Y(n_1199) );
BUFx2_ASAP7_75t_L g859 ( .A(n_860), .Y(n_859) );
INVx1_ASAP7_75t_L g1307 ( .A(n_860), .Y(n_1307) );
NAND2xp5_ASAP7_75t_L g1226 ( .A(n_872), .B(n_1227), .Y(n_1226) );
AOI22xp5_ASAP7_75t_L g1270 ( .A1(n_872), .A2(n_1271), .B1(n_1272), .B2(n_1273), .Y(n_1270) );
NAND2xp5_ASAP7_75t_L g873 ( .A(n_874), .B(n_875), .Y(n_873) );
XNOR2x1_ASAP7_75t_L g882 ( .A(n_883), .B(n_971), .Y(n_882) );
XNOR2x1_ASAP7_75t_L g883 ( .A(n_884), .B(n_970), .Y(n_883) );
OR2x2_ASAP7_75t_L g884 ( .A(n_885), .B(n_930), .Y(n_884) );
NAND3xp33_ASAP7_75t_SL g885 ( .A(n_886), .B(n_913), .C(n_925), .Y(n_885) );
AOI211xp5_ASAP7_75t_SL g886 ( .A1(n_887), .A2(n_890), .B(n_896), .C(n_905), .Y(n_886) );
INVxp67_ASAP7_75t_SL g892 ( .A(n_893), .Y(n_892) );
OAI21xp5_ASAP7_75t_L g1676 ( .A1(n_894), .A2(n_903), .B(n_1677), .Y(n_1676) );
INVx2_ASAP7_75t_L g894 ( .A(n_895), .Y(n_894) );
INVx1_ASAP7_75t_L g1016 ( .A(n_897), .Y(n_1016) );
INVx2_ASAP7_75t_SL g1673 ( .A(n_897), .Y(n_1673) );
NAND2x2_ASAP7_75t_L g897 ( .A(n_898), .B(n_900), .Y(n_897) );
INVx1_ASAP7_75t_L g904 ( .A(n_898), .Y(n_904) );
INVx2_ASAP7_75t_L g898 ( .A(n_899), .Y(n_898) );
INVx2_ASAP7_75t_SL g900 ( .A(n_901), .Y(n_900) );
INVx1_ASAP7_75t_SL g1671 ( .A(n_902), .Y(n_1671) );
CKINVDCx5p33_ASAP7_75t_R g1020 ( .A(n_903), .Y(n_1020) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
HB1xp67_ASAP7_75t_L g1007 ( .A(n_911), .Y(n_1007) );
NAND2xp5_ASAP7_75t_L g1667 ( .A(n_911), .B(n_1668), .Y(n_1667) );
AOI222xp33_ASAP7_75t_L g913 ( .A1(n_914), .A2(n_917), .B1(n_918), .B2(n_921), .C1(n_922), .C2(n_924), .Y(n_913) );
AOI21xp33_ASAP7_75t_SL g1018 ( .A1(n_914), .A2(n_1019), .B(n_1020), .Y(n_1018) );
AND2x4_ASAP7_75t_L g914 ( .A(n_915), .B(n_916), .Y(n_914) );
AOI222xp33_ASAP7_75t_L g1014 ( .A1(n_918), .A2(n_982), .B1(n_994), .B2(n_1015), .C1(n_1016), .C2(n_1017), .Y(n_1014) );
INVx1_ASAP7_75t_L g1685 ( .A(n_918), .Y(n_1685) );
INVx1_ASAP7_75t_L g919 ( .A(n_920), .Y(n_919) );
AOI211xp5_ASAP7_75t_L g949 ( .A1(n_921), .A2(n_950), .B(n_953), .C(n_961), .Y(n_949) );
AOI222xp33_ASAP7_75t_L g1002 ( .A1(n_922), .A2(n_983), .B1(n_1003), .B2(n_1007), .C1(n_1008), .C2(n_1011), .Y(n_1002) );
INVx2_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
NAND2xp5_ASAP7_75t_L g925 ( .A(n_926), .B(n_927), .Y(n_925) );
INVx1_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
INVx3_ASAP7_75t_L g928 ( .A(n_929), .Y(n_928) );
HB1xp67_ASAP7_75t_L g973 ( .A(n_929), .Y(n_973) );
A2O1A1Ixp33_ASAP7_75t_L g930 ( .A1(n_931), .A2(n_949), .B(n_967), .C(n_968), .Y(n_930) );
AOI221xp5_ASAP7_75t_L g931 ( .A1(n_932), .A2(n_935), .B1(n_936), .B2(n_940), .C(n_943), .Y(n_931) );
INVx2_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
OAI221xp5_ASAP7_75t_L g985 ( .A1(n_938), .A2(n_986), .B1(n_987), .B2(n_988), .C(n_989), .Y(n_985) );
OAI221xp5_ASAP7_75t_L g1648 ( .A1(n_938), .A2(n_959), .B1(n_1649), .B2(n_1650), .C(n_1651), .Y(n_1648) );
BUFx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx2_ASAP7_75t_L g944 ( .A(n_945), .Y(n_944) );
AOI22xp5_ASAP7_75t_L g993 ( .A1(n_945), .A2(n_948), .B1(n_974), .B2(n_994), .Y(n_993) );
INVx1_ASAP7_75t_L g947 ( .A(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g950 ( .A(n_951), .Y(n_950) );
INVx2_ASAP7_75t_L g951 ( .A(n_952), .Y(n_951) );
INVx4_ASAP7_75t_L g954 ( .A(n_955), .Y(n_954) );
AOI22xp33_ASAP7_75t_L g981 ( .A1(n_955), .A2(n_957), .B1(n_982), .B2(n_983), .Y(n_981) );
INVx2_ASAP7_75t_L g956 ( .A(n_957), .Y(n_956) );
OAI221xp5_ASAP7_75t_L g1643 ( .A1(n_958), .A2(n_1644), .B1(n_1648), .B2(n_1652), .C(n_1656), .Y(n_1643) );
OR2x6_ASAP7_75t_L g958 ( .A(n_959), .B(n_960), .Y(n_958) );
INVx2_ASAP7_75t_L g963 ( .A(n_964), .Y(n_963) );
HB1xp67_ASAP7_75t_L g1663 ( .A(n_964), .Y(n_1663) );
INVx3_ASAP7_75t_L g965 ( .A(n_966), .Y(n_965) );
HB1xp67_ASAP7_75t_L g1050 ( .A(n_967), .Y(n_1050) );
INVx1_ASAP7_75t_L g1364 ( .A(n_967), .Y(n_1364) );
AOI211x1_ASAP7_75t_L g972 ( .A1(n_973), .A2(n_974), .B(n_975), .C(n_1001), .Y(n_972) );
NAND2xp5_ASAP7_75t_L g975 ( .A(n_976), .B(n_978), .Y(n_975) );
NAND3xp33_ASAP7_75t_L g984 ( .A(n_985), .B(n_993), .C(n_995), .Y(n_984) );
INVx3_ASAP7_75t_L g991 ( .A(n_992), .Y(n_991) );
OAI211xp5_ASAP7_75t_L g995 ( .A1(n_996), .A2(n_997), .B(n_999), .C(n_1000), .Y(n_995) );
OAI21xp5_ASAP7_75t_SL g1656 ( .A1(n_997), .A2(n_1657), .B(n_1658), .Y(n_1656) );
INVx3_ASAP7_75t_L g997 ( .A(n_998), .Y(n_997) );
INVx2_ASAP7_75t_L g1258 ( .A(n_998), .Y(n_1258) );
NAND3xp33_ASAP7_75t_L g1001 ( .A(n_1002), .B(n_1014), .C(n_1018), .Y(n_1001) );
INVx1_ASAP7_75t_L g1012 ( .A(n_1013), .Y(n_1012) );
INVx2_ASAP7_75t_L g1021 ( .A(n_1022), .Y(n_1021) );
XNOR2x1_ASAP7_75t_L g1022 ( .A(n_1023), .B(n_1217), .Y(n_1022) );
XNOR2xp5_ASAP7_75t_L g1023 ( .A(n_1024), .B(n_1119), .Y(n_1023) );
INVx1_ASAP7_75t_L g1024 ( .A(n_1025), .Y(n_1024) );
OAI22xp33_ASAP7_75t_L g1025 ( .A1(n_1026), .A2(n_1073), .B1(n_1074), .B2(n_1118), .Y(n_1025) );
INVx2_ASAP7_75t_L g1118 ( .A(n_1026), .Y(n_1118) );
AOI21xp5_ASAP7_75t_L g1028 ( .A1(n_1029), .A2(n_1050), .B(n_1051), .Y(n_1028) );
NAND4xp25_ASAP7_75t_L g1029 ( .A(n_1030), .B(n_1032), .C(n_1041), .D(n_1046), .Y(n_1029) );
OAI22xp5_ASAP7_75t_SL g1055 ( .A1(n_1056), .A2(n_1057), .B1(n_1063), .B2(n_1064), .Y(n_1055) );
OAI221xp5_ASAP7_75t_L g1057 ( .A1(n_1058), .A2(n_1059), .B1(n_1060), .B2(n_1061), .C(n_1062), .Y(n_1057) );
OAI211xp5_ASAP7_75t_L g1277 ( .A1(n_1058), .A2(n_1278), .B(n_1279), .C(n_1280), .Y(n_1277) );
OAI22xp5_ASAP7_75t_L g1652 ( .A1(n_1058), .A2(n_1653), .B1(n_1654), .B2(n_1655), .Y(n_1652) );
INVx2_ASAP7_75t_L g1711 ( .A(n_1058), .Y(n_1711) );
OAI22xp5_ASAP7_75t_L g1251 ( .A1(n_1060), .A2(n_1085), .B1(n_1235), .B2(n_1252), .Y(n_1251) );
OAI22xp5_ASAP7_75t_L g1275 ( .A1(n_1063), .A2(n_1276), .B1(n_1277), .B2(n_1281), .Y(n_1275) );
NAND2xp5_ASAP7_75t_L g1068 ( .A(n_1069), .B(n_1070), .Y(n_1068) );
INVx2_ASAP7_75t_L g1073 ( .A(n_1074), .Y(n_1073) );
NAND3xp33_ASAP7_75t_L g1075 ( .A(n_1076), .B(n_1092), .C(n_1095), .Y(n_1075) );
NOR3xp33_ASAP7_75t_L g1076 ( .A(n_1077), .B(n_1089), .C(n_1091), .Y(n_1076) );
NAND2xp5_ASAP7_75t_L g1077 ( .A(n_1078), .B(n_1081), .Y(n_1077) );
INVx1_ASAP7_75t_L g1084 ( .A(n_1085), .Y(n_1084) );
NOR3xp33_ASAP7_75t_L g1368 ( .A(n_1091), .B(n_1369), .C(n_1381), .Y(n_1368) );
BUFx2_ASAP7_75t_L g1103 ( .A(n_1104), .Y(n_1103) );
HB1xp67_ASAP7_75t_L g1111 ( .A(n_1112), .Y(n_1111) );
HB1xp67_ASAP7_75t_L g1236 ( .A(n_1112), .Y(n_1236) );
INVx1_ASAP7_75t_L g1115 ( .A(n_1116), .Y(n_1115) );
AOI22xp5_ASAP7_75t_L g1119 ( .A1(n_1120), .A2(n_1121), .B1(n_1165), .B2(n_1216), .Y(n_1119) );
INVx1_ASAP7_75t_L g1120 ( .A(n_1121), .Y(n_1120) );
INVx2_ASAP7_75t_L g1121 ( .A(n_1122), .Y(n_1121) );
AO21x2_ASAP7_75t_L g1122 ( .A1(n_1123), .A2(n_1124), .B(n_1164), .Y(n_1122) );
NAND3xp33_ASAP7_75t_SL g1124 ( .A(n_1125), .B(n_1128), .C(n_1147), .Y(n_1124) );
OAI21xp5_ASAP7_75t_L g1128 ( .A1(n_1129), .A2(n_1138), .B(n_1146), .Y(n_1128) );
INVx1_ASAP7_75t_L g1135 ( .A(n_1136), .Y(n_1135) );
INVx1_ASAP7_75t_L g1145 ( .A(n_1136), .Y(n_1145) );
INVx2_ASAP7_75t_L g1140 ( .A(n_1141), .Y(n_1140) );
OAI31xp33_ASAP7_75t_L g1232 ( .A1(n_1146), .A2(n_1233), .A3(n_1239), .B(n_1245), .Y(n_1232) );
INVx1_ASAP7_75t_L g1148 ( .A(n_1149), .Y(n_1148) );
INVx1_ASAP7_75t_L g1155 ( .A(n_1156), .Y(n_1155) );
INVx1_ASAP7_75t_L g1259 ( .A(n_1158), .Y(n_1259) );
INVx1_ASAP7_75t_L g1287 ( .A(n_1162), .Y(n_1287) );
INVx2_ASAP7_75t_L g1216 ( .A(n_1165), .Y(n_1216) );
XOR2x2_ASAP7_75t_L g1165 ( .A(n_1166), .B(n_1215), .Y(n_1165) );
NAND2xp5_ASAP7_75t_SL g1166 ( .A(n_1167), .B(n_1194), .Y(n_1166) );
NAND2xp5_ASAP7_75t_L g1169 ( .A(n_1170), .B(n_1178), .Y(n_1169) );
NOR2xp33_ASAP7_75t_L g1170 ( .A(n_1171), .B(n_1175), .Y(n_1170) );
INVx2_ASAP7_75t_L g1180 ( .A(n_1181), .Y(n_1180) );
INVx1_ASAP7_75t_L g1187 ( .A(n_1188), .Y(n_1187) );
INVx1_ASAP7_75t_L g1188 ( .A(n_1189), .Y(n_1188) );
NAND3xp33_ASAP7_75t_SL g1195 ( .A(n_1196), .B(n_1197), .C(n_1204), .Y(n_1195) );
INVx1_ASAP7_75t_SL g1202 ( .A(n_1203), .Y(n_1202) );
INVx5_ASAP7_75t_L g1213 ( .A(n_1214), .Y(n_1213) );
INVx1_ASAP7_75t_L g1217 ( .A(n_1218), .Y(n_1217) );
AOI22xp5_ASAP7_75t_L g1218 ( .A1(n_1219), .A2(n_1220), .B1(n_1266), .B2(n_1340), .Y(n_1218) );
INVx2_ASAP7_75t_L g1219 ( .A(n_1220), .Y(n_1219) );
XNOR2x1_ASAP7_75t_L g1220 ( .A(n_1221), .B(n_1265), .Y(n_1220) );
NOR2x1_ASAP7_75t_L g1221 ( .A(n_1222), .B(n_1231), .Y(n_1221) );
NAND2xp5_ASAP7_75t_L g1231 ( .A(n_1232), .B(n_1247), .Y(n_1231) );
OAI22xp33_ASAP7_75t_L g1253 ( .A1(n_1242), .A2(n_1254), .B1(n_1257), .B2(n_1258), .Y(n_1253) );
AOI21xp5_ASAP7_75t_SL g1247 ( .A1(n_1248), .A2(n_1249), .B(n_1250), .Y(n_1247) );
INVx2_ASAP7_75t_L g1254 ( .A(n_1255), .Y(n_1254) );
INVx1_ASAP7_75t_L g1255 ( .A(n_1256), .Y(n_1255) );
OAI22xp5_ASAP7_75t_L g1644 ( .A1(n_1256), .A2(n_1645), .B1(n_1646), .B2(n_1647), .Y(n_1644) );
OAI221xp5_ASAP7_75t_L g1281 ( .A1(n_1262), .A2(n_1282), .B1(n_1283), .B2(n_1284), .C(n_1285), .Y(n_1281) );
INVx1_ASAP7_75t_L g1340 ( .A(n_1266), .Y(n_1340) );
XNOR2x1_ASAP7_75t_L g1266 ( .A(n_1267), .B(n_1311), .Y(n_1266) );
NAND4xp75_ASAP7_75t_L g1268 ( .A(n_1269), .B(n_1274), .C(n_1288), .D(n_1309), .Y(n_1268) );
NAND2xp5_ASAP7_75t_L g1289 ( .A(n_1290), .B(n_1294), .Y(n_1289) );
OAI221xp5_ASAP7_75t_L g1298 ( .A1(n_1299), .A2(n_1300), .B1(n_1301), .B2(n_1303), .C(n_1304), .Y(n_1298) );
BUFx3_ASAP7_75t_L g1301 ( .A(n_1302), .Y(n_1301) );
INVx2_ASAP7_75t_L g1305 ( .A(n_1306), .Y(n_1305) );
INVx1_ASAP7_75t_L g1306 ( .A(n_1307), .Y(n_1306) );
AND2x2_ASAP7_75t_L g1312 ( .A(n_1313), .B(n_1327), .Y(n_1312) );
AOI22xp5_ASAP7_75t_L g1320 ( .A1(n_1321), .A2(n_1323), .B1(n_1324), .B2(n_1326), .Y(n_1320) );
NAND3xp33_ASAP7_75t_L g1328 ( .A(n_1329), .B(n_1332), .C(n_1335), .Y(n_1328) );
INVx1_ASAP7_75t_L g1341 ( .A(n_1342), .Y(n_1341) );
NAND3xp33_ASAP7_75t_L g1343 ( .A(n_1344), .B(n_1365), .C(n_1368), .Y(n_1343) );
OAI31xp33_ASAP7_75t_L g1344 ( .A1(n_1345), .A2(n_1351), .A3(n_1362), .B(n_1363), .Y(n_1344) );
NAND2xp5_ASAP7_75t_L g1345 ( .A(n_1346), .B(n_1348), .Y(n_1345) );
OAI211xp5_ASAP7_75t_L g1352 ( .A1(n_1353), .A2(n_1354), .B(n_1355), .C(n_1356), .Y(n_1352) );
INVx1_ASAP7_75t_L g1363 ( .A(n_1364), .Y(n_1363) );
NAND2xp5_ASAP7_75t_L g1369 ( .A(n_1370), .B(n_1373), .Y(n_1369) );
INVx2_ASAP7_75t_L g1378 ( .A(n_1379), .Y(n_1378) );
INVx2_ASAP7_75t_L g1384 ( .A(n_1385), .Y(n_1384) );
OR2x2_ASAP7_75t_L g1385 ( .A(n_1386), .B(n_1392), .Y(n_1385) );
NOR2xp33_ASAP7_75t_L g1740 ( .A(n_1386), .B(n_1395), .Y(n_1740) );
INVx1_ASAP7_75t_L g1386 ( .A(n_1387), .Y(n_1386) );
NOR2xp33_ASAP7_75t_L g1387 ( .A(n_1388), .B(n_1390), .Y(n_1387) );
NOR2xp33_ASAP7_75t_L g1693 ( .A(n_1388), .B(n_1391), .Y(n_1693) );
INVx1_ASAP7_75t_L g1744 ( .A(n_1388), .Y(n_1744) );
HB1xp67_ASAP7_75t_L g1388 ( .A(n_1389), .Y(n_1388) );
INVx1_ASAP7_75t_L g1390 ( .A(n_1391), .Y(n_1390) );
NOR2xp33_ASAP7_75t_L g1746 ( .A(n_1391), .B(n_1744), .Y(n_1746) );
INVx1_ASAP7_75t_L g1392 ( .A(n_1393), .Y(n_1392) );
NAND2xp5_ASAP7_75t_L g1393 ( .A(n_1394), .B(n_1396), .Y(n_1393) );
INVx1_ASAP7_75t_L g1394 ( .A(n_1395), .Y(n_1394) );
AND2x4_ASAP7_75t_SL g1739 ( .A(n_1396), .B(n_1740), .Y(n_1739) );
INVx3_ASAP7_75t_L g1396 ( .A(n_1397), .Y(n_1396) );
OAI221xp5_ASAP7_75t_SL g1399 ( .A1(n_1400), .A2(n_1628), .B1(n_1632), .B2(n_1690), .C(n_1694), .Y(n_1399) );
AND5x1_ASAP7_75t_L g1400 ( .A(n_1401), .B(n_1542), .C(n_1589), .D(n_1611), .E(n_1624), .Y(n_1400) );
OAI31xp33_ASAP7_75t_L g1401 ( .A1(n_1402), .A2(n_1480), .A3(n_1519), .B(n_1533), .Y(n_1401) );
OAI221xp5_ASAP7_75t_L g1402 ( .A1(n_1403), .A2(n_1431), .B1(n_1442), .B2(n_1449), .C(n_1450), .Y(n_1402) );
NAND2x1_ASAP7_75t_L g1403 ( .A(n_1404), .B(n_1419), .Y(n_1403) );
NAND2xp5_ASAP7_75t_SL g1495 ( .A(n_1404), .B(n_1496), .Y(n_1495) );
CKINVDCx5p33_ASAP7_75t_R g1516 ( .A(n_1404), .Y(n_1516) );
OAI21xp33_ASAP7_75t_L g1556 ( .A1(n_1404), .A2(n_1469), .B(n_1557), .Y(n_1556) );
NOR2xp33_ASAP7_75t_L g1562 ( .A(n_1404), .B(n_1563), .Y(n_1562) );
AND2x2_ASAP7_75t_L g1566 ( .A(n_1404), .B(n_1472), .Y(n_1566) );
NOR2x1_ASAP7_75t_L g1571 ( .A(n_1404), .B(n_1572), .Y(n_1571) );
OAI22xp5_ASAP7_75t_SL g1594 ( .A1(n_1404), .A2(n_1550), .B1(n_1595), .B2(n_1599), .Y(n_1594) );
AND2x2_ASAP7_75t_L g1622 ( .A(n_1404), .B(n_1623), .Y(n_1622) );
INVx4_ASAP7_75t_L g1404 ( .A(n_1405), .Y(n_1404) );
INVx4_ASAP7_75t_L g1443 ( .A(n_1405), .Y(n_1443) );
OR2x2_ASAP7_75t_L g1476 ( .A(n_1405), .B(n_1420), .Y(n_1476) );
NAND2xp5_ASAP7_75t_SL g1478 ( .A(n_1405), .B(n_1420), .Y(n_1478) );
NOR2xp33_ASAP7_75t_L g1509 ( .A(n_1405), .B(n_1510), .Y(n_1509) );
NOR3xp33_ASAP7_75t_L g1530 ( .A(n_1405), .B(n_1531), .C(n_1532), .Y(n_1530) );
NOR2xp33_ASAP7_75t_L g1549 ( .A(n_1405), .B(n_1453), .Y(n_1549) );
NOR2xp33_ASAP7_75t_L g1574 ( .A(n_1405), .B(n_1575), .Y(n_1574) );
AND2x4_ASAP7_75t_SL g1405 ( .A(n_1406), .B(n_1414), .Y(n_1405) );
AND2x4_ASAP7_75t_L g1407 ( .A(n_1408), .B(n_1409), .Y(n_1407) );
AND2x6_ASAP7_75t_L g1412 ( .A(n_1408), .B(n_1413), .Y(n_1412) );
AND2x6_ASAP7_75t_L g1415 ( .A(n_1408), .B(n_1416), .Y(n_1415) );
AND2x2_ASAP7_75t_L g1417 ( .A(n_1408), .B(n_1418), .Y(n_1417) );
AND2x2_ASAP7_75t_L g1423 ( .A(n_1408), .B(n_1418), .Y(n_1423) );
AND2x2_ASAP7_75t_L g1436 ( .A(n_1408), .B(n_1418), .Y(n_1436) );
NAND2xp5_ASAP7_75t_L g1537 ( .A(n_1408), .B(n_1409), .Y(n_1537) );
AND2x2_ASAP7_75t_L g1409 ( .A(n_1410), .B(n_1411), .Y(n_1409) );
INVx2_ASAP7_75t_L g1539 ( .A(n_1412), .Y(n_1539) );
OAI21xp5_ASAP7_75t_L g1743 ( .A1(n_1418), .A2(n_1744), .B(n_1745), .Y(n_1743) );
AND2x2_ASAP7_75t_L g1419 ( .A(n_1420), .B(n_1424), .Y(n_1419) );
INVx1_ASAP7_75t_L g1446 ( .A(n_1420), .Y(n_1446) );
OR2x2_ASAP7_75t_L g1497 ( .A(n_1420), .B(n_1498), .Y(n_1497) );
OR2x2_ASAP7_75t_L g1554 ( .A(n_1420), .B(n_1425), .Y(n_1554) );
NAND2xp5_ASAP7_75t_L g1567 ( .A(n_1420), .B(n_1428), .Y(n_1567) );
OR2x2_ASAP7_75t_L g1575 ( .A(n_1420), .B(n_1465), .Y(n_1575) );
AND2x2_ASAP7_75t_L g1598 ( .A(n_1420), .B(n_1465), .Y(n_1598) );
AND2x2_ASAP7_75t_L g1420 ( .A(n_1421), .B(n_1422), .Y(n_1420) );
AND2x2_ASAP7_75t_L g1463 ( .A(n_1421), .B(n_1422), .Y(n_1463) );
INVx1_ASAP7_75t_L g1572 ( .A(n_1424), .Y(n_1572) );
AND2x2_ASAP7_75t_L g1588 ( .A(n_1424), .B(n_1525), .Y(n_1588) );
AND2x2_ASAP7_75t_L g1424 ( .A(n_1425), .B(n_1428), .Y(n_1424) );
NAND2xp5_ASAP7_75t_L g1447 ( .A(n_1425), .B(n_1448), .Y(n_1447) );
OR2x2_ASAP7_75t_L g1453 ( .A(n_1425), .B(n_1428), .Y(n_1453) );
INVx2_ASAP7_75t_L g1465 ( .A(n_1425), .Y(n_1465) );
AOI332xp33_ASAP7_75t_L g1508 ( .A1(n_1425), .A2(n_1463), .A3(n_1501), .B1(n_1509), .B2(n_1511), .B3(n_1514), .C1(n_1517), .C2(n_1518), .Y(n_1508) );
NAND2x1p5_ASAP7_75t_L g1425 ( .A(n_1426), .B(n_1427), .Y(n_1425) );
INVx1_ASAP7_75t_L g1448 ( .A(n_1428), .Y(n_1448) );
AND2x2_ASAP7_75t_L g1464 ( .A(n_1428), .B(n_1465), .Y(n_1464) );
INVx1_ASAP7_75t_L g1498 ( .A(n_1428), .Y(n_1498) );
OR2x2_ASAP7_75t_L g1563 ( .A(n_1428), .B(n_1463), .Y(n_1563) );
NAND3xp33_ASAP7_75t_L g1607 ( .A(n_1428), .B(n_1433), .C(n_1534), .Y(n_1607) );
AND2x2_ASAP7_75t_L g1428 ( .A(n_1429), .B(n_1430), .Y(n_1428) );
OAI21xp33_ASAP7_75t_L g1569 ( .A1(n_1431), .A2(n_1570), .B(n_1573), .Y(n_1569) );
INVx1_ASAP7_75t_L g1431 ( .A(n_1432), .Y(n_1431) );
AND2x2_ASAP7_75t_L g1432 ( .A(n_1433), .B(n_1437), .Y(n_1432) );
INVx3_ASAP7_75t_L g1456 ( .A(n_1433), .Y(n_1456) );
INVx1_ASAP7_75t_L g1515 ( .A(n_1433), .Y(n_1515) );
AND2x2_ASAP7_75t_L g1521 ( .A(n_1433), .B(n_1438), .Y(n_1521) );
OR2x2_ASAP7_75t_L g1532 ( .A(n_1433), .B(n_1438), .Y(n_1532) );
NOR2xp33_ASAP7_75t_SL g1583 ( .A(n_1433), .B(n_1535), .Y(n_1583) );
OAI322xp33_ASAP7_75t_L g1625 ( .A1(n_1433), .A2(n_1471), .A3(n_1474), .B1(n_1520), .B2(n_1554), .C1(n_1626), .C2(n_1627), .Y(n_1625) );
AND2x2_ASAP7_75t_L g1433 ( .A(n_1434), .B(n_1435), .Y(n_1433) );
HB1xp67_ASAP7_75t_L g1631 ( .A(n_1436), .Y(n_1631) );
INVx1_ASAP7_75t_L g1437 ( .A(n_1438), .Y(n_1437) );
INVx2_ASAP7_75t_L g1449 ( .A(n_1438), .Y(n_1449) );
OR2x2_ASAP7_75t_L g1457 ( .A(n_1438), .B(n_1458), .Y(n_1457) );
AND2x2_ASAP7_75t_L g1493 ( .A(n_1438), .B(n_1456), .Y(n_1493) );
AND2x2_ASAP7_75t_L g1501 ( .A(n_1438), .B(n_1472), .Y(n_1501) );
OR2x2_ASAP7_75t_L g1510 ( .A(n_1438), .B(n_1459), .Y(n_1510) );
INVx2_ASAP7_75t_L g1438 ( .A(n_1439), .Y(n_1438) );
OR2x2_ASAP7_75t_L g1470 ( .A(n_1439), .B(n_1458), .Y(n_1470) );
NAND2xp5_ASAP7_75t_L g1439 ( .A(n_1440), .B(n_1441), .Y(n_1439) );
NAND2xp5_ASAP7_75t_L g1442 ( .A(n_1443), .B(n_1444), .Y(n_1442) );
CKINVDCx5p33_ASAP7_75t_R g1468 ( .A(n_1443), .Y(n_1468) );
NOR2xp33_ASAP7_75t_L g1482 ( .A(n_1443), .B(n_1483), .Y(n_1482) );
AND2x2_ASAP7_75t_L g1579 ( .A(n_1443), .B(n_1488), .Y(n_1579) );
OR2x2_ASAP7_75t_L g1593 ( .A(n_1443), .B(n_1558), .Y(n_1593) );
INVx1_ASAP7_75t_L g1444 ( .A(n_1445), .Y(n_1444) );
OAI211xp5_ASAP7_75t_L g1590 ( .A1(n_1445), .A2(n_1527), .B(n_1548), .C(n_1591), .Y(n_1590) );
OR2x2_ASAP7_75t_L g1445 ( .A(n_1446), .B(n_1447), .Y(n_1445) );
AND2x2_ASAP7_75t_L g1451 ( .A(n_1446), .B(n_1452), .Y(n_1451) );
NOR2xp33_ASAP7_75t_L g1485 ( .A(n_1446), .B(n_1465), .Y(n_1485) );
AND2x2_ASAP7_75t_L g1517 ( .A(n_1446), .B(n_1464), .Y(n_1517) );
AND2x2_ASAP7_75t_L g1586 ( .A(n_1446), .B(n_1571), .Y(n_1586) );
OR2x2_ASAP7_75t_L g1618 ( .A(n_1446), .B(n_1453), .Y(n_1618) );
OR2x2_ASAP7_75t_L g1477 ( .A(n_1447), .B(n_1478), .Y(n_1477) );
NAND2xp5_ASAP7_75t_L g1512 ( .A(n_1447), .B(n_1513), .Y(n_1512) );
OR2x2_ASAP7_75t_L g1558 ( .A(n_1447), .B(n_1463), .Y(n_1558) );
INVx1_ASAP7_75t_L g1623 ( .A(n_1447), .Y(n_1623) );
INVx1_ASAP7_75t_L g1550 ( .A(n_1449), .Y(n_1550) );
NAND2xp5_ASAP7_75t_L g1597 ( .A(n_1449), .B(n_1534), .Y(n_1597) );
AOI221xp5_ASAP7_75t_L g1450 ( .A1(n_1451), .A2(n_1454), .B1(n_1462), .B2(n_1466), .C(n_1473), .Y(n_1450) );
AND2x2_ASAP7_75t_L g1528 ( .A(n_1451), .B(n_1468), .Y(n_1528) );
AND2x2_ASAP7_75t_L g1524 ( .A(n_1452), .B(n_1525), .Y(n_1524) );
INVx1_ASAP7_75t_L g1452 ( .A(n_1453), .Y(n_1452) );
OR2x2_ASAP7_75t_L g1503 ( .A(n_1453), .B(n_1476), .Y(n_1503) );
INVx1_ASAP7_75t_L g1454 ( .A(n_1455), .Y(n_1454) );
OR2x2_ASAP7_75t_L g1455 ( .A(n_1456), .B(n_1457), .Y(n_1455) );
NAND2xp5_ASAP7_75t_L g1471 ( .A(n_1456), .B(n_1472), .Y(n_1471) );
OR2x2_ASAP7_75t_L g1479 ( .A(n_1456), .B(n_1472), .Y(n_1479) );
AND2x2_ASAP7_75t_L g1487 ( .A(n_1456), .B(n_1488), .Y(n_1487) );
OR2x2_ASAP7_75t_L g1507 ( .A(n_1456), .B(n_1470), .Y(n_1507) );
CKINVDCx14_ASAP7_75t_R g1568 ( .A(n_1456), .Y(n_1568) );
OR2x2_ASAP7_75t_L g1610 ( .A(n_1456), .B(n_1492), .Y(n_1610) );
CKINVDCx5p33_ASAP7_75t_R g1488 ( .A(n_1457), .Y(n_1488) );
INVx1_ASAP7_75t_L g1492 ( .A(n_1458), .Y(n_1492) );
NOR2xp33_ASAP7_75t_L g1600 ( .A(n_1458), .B(n_1601), .Y(n_1600) );
INVx1_ASAP7_75t_L g1458 ( .A(n_1459), .Y(n_1458) );
INVx1_ASAP7_75t_L g1472 ( .A(n_1459), .Y(n_1472) );
NAND2xp5_ASAP7_75t_L g1459 ( .A(n_1460), .B(n_1461), .Y(n_1459) );
INVx1_ASAP7_75t_L g1531 ( .A(n_1462), .Y(n_1531) );
AOI22xp5_ASAP7_75t_L g1595 ( .A1(n_1462), .A2(n_1518), .B1(n_1596), .B2(n_1598), .Y(n_1595) );
AND2x2_ASAP7_75t_L g1462 ( .A(n_1463), .B(n_1464), .Y(n_1462) );
NAND2xp5_ASAP7_75t_L g1548 ( .A(n_1463), .B(n_1549), .Y(n_1548) );
NAND2xp5_ASAP7_75t_L g1474 ( .A(n_1464), .B(n_1475), .Y(n_1474) );
NAND2xp5_ASAP7_75t_L g1505 ( .A(n_1464), .B(n_1506), .Y(n_1505) );
INVx1_ASAP7_75t_L g1513 ( .A(n_1464), .Y(n_1513) );
OAI311xp33_ASAP7_75t_L g1544 ( .A1(n_1465), .A2(n_1468), .A3(n_1545), .B1(n_1546), .C1(n_1560), .Y(n_1544) );
NAND2xp5_ASAP7_75t_L g1466 ( .A(n_1467), .B(n_1471), .Y(n_1466) );
NAND2xp5_ASAP7_75t_L g1467 ( .A(n_1468), .B(n_1469), .Y(n_1467) );
AND2x2_ASAP7_75t_L g1606 ( .A(n_1468), .B(n_1488), .Y(n_1606) );
O2A1O1Ixp33_ASAP7_75t_L g1624 ( .A1(n_1469), .A2(n_1547), .B(n_1612), .C(n_1625), .Y(n_1624) );
CKINVDCx5p33_ASAP7_75t_R g1469 ( .A(n_1470), .Y(n_1469) );
INVx2_ASAP7_75t_L g1527 ( .A(n_1472), .Y(n_1527) );
AND2x2_ASAP7_75t_L g1555 ( .A(n_1472), .B(n_1516), .Y(n_1555) );
AOI21xp33_ASAP7_75t_L g1473 ( .A1(n_1474), .A2(n_1477), .B(n_1479), .Y(n_1473) );
INVx1_ASAP7_75t_L g1475 ( .A(n_1476), .Y(n_1475) );
NOR2xp33_ASAP7_75t_L g1581 ( .A(n_1477), .B(n_1527), .Y(n_1581) );
INVx1_ASAP7_75t_L g1525 ( .A(n_1478), .Y(n_1525) );
O2A1O1Ixp33_ASAP7_75t_L g1584 ( .A1(n_1479), .A2(n_1518), .B(n_1585), .C(n_1587), .Y(n_1584) );
INVx1_ASAP7_75t_L g1616 ( .A(n_1479), .Y(n_1616) );
OAI211xp5_ASAP7_75t_SL g1480 ( .A1(n_1481), .A2(n_1486), .B(n_1489), .C(n_1508), .Y(n_1480) );
INVx1_ASAP7_75t_L g1481 ( .A(n_1482), .Y(n_1481) );
INVx1_ASAP7_75t_L g1483 ( .A(n_1484), .Y(n_1483) );
HB1xp67_ASAP7_75t_L g1484 ( .A(n_1485), .Y(n_1484) );
INVx1_ASAP7_75t_L g1486 ( .A(n_1487), .Y(n_1486) );
AOI211xp5_ASAP7_75t_L g1489 ( .A1(n_1490), .A2(n_1494), .B(n_1499), .C(n_1504), .Y(n_1489) );
INVx1_ASAP7_75t_L g1490 ( .A(n_1491), .Y(n_1490) );
NAND2xp5_ASAP7_75t_L g1491 ( .A(n_1492), .B(n_1493), .Y(n_1491) );
INVx1_ASAP7_75t_L g1523 ( .A(n_1492), .Y(n_1523) );
O2A1O1Ixp33_ASAP7_75t_L g1580 ( .A1(n_1492), .A2(n_1549), .B(n_1557), .C(n_1581), .Y(n_1580) );
AOI211xp5_ASAP7_75t_L g1589 ( .A1(n_1493), .A2(n_1590), .B(n_1594), .C(n_1602), .Y(n_1589) );
INVxp67_ASAP7_75t_SL g1494 ( .A(n_1495), .Y(n_1494) );
INVx1_ASAP7_75t_L g1496 ( .A(n_1497), .Y(n_1496) );
INVxp67_ASAP7_75t_SL g1499 ( .A(n_1500), .Y(n_1499) );
NAND2xp5_ASAP7_75t_L g1500 ( .A(n_1501), .B(n_1502), .Y(n_1500) );
NAND2xp5_ASAP7_75t_L g1559 ( .A(n_1501), .B(n_1517), .Y(n_1559) );
INVx1_ASAP7_75t_L g1502 ( .A(n_1503), .Y(n_1502) );
INVx1_ASAP7_75t_L g1504 ( .A(n_1505), .Y(n_1504) );
INVx1_ASAP7_75t_L g1506 ( .A(n_1507), .Y(n_1506) );
AOI21xp33_ASAP7_75t_L g1619 ( .A1(n_1507), .A2(n_1620), .B(n_1621), .Y(n_1619) );
INVx1_ASAP7_75t_L g1626 ( .A(n_1509), .Y(n_1626) );
INVx1_ASAP7_75t_L g1518 ( .A(n_1510), .Y(n_1518) );
OR2x2_ASAP7_75t_L g1545 ( .A(n_1510), .B(n_1515), .Y(n_1545) );
INVx1_ASAP7_75t_L g1511 ( .A(n_1512), .Y(n_1511) );
AND2x2_ASAP7_75t_L g1514 ( .A(n_1515), .B(n_1516), .Y(n_1514) );
OAI21xp33_ASAP7_75t_SL g1613 ( .A1(n_1515), .A2(n_1614), .B(n_1615), .Y(n_1613) );
INVx1_ASAP7_75t_L g1603 ( .A(n_1517), .Y(n_1603) );
OAI21xp33_ASAP7_75t_L g1608 ( .A1(n_1518), .A2(n_1592), .B(n_1609), .Y(n_1608) );
OAI211xp5_ASAP7_75t_L g1519 ( .A1(n_1520), .A2(n_1522), .B(n_1526), .C(n_1529), .Y(n_1519) );
INVx1_ASAP7_75t_L g1520 ( .A(n_1521), .Y(n_1520) );
NAND2xp5_ASAP7_75t_L g1573 ( .A(n_1521), .B(n_1574), .Y(n_1573) );
NAND2xp5_ASAP7_75t_L g1522 ( .A(n_1523), .B(n_1524), .Y(n_1522) );
AND2x2_ASAP7_75t_L g1561 ( .A(n_1523), .B(n_1562), .Y(n_1561) );
NAND2xp5_ASAP7_75t_L g1587 ( .A(n_1523), .B(n_1588), .Y(n_1587) );
INVx1_ASAP7_75t_L g1601 ( .A(n_1524), .Y(n_1601) );
NAND2xp5_ASAP7_75t_L g1526 ( .A(n_1527), .B(n_1528), .Y(n_1526) );
NAND2xp5_ASAP7_75t_SL g1591 ( .A(n_1527), .B(n_1592), .Y(n_1591) );
OR2x2_ASAP7_75t_L g1604 ( .A(n_1527), .B(n_1532), .Y(n_1604) );
INVx1_ASAP7_75t_L g1620 ( .A(n_1528), .Y(n_1620) );
INVx1_ASAP7_75t_L g1529 ( .A(n_1530), .Y(n_1529) );
INVx1_ASAP7_75t_L g1543 ( .A(n_1533), .Y(n_1543) );
INVx2_ASAP7_75t_L g1533 ( .A(n_1534), .Y(n_1533) );
INVx1_ASAP7_75t_L g1534 ( .A(n_1535), .Y(n_1534) );
INVx1_ASAP7_75t_L g1535 ( .A(n_1536), .Y(n_1535) );
OAI221xp5_ASAP7_75t_L g1536 ( .A1(n_1537), .A2(n_1538), .B1(n_1539), .B2(n_1540), .C(n_1541), .Y(n_1536) );
AOI211xp5_ASAP7_75t_L g1542 ( .A1(n_1543), .A2(n_1544), .B(n_1576), .C(n_1584), .Y(n_1542) );
AOI221xp5_ASAP7_75t_L g1611 ( .A1(n_1543), .A2(n_1557), .B1(n_1612), .B2(n_1613), .C(n_1619), .Y(n_1611) );
INVx1_ASAP7_75t_L g1612 ( .A(n_1545), .Y(n_1612) );
AOI21xp5_ASAP7_75t_SL g1546 ( .A1(n_1547), .A2(n_1550), .B(n_1551), .Y(n_1546) );
INVx1_ASAP7_75t_L g1547 ( .A(n_1548), .Y(n_1547) );
NAND3xp33_ASAP7_75t_L g1552 ( .A(n_1550), .B(n_1553), .C(n_1555), .Y(n_1552) );
NAND3xp33_ASAP7_75t_SL g1551 ( .A(n_1552), .B(n_1556), .C(n_1559), .Y(n_1551) );
INVx1_ASAP7_75t_L g1553 ( .A(n_1554), .Y(n_1553) );
INVx1_ASAP7_75t_L g1557 ( .A(n_1558), .Y(n_1557) );
O2A1O1Ixp33_ASAP7_75t_L g1560 ( .A1(n_1561), .A2(n_1564), .B(n_1568), .C(n_1569), .Y(n_1560) );
INVxp67_ASAP7_75t_SL g1627 ( .A(n_1564), .Y(n_1627) );
NOR2xp33_ASAP7_75t_L g1564 ( .A(n_1565), .B(n_1567), .Y(n_1564) );
INVx1_ASAP7_75t_L g1565 ( .A(n_1566), .Y(n_1565) );
INVx1_ASAP7_75t_L g1577 ( .A(n_1567), .Y(n_1577) );
INVx1_ASAP7_75t_L g1570 ( .A(n_1571), .Y(n_1570) );
O2A1O1Ixp33_ASAP7_75t_SL g1576 ( .A1(n_1577), .A2(n_1578), .B(n_1580), .C(n_1582), .Y(n_1576) );
INVx1_ASAP7_75t_L g1578 ( .A(n_1579), .Y(n_1578) );
INVx1_ASAP7_75t_L g1582 ( .A(n_1583), .Y(n_1582) );
INVx1_ASAP7_75t_L g1585 ( .A(n_1586), .Y(n_1585) );
INVx1_ASAP7_75t_L g1614 ( .A(n_1588), .Y(n_1614) );
INVx1_ASAP7_75t_L g1592 ( .A(n_1593), .Y(n_1592) );
INVx1_ASAP7_75t_L g1596 ( .A(n_1597), .Y(n_1596) );
INVx1_ASAP7_75t_L g1599 ( .A(n_1600), .Y(n_1599) );
OAI221xp5_ASAP7_75t_L g1602 ( .A1(n_1603), .A2(n_1604), .B1(n_1605), .B2(n_1607), .C(n_1608), .Y(n_1602) );
INVx1_ASAP7_75t_L g1605 ( .A(n_1606), .Y(n_1605) );
INVx1_ASAP7_75t_L g1609 ( .A(n_1610), .Y(n_1609) );
NAND2xp5_ASAP7_75t_L g1615 ( .A(n_1616), .B(n_1617), .Y(n_1615) );
INVx1_ASAP7_75t_L g1617 ( .A(n_1618), .Y(n_1617) );
INVx1_ASAP7_75t_L g1621 ( .A(n_1622), .Y(n_1621) );
CKINVDCx20_ASAP7_75t_R g1628 ( .A(n_1629), .Y(n_1628) );
CKINVDCx20_ASAP7_75t_R g1629 ( .A(n_1630), .Y(n_1629) );
INVx4_ASAP7_75t_L g1630 ( .A(n_1631), .Y(n_1630) );
INVx1_ASAP7_75t_L g1634 ( .A(n_1635), .Y(n_1634) );
HB1xp67_ASAP7_75t_L g1635 ( .A(n_1636), .Y(n_1635) );
NOR2x1_ASAP7_75t_L g1636 ( .A(n_1637), .B(n_1664), .Y(n_1636) );
NAND2xp5_ASAP7_75t_L g1637 ( .A(n_1638), .B(n_1641), .Y(n_1637) );
OAI211xp5_ASAP7_75t_L g1677 ( .A1(n_1649), .A2(n_1678), .B(n_1680), .C(n_1681), .Y(n_1677) );
AOI22xp5_ASAP7_75t_L g1670 ( .A1(n_1661), .A2(n_1671), .B1(n_1672), .B2(n_1673), .Y(n_1670) );
INVx1_ASAP7_75t_L g1662 ( .A(n_1663), .Y(n_1662) );
NAND3xp33_ASAP7_75t_L g1664 ( .A(n_1665), .B(n_1682), .C(n_1686), .Y(n_1664) );
NOR3xp33_ASAP7_75t_SL g1665 ( .A(n_1666), .B(n_1674), .C(n_1676), .Y(n_1665) );
OAI21xp5_ASAP7_75t_SL g1666 ( .A1(n_1667), .A2(n_1669), .B(n_1670), .Y(n_1666) );
INVx2_ASAP7_75t_L g1678 ( .A(n_1679), .Y(n_1678) );
NAND2xp5_ASAP7_75t_L g1682 ( .A(n_1683), .B(n_1684), .Y(n_1682) );
NAND2xp5_ASAP7_75t_L g1686 ( .A(n_1687), .B(n_1688), .Y(n_1686) );
CKINVDCx5p33_ASAP7_75t_R g1690 ( .A(n_1691), .Y(n_1690) );
BUFx3_ASAP7_75t_L g1691 ( .A(n_1692), .Y(n_1691) );
BUFx3_ASAP7_75t_L g1692 ( .A(n_1693), .Y(n_1692) );
INVx1_ASAP7_75t_L g1695 ( .A(n_1696), .Y(n_1695) );
XNOR2x1_ASAP7_75t_L g1696 ( .A(n_1697), .B(n_1738), .Y(n_1696) );
OR2x2_ASAP7_75t_L g1697 ( .A(n_1698), .B(n_1713), .Y(n_1697) );
NAND4xp25_ASAP7_75t_SL g1698 ( .A(n_1699), .B(n_1703), .C(n_1705), .D(n_1709), .Y(n_1698) );
NAND3xp33_ASAP7_75t_SL g1713 ( .A(n_1714), .B(n_1717), .C(n_1719), .Y(n_1713) );
INVx2_ASAP7_75t_L g1724 ( .A(n_1725), .Y(n_1724) );
OAI21xp5_ASAP7_75t_SL g1726 ( .A1(n_1727), .A2(n_1728), .B(n_1731), .Y(n_1726) );
INVx1_ASAP7_75t_L g1741 ( .A(n_1742), .Y(n_1741) );
INVx1_ASAP7_75t_L g1742 ( .A(n_1743), .Y(n_1742) );
INVx1_ASAP7_75t_L g1745 ( .A(n_1746), .Y(n_1745) );
endmodule