module fake_jpeg_11494_n_438 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_438);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_438;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_396;
wire n_375;
wire n_186;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_10),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

HB1xp67_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_12),
.Y(n_22)
);

INVx11_ASAP7_75t_SL g23 ( 
.A(n_7),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_5),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_15),
.Y(n_27)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_9),
.Y(n_29)
);

INVx13_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVxp33_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_1),
.Y(n_33)
);

CKINVDCx16_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_1),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_4),
.Y(n_36)
);

BUFx3_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

BUFx12_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

BUFx3_ASAP7_75t_L g39 ( 
.A(n_1),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_2),
.Y(n_40)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_12),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_6),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_15),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_13),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_43),
.Y(n_47)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_38),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_48),
.B(n_55),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g49 ( 
.A(n_42),
.Y(n_49)
);

INVx5_ASAP7_75t_L g98 ( 
.A(n_49),
.Y(n_98)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_37),
.Y(n_50)
);

INVx3_ASAP7_75t_L g100 ( 
.A(n_50),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_16),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_51),
.Y(n_103)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_22),
.Y(n_52)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_52),
.Y(n_99)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_53),
.Y(n_131)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_16),
.Y(n_54)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_54),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_38),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_16),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_38),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_57),
.B(n_76),
.Y(n_115)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_22),
.Y(n_58)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx11_ASAP7_75t_L g59 ( 
.A(n_28),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g132 ( 
.A(n_59),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_16),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_60),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_17),
.Y(n_61)
);

INVx6_ASAP7_75t_L g96 ( 
.A(n_61),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_32),
.B(n_45),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_62),
.B(n_34),
.Y(n_95)
);

INVx5_ASAP7_75t_L g63 ( 
.A(n_37),
.Y(n_63)
);

BUFx2_ASAP7_75t_L g125 ( 
.A(n_63),
.Y(n_125)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx6_ASAP7_75t_L g142 ( 
.A(n_64),
.Y(n_142)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_17),
.Y(n_65)
);

INVx5_ASAP7_75t_L g144 ( 
.A(n_65),
.Y(n_144)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_66),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_17),
.Y(n_67)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_67),
.Y(n_111)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_45),
.Y(n_68)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_68),
.Y(n_114)
);

BUFx10_ASAP7_75t_L g69 ( 
.A(n_28),
.Y(n_69)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_69),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g70 ( 
.A(n_42),
.Y(n_70)
);

AND2x2_ASAP7_75t_L g116 ( 
.A(n_70),
.B(n_42),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_18),
.Y(n_71)
);

INVx4_ASAP7_75t_L g138 ( 
.A(n_71),
.Y(n_138)
);

BUFx6f_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_72),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_18),
.Y(n_73)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_73),
.Y(n_105)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_22),
.Y(n_74)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_74),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g75 ( 
.A(n_18),
.Y(n_75)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_75),
.Y(n_107)
);

CKINVDCx16_ASAP7_75t_R g76 ( 
.A(n_19),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_32),
.B(n_14),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_77),
.B(n_79),
.Y(n_97)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_78),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_34),
.B(n_14),
.Y(n_79)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_26),
.Y(n_80)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_80),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g81 ( 
.A(n_46),
.Y(n_81)
);

INVx2_ASAP7_75t_L g118 ( 
.A(n_81),
.Y(n_118)
);

BUFx12f_ASAP7_75t_L g82 ( 
.A(n_37),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_84),
.Y(n_126)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_46),
.Y(n_83)
);

INVx2_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_26),
.Y(n_84)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_46),
.Y(n_85)
);

INVx2_ASAP7_75t_L g128 ( 
.A(n_85),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g86 ( 
.A(n_38),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_86),
.B(n_82),
.Y(n_129)
);

INVx8_ASAP7_75t_L g87 ( 
.A(n_27),
.Y(n_87)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_87),
.Y(n_134)
);

BUFx10_ASAP7_75t_L g88 ( 
.A(n_28),
.Y(n_88)
);

INVx2_ASAP7_75t_L g139 ( 
.A(n_88),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_89),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_31),
.B(n_13),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_90),
.B(n_92),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g91 ( 
.A(n_27),
.Y(n_91)
);

INVx2_ASAP7_75t_L g141 ( 
.A(n_91),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_31),
.B(n_9),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_95),
.B(n_117),
.Y(n_166)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_52),
.B(n_19),
.C(n_41),
.Y(n_108)
);

AND2x2_ASAP7_75t_L g149 ( 
.A(n_108),
.B(n_116),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_58),
.B(n_20),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_110),
.B(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_74),
.B(n_20),
.Y(n_112)
);

AND2x2_ASAP7_75t_L g117 ( 
.A(n_70),
.B(n_26),
.Y(n_117)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_50),
.A2(n_41),
.B1(n_39),
.B2(n_33),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_119),
.A2(n_124),
.B1(n_87),
.B2(n_33),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_SL g120 ( 
.A(n_63),
.B(n_20),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g163 ( 
.A(n_120),
.B(n_130),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_89),
.A2(n_41),
.B1(n_44),
.B2(n_27),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_SL g167 ( 
.A1(n_122),
.A2(n_23),
.B1(n_83),
.B2(n_81),
.Y(n_167)
);

AOI22xp33_ASAP7_75t_SL g124 ( 
.A1(n_54),
.A2(n_39),
.B1(n_33),
.B2(n_42),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_129),
.B(n_133),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_82),
.B(n_40),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_49),
.B(n_40),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g135 ( 
.A(n_53),
.B(n_36),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_135),
.B(n_25),
.Y(n_180)
);

AOI22xp5_ASAP7_75t_SL g136 ( 
.A1(n_91),
.A2(n_39),
.B1(n_44),
.B2(n_23),
.Y(n_136)
);

OAI211xp5_ASAP7_75t_L g175 ( 
.A1(n_136),
.A2(n_69),
.B(n_30),
.C(n_21),
.Y(n_175)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_145),
.Y(n_146)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_146),
.Y(n_193)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_145),
.Y(n_147)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_147),
.Y(n_200)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_107),
.Y(n_148)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_148),
.Y(n_224)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_116),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_150),
.B(n_152),
.Y(n_209)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_151),
.A2(n_165),
.B1(n_175),
.B2(n_182),
.Y(n_195)
);

OAI32xp33_ASAP7_75t_L g152 ( 
.A1(n_97),
.A2(n_88),
.A3(n_69),
.B1(n_51),
.B2(n_56),
.Y(n_152)
);

INVx13_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

INVx2_ASAP7_75t_SL g227 ( 
.A(n_153),
.Y(n_227)
);

HAxp5_ASAP7_75t_SL g155 ( 
.A(n_117),
.B(n_88),
.CON(n_155),
.SN(n_155)
);

AND2x2_ASAP7_75t_L g228 ( 
.A(n_155),
.B(n_174),
.Y(n_228)
);

INVx2_ASAP7_75t_SL g156 ( 
.A(n_100),
.Y(n_156)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_156),
.Y(n_201)
);

BUFx2_ASAP7_75t_L g157 ( 
.A(n_98),
.Y(n_157)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_157),
.Y(n_216)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_113),
.Y(n_158)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_158),
.Y(n_205)
);

OAI21xp5_ASAP7_75t_L g159 ( 
.A1(n_115),
.A2(n_29),
.B(n_24),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g211 ( 
.A(n_159),
.B(n_177),
.C(n_123),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_143),
.B(n_35),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g202 ( 
.A(n_160),
.B(n_162),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g161 ( 
.A(n_94),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_161),
.B(n_169),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_108),
.B(n_35),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_93),
.B(n_29),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_164),
.B(n_179),
.Y(n_203)
);

AOI22xp33_ASAP7_75t_SL g165 ( 
.A1(n_125),
.A2(n_24),
.B1(n_21),
.B2(n_36),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g204 ( 
.A1(n_167),
.A2(n_173),
.B1(n_138),
.B2(n_111),
.Y(n_204)
);

HB1xp67_ASAP7_75t_L g168 ( 
.A(n_100),
.Y(n_168)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_168),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_126),
.Y(n_169)
);

INVx5_ASAP7_75t_L g170 ( 
.A(n_98),
.Y(n_170)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_170),
.Y(n_196)
);

INVx2_ASAP7_75t_L g171 ( 
.A(n_118),
.Y(n_171)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_171),
.Y(n_225)
);

INVx4_ASAP7_75t_L g172 ( 
.A(n_131),
.Y(n_172)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

AOI22xp33_ASAP7_75t_L g173 ( 
.A1(n_104),
.A2(n_85),
.B1(n_78),
.B2(n_75),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_101),
.A2(n_44),
.B1(n_72),
.B2(n_71),
.Y(n_177)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_121),
.Y(n_178)
);

INVx5_ASAP7_75t_L g206 ( 
.A(n_178),
.Y(n_206)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_105),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_SL g232 ( 
.A(n_180),
.B(n_0),
.Y(n_232)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_105),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_183),
.Y(n_207)
);

OA22x2_ASAP7_75t_L g182 ( 
.A1(n_136),
.A2(n_73),
.B1(n_67),
.B2(n_65),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_114),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_99),
.B(n_25),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_184),
.B(n_187),
.Y(n_222)
);

CKINVDCx20_ASAP7_75t_R g185 ( 
.A(n_137),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_L g217 ( 
.A(n_185),
.B(n_188),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_119),
.A2(n_44),
.B1(n_59),
.B2(n_60),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_SL g198 ( 
.A1(n_186),
.A2(n_142),
.B1(n_96),
.B2(n_131),
.Y(n_198)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_102),
.Y(n_187)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_144),
.Y(n_188)
);

INVx8_ASAP7_75t_L g189 ( 
.A(n_103),
.Y(n_189)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_189),
.Y(n_208)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_128),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_190),
.B(n_192),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_124),
.A2(n_64),
.B1(n_61),
.B2(n_30),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_132),
.B1(n_142),
.B2(n_96),
.Y(n_199)
);

CKINVDCx20_ASAP7_75t_R g192 ( 
.A(n_144),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g194 ( 
.A(n_162),
.B(n_106),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g243 ( 
.A(n_194),
.B(n_215),
.C(n_220),
.Y(n_243)
);

NOR2xp33_ASAP7_75t_SL g197 ( 
.A(n_166),
.B(n_127),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_197),
.B(n_213),
.Y(n_242)
);

INVxp67_ASAP7_75t_L g234 ( 
.A(n_198),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g262 ( 
.A1(n_199),
.A2(n_223),
.B1(n_178),
.B2(n_171),
.Y(n_262)
);

INVxp33_ASAP7_75t_L g266 ( 
.A(n_204),
.Y(n_266)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_154),
.A2(n_141),
.B1(n_140),
.B2(n_138),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_210),
.A2(n_218),
.B1(n_156),
.B2(n_182),
.Y(n_235)
);

AND2x2_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_172),
.Y(n_259)
);

INVx6_ASAP7_75t_L g212 ( 
.A(n_189),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g263 ( 
.A(n_212),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_161),
.B(n_127),
.Y(n_213)
);

MAJIxp5_ASAP7_75t_L g215 ( 
.A(n_149),
.B(n_134),
.C(n_139),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_167),
.A2(n_111),
.B1(n_123),
.B2(n_109),
.Y(n_218)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_149),
.B(n_109),
.C(n_103),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g223 ( 
.A1(n_149),
.A2(n_30),
.B1(n_38),
.B2(n_3),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_163),
.B(n_0),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_226),
.B(n_229),
.Y(n_251)
);

NOR2xp67_ASAP7_75t_L g229 ( 
.A(n_160),
.B(n_0),
.Y(n_229)
);

AOI22xp33_ASAP7_75t_SL g231 ( 
.A1(n_191),
.A2(n_182),
.B1(n_181),
.B2(n_174),
.Y(n_231)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_232),
.B(n_214),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_202),
.B(n_184),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_233),
.B(n_236),
.Y(n_275)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_235),
.B(n_265),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_202),
.B(n_194),
.Y(n_236)
);

AO21x2_ASAP7_75t_L g237 ( 
.A1(n_222),
.A2(n_203),
.B(n_207),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g281 ( 
.A(n_237),
.B(n_249),
.Y(n_281)
);

A2O1A1O1Ixp25_ASAP7_75t_L g238 ( 
.A1(n_209),
.A2(n_159),
.B(n_176),
.C(n_164),
.D(n_155),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_238),
.B(n_254),
.Y(n_276)
);

INVx1_ASAP7_75t_SL g239 ( 
.A(n_228),
.Y(n_239)
);

INVx2_ASAP7_75t_L g268 ( 
.A(n_239),
.Y(n_268)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_207),
.Y(n_240)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_240),
.Y(n_278)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_200),
.Y(n_241)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_241),
.Y(n_287)
);

OA21x2_ASAP7_75t_L g244 ( 
.A1(n_199),
.A2(n_204),
.B(n_228),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g271 ( 
.A(n_244),
.Y(n_271)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_211),
.A2(n_152),
.B1(n_185),
.B2(n_188),
.Y(n_245)
);

AOI21xp5_ASAP7_75t_L g290 ( 
.A1(n_245),
.A2(n_248),
.B(n_250),
.Y(n_290)
);

INVxp67_ASAP7_75t_SL g246 ( 
.A(n_201),
.Y(n_246)
);

INVxp33_ASAP7_75t_L g291 ( 
.A(n_246),
.Y(n_291)
);

BUFx2_ASAP7_75t_L g247 ( 
.A(n_208),
.Y(n_247)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_247),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_L g248 ( 
.A1(n_195),
.A2(n_177),
.B(n_156),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_222),
.B(n_183),
.Y(n_249)
);

OAI21xp5_ASAP7_75t_SL g250 ( 
.A1(n_228),
.A2(n_182),
.B(n_187),
.Y(n_250)
);

NOR2xp33_ASAP7_75t_SL g279 ( 
.A(n_252),
.B(n_251),
.Y(n_279)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_217),
.Y(n_253)
);

INVx1_ASAP7_75t_L g296 ( 
.A(n_253),
.Y(n_296)
);

INVx1_ASAP7_75t_L g254 ( 
.A(n_200),
.Y(n_254)
);

INVx11_ASAP7_75t_L g255 ( 
.A(n_227),
.Y(n_255)
);

CKINVDCx16_ASAP7_75t_R g284 ( 
.A(n_255),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g256 ( 
.A(n_219),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g280 ( 
.A(n_256),
.B(n_267),
.Y(n_280)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_218),
.A2(n_179),
.B1(n_192),
.B2(n_148),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_257),
.A2(n_224),
.B1(n_193),
.B2(n_216),
.Y(n_289)
);

XOR2xp5_ASAP7_75t_L g273 ( 
.A(n_259),
.B(n_221),
.Y(n_273)
);

AOI22x1_ASAP7_75t_SL g260 ( 
.A1(n_210),
.A2(n_147),
.B1(n_146),
.B2(n_190),
.Y(n_260)
);

AOI21xp5_ASAP7_75t_L g295 ( 
.A1(n_260),
.A2(n_206),
.B(n_230),
.Y(n_295)
);

AO21x2_ASAP7_75t_L g261 ( 
.A1(n_203),
.A2(n_157),
.B(n_170),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g286 ( 
.A(n_261),
.B(n_264),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_262),
.A2(n_225),
.B1(n_205),
.B2(n_224),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_220),
.B(n_215),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_201),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g267 ( 
.A(n_223),
.B(n_158),
.Y(n_267)
);

CKINVDCx20_ASAP7_75t_R g269 ( 
.A(n_255),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_269),
.B(n_270),
.Y(n_305)
);

CKINVDCx20_ASAP7_75t_R g270 ( 
.A(n_249),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g272 ( 
.A(n_236),
.B(n_221),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_272),
.B(n_273),
.C(n_297),
.Y(n_314)
);

CKINVDCx20_ASAP7_75t_R g274 ( 
.A(n_265),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_274),
.B(n_279),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_216),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_SL g308 ( 
.A(n_277),
.B(n_267),
.Y(n_308)
);

OAI22xp33_ASAP7_75t_L g318 ( 
.A1(n_282),
.A2(n_266),
.B1(n_235),
.B2(n_257),
.Y(n_318)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_244),
.A2(n_212),
.B1(n_208),
.B2(n_196),
.Y(n_283)
);

OAI22xp5_ASAP7_75t_SL g315 ( 
.A1(n_283),
.A2(n_261),
.B1(n_258),
.B2(n_248),
.Y(n_315)
);

XOR2x2_ASAP7_75t_L g285 ( 
.A(n_243),
.B(n_225),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g320 ( 
.A(n_285),
.B(n_298),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_289),
.B(n_294),
.Y(n_313)
);

CKINVDCx20_ASAP7_75t_R g292 ( 
.A(n_241),
.Y(n_292)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_292),
.B(n_260),
.Y(n_323)
);

OAI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_245),
.A2(n_196),
.B1(n_230),
.B2(n_193),
.Y(n_294)
);

INVxp67_ASAP7_75t_L g306 ( 
.A(n_295),
.Y(n_306)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_243),
.B(n_227),
.C(n_153),
.Y(n_297)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_264),
.B(n_206),
.Y(n_298)
);

XOR2xp5_ASAP7_75t_L g299 ( 
.A(n_233),
.B(n_227),
.Y(n_299)
);

NAND2xp5_ASAP7_75t_L g319 ( 
.A(n_299),
.B(n_237),
.Y(n_319)
);

AO21x1_ASAP7_75t_L g300 ( 
.A1(n_271),
.A2(n_259),
.B(n_258),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_300),
.Y(n_347)
);

INVx13_ASAP7_75t_L g301 ( 
.A(n_269),
.Y(n_301)
);

HB1xp67_ASAP7_75t_L g341 ( 
.A(n_301),
.Y(n_341)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_286),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_302),
.B(n_308),
.Y(n_342)
);

OA21x2_ASAP7_75t_SL g303 ( 
.A1(n_275),
.A2(n_238),
.B(n_240),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g336 ( 
.A(n_303),
.B(n_327),
.Y(n_336)
);

BUFx3_ASAP7_75t_L g304 ( 
.A(n_296),
.Y(n_304)
);

HB1xp67_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_307),
.Y(n_328)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_287),
.Y(n_309)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_309),
.Y(n_340)
);

BUFx3_ASAP7_75t_L g310 ( 
.A(n_296),
.Y(n_310)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_288),
.Y(n_311)
);

CKINVDCx16_ASAP7_75t_R g329 ( 
.A(n_311),
.Y(n_329)
);

OAI21xp33_ASAP7_75t_L g312 ( 
.A1(n_276),
.A2(n_259),
.B(n_239),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_SL g334 ( 
.A1(n_312),
.A2(n_315),
.B1(n_234),
.B2(n_293),
.Y(n_334)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_282),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g333 ( 
.A(n_316),
.B(n_317),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_270),
.B(n_237),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_318),
.A2(n_325),
.B1(n_293),
.B2(n_244),
.Y(n_331)
);

XNOR2xp5_ASAP7_75t_SL g337 ( 
.A(n_319),
.B(n_273),
.Y(n_337)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_286),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g339 ( 
.A(n_321),
.Y(n_339)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_323),
.B(n_324),
.Y(n_330)
);

INVx1_ASAP7_75t_L g324 ( 
.A(n_278),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g325 ( 
.A1(n_271),
.A2(n_237),
.B1(n_261),
.B2(n_234),
.Y(n_325)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_278),
.Y(n_326)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_326),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g327 ( 
.A(n_275),
.B(n_281),
.Y(n_327)
);

OAI22xp5_ASAP7_75t_L g354 ( 
.A1(n_331),
.A2(n_334),
.B1(n_344),
.B2(n_300),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g332 ( 
.A1(n_302),
.A2(n_293),
.B1(n_294),
.B2(n_281),
.Y(n_332)
);

OAI22xp5_ASAP7_75t_SL g361 ( 
.A1(n_332),
.A2(n_338),
.B1(n_261),
.B2(n_306),
.Y(n_361)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_314),
.B(n_285),
.C(n_298),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g360 ( 
.A(n_335),
.B(n_346),
.C(n_349),
.Y(n_360)
);

XNOR2xp5_ASAP7_75t_L g355 ( 
.A(n_337),
.B(n_327),
.Y(n_355)
);

AOI22xp5_ASAP7_75t_L g338 ( 
.A1(n_321),
.A2(n_266),
.B1(n_299),
.B2(n_290),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g343 ( 
.A1(n_317),
.A2(n_290),
.B1(n_283),
.B2(n_237),
.Y(n_343)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_343),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_300),
.A2(n_295),
.B1(n_261),
.B2(n_280),
.Y(n_344)
);

MAJIxp5_ASAP7_75t_L g346 ( 
.A(n_314),
.B(n_297),
.C(n_272),
.Y(n_346)
);

MAJIxp5_ASAP7_75t_L g349 ( 
.A(n_320),
.B(n_268),
.C(n_274),
.Y(n_349)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_320),
.B(n_268),
.C(n_291),
.Y(n_350)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_350),
.B(n_352),
.C(n_316),
.Y(n_363)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_319),
.B(n_284),
.C(n_250),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_303),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g381 ( 
.A(n_353),
.B(n_356),
.C(n_359),
.Y(n_381)
);

AOI22xp5_ASAP7_75t_L g382 ( 
.A1(n_354),
.A2(n_361),
.B1(n_343),
.B2(n_289),
.Y(n_382)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_355),
.B(n_364),
.Y(n_386)
);

XNOR2xp5_ASAP7_75t_L g356 ( 
.A(n_346),
.B(n_305),
.Y(n_356)
);

INVx1_ASAP7_75t_L g357 ( 
.A(n_328),
.Y(n_357)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_357),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_L g358 ( 
.A(n_336),
.B(n_322),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_SL g383 ( 
.A(n_358),
.B(n_366),
.Y(n_383)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_349),
.B(n_350),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_363),
.B(n_365),
.C(n_372),
.Y(n_384)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_340),
.Y(n_364)
);

XOR2xp5_ASAP7_75t_L g365 ( 
.A(n_337),
.B(n_325),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g366 ( 
.A(n_336),
.B(n_310),
.Y(n_366)
);

OA21x2_ASAP7_75t_SL g367 ( 
.A1(n_342),
.A2(n_324),
.B(n_326),
.Y(n_367)
);

CKINVDCx14_ASAP7_75t_R g374 ( 
.A(n_367),
.Y(n_374)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_341),
.Y(n_368)
);

INVx1_ASAP7_75t_SL g389 ( 
.A(n_368),
.Y(n_389)
);

INVxp67_ASAP7_75t_SL g369 ( 
.A(n_330),
.Y(n_369)
);

OAI22xp5_ASAP7_75t_L g378 ( 
.A1(n_369),
.A2(n_371),
.B1(n_373),
.B2(n_329),
.Y(n_378)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_333),
.Y(n_370)
);

INVxp67_ASAP7_75t_L g376 ( 
.A(n_370),
.Y(n_376)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_304),
.Y(n_371)
);

MAJIxp5_ASAP7_75t_SL g372 ( 
.A(n_352),
.B(n_313),
.C(n_315),
.Y(n_372)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_333),
.Y(n_373)
);

A2O1A1O1Ixp25_ASAP7_75t_L g377 ( 
.A1(n_362),
.A2(n_347),
.B(n_339),
.C(n_338),
.D(n_306),
.Y(n_377)
);

OAI21xp5_ASAP7_75t_SL g395 ( 
.A1(n_377),
.A2(n_301),
.B(n_353),
.Y(n_395)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_378),
.Y(n_399)
);

OAI321xp33_ASAP7_75t_L g379 ( 
.A1(n_362),
.A2(n_308),
.A3(n_313),
.B1(n_347),
.B2(n_334),
.C(n_344),
.Y(n_379)
);

OAI22xp5_ASAP7_75t_L g394 ( 
.A1(n_379),
.A2(n_382),
.B1(n_387),
.B2(n_355),
.Y(n_394)
);

OAI22xp5_ASAP7_75t_L g380 ( 
.A1(n_363),
.A2(n_331),
.B1(n_332),
.B2(n_307),
.Y(n_380)
);

NAND2xp5_ASAP7_75t_L g391 ( 
.A(n_380),
.B(n_385),
.Y(n_391)
);

MAJIxp5_ASAP7_75t_L g385 ( 
.A(n_360),
.B(n_351),
.C(n_348),
.Y(n_385)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_361),
.A2(n_309),
.B1(n_262),
.B2(n_288),
.Y(n_387)
);

MAJIxp5_ASAP7_75t_L g388 ( 
.A(n_360),
.B(n_247),
.C(n_301),
.Y(n_388)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_388),
.B(n_359),
.C(n_356),
.Y(n_390)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_390),
.B(n_389),
.C(n_382),
.Y(n_413)
);

XNOR2xp5_ASAP7_75t_L g392 ( 
.A(n_381),
.B(n_372),
.Y(n_392)
);

XNOR2xp5_ASAP7_75t_L g404 ( 
.A(n_392),
.B(n_397),
.Y(n_404)
);

XNOR2x1_ASAP7_75t_L g393 ( 
.A(n_384),
.B(n_365),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g406 ( 
.A(n_393),
.B(n_395),
.Y(n_406)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_394),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_L g396 ( 
.A1(n_374),
.A2(n_263),
.B1(n_2),
.B2(n_3),
.Y(n_396)
);

MAJIxp5_ASAP7_75t_L g412 ( 
.A(n_396),
.B(n_400),
.C(n_389),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g397 ( 
.A1(n_376),
.A2(n_263),
.B(n_2),
.Y(n_397)
);

OAI21xp5_ASAP7_75t_SL g398 ( 
.A1(n_377),
.A2(n_0),
.B(n_3),
.Y(n_398)
);

HB1xp67_ASAP7_75t_L g411 ( 
.A(n_398),
.Y(n_411)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_388),
.B(n_3),
.C(n_4),
.Y(n_400)
);

AOI21x1_ASAP7_75t_L g401 ( 
.A1(n_376),
.A2(n_4),
.B(n_5),
.Y(n_401)
);

XNOR2xp5_ASAP7_75t_L g405 ( 
.A(n_401),
.B(n_402),
.Y(n_405)
);

XNOR2xp5_ASAP7_75t_L g402 ( 
.A(n_381),
.B(n_4),
.Y(n_402)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_402),
.B(n_385),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g414 ( 
.A(n_407),
.B(n_410),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_391),
.B(n_383),
.Y(n_408)
);

NOR2xp33_ASAP7_75t_SL g417 ( 
.A(n_408),
.B(n_409),
.Y(n_417)
);

NOR2xp33_ASAP7_75t_SL g409 ( 
.A(n_392),
.B(n_386),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_390),
.B(n_384),
.Y(n_410)
);

NAND2xp5_ASAP7_75t_SL g415 ( 
.A(n_412),
.B(n_413),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g416 ( 
.A(n_413),
.B(n_393),
.C(n_399),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g428 ( 
.A(n_416),
.B(n_418),
.Y(n_428)
);

AOI22xp5_ASAP7_75t_L g418 ( 
.A1(n_403),
.A2(n_375),
.B1(n_401),
.B2(n_400),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_406),
.B(n_404),
.Y(n_419)
);

NAND2xp5_ASAP7_75t_SL g424 ( 
.A(n_419),
.B(n_420),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_L g420 ( 
.A1(n_411),
.A2(n_387),
.B1(n_398),
.B2(n_397),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g421 ( 
.A(n_411),
.B(n_5),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_SL g426 ( 
.A(n_421),
.B(n_8),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g422 ( 
.A(n_406),
.B(n_5),
.Y(n_422)
);

INVxp67_ASAP7_75t_L g425 ( 
.A(n_422),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g423 ( 
.A(n_414),
.B(n_405),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_SL g432 ( 
.A(n_423),
.B(n_426),
.Y(n_432)
);

XOR2xp5_ASAP7_75t_L g427 ( 
.A(n_415),
.B(n_6),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g430 ( 
.A(n_427),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_L g429 ( 
.A1(n_424),
.A2(n_417),
.B1(n_416),
.B2(n_422),
.Y(n_429)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_429),
.Y(n_433)
);

OAI21xp5_ASAP7_75t_L g431 ( 
.A1(n_428),
.A2(n_6),
.B(n_7),
.Y(n_431)
);

INVxp67_ASAP7_75t_L g434 ( 
.A(n_431),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_SL g435 ( 
.A1(n_433),
.A2(n_425),
.B1(n_432),
.B2(n_430),
.Y(n_435)
);

OAI221xp5_ASAP7_75t_L g436 ( 
.A1(n_435),
.A2(n_425),
.B1(n_434),
.B2(n_6),
.C(n_8),
.Y(n_436)
);

XOR2xp5_ASAP7_75t_L g437 ( 
.A(n_436),
.B(n_8),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_SL g438 ( 
.A(n_437),
.B(n_8),
.Y(n_438)
);


endmodule