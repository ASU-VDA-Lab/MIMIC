module fake_jpeg_26642_n_132 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_132);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_132;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_21;
wire n_57;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_107;
wire n_39;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_7),
.Y(n_15)
);

INVx2_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

BUFx12f_ASAP7_75t_L g17 ( 
.A(n_12),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_10),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_12),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_6),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_12),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_6),
.Y(n_22)
);

AND2x2_ASAP7_75t_L g23 ( 
.A(n_0),
.B(n_4),
.Y(n_23)
);

BUFx3_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_3),
.B(n_10),
.Y(n_28)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_17),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_29),
.Y(n_39)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_23),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_30),
.B(n_34),
.Y(n_48)
);

BUFx16f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_14),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_32),
.B(n_19),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g33 ( 
.A(n_24),
.Y(n_33)
);

BUFx2_ASAP7_75t_L g46 ( 
.A(n_33),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_0),
.Y(n_34)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_17),
.Y(n_35)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_35),
.Y(n_41)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_25),
.Y(n_36)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_36),
.Y(n_53)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_37),
.Y(n_47)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_38),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_40),
.B(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_28),
.Y(n_42)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_30),
.B(n_23),
.C(n_16),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_43),
.B(n_45),
.C(n_15),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVxp67_ASAP7_75t_L g55 ( 
.A(n_44),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g45 ( 
.A(n_30),
.B(n_28),
.Y(n_45)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_45),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g51 ( 
.A(n_29),
.Y(n_51)
);

INVx2_ASAP7_75t_L g58 ( 
.A(n_51),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_29),
.Y(n_52)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_52),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_32),
.B(n_34),
.Y(n_54)
);

INVxp67_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_53),
.A2(n_36),
.B1(n_37),
.B2(n_20),
.Y(n_56)
);

OAI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_56),
.A2(n_33),
.B1(n_38),
.B2(n_49),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_48),
.A2(n_36),
.B1(n_37),
.B2(n_34),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_62),
.B1(n_70),
.B2(n_33),
.Y(n_79)
);

AOI21xp5_ASAP7_75t_L g60 ( 
.A1(n_44),
.A2(n_33),
.B(n_31),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_SL g81 ( 
.A(n_60),
.B(n_69),
.C(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_48),
.B(n_20),
.Y(n_61)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_61),
.B(n_73),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_53),
.A2(n_36),
.B1(n_26),
.B2(n_29),
.Y(n_62)
);

CKINVDCx16_ASAP7_75t_R g63 ( 
.A(n_46),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_63),
.B(n_66),
.Y(n_80)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_46),
.Y(n_66)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

AND2x6_ASAP7_75t_L g69 ( 
.A(n_43),
.B(n_0),
.Y(n_69)
);

OAI22xp33_ASAP7_75t_SL g70 ( 
.A1(n_47),
.A2(n_38),
.B1(n_26),
.B2(n_35),
.Y(n_70)
);

INVx1_ASAP7_75t_L g71 ( 
.A(n_47),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g84 ( 
.A(n_72),
.B(n_18),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_41),
.B(n_15),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_61),
.B(n_41),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_75),
.B(n_77),
.Y(n_93)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_73),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_59),
.B(n_35),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_68),
.B(n_21),
.Y(n_78)
);

XNOR2x2_ASAP7_75t_SL g100 ( 
.A(n_81),
.B(n_24),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_67),
.B(n_18),
.Y(n_82)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_82),
.Y(n_95)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_70),
.Y(n_83)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_85),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_64),
.B(n_35),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_86),
.B(n_87),
.Y(n_94)
);

NOR2x1_ASAP7_75t_L g87 ( 
.A(n_57),
.B(n_31),
.Y(n_87)
);

XOR2xp5_ASAP7_75t_L g88 ( 
.A(n_72),
.B(n_31),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_89),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g89 ( 
.A(n_69),
.B(n_31),
.Y(n_89)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_60),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_90),
.B(n_35),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_SL g108 ( 
.A(n_91),
.B(n_99),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g92 ( 
.A(n_88),
.B(n_71),
.C(n_69),
.Y(n_92)
);

BUFx2_ASAP7_75t_L g96 ( 
.A(n_80),
.Y(n_96)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_74),
.B(n_66),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_97),
.B(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_86),
.B(n_63),
.Y(n_99)
);

AOI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_100),
.A2(n_27),
.B(n_19),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_74),
.B(n_65),
.Y(n_102)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_38),
.C(n_62),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_101),
.B(n_75),
.C(n_77),
.Y(n_104)
);

MAJIxp5_ASAP7_75t_L g114 ( 
.A(n_104),
.B(n_110),
.C(n_103),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g106 ( 
.A1(n_94),
.A2(n_81),
.B(n_87),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_106),
.A2(n_113),
.B1(n_22),
.B2(n_14),
.Y(n_118)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_95),
.B(n_76),
.Y(n_107)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_107),
.Y(n_119)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_98),
.A2(n_83),
.B1(n_79),
.B2(n_85),
.Y(n_109)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_58),
.B1(n_55),
.B2(n_27),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_92),
.C(n_97),
.Y(n_110)
);

XNOR2xp5_ASAP7_75t_L g112 ( 
.A(n_94),
.B(n_84),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_110),
.B(n_93),
.C(n_100),
.Y(n_115)
);

AO22x1_ASAP7_75t_L g116 ( 
.A1(n_106),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_117),
.A2(n_25),
.B1(n_2),
.B2(n_3),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_118),
.A2(n_22),
.B1(n_108),
.B2(n_105),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g126 ( 
.A(n_120),
.B(n_123),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_114),
.B(n_39),
.C(n_50),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_121),
.B(n_122),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_115),
.B(n_39),
.C(n_50),
.Y(n_122)
);

A2O1A1O1Ixp25_ASAP7_75t_L g124 ( 
.A1(n_116),
.A2(n_13),
.B(n_3),
.C(n_4),
.D(n_5),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_126),
.B(n_119),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_127),
.B(n_128),
.Y(n_129)
);

BUFx24_ASAP7_75t_SL g128 ( 
.A(n_125),
.Y(n_128)
);

AOI21x1_ASAP7_75t_L g130 ( 
.A1(n_129),
.A2(n_8),
.B(n_9),
.Y(n_130)
);

AOI32xp33_ASAP7_75t_L g131 ( 
.A1(n_130),
.A2(n_10),
.A3(n_11),
.B1(n_124),
.B2(n_78),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_131),
.Y(n_132)
);


endmodule