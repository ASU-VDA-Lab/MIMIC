module fake_ariane_2128_n_626 (n_83, n_8, n_56, n_60, n_64, n_38, n_47, n_18, n_86, n_75, n_67, n_34, n_69, n_74, n_33, n_19, n_40, n_12, n_53, n_21, n_66, n_71, n_24, n_7, n_49, n_20, n_17, n_50, n_62, n_51, n_76, n_79, n_26, n_3, n_46, n_0, n_84, n_36, n_72, n_44, n_30, n_82, n_31, n_42, n_57, n_70, n_10, n_85, n_6, n_48, n_4, n_2, n_32, n_37, n_58, n_65, n_9, n_45, n_11, n_52, n_73, n_77, n_15, n_23, n_61, n_22, n_43, n_1, n_81, n_87, n_13, n_27, n_29, n_41, n_55, n_28, n_80, n_14, n_88, n_68, n_78, n_39, n_59, n_63, n_16, n_5, n_35, n_54, n_25, n_626);

input n_83;
input n_8;
input n_56;
input n_60;
input n_64;
input n_38;
input n_47;
input n_18;
input n_86;
input n_75;
input n_67;
input n_34;
input n_69;
input n_74;
input n_33;
input n_19;
input n_40;
input n_12;
input n_53;
input n_21;
input n_66;
input n_71;
input n_24;
input n_7;
input n_49;
input n_20;
input n_17;
input n_50;
input n_62;
input n_51;
input n_76;
input n_79;
input n_26;
input n_3;
input n_46;
input n_0;
input n_84;
input n_36;
input n_72;
input n_44;
input n_30;
input n_82;
input n_31;
input n_42;
input n_57;
input n_70;
input n_10;
input n_85;
input n_6;
input n_48;
input n_4;
input n_2;
input n_32;
input n_37;
input n_58;
input n_65;
input n_9;
input n_45;
input n_11;
input n_52;
input n_73;
input n_77;
input n_15;
input n_23;
input n_61;
input n_22;
input n_43;
input n_1;
input n_81;
input n_87;
input n_13;
input n_27;
input n_29;
input n_41;
input n_55;
input n_28;
input n_80;
input n_14;
input n_88;
input n_68;
input n_78;
input n_39;
input n_59;
input n_63;
input n_16;
input n_5;
input n_35;
input n_54;
input n_25;

output n_626;

wire n_295;
wire n_356;
wire n_556;
wire n_170;
wire n_190;
wire n_160;
wire n_180;
wire n_119;
wire n_124;
wire n_386;
wire n_307;
wire n_516;
wire n_589;
wire n_332;
wire n_581;
wire n_294;
wire n_197;
wire n_463;
wire n_176;
wire n_404;
wire n_172;
wire n_347;
wire n_423;
wire n_183;
wire n_469;
wire n_479;
wire n_603;
wire n_373;
wire n_299;
wire n_541;
wire n_499;
wire n_564;
wire n_133;
wire n_610;
wire n_205;
wire n_341;
wire n_109;
wire n_245;
wire n_421;
wire n_96;
wire n_549;
wire n_522;
wire n_319;
wire n_591;
wire n_416;
wire n_283;
wire n_187;
wire n_525;
wire n_367;
wire n_598;
wire n_345;
wire n_374;
wire n_318;
wire n_103;
wire n_244;
wire n_226;
wire n_220;
wire n_261;
wire n_370;
wire n_189;
wire n_286;
wire n_443;
wire n_586;
wire n_605;
wire n_424;
wire n_528;
wire n_584;
wire n_387;
wire n_406;
wire n_117;
wire n_139;
wire n_524;
wire n_130;
wire n_349;
wire n_391;
wire n_466;
wire n_346;
wire n_214;
wire n_348;
wire n_552;
wire n_462;
wire n_607;
wire n_410;
wire n_379;
wire n_445;
wire n_515;
wire n_138;
wire n_162;
wire n_264;
wire n_137;
wire n_122;
wire n_198;
wire n_232;
wire n_441;
wire n_568;
wire n_385;
wire n_327;
wire n_372;
wire n_377;
wire n_396;
wire n_399;
wire n_554;
wire n_520;
wire n_279;
wire n_207;
wire n_363;
wire n_354;
wire n_140;
wire n_419;
wire n_151;
wire n_146;
wire n_230;
wire n_270;
wire n_194;
wire n_154;
wire n_338;
wire n_142;
wire n_285;
wire n_473;
wire n_186;
wire n_202;
wire n_145;
wire n_193;
wire n_500;
wire n_336;
wire n_315;
wire n_594;
wire n_311;
wire n_239;
wire n_402;
wire n_272;
wire n_339;
wire n_487;
wire n_167;
wire n_90;
wire n_422;
wire n_153;
wire n_269;
wire n_597;
wire n_158;
wire n_259;
wire n_95;
wire n_446;
wire n_553;
wire n_143;
wire n_566;
wire n_578;
wire n_625;
wire n_152;
wire n_405;
wire n_557;
wire n_120;
wire n_169;
wire n_106;
wire n_173;
wire n_242;
wire n_320;
wire n_309;
wire n_115;
wire n_331;
wire n_559;
wire n_401;
wire n_485;
wire n_267;
wire n_495;
wire n_504;
wire n_483;
wire n_335;
wire n_435;
wire n_350;
wire n_291;
wire n_344;
wire n_381;
wire n_426;
wire n_433;
wire n_481;
wire n_600;
wire n_398;
wire n_210;
wire n_200;
wire n_529;
wire n_502;
wire n_166;
wire n_253;
wire n_561;
wire n_218;
wire n_271;
wire n_465;
wire n_486;
wire n_507;
wire n_247;
wire n_569;
wire n_567;
wire n_91;
wire n_240;
wire n_369;
wire n_128;
wire n_224;
wire n_547;
wire n_420;
wire n_562;
wire n_518;
wire n_439;
wire n_604;
wire n_614;
wire n_222;
wire n_478;
wire n_510;
wire n_256;
wire n_326;
wire n_227;
wire n_188;
wire n_323;
wire n_550;
wire n_330;
wire n_400;
wire n_129;
wire n_126;
wire n_282;
wire n_328;
wire n_368;
wire n_590;
wire n_277;
wire n_248;
wire n_301;
wire n_467;
wire n_432;
wire n_545;
wire n_536;
wire n_293;
wire n_620;
wire n_228;
wire n_325;
wire n_276;
wire n_93;
wire n_427;
wire n_108;
wire n_587;
wire n_497;
wire n_303;
wire n_442;
wire n_168;
wire n_206;
wire n_352;
wire n_538;
wire n_576;
wire n_511;
wire n_611;
wire n_238;
wire n_365;
wire n_429;
wire n_455;
wire n_588;
wire n_136;
wire n_334;
wire n_192;
wire n_488;
wire n_300;
wire n_533;
wire n_505;
wire n_163;
wire n_141;
wire n_390;
wire n_498;
wire n_104;
wire n_501;
wire n_438;
wire n_314;
wire n_440;
wire n_273;
wire n_305;
wire n_539;
wire n_312;
wire n_233;
wire n_388;
wire n_333;
wire n_449;
wire n_612;
wire n_413;
wire n_392;
wire n_376;
wire n_512;
wire n_579;
wire n_459;
wire n_221;
wire n_321;
wire n_361;
wire n_458;
wire n_89;
wire n_149;
wire n_383;
wire n_623;
wire n_237;
wire n_175;
wire n_453;
wire n_491;
wire n_181;
wire n_617;
wire n_616;
wire n_570;
wire n_260;
wire n_362;
wire n_543;
wire n_310;
wire n_236;
wire n_601;
wire n_565;
wire n_281;
wire n_461;
wire n_209;
wire n_262;
wire n_490;
wire n_225;
wire n_235;
wire n_464;
wire n_575;
wire n_546;
wire n_297;
wire n_503;
wire n_290;
wire n_527;
wire n_371;
wire n_199;
wire n_107;
wire n_217;
wire n_452;
wire n_178;
wire n_551;
wire n_308;
wire n_417;
wire n_201;
wire n_572;
wire n_343;
wire n_414;
wire n_571;
wire n_287;
wire n_302;
wire n_380;
wire n_582;
wire n_94;
wire n_284;
wire n_448;
wire n_593;
wire n_249;
wire n_534;
wire n_123;
wire n_212;
wire n_355;
wire n_444;
wire n_609;
wire n_278;
wire n_255;
wire n_560;
wire n_450;
wire n_257;
wire n_148;
wire n_451;
wire n_613;
wire n_475;
wire n_135;
wire n_409;
wire n_171;
wire n_519;
wire n_384;
wire n_468;
wire n_526;
wire n_102;
wire n_182;
wire n_482;
wire n_316;
wire n_196;
wire n_125;
wire n_577;
wire n_407;
wire n_254;
wire n_596;
wire n_476;
wire n_460;
wire n_219;
wire n_535;
wire n_231;
wire n_366;
wire n_555;
wire n_234;
wire n_492;
wire n_574;
wire n_280;
wire n_215;
wire n_252;
wire n_161;
wire n_454;
wire n_298;
wire n_532;
wire n_415;
wire n_99;
wire n_544;
wire n_216;
wire n_540;
wire n_599;
wire n_514;
wire n_418;
wire n_537;
wire n_223;
wire n_403;
wire n_389;
wire n_513;
wire n_288;
wire n_179;
wire n_395;
wire n_621;
wire n_195;
wire n_606;
wire n_213;
wire n_110;
wire n_304;
wire n_509;
wire n_583;
wire n_306;
wire n_313;
wire n_92;
wire n_430;
wire n_493;
wire n_203;
wire n_378;
wire n_436;
wire n_150;
wire n_98;
wire n_375;
wire n_113;
wire n_114;
wire n_324;
wire n_585;
wire n_619;
wire n_337;
wire n_437;
wire n_111;
wire n_274;
wire n_622;
wire n_472;
wire n_296;
wire n_265;
wire n_208;
wire n_456;
wire n_156;
wire n_292;
wire n_174;
wire n_275;
wire n_100;
wire n_132;
wire n_147;
wire n_204;
wire n_615;
wire n_521;
wire n_496;
wire n_342;
wire n_246;
wire n_517;
wire n_530;
wire n_428;
wire n_159;
wire n_358;
wire n_105;
wire n_580;
wire n_608;
wire n_494;
wire n_131;
wire n_263;
wire n_434;
wire n_360;
wire n_563;
wire n_229;
wire n_394;
wire n_250;
wire n_165;
wire n_144;
wire n_317;
wire n_101;
wire n_243;
wire n_134;
wire n_329;
wire n_185;
wire n_340;
wire n_289;
wire n_112;
wire n_542;
wire n_548;
wire n_523;
wire n_268;
wire n_266;
wire n_470;
wire n_457;
wire n_164;
wire n_157;
wire n_184;
wire n_177;
wire n_477;
wire n_364;
wire n_258;
wire n_425;
wire n_431;
wire n_508;
wire n_624;
wire n_118;
wire n_121;
wire n_618;
wire n_411;
wire n_484;
wire n_353;
wire n_241;
wire n_357;
wire n_412;
wire n_447;
wire n_191;
wire n_382;
wire n_489;
wire n_480;
wire n_211;
wire n_97;
wire n_408;
wire n_595;
wire n_322;
wire n_251;
wire n_506;
wire n_602;
wire n_558;
wire n_592;
wire n_116;
wire n_397;
wire n_471;
wire n_351;
wire n_393;
wire n_474;
wire n_359;
wire n_155;
wire n_573;
wire n_127;
wire n_531;

HB1xp67_ASAP7_75t_L g89 ( 
.A(n_4),
.Y(n_89)
);

INVx1_ASAP7_75t_SL g90 ( 
.A(n_16),
.Y(n_90)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_49),
.Y(n_91)
);

BUFx3_ASAP7_75t_L g92 ( 
.A(n_54),
.Y(n_92)
);

HB1xp67_ASAP7_75t_L g93 ( 
.A(n_50),
.Y(n_93)
);

CKINVDCx5p33_ASAP7_75t_R g94 ( 
.A(n_67),
.Y(n_94)
);

INVxp33_ASAP7_75t_L g95 ( 
.A(n_76),
.Y(n_95)
);

NOR2xp67_ASAP7_75t_L g96 ( 
.A(n_82),
.B(n_2),
.Y(n_96)
);

CKINVDCx14_ASAP7_75t_R g97 ( 
.A(n_47),
.Y(n_97)
);

CKINVDCx5p33_ASAP7_75t_R g98 ( 
.A(n_20),
.Y(n_98)
);

BUFx5_ASAP7_75t_L g99 ( 
.A(n_68),
.Y(n_99)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_22),
.Y(n_100)
);

CKINVDCx5p33_ASAP7_75t_R g101 ( 
.A(n_79),
.Y(n_101)
);

INVx2_ASAP7_75t_L g102 ( 
.A(n_59),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_17),
.Y(n_103)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_7),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_13),
.Y(n_105)
);

CKINVDCx5p33_ASAP7_75t_R g106 ( 
.A(n_75),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g107 ( 
.A(n_13),
.Y(n_107)
);

NOR2xp67_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_32),
.Y(n_108)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_73),
.Y(n_109)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_1),
.Y(n_110)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_10),
.Y(n_111)
);

CKINVDCx5p33_ASAP7_75t_R g112 ( 
.A(n_12),
.Y(n_112)
);

BUFx2_ASAP7_75t_L g113 ( 
.A(n_57),
.Y(n_113)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_62),
.Y(n_114)
);

INVxp67_ASAP7_75t_SL g115 ( 
.A(n_19),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_39),
.Y(n_116)
);

CKINVDCx5p33_ASAP7_75t_R g117 ( 
.A(n_51),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_80),
.Y(n_118)
);

CKINVDCx5p33_ASAP7_75t_R g119 ( 
.A(n_26),
.Y(n_119)
);

CKINVDCx16_ASAP7_75t_R g120 ( 
.A(n_71),
.Y(n_120)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_83),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_69),
.Y(n_122)
);

INVxp67_ASAP7_75t_L g123 ( 
.A(n_81),
.Y(n_123)
);

CKINVDCx5p33_ASAP7_75t_R g124 ( 
.A(n_33),
.Y(n_124)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_21),
.Y(n_125)
);

INVx2_ASAP7_75t_L g126 ( 
.A(n_25),
.Y(n_126)
);

BUFx2_ASAP7_75t_L g127 ( 
.A(n_61),
.Y(n_127)
);

INVx1_ASAP7_75t_SL g128 ( 
.A(n_88),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_30),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_41),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_72),
.Y(n_131)
);

CKINVDCx20_ASAP7_75t_R g132 ( 
.A(n_52),
.Y(n_132)
);

INVx1_ASAP7_75t_SL g133 ( 
.A(n_5),
.Y(n_133)
);

CKINVDCx5p33_ASAP7_75t_R g134 ( 
.A(n_1),
.Y(n_134)
);

CKINVDCx5p33_ASAP7_75t_R g135 ( 
.A(n_8),
.Y(n_135)
);

HB1xp67_ASAP7_75t_L g136 ( 
.A(n_7),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_37),
.Y(n_137)
);

CKINVDCx5p33_ASAP7_75t_R g138 ( 
.A(n_65),
.Y(n_138)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_77),
.Y(n_139)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_6),
.Y(n_140)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_56),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_29),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_12),
.Y(n_143)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_2),
.Y(n_144)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_43),
.Y(n_145)
);

CKINVDCx16_ASAP7_75t_R g146 ( 
.A(n_3),
.Y(n_146)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_66),
.Y(n_147)
);

CKINVDCx5p33_ASAP7_75t_R g148 ( 
.A(n_48),
.Y(n_148)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_0),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_46),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_15),
.Y(n_151)
);

INVxp67_ASAP7_75t_SL g152 ( 
.A(n_11),
.Y(n_152)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_23),
.Y(n_153)
);

INVx2_ASAP7_75t_L g154 ( 
.A(n_74),
.Y(n_154)
);

CKINVDCx16_ASAP7_75t_R g155 ( 
.A(n_34),
.Y(n_155)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_9),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_63),
.Y(n_157)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_10),
.Y(n_158)
);

INVxp67_ASAP7_75t_SL g159 ( 
.A(n_6),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_31),
.Y(n_160)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_14),
.Y(n_161)
);

CKINVDCx5p33_ASAP7_75t_R g162 ( 
.A(n_87),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_3),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g164 ( 
.A(n_86),
.Y(n_164)
);

BUFx2_ASAP7_75t_L g165 ( 
.A(n_78),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_15),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_85),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_9),
.Y(n_168)
);

CKINVDCx5p33_ASAP7_75t_R g169 ( 
.A(n_4),
.Y(n_169)
);

INVx1_ASAP7_75t_L g170 ( 
.A(n_8),
.Y(n_170)
);

CKINVDCx5p33_ASAP7_75t_R g171 ( 
.A(n_36),
.Y(n_171)
);

INVx1_ASAP7_75t_L g172 ( 
.A(n_27),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_92),
.Y(n_173)
);

INVx1_ASAP7_75t_L g174 ( 
.A(n_104),
.Y(n_174)
);

AND2x4_ASAP7_75t_L g175 ( 
.A(n_110),
.B(n_0),
.Y(n_175)
);

INVx5_ASAP7_75t_L g176 ( 
.A(n_92),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_5),
.Y(n_177)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_105),
.Y(n_178)
);

INVx6_ASAP7_75t_L g179 ( 
.A(n_120),
.Y(n_179)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_111),
.Y(n_180)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_140),
.Y(n_181)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_100),
.Y(n_182)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_143),
.Y(n_183)
);

AND2x4_ASAP7_75t_L g184 ( 
.A(n_110),
.B(n_11),
.Y(n_184)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_149),
.B(n_14),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g186 ( 
.A(n_102),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_127),
.B(n_16),
.Y(n_187)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_144),
.Y(n_188)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_107),
.B(n_17),
.Y(n_189)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx6_ASAP7_75t_L g191 ( 
.A(n_131),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_95),
.B(n_18),
.Y(n_192)
);

INVx2_ASAP7_75t_L g193 ( 
.A(n_114),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_155),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g195 ( 
.A(n_102),
.Y(n_195)
);

INVx2_ASAP7_75t_L g196 ( 
.A(n_118),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g197 ( 
.A1(n_91),
.A2(n_18),
.B1(n_24),
.B2(n_28),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_91),
.A2(n_35),
.B1(n_38),
.B2(n_40),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g199 ( 
.A(n_165),
.B(n_42),
.Y(n_199)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

INVx2_ASAP7_75t_L g201 ( 
.A(n_121),
.Y(n_201)
);

INVx2_ASAP7_75t_L g202 ( 
.A(n_122),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_95),
.B(n_44),
.Y(n_203)
);

AND2x2_ASAP7_75t_L g204 ( 
.A(n_146),
.B(n_89),
.Y(n_204)
);

AND2x2_ASAP7_75t_L g205 ( 
.A(n_136),
.B(n_45),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g206 ( 
.A(n_151),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_156),
.Y(n_207)
);

AND2x4_ASAP7_75t_L g208 ( 
.A(n_126),
.B(n_53),
.Y(n_208)
);

INVx1_ASAP7_75t_L g209 ( 
.A(n_158),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_161),
.Y(n_210)
);

INVx5_ASAP7_75t_L g211 ( 
.A(n_157),
.Y(n_211)
);

INVx2_ASAP7_75t_L g212 ( 
.A(n_125),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g213 ( 
.A(n_126),
.Y(n_213)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_103),
.A2(n_55),
.B1(n_60),
.B2(n_64),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_SL g215 ( 
.A1(n_103),
.A2(n_70),
.B1(n_84),
.B2(n_132),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_129),
.Y(n_216)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_163),
.Y(n_217)
);

CKINVDCx8_ASAP7_75t_R g218 ( 
.A(n_164),
.Y(n_218)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_97),
.B(n_93),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_97),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_116),
.A2(n_132),
.B1(n_90),
.B2(n_133),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_116),
.A2(n_169),
.B1(n_135),
.B2(n_134),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_130),
.B(n_141),
.Y(n_223)
);

INVx1_ASAP7_75t_SL g224 ( 
.A(n_112),
.Y(n_224)
);

AND2x4_ASAP7_75t_L g225 ( 
.A(n_145),
.B(n_154),
.Y(n_225)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_168),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g227 ( 
.A(n_112),
.B(n_134),
.Y(n_227)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_170),
.Y(n_228)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_152),
.Y(n_229)
);

NOR2x1_ASAP7_75t_L g230 ( 
.A(n_137),
.B(n_139),
.Y(n_230)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_159),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_142),
.Y(n_232)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_147),
.Y(n_233)
);

INVx1_ASAP7_75t_L g234 ( 
.A(n_150),
.Y(n_234)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_153),
.Y(n_235)
);

BUFx3_ASAP7_75t_L g236 ( 
.A(n_160),
.Y(n_236)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_167),
.Y(n_237)
);

BUFx6f_ASAP7_75t_L g238 ( 
.A(n_145),
.Y(n_238)
);

BUFx6f_ASAP7_75t_L g239 ( 
.A(n_154),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_SL g240 ( 
.A1(n_135),
.A2(n_169),
.B1(n_166),
.B2(n_98),
.Y(n_240)
);

INVx2_ASAP7_75t_L g241 ( 
.A(n_172),
.Y(n_241)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_94),
.Y(n_242)
);

INVx3_ASAP7_75t_L g243 ( 
.A(n_171),
.Y(n_243)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_99),
.B(n_94),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g245 ( 
.A(n_98),
.Y(n_245)
);

INVx2_ASAP7_75t_L g246 ( 
.A(n_99),
.Y(n_246)
);

AND2x4_ASAP7_75t_L g247 ( 
.A(n_96),
.B(n_123),
.Y(n_247)
);

AND2x4_ASAP7_75t_L g248 ( 
.A(n_108),
.B(n_115),
.Y(n_248)
);

INVx4_ASAP7_75t_L g249 ( 
.A(n_176),
.Y(n_249)
);

BUFx10_ASAP7_75t_L g250 ( 
.A(n_179),
.Y(n_250)
);

HB1xp67_ASAP7_75t_L g251 ( 
.A(n_224),
.Y(n_251)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_186),
.Y(n_252)
);

NAND2xp5_ASAP7_75t_SL g253 ( 
.A(n_208),
.B(n_171),
.Y(n_253)
);

AO22x2_ASAP7_75t_L g254 ( 
.A1(n_208),
.A2(n_128),
.B1(n_99),
.B2(n_106),
.Y(n_254)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_186),
.Y(n_255)
);

INVx3_ASAP7_75t_L g256 ( 
.A(n_186),
.Y(n_256)
);

BUFx2_ASAP7_75t_L g257 ( 
.A(n_194),
.Y(n_257)
);

BUFx3_ASAP7_75t_L g258 ( 
.A(n_173),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_211),
.B(n_148),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_L g260 ( 
.A1(n_225),
.A2(n_101),
.B1(n_106),
.B2(n_117),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_211),
.B(n_148),
.Y(n_261)
);

INVx2_ASAP7_75t_SL g262 ( 
.A(n_211),
.Y(n_262)
);

INVx2_ASAP7_75t_SL g263 ( 
.A(n_211),
.Y(n_263)
);

INVx4_ASAP7_75t_L g264 ( 
.A(n_176),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_174),
.Y(n_265)
);

INVx1_ASAP7_75t_L g266 ( 
.A(n_178),
.Y(n_266)
);

BUFx3_ASAP7_75t_L g267 ( 
.A(n_173),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_180),
.Y(n_268)
);

INVx4_ASAP7_75t_L g269 ( 
.A(n_176),
.Y(n_269)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_219),
.B(n_119),
.Y(n_270)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_176),
.Y(n_271)
);

BUFx6f_ASAP7_75t_L g272 ( 
.A(n_186),
.Y(n_272)
);

INVx4_ASAP7_75t_SL g273 ( 
.A(n_208),
.Y(n_273)
);

INVx6_ASAP7_75t_L g274 ( 
.A(n_173),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_242),
.B(n_124),
.Y(n_275)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

OAI22xp33_ASAP7_75t_L g277 ( 
.A1(n_221),
.A2(n_222),
.B1(n_197),
.B2(n_198),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_195),
.Y(n_278)
);

OR2x6_ASAP7_75t_L g279 ( 
.A(n_215),
.B(n_101),
.Y(n_279)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_181),
.Y(n_280)
);

INVx3_ASAP7_75t_L g281 ( 
.A(n_195),
.Y(n_281)
);

INVx2_ASAP7_75t_SL g282 ( 
.A(n_179),
.Y(n_282)
);

OR2x2_ASAP7_75t_L g283 ( 
.A(n_204),
.B(n_117),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g284 ( 
.A1(n_225),
.A2(n_138),
.B1(n_162),
.B2(n_99),
.Y(n_284)
);

AO21x2_ASAP7_75t_L g285 ( 
.A1(n_199),
.A2(n_138),
.B(n_99),
.Y(n_285)
);

INVx2_ASAP7_75t_L g286 ( 
.A(n_246),
.Y(n_286)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_243),
.B(n_99),
.Y(n_287)
);

BUFx3_ASAP7_75t_L g288 ( 
.A(n_173),
.Y(n_288)
);

OR2x2_ASAP7_75t_L g289 ( 
.A(n_227),
.B(n_99),
.Y(n_289)
);

AND2x4_ASAP7_75t_L g290 ( 
.A(n_248),
.B(n_247),
.Y(n_290)
);

CKINVDCx5p33_ASAP7_75t_R g291 ( 
.A(n_220),
.Y(n_291)
);

AND2x2_ASAP7_75t_L g292 ( 
.A(n_206),
.B(n_200),
.Y(n_292)
);

AND2x4_ASAP7_75t_L g293 ( 
.A(n_248),
.B(n_247),
.Y(n_293)
);

BUFx2_ASAP7_75t_L g294 ( 
.A(n_194),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g295 ( 
.A(n_243),
.B(n_220),
.Y(n_295)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_195),
.Y(n_296)
);

INVx2_ASAP7_75t_L g297 ( 
.A(n_195),
.Y(n_297)
);

OAI21xp5_ASAP7_75t_L g298 ( 
.A1(n_244),
.A2(n_248),
.B(n_230),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_245),
.B(n_247),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g300 ( 
.A(n_179),
.Y(n_300)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_245),
.B(n_232),
.Y(n_301)
);

INVxp33_ASAP7_75t_SL g302 ( 
.A(n_240),
.Y(n_302)
);

INVx4_ASAP7_75t_L g303 ( 
.A(n_213),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_183),
.Y(n_304)
);

AND2x6_ASAP7_75t_L g305 ( 
.A(n_205),
.B(n_175),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_188),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_245),
.B(n_235),
.Y(n_307)
);

AND2x2_ASAP7_75t_L g308 ( 
.A(n_206),
.B(n_200),
.Y(n_308)
);

INVx2_ASAP7_75t_SL g309 ( 
.A(n_191),
.Y(n_309)
);

BUFx2_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

HB1xp67_ASAP7_75t_L g311 ( 
.A(n_300),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_189),
.B1(n_192),
.B2(n_203),
.Y(n_312)
);

AND2x4_ASAP7_75t_L g313 ( 
.A(n_290),
.B(n_175),
.Y(n_313)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_265),
.Y(n_314)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_298),
.B(n_290),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_L g316 ( 
.A(n_290),
.B(n_245),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_L g317 ( 
.A(n_293),
.B(n_191),
.Y(n_317)
);

NOR2xp67_ASAP7_75t_L g318 ( 
.A(n_291),
.B(n_234),
.Y(n_318)
);

INVx2_ASAP7_75t_SL g319 ( 
.A(n_250),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_266),
.Y(n_320)
);

AOI22xp33_ASAP7_75t_L g321 ( 
.A1(n_254),
.A2(n_225),
.B1(n_185),
.B2(n_184),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_293),
.B(n_191),
.Y(n_322)
);

AOI22xp5_ASAP7_75t_L g323 ( 
.A1(n_305),
.A2(n_192),
.B1(n_203),
.B2(n_177),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_293),
.B(n_236),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_275),
.B(n_187),
.Y(n_325)
);

BUFx3_ASAP7_75t_L g326 ( 
.A(n_258),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_268),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_253),
.B(n_299),
.Y(n_328)
);

NAND2xp5_ASAP7_75t_L g329 ( 
.A(n_253),
.B(n_262),
.Y(n_329)
);

NAND2xp5_ASAP7_75t_SL g330 ( 
.A(n_273),
.B(n_289),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_262),
.B(n_236),
.Y(n_331)
);

NAND2xp5_ASAP7_75t_L g332 ( 
.A(n_263),
.B(n_241),
.Y(n_332)
);

AO22x1_ASAP7_75t_L g333 ( 
.A1(n_302),
.A2(n_175),
.B1(n_184),
.B2(n_185),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_263),
.B(n_182),
.Y(n_334)
);

INVx2_ASAP7_75t_L g335 ( 
.A(n_276),
.Y(n_335)
);

OR2x2_ASAP7_75t_L g336 ( 
.A(n_283),
.B(n_257),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g337 ( 
.A(n_273),
.B(n_184),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_273),
.B(n_185),
.Y(n_338)
);

INVx1_ASAP7_75t_L g339 ( 
.A(n_280),
.Y(n_339)
);

AND2x2_ASAP7_75t_L g340 ( 
.A(n_292),
.B(n_218),
.Y(n_340)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_276),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g342 ( 
.A(n_270),
.B(n_182),
.Y(n_342)
);

BUFx6f_ASAP7_75t_SL g343 ( 
.A(n_250),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_295),
.B(n_190),
.Y(n_344)
);

AOI22xp33_ASAP7_75t_L g345 ( 
.A1(n_254),
.A2(n_223),
.B1(n_231),
.B2(n_229),
.Y(n_345)
);

AOI22xp33_ASAP7_75t_L g346 ( 
.A1(n_254),
.A2(n_190),
.B1(n_193),
.B2(n_196),
.Y(n_346)
);

BUFx12f_ASAP7_75t_L g347 ( 
.A(n_250),
.Y(n_347)
);

NOR2xp33_ASAP7_75t_L g348 ( 
.A(n_289),
.B(n_193),
.Y(n_348)
);

NOR3xp33_ASAP7_75t_L g349 ( 
.A(n_277),
.B(n_214),
.C(n_226),
.Y(n_349)
);

NOR2xp33_ASAP7_75t_L g350 ( 
.A(n_301),
.B(n_196),
.Y(n_350)
);

NAND2xp5_ASAP7_75t_SL g351 ( 
.A(n_273),
.B(n_239),
.Y(n_351)
);

AOI22xp33_ASAP7_75t_L g352 ( 
.A1(n_254),
.A2(n_201),
.B1(n_202),
.B2(n_241),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g353 ( 
.A1(n_305),
.A2(n_201),
.B1(n_202),
.B2(n_237),
.Y(n_353)
);

AOI22xp33_ASAP7_75t_L g354 ( 
.A1(n_305),
.A2(n_237),
.B1(n_212),
.B2(n_216),
.Y(n_354)
);

AOI22xp5_ASAP7_75t_L g355 ( 
.A1(n_305),
.A2(n_216),
.B1(n_233),
.B2(n_212),
.Y(n_355)
);

OR2x6_ASAP7_75t_L g356 ( 
.A(n_279),
.B(n_233),
.Y(n_356)
);

INVx2_ASAP7_75t_L g357 ( 
.A(n_286),
.Y(n_357)
);

AOI22xp33_ASAP7_75t_L g358 ( 
.A1(n_305),
.A2(n_239),
.B1(n_238),
.B2(n_213),
.Y(n_358)
);

NAND2xp5_ASAP7_75t_L g359 ( 
.A(n_259),
.B(n_261),
.Y(n_359)
);

NOR2xp67_ASAP7_75t_L g360 ( 
.A(n_291),
.B(n_207),
.Y(n_360)
);

AOI22xp33_ASAP7_75t_SL g361 ( 
.A1(n_302),
.A2(n_209),
.B1(n_210),
.B2(n_217),
.Y(n_361)
);

INVx2_ASAP7_75t_SL g362 ( 
.A(n_283),
.Y(n_362)
);

NAND2xp5_ASAP7_75t_L g363 ( 
.A(n_307),
.B(n_213),
.Y(n_363)
);

INVx1_ASAP7_75t_L g364 ( 
.A(n_304),
.Y(n_364)
);

CKINVDCx5p33_ASAP7_75t_R g365 ( 
.A(n_294),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_306),
.Y(n_366)
);

INVx1_ASAP7_75t_L g367 ( 
.A(n_314),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g368 ( 
.A(n_310),
.B(n_292),
.Y(n_368)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_335),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g370 ( 
.A(n_348),
.B(n_325),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_320),
.Y(n_371)
);

AND2x2_ASAP7_75t_L g372 ( 
.A(n_311),
.B(n_308),
.Y(n_372)
);

NOR2xp33_ASAP7_75t_L g373 ( 
.A(n_325),
.B(n_309),
.Y(n_373)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_348),
.B(n_286),
.Y(n_374)
);

INVx1_ASAP7_75t_L g375 ( 
.A(n_327),
.Y(n_375)
);

AOI21xp5_ASAP7_75t_L g376 ( 
.A1(n_359),
.A2(n_344),
.B(n_342),
.Y(n_376)
);

INVx1_ASAP7_75t_SL g377 ( 
.A(n_340),
.Y(n_377)
);

AOI21xp5_ASAP7_75t_L g378 ( 
.A1(n_328),
.A2(n_316),
.B(n_330),
.Y(n_378)
);

NAND2xp33_ASAP7_75t_L g379 ( 
.A(n_319),
.B(n_287),
.Y(n_379)
);

AOI21xp5_ASAP7_75t_L g380 ( 
.A1(n_330),
.A2(n_285),
.B(n_282),
.Y(n_380)
);

OR2x2_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_309),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_SL g382 ( 
.A(n_318),
.B(n_260),
.Y(n_382)
);

AOI21xp5_ASAP7_75t_L g383 ( 
.A1(n_329),
.A2(n_285),
.B(n_282),
.Y(n_383)
);

BUFx4f_ASAP7_75t_L g384 ( 
.A(n_347),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_360),
.B(n_284),
.Y(n_385)
);

NOR2xp33_ASAP7_75t_L g386 ( 
.A(n_362),
.B(n_315),
.Y(n_386)
);

INVx2_ASAP7_75t_L g387 ( 
.A(n_335),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_339),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_313),
.B(n_285),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g390 ( 
.A(n_326),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_SL g391 ( 
.A(n_313),
.B(n_308),
.Y(n_391)
);

BUFx6f_ASAP7_75t_L g392 ( 
.A(n_326),
.Y(n_392)
);

BUFx6f_ASAP7_75t_L g393 ( 
.A(n_313),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g394 ( 
.A1(n_361),
.A2(n_279),
.B1(n_356),
.B2(n_365),
.Y(n_394)
);

CKINVDCx16_ASAP7_75t_R g395 ( 
.A(n_347),
.Y(n_395)
);

AO32x1_ASAP7_75t_L g396 ( 
.A1(n_341),
.A2(n_303),
.A3(n_297),
.B1(n_296),
.B2(n_228),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g397 ( 
.A(n_350),
.B(n_303),
.Y(n_397)
);

NOR3xp33_ASAP7_75t_L g398 ( 
.A(n_365),
.B(n_279),
.C(n_303),
.Y(n_398)
);

NAND2xp5_ASAP7_75t_L g399 ( 
.A(n_350),
.B(n_252),
.Y(n_399)
);

BUFx2_ASAP7_75t_L g400 ( 
.A(n_362),
.Y(n_400)
);

BUFx3_ASAP7_75t_L g401 ( 
.A(n_364),
.Y(n_401)
);

INVx2_ASAP7_75t_L g402 ( 
.A(n_341),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_366),
.Y(n_403)
);

A2O1A1Ixp33_ASAP7_75t_L g404 ( 
.A1(n_312),
.A2(n_252),
.B(n_256),
.C(n_278),
.Y(n_404)
);

NOR2xp33_ASAP7_75t_L g405 ( 
.A(n_317),
.B(n_279),
.Y(n_405)
);

AOI22xp5_ASAP7_75t_L g406 ( 
.A1(n_349),
.A2(n_267),
.B1(n_288),
.B2(n_258),
.Y(n_406)
);

INVx1_ASAP7_75t_L g407 ( 
.A(n_363),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_SL g408 ( 
.A(n_323),
.B(n_288),
.Y(n_408)
);

INVx2_ASAP7_75t_L g409 ( 
.A(n_357),
.Y(n_409)
);

NAND2xp5_ASAP7_75t_L g410 ( 
.A(n_333),
.B(n_281),
.Y(n_410)
);

BUFx2_ASAP7_75t_L g411 ( 
.A(n_356),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_SL g412 ( 
.A(n_356),
.B(n_271),
.Y(n_412)
);

NAND2xp33_ASAP7_75t_L g413 ( 
.A(n_354),
.B(n_272),
.Y(n_413)
);

INVx2_ASAP7_75t_L g414 ( 
.A(n_357),
.Y(n_414)
);

AND2x2_ASAP7_75t_L g415 ( 
.A(n_322),
.B(n_324),
.Y(n_415)
);

CKINVDCx5p33_ASAP7_75t_R g416 ( 
.A(n_343),
.Y(n_416)
);

OR2x6_ASAP7_75t_L g417 ( 
.A(n_356),
.B(n_338),
.Y(n_417)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_337),
.A2(n_297),
.B(n_296),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g419 ( 
.A(n_346),
.B(n_278),
.Y(n_419)
);

NAND2x1p5_ASAP7_75t_L g420 ( 
.A(n_337),
.B(n_267),
.Y(n_420)
);

INVx2_ASAP7_75t_L g421 ( 
.A(n_332),
.Y(n_421)
);

INVx1_ASAP7_75t_L g422 ( 
.A(n_334),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g423 ( 
.A(n_352),
.B(n_281),
.Y(n_423)
);

INVx2_ASAP7_75t_L g424 ( 
.A(n_351),
.Y(n_424)
);

BUFx6f_ASAP7_75t_L g425 ( 
.A(n_351),
.Y(n_425)
);

INVx2_ASAP7_75t_L g426 ( 
.A(n_338),
.Y(n_426)
);

AND2x2_ASAP7_75t_SL g427 ( 
.A(n_321),
.B(n_264),
.Y(n_427)
);

AND2x2_ASAP7_75t_L g428 ( 
.A(n_345),
.B(n_281),
.Y(n_428)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_353),
.Y(n_429)
);

OR2x2_ASAP7_75t_L g430 ( 
.A(n_331),
.B(n_256),
.Y(n_430)
);

AOI21xp5_ASAP7_75t_L g431 ( 
.A1(n_355),
.A2(n_256),
.B(n_278),
.Y(n_431)
);

BUFx6f_ASAP7_75t_L g432 ( 
.A(n_358),
.Y(n_432)
);

AND2x2_ASAP7_75t_L g433 ( 
.A(n_310),
.B(n_252),
.Y(n_433)
);

AOI22xp33_ASAP7_75t_SL g434 ( 
.A1(n_356),
.A2(n_213),
.B1(n_238),
.B2(n_239),
.Y(n_434)
);

BUFx6f_ASAP7_75t_L g435 ( 
.A(n_326),
.Y(n_435)
);

BUFx2_ASAP7_75t_L g436 ( 
.A(n_310),
.Y(n_436)
);

NOR2xp33_ASAP7_75t_L g437 ( 
.A(n_325),
.B(n_274),
.Y(n_437)
);

AO31x2_ASAP7_75t_L g438 ( 
.A1(n_404),
.A2(n_269),
.A3(n_249),
.B(n_271),
.Y(n_438)
);

AOI221xp5_ASAP7_75t_L g439 ( 
.A1(n_394),
.A2(n_238),
.B1(n_272),
.B2(n_255),
.C(n_264),
.Y(n_439)
);

A2O1A1Ixp33_ASAP7_75t_L g440 ( 
.A1(n_386),
.A2(n_255),
.B(n_272),
.C(n_274),
.Y(n_440)
);

OAI21xp5_ASAP7_75t_L g441 ( 
.A1(n_378),
.A2(n_249),
.B(n_264),
.Y(n_441)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_367),
.Y(n_442)
);

AO32x2_ASAP7_75t_L g443 ( 
.A1(n_396),
.A2(n_249),
.A3(n_269),
.B1(n_271),
.B2(n_255),
.Y(n_443)
);

BUFx3_ASAP7_75t_L g444 ( 
.A(n_436),
.Y(n_444)
);

INVx4_ASAP7_75t_L g445 ( 
.A(n_384),
.Y(n_445)
);

OAI21xp5_ASAP7_75t_L g446 ( 
.A1(n_378),
.A2(n_269),
.B(n_376),
.Y(n_446)
);

O2A1O1Ixp33_ASAP7_75t_L g447 ( 
.A1(n_370),
.A2(n_373),
.B(n_391),
.C(n_408),
.Y(n_447)
);

OAI21x1_ASAP7_75t_L g448 ( 
.A1(n_380),
.A2(n_418),
.B(n_431),
.Y(n_448)
);

OAI21x1_ASAP7_75t_L g449 ( 
.A1(n_431),
.A2(n_383),
.B(n_389),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_371),
.Y(n_450)
);

OAI211xp5_ASAP7_75t_L g451 ( 
.A1(n_400),
.A2(n_370),
.B(n_381),
.C(n_382),
.Y(n_451)
);

A2O1A1Ixp33_ASAP7_75t_L g452 ( 
.A1(n_405),
.A2(n_385),
.B(n_415),
.C(n_437),
.Y(n_452)
);

INVxp67_ASAP7_75t_L g453 ( 
.A(n_368),
.Y(n_453)
);

OAI21xp5_ASAP7_75t_L g454 ( 
.A1(n_397),
.A2(n_389),
.B(n_399),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g455 ( 
.A(n_372),
.Y(n_455)
);

AO31x2_ASAP7_75t_L g456 ( 
.A1(n_419),
.A2(n_423),
.A3(n_374),
.B(n_402),
.Y(n_456)
);

BUFx10_ASAP7_75t_L g457 ( 
.A(n_416),
.Y(n_457)
);

BUFx2_ASAP7_75t_L g458 ( 
.A(n_411),
.Y(n_458)
);

AOI22xp5_ASAP7_75t_L g459 ( 
.A1(n_393),
.A2(n_398),
.B1(n_377),
.B2(n_412),
.Y(n_459)
);

AOI22xp33_ASAP7_75t_L g460 ( 
.A1(n_428),
.A2(n_427),
.B1(n_401),
.B2(n_432),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_369),
.Y(n_461)
);

A2O1A1Ixp33_ASAP7_75t_L g462 ( 
.A1(n_426),
.A2(n_429),
.B(n_375),
.C(n_403),
.Y(n_462)
);

AOI21xp33_ASAP7_75t_L g463 ( 
.A1(n_410),
.A2(n_423),
.B(n_419),
.Y(n_463)
);

BUFx2_ASAP7_75t_R g464 ( 
.A(n_410),
.Y(n_464)
);

A2O1A1Ixp33_ASAP7_75t_L g465 ( 
.A1(n_388),
.A2(n_422),
.B(n_407),
.C(n_374),
.Y(n_465)
);

NAND2x1p5_ASAP7_75t_L g466 ( 
.A(n_393),
.B(n_384),
.Y(n_466)
);

CKINVDCx20_ASAP7_75t_R g467 ( 
.A(n_395),
.Y(n_467)
);

OAI22xp5_ASAP7_75t_L g468 ( 
.A1(n_393),
.A2(n_397),
.B1(n_417),
.B2(n_399),
.Y(n_468)
);

INVx3_ASAP7_75t_L g469 ( 
.A(n_390),
.Y(n_469)
);

A2O1A1Ixp33_ASAP7_75t_L g470 ( 
.A1(n_421),
.A2(n_406),
.B(n_424),
.C(n_412),
.Y(n_470)
);

INVx1_ASAP7_75t_L g471 ( 
.A(n_387),
.Y(n_471)
);

OAI22x1_ASAP7_75t_L g472 ( 
.A1(n_433),
.A2(n_420),
.B1(n_417),
.B2(n_430),
.Y(n_472)
);

AO31x2_ASAP7_75t_L g473 ( 
.A1(n_409),
.A2(n_414),
.A3(n_396),
.B(n_413),
.Y(n_473)
);

OR2x6_ASAP7_75t_L g474 ( 
.A(n_390),
.B(n_435),
.Y(n_474)
);

AOI21xp5_ASAP7_75t_L g475 ( 
.A1(n_379),
.A2(n_420),
.B(n_396),
.Y(n_475)
);

AOI22xp33_ASAP7_75t_L g476 ( 
.A1(n_432),
.A2(n_425),
.B1(n_434),
.B2(n_392),
.Y(n_476)
);

AOI21xp5_ASAP7_75t_L g477 ( 
.A1(n_425),
.A2(n_370),
.B(n_376),
.Y(n_477)
);

AO31x2_ASAP7_75t_L g478 ( 
.A1(n_432),
.A2(n_404),
.A3(n_383),
.B(n_380),
.Y(n_478)
);

AND2x4_ASAP7_75t_L g479 ( 
.A(n_436),
.B(n_311),
.Y(n_479)
);

AOI21xp5_ASAP7_75t_L g480 ( 
.A1(n_370),
.A2(n_376),
.B(n_359),
.Y(n_480)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_386),
.A2(n_349),
.B1(n_405),
.B2(n_394),
.Y(n_481)
);

O2A1O1Ixp33_ASAP7_75t_SL g482 ( 
.A1(n_370),
.A2(n_404),
.B(n_359),
.C(n_373),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_L g483 ( 
.A(n_370),
.B(n_251),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_370),
.B(n_373),
.Y(n_484)
);

O2A1O1Ixp33_ASAP7_75t_L g485 ( 
.A1(n_370),
.A2(n_373),
.B(n_362),
.C(n_386),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g486 ( 
.A(n_370),
.B(n_373),
.Y(n_486)
);

AOI21xp5_ASAP7_75t_L g487 ( 
.A1(n_370),
.A2(n_376),
.B(n_359),
.Y(n_487)
);

NAND2xp5_ASAP7_75t_L g488 ( 
.A(n_370),
.B(n_373),
.Y(n_488)
);

AND2x4_ASAP7_75t_L g489 ( 
.A(n_417),
.B(n_393),
.Y(n_489)
);

AO32x2_ASAP7_75t_L g490 ( 
.A1(n_394),
.A2(n_396),
.A3(n_303),
.B1(n_362),
.B2(n_214),
.Y(n_490)
);

INVxp67_ASAP7_75t_SL g491 ( 
.A(n_393),
.Y(n_491)
);

O2A1O1Ixp33_ASAP7_75t_SL g492 ( 
.A1(n_370),
.A2(n_404),
.B(n_359),
.C(n_373),
.Y(n_492)
);

AOI21xp5_ASAP7_75t_L g493 ( 
.A1(n_370),
.A2(n_376),
.B(n_359),
.Y(n_493)
);

AOI21xp5_ASAP7_75t_L g494 ( 
.A1(n_370),
.A2(n_376),
.B(n_359),
.Y(n_494)
);

INVx1_ASAP7_75t_L g495 ( 
.A(n_367),
.Y(n_495)
);

O2A1O1Ixp33_ASAP7_75t_SL g496 ( 
.A1(n_370),
.A2(n_404),
.B(n_359),
.C(n_373),
.Y(n_496)
);

AO32x2_ASAP7_75t_L g497 ( 
.A1(n_394),
.A2(n_396),
.A3(n_303),
.B1(n_362),
.B2(n_214),
.Y(n_497)
);

INVx1_ASAP7_75t_L g498 ( 
.A(n_367),
.Y(n_498)
);

INVx1_ASAP7_75t_L g499 ( 
.A(n_367),
.Y(n_499)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_499),
.Y(n_500)
);

BUFx3_ASAP7_75t_L g501 ( 
.A(n_444),
.Y(n_501)
);

OR2x6_ASAP7_75t_L g502 ( 
.A(n_489),
.B(n_466),
.Y(n_502)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_442),
.Y(n_503)
);

AOI22xp5_ASAP7_75t_L g504 ( 
.A1(n_483),
.A2(n_481),
.B1(n_479),
.B2(n_484),
.Y(n_504)
);

AOI21xp5_ASAP7_75t_L g505 ( 
.A1(n_480),
.A2(n_493),
.B(n_494),
.Y(n_505)
);

BUFx3_ASAP7_75t_L g506 ( 
.A(n_467),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g507 ( 
.A(n_486),
.B(n_488),
.Y(n_507)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_450),
.Y(n_508)
);

AOI21xp33_ASAP7_75t_L g509 ( 
.A1(n_451),
.A2(n_453),
.B(n_472),
.Y(n_509)
);

AND2x2_ASAP7_75t_L g510 ( 
.A(n_455),
.B(n_458),
.Y(n_510)
);

OR2x2_ASAP7_75t_L g511 ( 
.A(n_495),
.B(n_498),
.Y(n_511)
);

OAI21x1_ASAP7_75t_L g512 ( 
.A1(n_449),
.A2(n_448),
.B(n_446),
.Y(n_512)
);

AND2x2_ASAP7_75t_L g513 ( 
.A(n_464),
.B(n_460),
.Y(n_513)
);

AOI22xp33_ASAP7_75t_L g514 ( 
.A1(n_439),
.A2(n_463),
.B1(n_454),
.B2(n_471),
.Y(n_514)
);

OA21x2_ASAP7_75t_L g515 ( 
.A1(n_475),
.A2(n_487),
.B(n_477),
.Y(n_515)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_462),
.Y(n_516)
);

BUFx2_ASAP7_75t_L g517 ( 
.A(n_474),
.Y(n_517)
);

AOI22xp33_ASAP7_75t_L g518 ( 
.A1(n_468),
.A2(n_459),
.B1(n_476),
.B2(n_491),
.Y(n_518)
);

OAI21xp5_ASAP7_75t_L g519 ( 
.A1(n_447),
.A2(n_465),
.B(n_485),
.Y(n_519)
);

AOI222xp33_ASAP7_75t_L g520 ( 
.A1(n_452),
.A2(n_445),
.B1(n_497),
.B2(n_490),
.C1(n_470),
.C2(n_469),
.Y(n_520)
);

OA21x2_ASAP7_75t_L g521 ( 
.A1(n_440),
.A2(n_441),
.B(n_443),
.Y(n_521)
);

AOI21xp5_ASAP7_75t_L g522 ( 
.A1(n_482),
.A2(n_496),
.B(n_492),
.Y(n_522)
);

OAI221xp5_ASAP7_75t_L g523 ( 
.A1(n_457),
.A2(n_443),
.B1(n_438),
.B2(n_478),
.C(n_456),
.Y(n_523)
);

BUFx8_ASAP7_75t_L g524 ( 
.A(n_443),
.Y(n_524)
);

AOI211xp5_ASAP7_75t_L g525 ( 
.A1(n_438),
.A2(n_478),
.B(n_473),
.C(n_456),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_473),
.B(n_483),
.Y(n_526)
);

AO31x2_ASAP7_75t_L g527 ( 
.A1(n_475),
.A2(n_404),
.A3(n_470),
.B(n_452),
.Y(n_527)
);

AOI221xp5_ASAP7_75t_L g528 ( 
.A1(n_483),
.A2(n_349),
.B1(n_302),
.B2(n_277),
.C(n_394),
.Y(n_528)
);

OAI22xp5_ASAP7_75t_L g529 ( 
.A1(n_484),
.A2(n_488),
.B1(n_486),
.B2(n_370),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_484),
.Y(n_530)
);

INVx1_ASAP7_75t_L g531 ( 
.A(n_499),
.Y(n_531)
);

INVx4_ASAP7_75t_L g532 ( 
.A(n_445),
.Y(n_532)
);

NAND2xp5_ASAP7_75t_L g533 ( 
.A(n_483),
.B(n_484),
.Y(n_533)
);

A2O1A1Ixp33_ASAP7_75t_L g534 ( 
.A1(n_483),
.A2(n_486),
.B(n_488),
.C(n_484),
.Y(n_534)
);

OAI22xp5_ASAP7_75t_L g535 ( 
.A1(n_484),
.A2(n_488),
.B1(n_486),
.B2(n_370),
.Y(n_535)
);

INVx2_ASAP7_75t_L g536 ( 
.A(n_461),
.Y(n_536)
);

AOI21xp5_ASAP7_75t_L g537 ( 
.A1(n_480),
.A2(n_370),
.B(n_487),
.Y(n_537)
);

INVx1_ASAP7_75t_L g538 ( 
.A(n_516),
.Y(n_538)
);

AND2x2_ASAP7_75t_L g539 ( 
.A(n_519),
.B(n_520),
.Y(n_539)
);

INVx2_ASAP7_75t_L g540 ( 
.A(n_512),
.Y(n_540)
);

BUFx2_ASAP7_75t_L g541 ( 
.A(n_524),
.Y(n_541)
);

OR2x2_ASAP7_75t_SL g542 ( 
.A(n_524),
.B(n_530),
.Y(n_542)
);

OAI21xp5_ASAP7_75t_L g543 ( 
.A1(n_534),
.A2(n_535),
.B(n_529),
.Y(n_543)
);

INVx1_ASAP7_75t_L g544 ( 
.A(n_525),
.Y(n_544)
);

INVx4_ASAP7_75t_L g545 ( 
.A(n_502),
.Y(n_545)
);

OR2x2_ASAP7_75t_L g546 ( 
.A(n_526),
.B(n_504),
.Y(n_546)
);

INVx1_ASAP7_75t_L g547 ( 
.A(n_523),
.Y(n_547)
);

BUFx12f_ASAP7_75t_L g548 ( 
.A(n_532),
.Y(n_548)
);

BUFx3_ASAP7_75t_L g549 ( 
.A(n_524),
.Y(n_549)
);

AO21x2_ASAP7_75t_L g550 ( 
.A1(n_505),
.A2(n_537),
.B(n_522),
.Y(n_550)
);

NOR2xp33_ASAP7_75t_L g551 ( 
.A(n_533),
.B(n_507),
.Y(n_551)
);

AND2x2_ASAP7_75t_L g552 ( 
.A(n_534),
.B(n_507),
.Y(n_552)
);

BUFx2_ASAP7_75t_L g553 ( 
.A(n_521),
.Y(n_553)
);

OAI21xp5_ASAP7_75t_L g554 ( 
.A1(n_514),
.A2(n_521),
.B(n_528),
.Y(n_554)
);

AO21x2_ASAP7_75t_L g555 ( 
.A1(n_509),
.A2(n_515),
.B(n_521),
.Y(n_555)
);

OAI211xp5_ASAP7_75t_L g556 ( 
.A1(n_514),
.A2(n_518),
.B(n_510),
.C(n_503),
.Y(n_556)
);

AND2x2_ASAP7_75t_L g557 ( 
.A(n_527),
.B(n_518),
.Y(n_557)
);

AO21x2_ASAP7_75t_L g558 ( 
.A1(n_515),
.A2(n_536),
.B(n_500),
.Y(n_558)
);

OAI21xp5_ASAP7_75t_L g559 ( 
.A1(n_508),
.A2(n_531),
.B(n_511),
.Y(n_559)
);

INVxp67_ASAP7_75t_L g560 ( 
.A(n_559),
.Y(n_560)
);

AND2x2_ASAP7_75t_L g561 ( 
.A(n_557),
.B(n_527),
.Y(n_561)
);

AND2x2_ASAP7_75t_L g562 ( 
.A(n_557),
.B(n_513),
.Y(n_562)
);

BUFx3_ASAP7_75t_L g563 ( 
.A(n_542),
.Y(n_563)
);

INVxp67_ASAP7_75t_L g564 ( 
.A(n_559),
.Y(n_564)
);

INVx3_ASAP7_75t_L g565 ( 
.A(n_550),
.Y(n_565)
);

AOI22xp5_ASAP7_75t_L g566 ( 
.A1(n_539),
.A2(n_551),
.B1(n_552),
.B2(n_556),
.Y(n_566)
);

BUFx3_ASAP7_75t_L g567 ( 
.A(n_542),
.Y(n_567)
);

BUFx3_ASAP7_75t_L g568 ( 
.A(n_542),
.Y(n_568)
);

INVx3_ASAP7_75t_L g569 ( 
.A(n_550),
.Y(n_569)
);

AOI22xp33_ASAP7_75t_L g570 ( 
.A1(n_539),
.A2(n_506),
.B1(n_517),
.B2(n_501),
.Y(n_570)
);

AND2x2_ASAP7_75t_L g571 ( 
.A(n_553),
.B(n_501),
.Y(n_571)
);

OR2x2_ASAP7_75t_L g572 ( 
.A(n_546),
.B(n_506),
.Y(n_572)
);

AND2x4_ASAP7_75t_L g573 ( 
.A(n_563),
.B(n_549),
.Y(n_573)
);

OR2x2_ASAP7_75t_L g574 ( 
.A(n_561),
.B(n_546),
.Y(n_574)
);

BUFx2_ASAP7_75t_L g575 ( 
.A(n_571),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g576 ( 
.A(n_566),
.B(n_551),
.Y(n_576)
);

NAND2x1p5_ASAP7_75t_L g577 ( 
.A(n_572),
.B(n_545),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_572),
.Y(n_578)
);

AND2x2_ASAP7_75t_L g579 ( 
.A(n_561),
.B(n_553),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_566),
.B(n_552),
.Y(n_580)
);

NAND2xp5_ASAP7_75t_L g581 ( 
.A(n_560),
.B(n_543),
.Y(n_581)
);

NAND2x1_ASAP7_75t_SL g582 ( 
.A(n_571),
.B(n_539),
.Y(n_582)
);

NAND2xp5_ASAP7_75t_L g583 ( 
.A(n_560),
.B(n_543),
.Y(n_583)
);

NAND2xp5_ASAP7_75t_L g584 ( 
.A(n_564),
.B(n_546),
.Y(n_584)
);

INVx1_ASAP7_75t_L g585 ( 
.A(n_578),
.Y(n_585)
);

INVx1_ASAP7_75t_L g586 ( 
.A(n_574),
.Y(n_586)
);

NAND2xp5_ASAP7_75t_L g587 ( 
.A(n_581),
.B(n_564),
.Y(n_587)
);

NAND2xp33_ASAP7_75t_R g588 ( 
.A(n_573),
.B(n_541),
.Y(n_588)
);

INVx1_ASAP7_75t_L g589 ( 
.A(n_574),
.Y(n_589)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_584),
.Y(n_590)
);

INVx2_ASAP7_75t_SL g591 ( 
.A(n_582),
.Y(n_591)
);

AOI22xp5_ASAP7_75t_L g592 ( 
.A1(n_576),
.A2(n_556),
.B1(n_554),
.B2(n_570),
.Y(n_592)
);

NAND2xp5_ASAP7_75t_L g593 ( 
.A(n_583),
.B(n_572),
.Y(n_593)
);

AND2x2_ASAP7_75t_L g594 ( 
.A(n_575),
.B(n_571),
.Y(n_594)
);

NAND2xp5_ASAP7_75t_L g595 ( 
.A(n_590),
.B(n_580),
.Y(n_595)
);

INVx2_ASAP7_75t_L g596 ( 
.A(n_585),
.Y(n_596)
);

INVx2_ASAP7_75t_L g597 ( 
.A(n_586),
.Y(n_597)
);

NAND2xp5_ASAP7_75t_L g598 ( 
.A(n_587),
.B(n_579),
.Y(n_598)
);

NOR2xp67_ASAP7_75t_SL g599 ( 
.A(n_591),
.B(n_548),
.Y(n_599)
);

NAND2xp5_ASAP7_75t_L g600 ( 
.A(n_593),
.B(n_579),
.Y(n_600)
);

INVxp67_ASAP7_75t_L g601 ( 
.A(n_589),
.Y(n_601)
);

AND2x2_ASAP7_75t_L g602 ( 
.A(n_594),
.B(n_573),
.Y(n_602)
);

AND2x2_ASAP7_75t_L g603 ( 
.A(n_591),
.B(n_573),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_596),
.Y(n_604)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_598),
.B(n_592),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_598),
.B(n_600),
.Y(n_606)
);

INVx1_ASAP7_75t_L g607 ( 
.A(n_597),
.Y(n_607)
);

OAI22xp5_ASAP7_75t_L g608 ( 
.A1(n_601),
.A2(n_570),
.B1(n_567),
.B2(n_568),
.Y(n_608)
);

O2A1O1Ixp33_ASAP7_75t_L g609 ( 
.A1(n_605),
.A2(n_608),
.B(n_554),
.C(n_595),
.Y(n_609)
);

OAI21xp33_ASAP7_75t_L g610 ( 
.A1(n_606),
.A2(n_595),
.B(n_602),
.Y(n_610)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_604),
.Y(n_611)
);

AOI221xp5_ASAP7_75t_L g612 ( 
.A1(n_609),
.A2(n_607),
.B1(n_562),
.B2(n_547),
.C(n_544),
.Y(n_612)
);

OAI211xp5_ASAP7_75t_L g613 ( 
.A1(n_610),
.A2(n_565),
.B(n_569),
.C(n_541),
.Y(n_613)
);

OAI221xp5_ASAP7_75t_L g614 ( 
.A1(n_612),
.A2(n_611),
.B1(n_588),
.B2(n_599),
.C(n_547),
.Y(n_614)
);

NAND3xp33_ASAP7_75t_SL g615 ( 
.A(n_613),
.B(n_603),
.C(n_577),
.Y(n_615)
);

OAI211xp5_ASAP7_75t_L g616 ( 
.A1(n_615),
.A2(n_565),
.B(n_532),
.C(n_569),
.Y(n_616)
);

INVx2_ASAP7_75t_L g617 ( 
.A(n_614),
.Y(n_617)
);

INVx2_ASAP7_75t_L g618 ( 
.A(n_617),
.Y(n_618)
);

NOR4xp25_ASAP7_75t_L g619 ( 
.A(n_616),
.B(n_565),
.C(n_569),
.D(n_547),
.Y(n_619)
);

INVx1_ASAP7_75t_L g620 ( 
.A(n_618),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_R g621 ( 
.A(n_619),
.B(n_548),
.Y(n_621)
);

NOR2x1_ASAP7_75t_L g622 ( 
.A(n_620),
.B(n_548),
.Y(n_622)
);

AOI222xp33_ASAP7_75t_SL g623 ( 
.A1(n_622),
.A2(n_621),
.B1(n_565),
.B2(n_569),
.C1(n_541),
.C2(n_540),
.Y(n_623)
);

OAI22xp5_ASAP7_75t_L g624 ( 
.A1(n_623),
.A2(n_548),
.B1(n_565),
.B2(n_569),
.Y(n_624)
);

AO21x2_ASAP7_75t_L g625 ( 
.A1(n_624),
.A2(n_550),
.B(n_544),
.Y(n_625)
);

AOI22xp33_ASAP7_75t_L g626 ( 
.A1(n_625),
.A2(n_558),
.B1(n_555),
.B2(n_538),
.Y(n_626)
);


endmodule