module real_jpeg_26028_n_16 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_349, n_6, n_7, n_3, n_10, n_9, n_16);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_349;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_16;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_332;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_216;
wire n_202;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_345;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_337;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_335;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_334;
wire n_17;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_341;
wire n_331;
wire n_49;
wire n_68;
wire n_146;
wire n_286;
wire n_215;
wire n_166;
wire n_176;
wire n_323;
wire n_312;
wire n_325;
wire n_316;
wire n_307;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_342;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_336;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_343;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_324;
wire n_86;
wire n_261;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

AOI22xp33_ASAP7_75t_SL g117 ( 
.A1(n_2),
.A2(n_25),
.B1(n_28),
.B2(n_118),
.Y(n_117)
);

CKINVDCx20_ASAP7_75t_R g118 ( 
.A(n_2),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_L g137 ( 
.A1(n_2),
.A2(n_58),
.B1(n_70),
.B2(n_118),
.Y(n_137)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_2),
.A2(n_31),
.B1(n_32),
.B2(n_118),
.Y(n_177)
);

AOI22xp33_ASAP7_75t_L g216 ( 
.A1(n_2),
.A2(n_47),
.B1(n_48),
.B2(n_118),
.Y(n_216)
);

BUFx12f_ASAP7_75t_L g48 ( 
.A(n_3),
.Y(n_48)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_4),
.A2(n_70),
.B(n_125),
.Y(n_124)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_4),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_4),
.B(n_61),
.Y(n_158)
);

OAI22xp33_ASAP7_75t_L g197 ( 
.A1(n_4),
.A2(n_31),
.B1(n_32),
.B2(n_127),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_4),
.B(n_43),
.C(n_48),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_4),
.B(n_29),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_4),
.A2(n_99),
.B1(n_225),
.B2(n_230),
.Y(n_229)
);

INVx8_ASAP7_75t_SL g62 ( 
.A(n_5),
.Y(n_62)
);

AOI22xp33_ASAP7_75t_SL g119 ( 
.A1(n_6),
.A2(n_25),
.B1(n_28),
.B2(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_6),
.Y(n_120)
);

OAI22xp5_ASAP7_75t_L g179 ( 
.A1(n_6),
.A2(n_31),
.B1(n_32),
.B2(n_120),
.Y(n_179)
);

AOI22xp33_ASAP7_75t_L g208 ( 
.A1(n_6),
.A2(n_47),
.B1(n_48),
.B2(n_120),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_L g265 ( 
.A1(n_6),
.A2(n_54),
.B1(n_69),
.B2(n_120),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_SL g129 ( 
.A1(n_7),
.A2(n_58),
.B1(n_65),
.B2(n_130),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g130 ( 
.A(n_7),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_7),
.A2(n_25),
.B1(n_28),
.B2(n_130),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_7),
.A2(n_31),
.B1(n_32),
.B2(n_130),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_SL g225 ( 
.A1(n_7),
.A2(n_47),
.B1(n_48),
.B2(n_130),
.Y(n_225)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_8),
.A2(n_56),
.B1(n_68),
.B2(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_8),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_8),
.A2(n_47),
.B1(n_48),
.B2(n_68),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_8),
.A2(n_31),
.B1(n_32),
.B2(n_68),
.Y(n_259)
);

AOI22xp33_ASAP7_75t_SL g304 ( 
.A1(n_8),
.A2(n_25),
.B1(n_28),
.B2(n_68),
.Y(n_304)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_9),
.A2(n_54),
.B1(n_57),
.B2(n_58),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_9),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g94 ( 
.A1(n_9),
.A2(n_31),
.B1(n_32),
.B2(n_57),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_SL g146 ( 
.A1(n_9),
.A2(n_47),
.B1(n_48),
.B2(n_57),
.Y(n_146)
);

AOI22xp33_ASAP7_75t_SL g290 ( 
.A1(n_9),
.A2(n_25),
.B1(n_28),
.B2(n_57),
.Y(n_290)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_11),
.A2(n_25),
.B1(n_28),
.B2(n_38),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

AOI22xp33_ASAP7_75t_L g76 ( 
.A1(n_11),
.A2(n_38),
.B1(n_56),
.B2(n_58),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_11),
.A2(n_31),
.B1(n_32),
.B2(n_38),
.Y(n_97)
);

OAI22xp5_ASAP7_75t_L g106 ( 
.A1(n_11),
.A2(n_38),
.B1(n_47),
.B2(n_48),
.Y(n_106)
);

INVx13_ASAP7_75t_L g56 ( 
.A(n_12),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g32 ( 
.A(n_13),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_14),
.A2(n_25),
.B1(n_27),
.B2(n_28),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_14),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_14),
.A2(n_27),
.B1(n_31),
.B2(n_32),
.Y(n_50)
);

AOI22xp33_ASAP7_75t_L g82 ( 
.A1(n_14),
.A2(n_27),
.B1(n_58),
.B2(n_70),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_14),
.A2(n_27),
.B1(n_47),
.B2(n_48),
.Y(n_174)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_15),
.Y(n_102)
);

INVx6_ASAP7_75t_L g110 ( 
.A(n_15),
.Y(n_110)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_15),
.Y(n_211)
);

INVx3_ASAP7_75t_L g230 ( 
.A(n_15),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_84),
.Y(n_16)
);

NAND2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_83),
.Y(n_17)
);

OR2x2_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_77),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_19),
.B(n_77),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_72),
.C(n_73),
.Y(n_19)
);

XNOR2xp5_ASAP7_75t_L g343 ( 
.A(n_20),
.B(n_344),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_39),
.C(n_51),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g333 ( 
.A1(n_21),
.A2(n_22),
.B1(n_39),
.B2(n_328),
.Y(n_333)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_22),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_34),
.Y(n_22)
);

OAI21xp33_ASAP7_75t_L g139 ( 
.A1(n_23),
.A2(n_116),
.B(n_119),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g23 ( 
.A(n_24),
.B(n_29),
.Y(n_23)
);

OAI21xp5_ASAP7_75t_L g72 ( 
.A1(n_24),
.A2(n_29),
.B(n_35),
.Y(n_72)
);

INVxp67_ASAP7_75t_L g268 ( 
.A(n_24),
.Y(n_268)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_25),
.Y(n_28)
);

AOI22xp33_ASAP7_75t_L g36 ( 
.A1(n_25),
.A2(n_28),
.B1(n_30),
.B2(n_33),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_25),
.A2(n_28),
.B1(n_62),
.B2(n_63),
.Y(n_61)
);

A2O1A1Ixp33_ASAP7_75t_L g141 ( 
.A1(n_25),
.A2(n_63),
.B(n_126),
.C(n_142),
.Y(n_141)
);

HAxp5_ASAP7_75t_SL g170 ( 
.A(n_25),
.B(n_127),
.CON(n_170),
.SN(n_170)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND3xp33_ASAP7_75t_L g142 ( 
.A(n_28),
.B(n_55),
.C(n_62),
.Y(n_142)
);

OAI32xp33_ASAP7_75t_L g169 ( 
.A1(n_28),
.A2(n_30),
.A3(n_32),
.B1(n_170),
.B2(n_171),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_29),
.B(n_36),
.Y(n_35)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_29),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_29),
.A2(n_35),
.B1(n_161),
.B2(n_170),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g269 ( 
.A(n_29),
.B(n_37),
.Y(n_269)
);

AO22x1_ASAP7_75t_L g29 ( 
.A1(n_30),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_29)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_30),
.Y(n_33)
);

OAI22xp33_ASAP7_75t_L g42 ( 
.A1(n_31),
.A2(n_32),
.B1(n_43),
.B2(n_45),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_31),
.B(n_33),
.Y(n_171)
);

INVx2_ASAP7_75t_SL g31 ( 
.A(n_32),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_SL g199 ( 
.A(n_32),
.B(n_200),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g289 ( 
.A1(n_34),
.A2(n_121),
.B(n_290),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g34 ( 
.A(n_35),
.B(n_37),
.Y(n_34)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_35),
.Y(n_116)
);

AOI21xp5_ASAP7_75t_L g325 ( 
.A1(n_35),
.A2(n_326),
.B(n_327),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g323 ( 
.A1(n_39),
.A2(n_324),
.B1(n_325),
.B2(n_328),
.Y(n_323)
);

CKINVDCx20_ASAP7_75t_R g328 ( 
.A(n_39),
.Y(n_328)
);

AOI21xp5_ASAP7_75t_L g39 ( 
.A1(n_40),
.A2(n_46),
.B(n_49),
.Y(n_39)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_41),
.B(n_96),
.Y(n_95)
);

AOI21xp5_ASAP7_75t_L g113 ( 
.A1(n_41),
.A2(n_50),
.B(n_114),
.Y(n_113)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_41),
.A2(n_177),
.B1(n_178),
.B2(n_179),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g189 ( 
.A1(n_41),
.A2(n_179),
.B(n_190),
.Y(n_189)
);

AOI22xp5_ASAP7_75t_L g196 ( 
.A1(n_41),
.A2(n_178),
.B1(n_197),
.B2(n_198),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_41),
.A2(n_177),
.B1(n_178),
.B2(n_198),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_41),
.A2(n_178),
.B1(n_258),
.B2(n_259),
.Y(n_257)
);

AOI21xp5_ASAP7_75t_L g280 ( 
.A1(n_41),
.A2(n_114),
.B(n_259),
.Y(n_280)
);

AND2x2_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_46),
.Y(n_41)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_43),
.A2(n_45),
.B1(n_47),
.B2(n_48),
.Y(n_46)
);

BUFx24_ASAP7_75t_L g43 ( 
.A(n_44),
.Y(n_43)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_46),
.A2(n_94),
.B(n_95),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_46),
.B(n_97),
.Y(n_114)
);

INVx1_ASAP7_75t_L g178 ( 
.A(n_46),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g190 ( 
.A(n_46),
.B(n_49),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_SL g223 ( 
.A(n_46),
.B(n_127),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g100 ( 
.A(n_47),
.B(n_101),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_SL g231 ( 
.A(n_47),
.B(n_232),
.Y(n_231)
);

INVx6_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

XNOR2xp5_ASAP7_75t_SL g332 ( 
.A(n_51),
.B(n_333),
.Y(n_332)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_59),
.B1(n_61),
.B2(n_67),
.Y(n_51)
);

CKINVDCx20_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_53),
.A2(n_60),
.B(n_78),
.Y(n_321)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_55),
.B(n_127),
.Y(n_126)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx11_ASAP7_75t_L g58 ( 
.A(n_56),
.Y(n_58)
);

INVx8_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

INVx6_ASAP7_75t_L g71 ( 
.A(n_56),
.Y(n_71)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g74 ( 
.A1(n_59),
.A2(n_67),
.B(n_75),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_59),
.B(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_59),
.Y(n_123)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_59),
.A2(n_61),
.B1(n_129),
.B2(n_137),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_59),
.A2(n_61),
.B1(n_137),
.B2(n_265),
.Y(n_264)
);

AOI21xp5_ASAP7_75t_L g287 ( 
.A1(n_59),
.A2(n_81),
.B(n_265),
.Y(n_287)
);

AOI21xp5_ASAP7_75t_L g308 ( 
.A1(n_59),
.A2(n_75),
.B(n_309),
.Y(n_308)
);

AND2x2_ASAP7_75t_SL g59 ( 
.A(n_60),
.B(n_64),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_60),
.B(n_76),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_60),
.B(n_82),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_SL g122 ( 
.A1(n_60),
.A2(n_123),
.B1(n_124),
.B2(n_128),
.Y(n_122)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_62),
.A2(n_63),
.B1(n_65),
.B2(n_66),
.Y(n_64)
);

INVx8_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

INVx8_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_72),
.A2(n_73),
.B1(n_74),
.B2(n_345),
.Y(n_344)
);

CKINVDCx20_ASAP7_75t_R g345 ( 
.A(n_72),
.Y(n_345)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_74),
.Y(n_73)
);

INVxp67_ASAP7_75t_L g79 ( 
.A(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

CKINVDCx14_ASAP7_75t_R g80 ( 
.A(n_81),
.Y(n_80)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_82),
.Y(n_309)
);

AOI21xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_341),
.B(n_346),
.Y(n_84)
);

OAI321xp33_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_317),
.A3(n_336),
.B1(n_339),
.B2(n_340),
.C(n_349),
.Y(n_85)
);

AOI21xp5_ASAP7_75t_L g86 ( 
.A1(n_87),
.A2(n_295),
.B(n_316),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g87 ( 
.A1(n_88),
.A2(n_274),
.B(n_294),
.Y(n_87)
);

O2A1O1Ixp33_ASAP7_75t_SL g88 ( 
.A1(n_89),
.A2(n_162),
.B(n_249),
.C(n_273),
.Y(n_88)
);

AND2x2_ASAP7_75t_L g89 ( 
.A(n_90),
.B(n_147),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_90),
.B(n_147),
.Y(n_163)
);

XNOR2xp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_133),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g91 ( 
.A1(n_92),
.A2(n_111),
.B1(n_131),
.B2(n_132),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g131 ( 
.A(n_92),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_92),
.B(n_132),
.C(n_133),
.Y(n_250)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_98),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_93),
.B(n_98),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_94),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_95),
.B(n_302),
.Y(n_301)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_L g98 ( 
.A1(n_99),
.A2(n_103),
.B(n_105),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g172 ( 
.A1(n_99),
.A2(n_105),
.B(n_173),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_L g207 ( 
.A1(n_99),
.A2(n_208),
.B(n_209),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_99),
.A2(n_216),
.B1(n_225),
.B2(n_226),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g282 ( 
.A1(n_99),
.A2(n_173),
.B(n_226),
.Y(n_282)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_100),
.A2(n_104),
.B1(n_109),
.B2(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_100),
.B(n_106),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_100),
.A2(n_215),
.B1(n_217),
.B2(n_218),
.Y(n_214)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_101),
.Y(n_155)
);

INVx5_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_102),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_104),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_106),
.B(n_107),
.Y(n_105)
);

INVx3_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

INVx5_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_110),
.Y(n_109)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_110),
.Y(n_234)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_111),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g111 ( 
.A(n_112),
.B(n_115),
.C(n_122),
.Y(n_111)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_112),
.A2(n_113),
.B1(n_115),
.B2(n_150),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_115),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_121),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g159 ( 
.A1(n_116),
.A2(n_117),
.B1(n_121),
.B2(n_160),
.Y(n_159)
);

OAI21xp5_ASAP7_75t_L g267 ( 
.A1(n_116),
.A2(n_268),
.B(n_269),
.Y(n_267)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_116),
.A2(n_121),
.B1(n_290),
.B2(n_304),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_SL g148 ( 
.A(n_122),
.B(n_149),
.Y(n_148)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_127),
.B(n_233),
.Y(n_232)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g133 ( 
.A(n_134),
.B(n_140),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_135),
.A2(n_136),
.B1(n_138),
.B2(n_139),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_136),
.B(n_138),
.C(n_140),
.Y(n_271)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_141),
.B(n_143),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_141),
.A2(n_143),
.B1(n_144),
.B2(n_152),
.Y(n_151)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_141),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_144),
.Y(n_143)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g154 ( 
.A1(n_146),
.A2(n_155),
.B(n_156),
.Y(n_154)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_151),
.C(n_153),
.Y(n_147)
);

XNOR2xp5_ASAP7_75t_L g246 ( 
.A(n_148),
.B(n_247),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_151),
.B(n_153),
.Y(n_247)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_159),
.Y(n_153)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_154),
.A2(n_157),
.B1(n_158),
.B2(n_184),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_154),
.Y(n_184)
);

AND2x2_ASAP7_75t_L g256 ( 
.A(n_156),
.B(n_209),
.Y(n_256)
);

CKINVDCx16_ASAP7_75t_R g157 ( 
.A(n_158),
.Y(n_157)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_183),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g160 ( 
.A(n_161),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_163),
.B(n_164),
.Y(n_162)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_165),
.A2(n_244),
.B(n_248),
.Y(n_164)
);

OAI21xp5_ASAP7_75t_L g165 ( 
.A1(n_166),
.A2(n_192),
.B(n_243),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_167),
.B(n_180),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g243 ( 
.A(n_167),
.B(n_180),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_175),
.C(n_176),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g240 ( 
.A(n_168),
.B(n_241),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_SL g168 ( 
.A(n_169),
.B(n_172),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_169),
.B(n_172),
.Y(n_187)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_210),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g241 ( 
.A(n_175),
.B(n_176),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g180 ( 
.A1(n_181),
.A2(n_182),
.B1(n_185),
.B2(n_186),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g245 ( 
.A(n_181),
.B(n_188),
.C(n_191),
.Y(n_245)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_186),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g186 ( 
.A1(n_187),
.A2(n_188),
.B1(n_189),
.B2(n_191),
.Y(n_186)
);

CKINVDCx16_ASAP7_75t_R g191 ( 
.A(n_187),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g188 ( 
.A(n_189),
.Y(n_188)
);

INVxp67_ASAP7_75t_L g302 ( 
.A(n_190),
.Y(n_302)
);

AOI21xp5_ASAP7_75t_L g192 ( 
.A1(n_193),
.A2(n_238),
.B(n_242),
.Y(n_192)
);

OAI21xp5_ASAP7_75t_SL g193 ( 
.A1(n_194),
.A2(n_212),
.B(n_237),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g194 ( 
.A(n_195),
.B(n_201),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_195),
.B(n_201),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g195 ( 
.A(n_196),
.B(n_199),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g220 ( 
.A(n_196),
.B(n_199),
.Y(n_220)
);

XNOR2xp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_207),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g202 ( 
.A1(n_203),
.A2(n_204),
.B1(n_205),
.B2(n_206),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_203),
.B(n_206),
.C(n_207),
.Y(n_239)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_204),
.Y(n_203)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_205),
.Y(n_206)
);

INVxp67_ASAP7_75t_L g217 ( 
.A(n_208),
.Y(n_217)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

BUFx2_ASAP7_75t_L g219 ( 
.A(n_211),
.Y(n_219)
);

AOI21xp33_ASAP7_75t_L g212 ( 
.A1(n_213),
.A2(n_221),
.B(n_236),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g213 ( 
.A(n_214),
.B(n_220),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g236 ( 
.A(n_214),
.B(n_220),
.Y(n_236)
);

CKINVDCx14_ASAP7_75t_R g215 ( 
.A(n_216),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g218 ( 
.A(n_219),
.Y(n_218)
);

OAI21xp5_ASAP7_75t_SL g221 ( 
.A1(n_222),
.A2(n_228),
.B(n_235),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g235 ( 
.A(n_223),
.B(n_224),
.Y(n_235)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

INVx2_ASAP7_75t_L g233 ( 
.A(n_234),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_239),
.B(n_240),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g242 ( 
.A(n_239),
.B(n_240),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_245),
.B(n_246),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_SL g248 ( 
.A(n_245),
.B(n_246),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_251),
.Y(n_249)
);

NOR2xp33_ASAP7_75t_L g273 ( 
.A(n_250),
.B(n_251),
.Y(n_273)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_252),
.A2(n_253),
.B1(n_271),
.B2(n_272),
.Y(n_251)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_253),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g253 ( 
.A(n_254),
.B(n_261),
.Y(n_253)
);

MAJIxp5_ASAP7_75t_L g275 ( 
.A(n_254),
.B(n_261),
.C(n_272),
.Y(n_275)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_255),
.A2(n_256),
.B1(n_257),
.B2(n_260),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_L g284 ( 
.A(n_255),
.B(n_260),
.Y(n_284)
);

CKINVDCx20_ASAP7_75t_R g255 ( 
.A(n_256),
.Y(n_255)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_257),
.Y(n_260)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_262),
.B(n_270),
.Y(n_261)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_263),
.A2(n_264),
.B1(n_266),
.B2(n_267),
.Y(n_262)
);

CKINVDCx14_ASAP7_75t_R g263 ( 
.A(n_264),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_264),
.B(n_266),
.C(n_270),
.Y(n_293)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_267),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g327 ( 
.A(n_269),
.Y(n_327)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_271),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_276),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g294 ( 
.A(n_275),
.B(n_276),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_293),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g277 ( 
.A1(n_278),
.A2(n_283),
.B1(n_291),
.B2(n_292),
.Y(n_277)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_278),
.Y(n_291)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_278),
.B(n_292),
.C(n_293),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_279),
.A2(n_280),
.B1(n_281),
.B2(n_282),
.Y(n_278)
);

CKINVDCx20_ASAP7_75t_R g279 ( 
.A(n_280),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_280),
.B(n_281),
.Y(n_311)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_281),
.A2(n_282),
.B1(n_308),
.B2(n_310),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_L g329 ( 
.A1(n_281),
.A2(n_310),
.B(n_311),
.Y(n_329)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_282),
.Y(n_281)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_283),
.Y(n_292)
);

XNOR2xp5_ASAP7_75t_SL g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g314 ( 
.A(n_284),
.B(n_287),
.C(n_288),
.Y(n_314)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_286),
.A2(n_287),
.B1(n_288),
.B2(n_289),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_287),
.Y(n_286)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_289),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_297),
.Y(n_295)
);

NOR2xp33_ASAP7_75t_SL g316 ( 
.A(n_296),
.B(n_297),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_298),
.A2(n_299),
.B1(n_314),
.B2(n_315),
.Y(n_297)
);

INVx1_ASAP7_75t_L g298 ( 
.A(n_299),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g299 ( 
.A1(n_300),
.A2(n_306),
.B1(n_312),
.B2(n_313),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_300),
.Y(n_312)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_300),
.B(n_313),
.C(n_315),
.Y(n_337)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_301),
.A2(n_303),
.B(n_305),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_301),
.B(n_303),
.Y(n_305)
);

INVxp67_ASAP7_75t_L g326 ( 
.A(n_304),
.Y(n_326)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_305),
.B(n_319),
.C(n_329),
.Y(n_318)
);

FAx1_ASAP7_75t_SL g338 ( 
.A(n_305),
.B(n_319),
.CI(n_329),
.CON(n_338),
.SN(n_338)
);

INVx1_ASAP7_75t_L g313 ( 
.A(n_306),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_SL g306 ( 
.A(n_307),
.B(n_311),
.Y(n_306)
);

CKINVDCx16_ASAP7_75t_R g310 ( 
.A(n_308),
.Y(n_310)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_314),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g317 ( 
.A(n_318),
.B(n_330),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g340 ( 
.A(n_318),
.B(n_330),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_320),
.A2(n_321),
.B1(n_322),
.B2(n_323),
.Y(n_319)
);

AOI22xp5_ASAP7_75t_L g331 ( 
.A1(n_320),
.A2(n_321),
.B1(n_332),
.B2(n_334),
.Y(n_331)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_321),
.B(n_325),
.C(n_328),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_334),
.C(n_335),
.Y(n_342)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_323),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g324 ( 
.A(n_325),
.Y(n_324)
);

XNOR2xp5_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_335),
.Y(n_330)
);

INVx1_ASAP7_75t_L g334 ( 
.A(n_332),
.Y(n_334)
);

NOR2xp33_ASAP7_75t_L g336 ( 
.A(n_337),
.B(n_338),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_SL g339 ( 
.A(n_337),
.B(n_338),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g347 ( 
.A(n_338),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_SL g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g346 ( 
.A(n_342),
.B(n_343),
.Y(n_346)
);


endmodule