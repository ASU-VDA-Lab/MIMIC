module fake_netlist_1_12409_n_29 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_29);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_29;
wire n_20;
wire n_23;
wire n_28;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_27;
INVx2_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
NOR2xp33_ASAP7_75t_L g13 ( .A(n_9), .B(n_6), .Y(n_13) );
AND2x2_ASAP7_75t_L g14 ( .A(n_0), .B(n_3), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_11), .Y(n_15) );
INVx1_ASAP7_75t_L g16 ( .A(n_2), .Y(n_16) );
CKINVDCx20_ASAP7_75t_R g17 ( .A(n_8), .Y(n_17) );
INVx2_ASAP7_75t_L g18 ( .A(n_12), .Y(n_18) );
NAND2xp5_ASAP7_75t_L g19 ( .A(n_15), .B(n_0), .Y(n_19) );
INVx2_ASAP7_75t_SL g20 ( .A(n_18), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_17), .B1(n_16), .B2(n_14), .Y(n_21) );
OAI211xp5_ASAP7_75t_L g22 ( .A1(n_21), .A2(n_13), .B(n_1), .C(n_4), .Y(n_22) );
INVx1_ASAP7_75t_L g23 ( .A(n_22), .Y(n_23) );
NAND2xp5_ASAP7_75t_L g24 ( .A(n_23), .B(n_20), .Y(n_24) );
XNOR2x1_ASAP7_75t_L g25 ( .A(n_24), .B(n_1), .Y(n_25) );
NOR2x1_ASAP7_75t_L g26 ( .A(n_24), .B(n_13), .Y(n_26) );
INVx1_ASAP7_75t_SL g27 ( .A(n_25), .Y(n_27) );
BUFx2_ASAP7_75t_L g28 ( .A(n_27), .Y(n_28) );
OAI22xp5_ASAP7_75t_L g29 ( .A1(n_28), .A2(n_26), .B1(n_5), .B2(n_7), .Y(n_29) );
endmodule