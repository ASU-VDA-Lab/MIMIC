module fake_jpeg_12672_n_104 (n_3, n_2, n_1, n_0, n_4, n_8, n_9, n_6, n_5, n_7, n_104);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_104;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_42;
wire n_49;
wire n_16;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_30;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_11;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_7),
.Y(n_10)
);

INVx3_ASAP7_75t_L g11 ( 
.A(n_7),
.Y(n_11)
);

INVx1_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

BUFx10_ASAP7_75t_L g13 ( 
.A(n_2),
.Y(n_13)
);

INVx3_ASAP7_75t_L g14 ( 
.A(n_8),
.Y(n_14)
);

BUFx8_ASAP7_75t_L g15 ( 
.A(n_1),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_2),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

BUFx6f_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_3),
.Y(n_19)
);

INVx6_ASAP7_75t_L g20 ( 
.A(n_18),
.Y(n_20)
);

INVx6_ASAP7_75t_L g32 ( 
.A(n_20),
.Y(n_32)
);

INVx4_ASAP7_75t_L g21 ( 
.A(n_13),
.Y(n_21)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_21),
.Y(n_34)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_15),
.Y(n_22)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_22),
.Y(n_31)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g27 ( 
.A(n_23),
.B(n_26),
.Y(n_27)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx6p67_ASAP7_75t_R g29 ( 
.A(n_24),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_13),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_25),
.B(n_13),
.Y(n_33)
);

INVx3_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

INVx8_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_23),
.B(n_10),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_30),
.B(n_36),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_19),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_L g35 ( 
.A1(n_20),
.A2(n_25),
.B1(n_13),
.B2(n_11),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_35),
.A2(n_26),
.B1(n_24),
.B2(n_21),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g36 ( 
.A(n_22),
.B(n_10),
.Y(n_36)
);

BUFx12f_ASAP7_75t_L g37 ( 
.A(n_29),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_37),
.B(n_41),
.Y(n_46)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_40),
.A2(n_29),
.B1(n_31),
.B2(n_28),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_30),
.Y(n_41)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_27),
.B(n_24),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_42),
.B(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_27),
.B(n_19),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_43),
.B(n_44),
.Y(n_47)
);

AND2x6_ASAP7_75t_L g45 ( 
.A(n_29),
.B(n_9),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_45),
.B(n_8),
.Y(n_52)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_39),
.Y(n_48)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_48),
.Y(n_59)
);

OAI21xp33_ASAP7_75t_L g57 ( 
.A1(n_49),
.A2(n_37),
.B(n_29),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_35),
.Y(n_50)
);

XNOR2xp5_ASAP7_75t_L g55 ( 
.A(n_50),
.B(n_40),
.Y(n_55)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_51),
.B(n_52),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g58 ( 
.A1(n_53),
.A2(n_28),
.B1(n_32),
.B2(n_34),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_14),
.Y(n_54)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_37),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_55),
.B(n_60),
.C(n_18),
.Y(n_72)
);

OAI21x1_ASAP7_75t_L g56 ( 
.A1(n_47),
.A2(n_42),
.B(n_45),
.Y(n_56)
);

NOR3xp33_ASAP7_75t_L g66 ( 
.A(n_56),
.B(n_57),
.C(n_61),
.Y(n_66)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_34),
.C(n_14),
.Y(n_60)
);

OAI21xp5_ASAP7_75t_L g61 ( 
.A1(n_46),
.A2(n_16),
.B(n_12),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_50),
.A2(n_32),
.B1(n_16),
.B2(n_11),
.Y(n_63)
);

AOI22xp5_ASAP7_75t_L g68 ( 
.A1(n_63),
.A2(n_53),
.B1(n_32),
.B2(n_14),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_64),
.B(n_48),
.Y(n_67)
);

CKINVDCx14_ASAP7_75t_R g77 ( 
.A(n_67),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_68),
.B(n_70),
.Y(n_76)
);

BUFx3_ASAP7_75t_L g69 ( 
.A(n_58),
.Y(n_69)
);

INVx1_ASAP7_75t_SL g81 ( 
.A(n_69),
.Y(n_81)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_59),
.Y(n_70)
);

MAJIxp5_ASAP7_75t_L g71 ( 
.A(n_60),
.B(n_11),
.C(n_18),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g75 ( 
.A(n_71),
.B(n_61),
.C(n_15),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_72),
.B(n_55),
.Y(n_74)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_59),
.Y(n_73)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_73),
.Y(n_80)
);

NAND3xp33_ASAP7_75t_L g86 ( 
.A(n_74),
.B(n_66),
.C(n_5),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g84 ( 
.A(n_75),
.B(n_15),
.Y(n_84)
);

INVxp33_ASAP7_75t_L g78 ( 
.A(n_69),
.Y(n_78)
);

OAI21xp5_ASAP7_75t_L g82 ( 
.A1(n_78),
.A2(n_79),
.B(n_81),
.Y(n_82)
);

OAI21xp5_ASAP7_75t_L g79 ( 
.A1(n_72),
.A2(n_62),
.B(n_17),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g93 ( 
.A(n_82),
.B(n_86),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_80),
.B(n_66),
.C(n_65),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g91 ( 
.A(n_83),
.B(n_84),
.C(n_88),
.Y(n_91)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_76),
.Y(n_85)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_85),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g87 ( 
.A1(n_77),
.A2(n_17),
.B1(n_1),
.B2(n_2),
.Y(n_87)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_87),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_17),
.C(n_4),
.Y(n_88)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_90),
.B(n_78),
.Y(n_94)
);

OAI221xp5_ASAP7_75t_L g99 ( 
.A1(n_94),
.A2(n_95),
.B1(n_96),
.B2(n_97),
.C(n_6),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_89),
.B(n_4),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_93),
.B(n_9),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_91),
.B(n_92),
.Y(n_97)
);

NOR2xp67_ASAP7_75t_L g98 ( 
.A(n_94),
.B(n_91),
.Y(n_98)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_98),
.A2(n_100),
.B(n_0),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g102 ( 
.A(n_99),
.B(n_3),
.Y(n_102)
);

NOR2x1_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_0),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_101),
.Y(n_103)
);

XOR2xp5_ASAP7_75t_L g104 ( 
.A(n_103),
.B(n_102),
.Y(n_104)
);


endmodule