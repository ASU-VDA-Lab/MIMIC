module fake_jpeg_27488_n_59 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_59);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_59;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_45;
wire n_23;
wire n_27;
wire n_55;
wire n_22;
wire n_47;
wire n_51;
wire n_40;
wire n_35;
wire n_48;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_38;
wire n_44;
wire n_26;
wire n_36;
wire n_31;
wire n_25;
wire n_56;
wire n_29;
wire n_43;
wire n_37;
wire n_50;
wire n_32;

AND2x2_ASAP7_75t_L g22 ( 
.A(n_5),
.B(n_1),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_2),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_14),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_20),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_4),
.B(n_12),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_11),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g28 ( 
.A(n_1),
.B(n_5),
.Y(n_28)
);

CKINVDCx16_ASAP7_75t_R g29 ( 
.A(n_22),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_29),
.B(n_30),
.Y(n_37)
);

INVx4_ASAP7_75t_SL g30 ( 
.A(n_23),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_24),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_31),
.B(n_32),
.Y(n_36)
);

INVx2_ASAP7_75t_R g32 ( 
.A(n_23),
.Y(n_32)
);

OR2x2_ASAP7_75t_L g33 ( 
.A(n_22),
.B(n_0),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_33),
.B(n_34),
.Y(n_39)
);

NAND2xp5_ASAP7_75t_L g34 ( 
.A(n_22),
.B(n_0),
.Y(n_34)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_2),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_28),
.Y(n_41)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_38),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_34),
.A2(n_27),
.B1(n_25),
.B2(n_24),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_40),
.A2(n_44),
.B1(n_6),
.B2(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_41),
.B(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_35),
.Y(n_42)
);

OAI21xp5_ASAP7_75t_SL g43 ( 
.A1(n_33),
.A2(n_25),
.B(n_26),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g48 ( 
.A(n_43),
.B(n_3),
.C(n_6),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g44 ( 
.A1(n_30),
.A2(n_27),
.B1(n_13),
.B2(n_15),
.Y(n_44)
);

XNOR2xp5_ASAP7_75t_L g46 ( 
.A(n_39),
.B(n_10),
.Y(n_46)
);

MAJIxp5_ASAP7_75t_L g54 ( 
.A(n_46),
.B(n_47),
.C(n_48),
.Y(n_54)
);

OAI21xp5_ASAP7_75t_SL g47 ( 
.A1(n_37),
.A2(n_3),
.B(n_4),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_16),
.C(n_19),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_49),
.B(n_50),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_45),
.A2(n_36),
.B(n_38),
.C(n_44),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g55 ( 
.A(n_52),
.B(n_51),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g57 ( 
.A(n_55),
.B(n_56),
.Y(n_57)
);

MAJIxp5_ASAP7_75t_L g56 ( 
.A(n_53),
.B(n_51),
.C(n_43),
.Y(n_56)
);

AOI322xp5_ASAP7_75t_L g58 ( 
.A1(n_57),
.A2(n_54),
.A3(n_9),
.B1(n_17),
.B2(n_18),
.C1(n_21),
.C2(n_8),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_L g59 ( 
.A1(n_58),
.A2(n_7),
.B(n_8),
.Y(n_59)
);


endmodule