module real_aes_1814_n_99 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_753, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_43, n_96, n_54, n_35, n_42, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_754, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_99);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_753;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_754;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_99;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_100;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_744;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_656;
wire n_532;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_455;
wire n_310;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_449;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_434;
wire n_527;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_501;
wire n_488;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_430;
wire n_269;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_358;
wire n_275;
wire n_214;
wire n_385;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_720;
wire n_265;
wire n_354;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_101;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_633;
wire n_520;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_420;
wire n_336;
wire n_349;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_717;
wire n_456;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_524;
wire n_219;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_103;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_674;
wire n_644;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND2xp5_ASAP7_75t_L g162 ( .A(n_0), .B(n_136), .Y(n_162) );
NAND2xp5_ASAP7_75t_L g106 ( .A(n_1), .B(n_107), .Y(n_106) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_2), .B(n_120), .Y(n_526) );
NAND2xp5_ASAP7_75t_L g453 ( .A(n_3), .B(n_138), .Y(n_453) );
INVx1_ASAP7_75t_L g127 ( .A(n_4), .Y(n_127) );
NAND2xp5_ASAP7_75t_L g189 ( .A(n_5), .B(n_120), .Y(n_189) );
NAND2xp33_ASAP7_75t_SL g232 ( .A(n_6), .B(n_126), .Y(n_232) );
INVx1_ASAP7_75t_L g224 ( .A(n_7), .Y(n_224) );
CKINVDCx16_ASAP7_75t_R g107 ( .A(n_8), .Y(n_107) );
AND2x2_ASAP7_75t_L g187 ( .A(n_9), .B(n_144), .Y(n_187) );
AND2x2_ASAP7_75t_L g455 ( .A(n_10), .B(n_140), .Y(n_455) );
AND2x2_ASAP7_75t_L g465 ( .A(n_11), .B(n_230), .Y(n_465) );
INVx2_ASAP7_75t_L g142 ( .A(n_12), .Y(n_142) );
NAND2xp5_ASAP7_75t_L g505 ( .A(n_13), .B(n_138), .Y(n_505) );
CKINVDCx16_ASAP7_75t_R g108 ( .A(n_14), .Y(n_108) );
AOI221x1_ASAP7_75t_L g227 ( .A1(n_15), .A2(n_129), .B1(n_228), .B2(n_230), .C(n_231), .Y(n_227) );
NAND2xp5_ASAP7_75t_SL g119 ( .A(n_16), .B(n_120), .Y(n_119) );
NAND2xp5_ASAP7_75t_SL g510 ( .A(n_17), .B(n_120), .Y(n_510) );
INVx1_ASAP7_75t_L g104 ( .A(n_18), .Y(n_104) );
AOI22xp33_ASAP7_75t_L g469 ( .A1(n_19), .A2(n_88), .B1(n_120), .B2(n_173), .Y(n_469) );
AOI221xp5_ASAP7_75t_SL g151 ( .A1(n_20), .A2(n_37), .B1(n_120), .B2(n_129), .C(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g190 ( .A1(n_21), .A2(n_129), .B(n_191), .Y(n_190) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_22), .B(n_136), .Y(n_192) );
OA21x2_ASAP7_75t_L g141 ( .A1(n_23), .A2(n_87), .B(n_142), .Y(n_141) );
OR2x2_ASAP7_75t_L g145 ( .A(n_23), .B(n_87), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_24), .B(n_138), .Y(n_137) );
INVxp67_ASAP7_75t_L g226 ( .A(n_25), .Y(n_226) );
AND2x2_ASAP7_75t_L g213 ( .A(n_26), .B(n_150), .Y(n_213) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_27), .Y(n_750) );
AOI21xp5_ASAP7_75t_L g160 ( .A1(n_28), .A2(n_129), .B(n_161), .Y(n_160) );
AO21x2_ASAP7_75t_L g500 ( .A1(n_29), .A2(n_230), .B(n_501), .Y(n_500) );
CKINVDCx20_ASAP7_75t_R g727 ( .A(n_30), .Y(n_727) );
NAND2xp5_ASAP7_75t_L g153 ( .A(n_31), .B(n_138), .Y(n_153) );
OAI22xp5_ASAP7_75t_L g743 ( .A1(n_32), .A2(n_744), .B1(n_745), .B2(n_746), .Y(n_743) );
CKINVDCx20_ASAP7_75t_R g744 ( .A(n_32), .Y(n_744) );
AOI21xp5_ASAP7_75t_L g450 ( .A1(n_33), .A2(n_129), .B(n_451), .Y(n_450) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_34), .B(n_138), .Y(n_525) );
AND2x2_ASAP7_75t_L g126 ( .A(n_35), .B(n_127), .Y(n_126) );
AND2x2_ASAP7_75t_L g130 ( .A(n_35), .B(n_131), .Y(n_130) );
INVx1_ASAP7_75t_L g181 ( .A(n_35), .Y(n_181) );
NOR3xp33_ASAP7_75t_L g105 ( .A(n_36), .B(n_106), .C(n_108), .Y(n_105) );
OR2x6_ASAP7_75t_L g427 ( .A(n_36), .B(n_428), .Y(n_427) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_38), .B(n_120), .Y(n_454) );
AOI22xp5_ASAP7_75t_L g178 ( .A1(n_39), .A2(n_79), .B1(n_129), .B2(n_179), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g497 ( .A(n_40), .B(n_138), .Y(n_497) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_41), .B(n_120), .Y(n_441) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_42), .B(n_136), .Y(n_211) );
AOI21xp5_ASAP7_75t_L g460 ( .A1(n_43), .A2(n_129), .B(n_461), .Y(n_460) );
AND2x2_ASAP7_75t_L g165 ( .A(n_44), .B(n_150), .Y(n_165) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_45), .B(n_136), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g155 ( .A(n_46), .B(n_150), .Y(n_155) );
NAND2xp5_ASAP7_75t_SL g502 ( .A(n_47), .B(n_120), .Y(n_502) );
INVx1_ASAP7_75t_L g123 ( .A(n_48), .Y(n_123) );
INVx1_ASAP7_75t_L g133 ( .A(n_48), .Y(n_133) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_49), .B(n_138), .Y(n_463) );
AND2x2_ASAP7_75t_L g492 ( .A(n_50), .B(n_150), .Y(n_492) );
NAND2xp5_ASAP7_75t_SL g212 ( .A(n_51), .B(n_120), .Y(n_212) );
NAND2xp5_ASAP7_75t_L g462 ( .A(n_52), .B(n_136), .Y(n_462) );
NAND2xp5_ASAP7_75t_L g524 ( .A(n_53), .B(n_136), .Y(n_524) );
AND2x2_ASAP7_75t_L g204 ( .A(n_54), .B(n_150), .Y(n_204) );
NAND2xp5_ASAP7_75t_SL g464 ( .A(n_55), .B(n_120), .Y(n_464) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_56), .B(n_138), .Y(n_163) );
NAND2xp5_ASAP7_75t_SL g494 ( .A(n_57), .B(n_120), .Y(n_494) );
AOI21xp5_ASAP7_75t_L g522 ( .A1(n_58), .A2(n_129), .B(n_523), .Y(n_522) );
AND2x2_ASAP7_75t_SL g143 ( .A(n_59), .B(n_144), .Y(n_143) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_60), .B(n_136), .Y(n_201) );
AND2x2_ASAP7_75t_L g516 ( .A(n_61), .B(n_144), .Y(n_516) );
AOI21xp5_ASAP7_75t_L g208 ( .A1(n_62), .A2(n_129), .B(n_209), .Y(n_208) );
NAND2xp5_ASAP7_75t_L g193 ( .A(n_63), .B(n_138), .Y(n_193) );
AND2x2_ASAP7_75t_SL g184 ( .A(n_64), .B(n_140), .Y(n_184) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_65), .B(n_136), .Y(n_498) );
NAND2xp5_ASAP7_75t_L g506 ( .A(n_66), .B(n_136), .Y(n_506) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_67), .A2(n_90), .B1(n_129), .B2(n_179), .Y(n_470) );
NAND2xp5_ASAP7_75t_L g513 ( .A(n_68), .B(n_138), .Y(n_513) );
INVx1_ASAP7_75t_L g125 ( .A(n_69), .Y(n_125) );
INVx1_ASAP7_75t_L g131 ( .A(n_69), .Y(n_131) );
NAND2xp5_ASAP7_75t_L g452 ( .A(n_70), .B(n_136), .Y(n_452) );
OAI222xp33_ASAP7_75t_L g110 ( .A1(n_71), .A2(n_111), .B1(n_717), .B2(n_718), .C1(n_724), .C2(n_727), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g717 ( .A(n_71), .Y(n_717) );
AOI21xp5_ASAP7_75t_L g495 ( .A1(n_72), .A2(n_129), .B(n_496), .Y(n_495) );
AOI21xp5_ASAP7_75t_L g442 ( .A1(n_73), .A2(n_129), .B(n_443), .Y(n_442) );
AOI21xp5_ASAP7_75t_L g503 ( .A1(n_74), .A2(n_129), .B(n_504), .Y(n_503) );
AND2x2_ASAP7_75t_L g527 ( .A(n_75), .B(n_144), .Y(n_527) );
NAND2xp5_ASAP7_75t_SL g467 ( .A(n_76), .B(n_150), .Y(n_467) );
AOI22xp5_ASAP7_75t_L g172 ( .A1(n_77), .A2(n_81), .B1(n_120), .B2(n_173), .Y(n_172) );
NAND2xp5_ASAP7_75t_SL g202 ( .A(n_78), .B(n_120), .Y(n_202) );
NOR2xp33_ASAP7_75t_L g103 ( .A(n_80), .B(n_104), .Y(n_103) );
INVx1_ASAP7_75t_L g429 ( .A(n_80), .Y(n_429) );
NAND2xp5_ASAP7_75t_L g135 ( .A(n_82), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_83), .B(n_136), .Y(n_154) );
AND2x2_ASAP7_75t_L g446 ( .A(n_84), .B(n_140), .Y(n_446) );
CKINVDCx20_ASAP7_75t_R g738 ( .A(n_85), .Y(n_738) );
AOI21xp5_ASAP7_75t_L g198 ( .A1(n_86), .A2(n_129), .B(n_199), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g200 ( .A(n_89), .B(n_138), .Y(n_200) );
AOI21xp5_ASAP7_75t_L g511 ( .A1(n_91), .A2(n_129), .B(n_512), .Y(n_511) );
NAND2xp5_ASAP7_75t_L g444 ( .A(n_92), .B(n_138), .Y(n_444) );
NAND2xp5_ASAP7_75t_L g164 ( .A(n_93), .B(n_120), .Y(n_164) );
INVxp67_ASAP7_75t_L g229 ( .A(n_94), .Y(n_229) );
NAND2xp5_ASAP7_75t_L g210 ( .A(n_95), .B(n_138), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g128 ( .A1(n_96), .A2(n_129), .B(n_134), .Y(n_128) );
BUFx2_ASAP7_75t_L g515 ( .A(n_97), .Y(n_515) );
BUFx2_ASAP7_75t_L g732 ( .A(n_98), .Y(n_732) );
BUFx2_ASAP7_75t_SL g741 ( .A(n_98), .Y(n_741) );
AOI21xp33_ASAP7_75t_SL g99 ( .A1(n_100), .A2(n_109), .B(n_749), .Y(n_99) );
INVx2_ASAP7_75t_L g100 ( .A(n_101), .Y(n_100) );
INVx1_ASAP7_75t_SL g751 ( .A(n_101), .Y(n_751) );
INVx3_ASAP7_75t_SL g101 ( .A(n_102), .Y(n_101) );
AND2x2_ASAP7_75t_SL g102 ( .A(n_103), .B(n_105), .Y(n_102) );
NAND2xp5_ASAP7_75t_L g428 ( .A(n_104), .B(n_429), .Y(n_428) );
AND2x6_ASAP7_75t_SL g426 ( .A(n_108), .B(n_427), .Y(n_426) );
OR2x6_ASAP7_75t_SL g715 ( .A(n_108), .B(n_716), .Y(n_715) );
OR2x2_ASAP7_75t_L g726 ( .A(n_108), .B(n_427), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_108), .B(n_716), .Y(n_737) );
OA21x2_ASAP7_75t_L g109 ( .A1(n_110), .A2(n_728), .B(n_739), .Y(n_109) );
AOI22xp5_ASAP7_75t_SL g111 ( .A1(n_112), .A2(n_426), .B1(n_430), .B2(n_714), .Y(n_111) );
OAI22xp5_ASAP7_75t_L g719 ( .A1(n_112), .A2(n_430), .B1(n_720), .B2(n_723), .Y(n_719) );
INVx3_ASAP7_75t_SL g745 ( .A(n_112), .Y(n_745) );
HB1xp67_ASAP7_75t_L g746 ( .A(n_112), .Y(n_746) );
AND2x4_ASAP7_75t_L g112 ( .A(n_113), .B(n_318), .Y(n_112) );
NOR3xp33_ASAP7_75t_L g113 ( .A(n_114), .B(n_246), .C(n_296), .Y(n_113) );
OAI211xp5_ASAP7_75t_SL g114 ( .A1(n_115), .A2(n_166), .B(n_214), .C(n_235), .Y(n_114) );
OR2x2_ASAP7_75t_L g115 ( .A(n_116), .B(n_146), .Y(n_115) );
AND2x2_ASAP7_75t_L g245 ( .A(n_116), .B(n_147), .Y(n_245) );
INVx1_ASAP7_75t_L g376 ( .A(n_116), .Y(n_376) );
NOR2x1p5_ASAP7_75t_L g408 ( .A(n_116), .B(n_409), .Y(n_408) );
INVx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AND2x2_ASAP7_75t_L g219 ( .A(n_117), .B(n_220), .Y(n_219) );
INVx2_ASAP7_75t_L g267 ( .A(n_117), .Y(n_267) );
OR2x2_ASAP7_75t_L g271 ( .A(n_117), .B(n_272), .Y(n_271) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_117), .B(n_149), .Y(n_283) );
OR2x2_ASAP7_75t_L g305 ( .A(n_117), .B(n_149), .Y(n_305) );
AND2x4_ASAP7_75t_L g311 ( .A(n_117), .B(n_275), .Y(n_311) );
OR2x2_ASAP7_75t_L g328 ( .A(n_117), .B(n_221), .Y(n_328) );
INVx1_ASAP7_75t_L g363 ( .A(n_117), .Y(n_363) );
HB1xp67_ASAP7_75t_L g385 ( .A(n_117), .Y(n_385) );
OR2x2_ASAP7_75t_L g399 ( .A(n_117), .B(n_332), .Y(n_399) );
AND2x4_ASAP7_75t_SL g403 ( .A(n_117), .B(n_221), .Y(n_403) );
OR2x6_ASAP7_75t_L g117 ( .A(n_118), .B(n_143), .Y(n_117) );
AOI21xp5_ASAP7_75t_L g118 ( .A1(n_119), .A2(n_128), .B(n_140), .Y(n_118) );
AND2x4_ASAP7_75t_L g120 ( .A(n_121), .B(n_126), .Y(n_120) );
INVx1_ASAP7_75t_L g233 ( .A(n_121), .Y(n_233) );
AND2x4_ASAP7_75t_L g121 ( .A(n_122), .B(n_124), .Y(n_121) );
AND2x6_ASAP7_75t_L g136 ( .A(n_122), .B(n_131), .Y(n_136) );
INVx2_ASAP7_75t_L g122 ( .A(n_123), .Y(n_122) );
AND2x4_ASAP7_75t_L g138 ( .A(n_124), .B(n_133), .Y(n_138) );
INVx2_ASAP7_75t_L g124 ( .A(n_125), .Y(n_124) );
INVx5_ASAP7_75t_L g139 ( .A(n_126), .Y(n_139) );
AND2x2_ASAP7_75t_L g132 ( .A(n_127), .B(n_133), .Y(n_132) );
HB1xp67_ASAP7_75t_L g176 ( .A(n_127), .Y(n_176) );
AND2x6_ASAP7_75t_L g129 ( .A(n_130), .B(n_132), .Y(n_129) );
BUFx3_ASAP7_75t_L g177 ( .A(n_130), .Y(n_177) );
INVx2_ASAP7_75t_L g183 ( .A(n_131), .Y(n_183) );
AND2x4_ASAP7_75t_L g179 ( .A(n_132), .B(n_180), .Y(n_179) );
INVx2_ASAP7_75t_L g175 ( .A(n_133), .Y(n_175) );
AOI21xp5_ASAP7_75t_L g134 ( .A1(n_135), .A2(n_137), .B(n_139), .Y(n_134) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_136), .B(n_515), .Y(n_514) );
AOI21xp5_ASAP7_75t_L g152 ( .A1(n_139), .A2(n_153), .B(n_154), .Y(n_152) );
AOI21xp5_ASAP7_75t_L g161 ( .A1(n_139), .A2(n_162), .B(n_163), .Y(n_161) );
AOI21xp5_ASAP7_75t_L g191 ( .A1(n_139), .A2(n_192), .B(n_193), .Y(n_191) );
AOI21xp5_ASAP7_75t_L g199 ( .A1(n_139), .A2(n_200), .B(n_201), .Y(n_199) );
AOI21xp5_ASAP7_75t_L g209 ( .A1(n_139), .A2(n_210), .B(n_211), .Y(n_209) );
AOI21xp5_ASAP7_75t_L g443 ( .A1(n_139), .A2(n_444), .B(n_445), .Y(n_443) );
AOI21xp5_ASAP7_75t_L g451 ( .A1(n_139), .A2(n_452), .B(n_453), .Y(n_451) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_139), .A2(n_462), .B(n_463), .Y(n_461) );
AOI21xp5_ASAP7_75t_L g496 ( .A1(n_139), .A2(n_497), .B(n_498), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g504 ( .A1(n_139), .A2(n_505), .B(n_506), .Y(n_504) );
AOI21xp5_ASAP7_75t_L g512 ( .A1(n_139), .A2(n_513), .B(n_514), .Y(n_512) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_139), .A2(n_524), .B(n_525), .Y(n_523) );
INVx2_ASAP7_75t_SL g170 ( .A(n_140), .Y(n_170) );
AOI21xp5_ASAP7_75t_L g509 ( .A1(n_140), .A2(n_510), .B(n_511), .Y(n_509) );
BUFx4f_ASAP7_75t_L g140 ( .A(n_141), .Y(n_140) );
INVx3_ASAP7_75t_L g158 ( .A(n_141), .Y(n_158) );
AND2x2_ASAP7_75t_SL g144 ( .A(n_142), .B(n_145), .Y(n_144) );
AND2x4_ASAP7_75t_L g194 ( .A(n_142), .B(n_145), .Y(n_194) );
BUFx6f_ASAP7_75t_L g150 ( .A(n_144), .Y(n_150) );
INVx1_ASAP7_75t_L g146 ( .A(n_147), .Y(n_146) );
AND2x2_ASAP7_75t_L g355 ( .A(n_147), .B(n_311), .Y(n_355) );
AND2x2_ASAP7_75t_L g402 ( .A(n_147), .B(n_403), .Y(n_402) );
AND2x2_ASAP7_75t_L g147 ( .A(n_148), .B(n_156), .Y(n_147) );
INVx2_ASAP7_75t_L g148 ( .A(n_149), .Y(n_148) );
INVx1_ASAP7_75t_L g218 ( .A(n_149), .Y(n_218) );
AND2x2_ASAP7_75t_L g265 ( .A(n_149), .B(n_156), .Y(n_265) );
INVx2_ASAP7_75t_L g272 ( .A(n_149), .Y(n_272) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_149), .Y(n_393) );
BUFx3_ASAP7_75t_L g409 ( .A(n_149), .Y(n_409) );
OA21x2_ASAP7_75t_L g149 ( .A1(n_150), .A2(n_151), .B(n_155), .Y(n_149) );
CKINVDCx5p33_ASAP7_75t_R g203 ( .A(n_150), .Y(n_203) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_150), .A2(n_441), .B(n_442), .Y(n_440) );
AO21x2_ASAP7_75t_L g468 ( .A1(n_150), .A2(n_469), .B(n_470), .Y(n_468) );
INVx2_ASAP7_75t_L g234 ( .A(n_156), .Y(n_234) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_156), .B(n_275), .Y(n_274) );
OR2x2_ASAP7_75t_L g332 ( .A(n_156), .B(n_272), .Y(n_332) );
INVx1_ASAP7_75t_L g350 ( .A(n_156), .Y(n_350) );
HB1xp67_ASAP7_75t_L g366 ( .A(n_156), .Y(n_366) );
INVx1_ASAP7_75t_L g388 ( .A(n_156), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_156), .B(n_267), .Y(n_415) );
NAND2xp5_ASAP7_75t_L g425 ( .A(n_156), .B(n_221), .Y(n_425) );
INVx3_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AOI21x1_ASAP7_75t_L g157 ( .A1(n_158), .A2(n_159), .B(n_165), .Y(n_157) );
INVx4_ASAP7_75t_L g230 ( .A(n_158), .Y(n_230) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_158), .A2(n_459), .B(n_465), .Y(n_458) );
NAND2xp5_ASAP7_75t_L g159 ( .A(n_160), .B(n_164), .Y(n_159) );
INVx1_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_185), .Y(n_167) );
AND2x4_ASAP7_75t_L g239 ( .A(n_168), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g250 ( .A(n_168), .Y(n_250) );
AND2x2_ASAP7_75t_L g255 ( .A(n_168), .B(n_256), .Y(n_255) );
AND2x2_ASAP7_75t_L g290 ( .A(n_168), .B(n_195), .Y(n_290) );
AND2x2_ASAP7_75t_L g300 ( .A(n_168), .B(n_196), .Y(n_300) );
OR2x2_ASAP7_75t_L g380 ( .A(n_168), .B(n_295), .Y(n_380) );
OAI322xp33_ASAP7_75t_L g410 ( .A1(n_168), .A2(n_323), .A3(n_362), .B1(n_395), .B2(n_411), .C1(n_412), .C2(n_413), .Y(n_410) );
OR2x2_ASAP7_75t_L g411 ( .A(n_168), .B(n_393), .Y(n_411) );
BUFx6f_ASAP7_75t_L g168 ( .A(n_169), .Y(n_168) );
INVx2_ASAP7_75t_L g244 ( .A(n_169), .Y(n_244) );
AOI21x1_ASAP7_75t_L g169 ( .A1(n_170), .A2(n_171), .B(n_184), .Y(n_169) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_178), .Y(n_171) );
AOI22xp5_ASAP7_75t_L g222 ( .A1(n_173), .A2(n_179), .B1(n_223), .B2(n_225), .Y(n_222) );
AND2x4_ASAP7_75t_L g173 ( .A(n_174), .B(n_177), .Y(n_173) );
AND2x2_ASAP7_75t_L g174 ( .A(n_175), .B(n_176), .Y(n_174) );
NOR2x1p5_ASAP7_75t_L g180 ( .A(n_181), .B(n_182), .Y(n_180) );
INVx3_ASAP7_75t_L g182 ( .A(n_183), .Y(n_182) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_185), .A2(n_357), .B1(n_361), .B2(n_364), .Y(n_356) );
AOI211xp5_ASAP7_75t_L g416 ( .A1(n_185), .A2(n_417), .B(n_418), .C(n_421), .Y(n_416) );
AND2x4_ASAP7_75t_SL g185 ( .A(n_186), .B(n_195), .Y(n_185) );
AND2x4_ASAP7_75t_L g238 ( .A(n_186), .B(n_206), .Y(n_238) );
HB1xp67_ASAP7_75t_L g242 ( .A(n_186), .Y(n_242) );
INVx5_ASAP7_75t_L g254 ( .A(n_186), .Y(n_254) );
INVx2_ASAP7_75t_L g263 ( .A(n_186), .Y(n_263) );
AND2x2_ASAP7_75t_L g286 ( .A(n_186), .B(n_196), .Y(n_286) );
AND2x2_ASAP7_75t_L g315 ( .A(n_186), .B(n_205), .Y(n_315) );
OR2x2_ASAP7_75t_L g324 ( .A(n_186), .B(n_244), .Y(n_324) );
OR2x2_ASAP7_75t_L g339 ( .A(n_186), .B(n_253), .Y(n_339) );
OR2x6_ASAP7_75t_L g186 ( .A(n_187), .B(n_188), .Y(n_186) );
AOI21xp5_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_194), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_194), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g225 ( .A(n_194), .B(n_226), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g228 ( .A(n_194), .B(n_229), .Y(n_228) );
NOR3xp33_ASAP7_75t_L g231 ( .A(n_194), .B(n_232), .C(n_233), .Y(n_231) );
AOI21xp5_ASAP7_75t_L g493 ( .A1(n_194), .A2(n_494), .B(n_495), .Y(n_493) );
AOI21xp5_ASAP7_75t_L g501 ( .A1(n_194), .A2(n_502), .B(n_503), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_195), .B(n_215), .Y(n_214) );
INVx3_ASAP7_75t_SL g323 ( .A(n_195), .Y(n_323) );
AND2x2_ASAP7_75t_L g346 ( .A(n_195), .B(n_254), .Y(n_346) );
AND2x4_ASAP7_75t_L g195 ( .A(n_196), .B(n_205), .Y(n_195) );
INVx2_ASAP7_75t_L g240 ( .A(n_196), .Y(n_240) );
AND2x2_ASAP7_75t_L g243 ( .A(n_196), .B(n_244), .Y(n_243) );
OR2x2_ASAP7_75t_L g257 ( .A(n_196), .B(n_206), .Y(n_257) );
INVx1_ASAP7_75t_L g261 ( .A(n_196), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g295 ( .A(n_196), .B(n_206), .Y(n_295) );
HB1xp67_ASAP7_75t_L g359 ( .A(n_196), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g370 ( .A(n_196), .B(n_254), .Y(n_370) );
AO21x2_ASAP7_75t_L g196 ( .A1(n_197), .A2(n_203), .B(n_204), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g197 ( .A(n_198), .B(n_202), .Y(n_197) );
AO21x2_ASAP7_75t_L g206 ( .A1(n_203), .A2(n_207), .B(n_213), .Y(n_206) );
AO21x2_ASAP7_75t_L g253 ( .A1(n_203), .A2(n_207), .B(n_213), .Y(n_253) );
AOI21x1_ASAP7_75t_L g448 ( .A1(n_203), .A2(n_449), .B(n_455), .Y(n_448) );
INVx2_ASAP7_75t_L g205 ( .A(n_206), .Y(n_205) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_206), .Y(n_276) );
AND2x2_ASAP7_75t_L g360 ( .A(n_206), .B(n_244), .Y(n_360) );
NAND2xp5_ASAP7_75t_L g207 ( .A(n_208), .B(n_212), .Y(n_207) );
AND2x2_ASAP7_75t_L g215 ( .A(n_216), .B(n_219), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g326 ( .A(n_216), .B(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
OR2x6_ASAP7_75t_SL g424 ( .A(n_217), .B(n_425), .Y(n_424) );
INVxp67_ASAP7_75t_SL g217 ( .A(n_218), .Y(n_217) );
HB1xp67_ASAP7_75t_L g310 ( .A(n_218), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g349 ( .A(n_218), .B(n_350), .Y(n_349) );
INVx1_ASAP7_75t_L g372 ( .A(n_218), .Y(n_372) );
AOI22xp5_ASAP7_75t_L g280 ( .A1(n_219), .A2(n_281), .B1(n_284), .B2(n_291), .Y(n_280) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_220), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g316 ( .A(n_220), .B(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g362 ( .A(n_220), .B(n_363), .Y(n_362) );
AND2x2_ASAP7_75t_SL g371 ( .A(n_220), .B(n_372), .Y(n_371) );
AND2x4_ASAP7_75t_L g220 ( .A(n_221), .B(n_234), .Y(n_220) );
AND2x2_ASAP7_75t_L g266 ( .A(n_221), .B(n_267), .Y(n_266) );
INVx3_ASAP7_75t_L g275 ( .A(n_221), .Y(n_275) );
OAI22xp33_ASAP7_75t_L g333 ( .A1(n_221), .A2(n_282), .B1(n_334), .B2(n_336), .Y(n_333) );
INVx1_ASAP7_75t_L g341 ( .A(n_221), .Y(n_341) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_221), .B(n_335), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g396 ( .A(n_221), .B(n_265), .Y(n_396) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_221), .B(n_272), .Y(n_414) );
AND2x4_ASAP7_75t_L g221 ( .A(n_222), .B(n_227), .Y(n_221) );
INVx3_ASAP7_75t_L g520 ( .A(n_230), .Y(n_520) );
OAI21xp33_ASAP7_75t_L g235 ( .A1(n_236), .A2(n_241), .B(n_245), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_237), .B(n_239), .Y(n_236) );
NAND4xp25_ASAP7_75t_SL g284 ( .A(n_237), .B(n_285), .C(n_287), .D(n_289), .Y(n_284) );
INVx2_ASAP7_75t_SL g237 ( .A(n_238), .Y(n_237) );
NAND2xp5_ASAP7_75t_L g374 ( .A(n_238), .B(n_345), .Y(n_374) );
AND2x2_ASAP7_75t_L g401 ( .A(n_238), .B(n_239), .Y(n_401) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_238), .B(n_261), .Y(n_412) );
INVx1_ASAP7_75t_L g277 ( .A(n_239), .Y(n_277) );
AOI22xp5_ASAP7_75t_L g312 ( .A1(n_239), .A2(n_302), .B1(n_313), .B2(n_316), .Y(n_312) );
NAND3xp33_ASAP7_75t_L g334 ( .A(n_239), .B(n_252), .C(n_335), .Y(n_334) );
NAND2xp5_ASAP7_75t_L g353 ( .A(n_239), .B(n_254), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_239), .B(n_262), .Y(n_405) );
AND2x2_ASAP7_75t_L g337 ( .A(n_240), .B(n_244), .Y(n_337) );
HB1xp67_ASAP7_75t_L g398 ( .A(n_240), .Y(n_398) );
AND2x2_ASAP7_75t_L g241 ( .A(n_242), .B(n_243), .Y(n_241) );
INVx1_ASAP7_75t_L g293 ( .A(n_242), .Y(n_293) );
INVx1_ASAP7_75t_L g383 ( .A(n_243), .Y(n_383) );
AND2x2_ASAP7_75t_L g390 ( .A(n_243), .B(n_254), .Y(n_390) );
BUFx2_ASAP7_75t_L g345 ( .A(n_244), .Y(n_345) );
NAND3xp33_ASAP7_75t_SL g246 ( .A(n_247), .B(n_268), .C(n_280), .Y(n_246) );
OAI31xp33_ASAP7_75t_L g247 ( .A1(n_248), .A2(n_255), .A3(n_258), .B(n_264), .Y(n_247) );
AOI22xp5_ASAP7_75t_L g301 ( .A1(n_248), .A2(n_302), .B1(n_306), .B2(n_307), .Y(n_301) );
INVx1_ASAP7_75t_L g248 ( .A(n_249), .Y(n_248) );
OR2x2_ASAP7_75t_L g249 ( .A(n_250), .B(n_251), .Y(n_249) );
OR2x2_ASAP7_75t_L g287 ( .A(n_250), .B(n_288), .Y(n_287) );
NOR2x1_ASAP7_75t_L g313 ( .A(n_250), .B(n_314), .Y(n_313) );
O2A1O1Ixp33_ASAP7_75t_L g382 ( .A1(n_251), .A2(n_353), .B(n_383), .C(n_384), .Y(n_382) );
INVx2_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_252), .B(n_398), .Y(n_397) );
AND2x4_ASAP7_75t_L g252 ( .A(n_253), .B(n_254), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_253), .B(n_261), .Y(n_288) );
AND2x2_ASAP7_75t_L g306 ( .A(n_253), .B(n_286), .Y(n_306) );
AND2x2_ASAP7_75t_L g423 ( .A(n_256), .B(n_345), .Y(n_423) );
INVx2_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g279 ( .A(n_257), .B(n_263), .Y(n_279) );
NOR2xp33_ASAP7_75t_L g258 ( .A(n_259), .B(n_262), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_260), .Y(n_259) );
HB1xp67_ASAP7_75t_L g260 ( .A(n_261), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g299 ( .A(n_262), .B(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g354 ( .A(n_262), .B(n_337), .Y(n_354) );
INVx2_ASAP7_75t_L g262 ( .A(n_263), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g343 ( .A(n_263), .B(n_337), .Y(n_343) );
AND2x2_ASAP7_75t_L g264 ( .A(n_265), .B(n_266), .Y(n_264) );
INVx2_ASAP7_75t_L g335 ( .A(n_265), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_266), .B(n_366), .Y(n_365) );
AOI32xp33_ASAP7_75t_L g268 ( .A1(n_269), .A2(n_276), .A3(n_277), .B1(n_278), .B2(n_753), .Y(n_268) );
AOI221xp5_ASAP7_75t_L g389 ( .A1(n_269), .A2(n_354), .B1(n_390), .B2(n_391), .C(n_394), .Y(n_389) );
AND2x4_ASAP7_75t_L g269 ( .A(n_270), .B(n_273), .Y(n_269) );
INVx2_ASAP7_75t_L g270 ( .A(n_271), .Y(n_270) );
HB1xp67_ASAP7_75t_L g317 ( .A(n_272), .Y(n_317) );
INVx1_ASAP7_75t_L g273 ( .A(n_274), .Y(n_273) );
OR2x2_ASAP7_75t_L g282 ( .A(n_274), .B(n_283), .Y(n_282) );
AND2x2_ASAP7_75t_L g387 ( .A(n_275), .B(n_388), .Y(n_387) );
NAND2xp5_ASAP7_75t_SL g297 ( .A(n_276), .B(n_298), .Y(n_297) );
AOI221xp5_ASAP7_75t_L g320 ( .A1(n_278), .A2(n_321), .B1(n_325), .B2(n_329), .C(n_333), .Y(n_320) );
INVx1_ASAP7_75t_L g278 ( .A(n_279), .Y(n_278) );
INVx2_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OAI211xp5_ASAP7_75t_L g296 ( .A1(n_283), .A2(n_297), .B(n_301), .C(n_312), .Y(n_296) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
OAI322xp33_ASAP7_75t_L g394 ( .A1(n_289), .A2(n_299), .A3(n_348), .B1(n_395), .B2(n_396), .C1(n_397), .C2(n_399), .Y(n_394) );
INVx2_ASAP7_75t_L g289 ( .A(n_290), .Y(n_289) );
INVx2_ASAP7_75t_L g291 ( .A(n_292), .Y(n_291) );
AOI21xp33_ASAP7_75t_L g421 ( .A1(n_292), .A2(n_422), .B(n_424), .Y(n_421) );
NAND2xp5_ASAP7_75t_SL g292 ( .A(n_293), .B(n_294), .Y(n_292) );
INVx1_ASAP7_75t_L g294 ( .A(n_295), .Y(n_294) );
O2A1O1Ixp33_ASAP7_75t_L g378 ( .A1(n_298), .A2(n_379), .B(n_381), .C(n_382), .Y(n_378) );
INVx1_ASAP7_75t_L g298 ( .A(n_299), .Y(n_298) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVx1_ASAP7_75t_SL g304 ( .A(n_305), .Y(n_304) );
OR2x2_ASAP7_75t_L g420 ( .A(n_305), .B(n_386), .Y(n_420) );
INVx1_ASAP7_75t_L g307 ( .A(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g308 ( .A(n_309), .B(n_311), .Y(n_308) );
INVxp67_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_311), .B(n_331), .Y(n_330) );
INVx1_ASAP7_75t_L g395 ( .A(n_311), .Y(n_395) );
INVx2_ASAP7_75t_L g314 ( .A(n_315), .Y(n_314) );
OAI31xp33_ASAP7_75t_L g351 ( .A1(n_315), .A2(n_352), .A3(n_354), .B(n_355), .Y(n_351) );
NOR2x1_ASAP7_75t_L g318 ( .A(n_319), .B(n_377), .Y(n_318) );
NAND5xp2_ASAP7_75t_L g319 ( .A(n_320), .B(n_340), .C(n_351), .D(n_356), .E(n_367), .Y(n_319) );
INVx1_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
OR2x2_ASAP7_75t_L g322 ( .A(n_323), .B(n_324), .Y(n_322) );
AOI21xp33_ASAP7_75t_L g418 ( .A1(n_323), .A2(n_419), .B(n_420), .Y(n_418) );
INVx1_ASAP7_75t_SL g325 ( .A(n_326), .Y(n_325) );
AND2x2_ASAP7_75t_L g391 ( .A(n_327), .B(n_392), .Y(n_391) );
INVx1_ASAP7_75t_SL g327 ( .A(n_328), .Y(n_327) );
INVx1_ASAP7_75t_L g329 ( .A(n_330), .Y(n_329) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
INVx1_ASAP7_75t_SL g338 ( .A(n_339), .Y(n_338) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_342), .B(n_344), .C(n_347), .Y(n_340) );
INVxp33_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g344 ( .A(n_345), .B(n_346), .Y(n_344) );
OR2x2_ASAP7_75t_L g369 ( .A(n_345), .B(n_370), .Y(n_369) );
HB1xp67_ASAP7_75t_L g347 ( .A(n_348), .Y(n_347) );
NAND2xp5_ASAP7_75t_L g375 ( .A(n_348), .B(n_376), .Y(n_375) );
INVx1_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AND2x2_ASAP7_75t_SL g357 ( .A(n_358), .B(n_360), .Y(n_357) );
INVx1_ASAP7_75t_L g358 ( .A(n_359), .Y(n_358) );
INVx1_ASAP7_75t_L g419 ( .A(n_360), .Y(n_419) );
INVx1_ASAP7_75t_SL g361 ( .A(n_362), .Y(n_361) );
INVx1_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
AOI21xp5_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_371), .B(n_373), .Y(n_367) );
INVx1_ASAP7_75t_L g368 ( .A(n_369), .Y(n_368) );
AOI21xp33_ASAP7_75t_L g373 ( .A1(n_369), .A2(n_374), .B(n_375), .Y(n_373) );
NAND4xp25_ASAP7_75t_L g377 ( .A(n_378), .B(n_389), .C(n_400), .D(n_416), .Y(n_377) );
INVx1_ASAP7_75t_SL g379 ( .A(n_380), .Y(n_379) );
OR2x2_ASAP7_75t_L g384 ( .A(n_385), .B(n_386), .Y(n_384) );
INVx1_ASAP7_75t_SL g386 ( .A(n_387), .Y(n_386) );
NAND2xp5_ASAP7_75t_L g407 ( .A(n_387), .B(n_408), .Y(n_407) );
HB1xp67_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
INVx1_ASAP7_75t_L g417 ( .A(n_399), .Y(n_417) );
AOI221xp5_ASAP7_75t_L g400 ( .A1(n_401), .A2(n_402), .B1(n_404), .B2(n_406), .C(n_410), .Y(n_400) );
INVx1_ASAP7_75t_L g404 ( .A(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g406 ( .A(n_407), .Y(n_406) );
OR2x2_ASAP7_75t_L g413 ( .A(n_414), .B(n_415), .Y(n_413) );
INVx2_ASAP7_75t_L g422 ( .A(n_423), .Y(n_422) );
CKINVDCx5p33_ASAP7_75t_R g722 ( .A(n_426), .Y(n_722) );
CKINVDCx5p33_ASAP7_75t_R g716 ( .A(n_427), .Y(n_716) );
AND2x4_ASAP7_75t_L g430 ( .A(n_431), .B(n_627), .Y(n_430) );
NOR4xp75_ASAP7_75t_L g431 ( .A(n_432), .B(n_550), .C(n_575), .D(n_602), .Y(n_431) );
OAI21xp5_ASAP7_75t_L g432 ( .A1(n_433), .A2(n_487), .B(n_528), .Y(n_432) );
NOR4xp25_ASAP7_75t_L g433 ( .A(n_434), .B(n_471), .C(n_478), .D(n_482), .Y(n_433) );
INVx1_ASAP7_75t_SL g434 ( .A(n_435), .Y(n_434) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_436), .B(n_456), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_437), .Y(n_436) );
NAND2xp5_ASAP7_75t_L g437 ( .A(n_438), .B(n_447), .Y(n_437) );
NAND2x1p5_ASAP7_75t_L g590 ( .A(n_438), .B(n_591), .Y(n_590) );
NAND2xp5_ASAP7_75t_L g621 ( .A(n_438), .B(n_475), .Y(n_621) );
AND2x2_ASAP7_75t_L g646 ( .A(n_438), .B(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g671 ( .A(n_438), .B(n_466), .Y(n_671) );
AND2x2_ASAP7_75t_L g712 ( .A(n_438), .B(n_480), .Y(n_712) );
INVx4_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
AND2x4_ASAP7_75t_SL g484 ( .A(n_439), .B(n_477), .Y(n_484) );
AND2x2_ASAP7_75t_L g486 ( .A(n_439), .B(n_458), .Y(n_486) );
NOR2x1_ASAP7_75t_L g536 ( .A(n_439), .B(n_537), .Y(n_536) );
INVx1_ASAP7_75t_L g547 ( .A(n_439), .Y(n_547) );
AND2x2_ASAP7_75t_L g553 ( .A(n_439), .B(n_480), .Y(n_553) );
BUFx2_ASAP7_75t_L g566 ( .A(n_439), .Y(n_566) );
AND2x4_ASAP7_75t_L g597 ( .A(n_439), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g644 ( .A(n_439), .B(n_645), .Y(n_644) );
OR2x6_ASAP7_75t_L g439 ( .A(n_440), .B(n_446), .Y(n_439) );
INVx1_ASAP7_75t_L g638 ( .A(n_447), .Y(n_638) );
HB1xp67_ASAP7_75t_L g447 ( .A(n_448), .Y(n_447) );
INVx3_ASAP7_75t_L g477 ( .A(n_448), .Y(n_477) );
AND2x2_ASAP7_75t_L g480 ( .A(n_448), .B(n_458), .Y(n_480) );
NAND2xp5_ASAP7_75t_L g449 ( .A(n_450), .B(n_454), .Y(n_449) );
NAND2xp5_ASAP7_75t_L g709 ( .A(n_456), .B(n_656), .Y(n_709) );
INVx2_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
OR2x2_ASAP7_75t_L g546 ( .A(n_457), .B(n_547), .Y(n_546) );
OR2x2_ASAP7_75t_L g457 ( .A(n_458), .B(n_466), .Y(n_457) );
INVx2_ASAP7_75t_L g476 ( .A(n_458), .Y(n_476) );
INVx2_ASAP7_75t_L g537 ( .A(n_458), .Y(n_537) );
AND2x2_ASAP7_75t_L g647 ( .A(n_458), .B(n_477), .Y(n_647) );
NAND2xp5_ASAP7_75t_L g459 ( .A(n_460), .B(n_464), .Y(n_459) );
INVx2_ASAP7_75t_L g535 ( .A(n_466), .Y(n_535) );
BUFx3_ASAP7_75t_L g552 ( .A(n_466), .Y(n_552) );
AND2x2_ASAP7_75t_L g579 ( .A(n_466), .B(n_580), .Y(n_579) );
AND2x4_ASAP7_75t_L g466 ( .A(n_467), .B(n_468), .Y(n_466) );
AND2x4_ASAP7_75t_L g473 ( .A(n_467), .B(n_468), .Y(n_473) );
NOR2x1_ASAP7_75t_L g471 ( .A(n_472), .B(n_474), .Y(n_471) );
INVx2_ASAP7_75t_L g481 ( .A(n_472), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g637 ( .A(n_472), .B(n_638), .Y(n_637) );
OR2x2_ASAP7_75t_L g650 ( .A(n_472), .B(n_590), .Y(n_650) );
AND2x2_ASAP7_75t_L g674 ( .A(n_472), .B(n_484), .Y(n_674) );
INVx3_ASAP7_75t_L g472 ( .A(n_473), .Y(n_472) );
AND2x2_ASAP7_75t_L g570 ( .A(n_473), .B(n_476), .Y(n_570) );
AND2x2_ASAP7_75t_L g652 ( .A(n_473), .B(n_645), .Y(n_652) );
INVx1_ASAP7_75t_L g474 ( .A(n_475), .Y(n_474) );
INVx1_ASAP7_75t_SL g695 ( .A(n_475), .Y(n_695) );
AND2x2_ASAP7_75t_L g475 ( .A(n_476), .B(n_477), .Y(n_475) );
INVx1_ASAP7_75t_L g580 ( .A(n_476), .Y(n_580) );
HB1xp67_ASAP7_75t_L g584 ( .A(n_477), .Y(n_584) );
INVx2_ASAP7_75t_L g592 ( .A(n_477), .Y(n_592) );
INVx1_ASAP7_75t_L g598 ( .A(n_477), .Y(n_598) );
AOI222xp33_ASAP7_75t_SL g528 ( .A1(n_478), .A2(n_529), .B1(n_533), .B2(n_538), .C1(n_545), .C2(n_548), .Y(n_528) );
INVx1_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
INVx1_ASAP7_75t_L g605 ( .A(n_480), .Y(n_605) );
BUFx2_ASAP7_75t_L g634 ( .A(n_480), .Y(n_634) );
OAI211xp5_ASAP7_75t_L g628 ( .A1(n_481), .A2(n_629), .B(n_633), .C(n_641), .Y(n_628) );
OR2x2_ASAP7_75t_L g699 ( .A(n_481), .B(n_700), .Y(n_699) );
AND2x2_ASAP7_75t_L g707 ( .A(n_481), .B(n_612), .Y(n_707) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_485), .Y(n_482) );
INVx2_ASAP7_75t_SL g483 ( .A(n_484), .Y(n_483) );
AND2x2_ASAP7_75t_SL g664 ( .A(n_484), .B(n_665), .Y(n_664) );
AND2x2_ASAP7_75t_L g682 ( .A(n_484), .B(n_570), .Y(n_682) );
NAND2xp5_ASAP7_75t_L g689 ( .A(n_484), .B(n_662), .Y(n_689) );
OR2x2_ASAP7_75t_L g690 ( .A(n_485), .B(n_552), .Y(n_690) );
INVx1_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
AND2x2_ASAP7_75t_L g612 ( .A(n_486), .B(n_584), .Y(n_612) );
INVx1_ASAP7_75t_L g487 ( .A(n_488), .Y(n_487) );
AND2x2_ASAP7_75t_L g488 ( .A(n_489), .B(n_507), .Y(n_488) );
INVx1_ASAP7_75t_L g706 ( .A(n_489), .Y(n_706) );
NOR2xp67_ASAP7_75t_L g489 ( .A(n_490), .B(n_499), .Y(n_489) );
AND2x2_ASAP7_75t_L g549 ( .A(n_490), .B(n_508), .Y(n_549) );
INVx1_ASAP7_75t_L g626 ( .A(n_490), .Y(n_626) );
OR2x2_ASAP7_75t_L g685 ( .A(n_490), .B(n_508), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_490), .B(n_557), .Y(n_691) );
INVx4_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
INVx2_ASAP7_75t_L g532 ( .A(n_491), .Y(n_532) );
OR2x2_ASAP7_75t_L g564 ( .A(n_491), .B(n_518), .Y(n_564) );
AND2x2_ASAP7_75t_L g573 ( .A(n_491), .B(n_500), .Y(n_573) );
NAND2x1_ASAP7_75t_L g601 ( .A(n_491), .B(n_508), .Y(n_601) );
AND2x2_ASAP7_75t_L g648 ( .A(n_491), .B(n_543), .Y(n_648) );
OR2x6_ASAP7_75t_L g491 ( .A(n_492), .B(n_493), .Y(n_491) );
HB1xp67_ASAP7_75t_L g499 ( .A(n_500), .Y(n_499) );
INVx1_ASAP7_75t_L g531 ( .A(n_500), .Y(n_531) );
INVx1_ASAP7_75t_L g541 ( .A(n_500), .Y(n_541) );
AND2x2_ASAP7_75t_L g557 ( .A(n_500), .B(n_544), .Y(n_557) );
INVx2_ASAP7_75t_L g562 ( .A(n_500), .Y(n_562) );
OR2x2_ASAP7_75t_L g658 ( .A(n_500), .B(n_508), .Y(n_658) );
AND2x2_ASAP7_75t_L g507 ( .A(n_508), .B(n_517), .Y(n_507) );
NOR2x1_ASAP7_75t_SL g543 ( .A(n_508), .B(n_544), .Y(n_543) );
AND2x2_ASAP7_75t_L g561 ( .A(n_508), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g574 ( .A(n_508), .B(n_518), .Y(n_574) );
BUFx2_ASAP7_75t_L g593 ( .A(n_508), .Y(n_593) );
INVx2_ASAP7_75t_SL g620 ( .A(n_508), .Y(n_620) );
OR2x6_ASAP7_75t_L g508 ( .A(n_509), .B(n_516), .Y(n_508) );
INVx2_ASAP7_75t_L g517 ( .A(n_518), .Y(n_517) );
AND2x2_ASAP7_75t_L g530 ( .A(n_518), .B(n_531), .Y(n_530) );
AND2x2_ASAP7_75t_L g676 ( .A(n_518), .B(n_618), .Y(n_676) );
INVx3_ASAP7_75t_L g518 ( .A(n_519), .Y(n_518) );
AO21x2_ASAP7_75t_L g519 ( .A1(n_520), .A2(n_521), .B(n_527), .Y(n_519) );
AO21x1_ASAP7_75t_SL g544 ( .A1(n_520), .A2(n_521), .B(n_527), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g521 ( .A(n_522), .B(n_526), .Y(n_521) );
AOI211xp5_ASAP7_75t_L g692 ( .A1(n_529), .A2(n_553), .B(n_693), .C(n_697), .Y(n_692) );
AND2x2_ASAP7_75t_L g529 ( .A(n_530), .B(n_532), .Y(n_529) );
NAND2xp5_ASAP7_75t_L g643 ( .A(n_530), .B(n_608), .Y(n_643) );
BUFx2_ASAP7_75t_L g607 ( .A(n_531), .Y(n_607) );
OR2x2_ASAP7_75t_L g555 ( .A(n_532), .B(n_556), .Y(n_555) );
AND2x2_ASAP7_75t_L g640 ( .A(n_532), .B(n_574), .Y(n_640) );
AND2x2_ASAP7_75t_L g661 ( .A(n_532), .B(n_617), .Y(n_661) );
INVx2_ASAP7_75t_L g668 ( .A(n_532), .Y(n_668) );
OAI21xp5_ASAP7_75t_SL g673 ( .A1(n_533), .A2(n_674), .B(n_675), .Y(n_673) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_536), .Y(n_533) );
AND2x2_ASAP7_75t_L g615 ( .A(n_534), .B(n_597), .Y(n_615) );
OR2x2_ASAP7_75t_L g694 ( .A(n_534), .B(n_695), .Y(n_694) );
INVx2_ASAP7_75t_L g534 ( .A(n_535), .Y(n_534) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_535), .B(n_568), .Y(n_567) );
INVx1_ASAP7_75t_L g568 ( .A(n_537), .Y(n_568) );
AND2x2_ASAP7_75t_L g645 ( .A(n_537), .B(n_592), .Y(n_645) );
INVx1_ASAP7_75t_L g538 ( .A(n_539), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_540), .B(n_542), .Y(n_539) );
AND2x2_ASAP7_75t_L g630 ( .A(n_540), .B(n_631), .Y(n_630) );
AND2x4_ASAP7_75t_SL g639 ( .A(n_540), .B(n_640), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g672 ( .A(n_540), .B(n_549), .Y(n_672) );
INVx3_ASAP7_75t_L g540 ( .A(n_541), .Y(n_540) );
AND2x2_ASAP7_75t_L g548 ( .A(n_541), .B(n_549), .Y(n_548) );
OR2x2_ASAP7_75t_L g667 ( .A(n_542), .B(n_668), .Y(n_667) );
INVx2_ASAP7_75t_L g542 ( .A(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g617 ( .A(n_543), .B(n_618), .Y(n_617) );
AND2x2_ASAP7_75t_L g587 ( .A(n_544), .B(n_562), .Y(n_587) );
OAI31xp33_ASAP7_75t_L g594 ( .A1(n_545), .A2(n_595), .A3(n_597), .B(n_599), .Y(n_594) );
INVx1_ASAP7_75t_L g545 ( .A(n_546), .Y(n_545) );
NAND2xp5_ASAP7_75t_SL g596 ( .A(n_547), .B(n_570), .Y(n_596) );
AO21x1_ASAP7_75t_L g550 ( .A1(n_551), .A2(n_554), .B(n_558), .Y(n_550) );
AND2x2_ASAP7_75t_L g551 ( .A(n_552), .B(n_553), .Y(n_551) );
OR2x2_ASAP7_75t_L g606 ( .A(n_552), .B(n_607), .Y(n_606) );
INVx1_ASAP7_75t_L g711 ( .A(n_552), .Y(n_711) );
INVx2_ASAP7_75t_SL g696 ( .A(n_553), .Y(n_696) );
INVx1_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
OR2x2_ASAP7_75t_L g600 ( .A(n_556), .B(n_601), .Y(n_600) );
OR2x2_ASAP7_75t_L g684 ( .A(n_556), .B(n_685), .Y(n_684) );
INVx2_ASAP7_75t_SL g556 ( .A(n_557), .Y(n_556) );
NAND2xp5_ASAP7_75t_L g701 ( .A(n_557), .B(n_620), .Y(n_701) );
OAI22xp5_ASAP7_75t_L g558 ( .A1(n_559), .A2(n_565), .B1(n_569), .B2(n_571), .Y(n_558) );
AOI21xp33_ASAP7_75t_L g677 ( .A1(n_559), .A2(n_678), .B(n_679), .Y(n_677) );
INVx3_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
AND2x4_ASAP7_75t_L g560 ( .A(n_561), .B(n_563), .Y(n_560) );
INVx1_ASAP7_75t_L g618 ( .A(n_562), .Y(n_618) );
INVx1_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
OR2x2_ASAP7_75t_L g632 ( .A(n_564), .B(n_593), .Y(n_632) );
OR2x2_ASAP7_75t_L g657 ( .A(n_564), .B(n_658), .Y(n_657) );
OR2x2_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NAND2xp5_ASAP7_75t_L g569 ( .A(n_566), .B(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_L g578 ( .A(n_566), .B(n_579), .Y(n_578) );
INVx2_ASAP7_75t_L g656 ( .A(n_566), .Y(n_656) );
INVx2_ASAP7_75t_L g585 ( .A(n_567), .Y(n_585) );
INVx1_ASAP7_75t_L g665 ( .A(n_568), .Y(n_665) );
AND2x2_ASAP7_75t_L g588 ( .A(n_570), .B(n_589), .Y(n_588) );
INVx1_ASAP7_75t_L g662 ( .A(n_570), .Y(n_662) );
INVx2_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
AND2x2_ASAP7_75t_L g572 ( .A(n_573), .B(n_574), .Y(n_572) );
NAND2xp5_ASAP7_75t_SL g575 ( .A(n_576), .B(n_594), .Y(n_575) );
OAI321xp33_ASAP7_75t_L g576 ( .A1(n_577), .A2(n_581), .A3(n_586), .B1(n_587), .B2(n_588), .C(n_593), .Y(n_576) );
AOI322xp5_ASAP7_75t_L g702 ( .A1(n_577), .A2(n_608), .A3(n_703), .B1(n_705), .B2(n_707), .C1(n_708), .C2(n_713), .Y(n_702) );
INVx1_ASAP7_75t_L g577 ( .A(n_578), .Y(n_577) );
BUFx2_ASAP7_75t_L g655 ( .A(n_580), .Y(n_655) );
AND2x2_ASAP7_75t_L g581 ( .A(n_582), .B(n_585), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_582), .B(n_662), .Y(n_679) );
INVx2_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
INVx1_ASAP7_75t_L g687 ( .A(n_585), .Y(n_687) );
INVx1_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp33_ASAP7_75t_SL g619 ( .A(n_587), .B(n_620), .Y(n_619) );
INVx1_ASAP7_75t_L g589 ( .A(n_590), .Y(n_589) );
OAI21xp33_ASAP7_75t_SL g686 ( .A1(n_590), .A2(n_596), .B(n_687), .Y(n_686) );
INVx1_ASAP7_75t_SL g591 ( .A(n_592), .Y(n_591) );
INVx1_ASAP7_75t_L g595 ( .A(n_596), .Y(n_595) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
INVx3_ASAP7_75t_L g608 ( .A(n_601), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g602 ( .A(n_603), .B(n_622), .Y(n_602) );
AOI221xp5_ASAP7_75t_L g603 ( .A1(n_604), .A2(n_608), .B1(n_609), .B2(n_610), .C(n_613), .Y(n_603) );
NOR2xp33_ASAP7_75t_L g604 ( .A(n_605), .B(n_606), .Y(n_604) );
HB1xp67_ASAP7_75t_L g624 ( .A(n_605), .Y(n_624) );
AND2x2_ASAP7_75t_L g609 ( .A(n_607), .B(n_608), .Y(n_609) );
INVx2_ASAP7_75t_L g610 ( .A(n_611), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
OAI22xp33_ASAP7_75t_SL g613 ( .A1(n_614), .A2(n_616), .B1(n_619), .B2(n_621), .Y(n_613) );
INVx1_ASAP7_75t_L g614 ( .A(n_615), .Y(n_614) );
INVx1_ASAP7_75t_L g616 ( .A(n_617), .Y(n_616) );
AND2x2_ASAP7_75t_L g625 ( .A(n_617), .B(n_626), .Y(n_625) );
OAI21xp33_ASAP7_75t_L g708 ( .A1(n_620), .A2(n_709), .B(n_710), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_623), .B(n_625), .Y(n_622) );
INVx1_ASAP7_75t_L g623 ( .A(n_624), .Y(n_623) );
NOR3xp33_ASAP7_75t_SL g627 ( .A(n_628), .B(n_659), .C(n_680), .Y(n_627) );
INVx1_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
INVx1_ASAP7_75t_SL g631 ( .A(n_632), .Y(n_631) );
OAI22xp5_ASAP7_75t_L g693 ( .A1(n_632), .A2(n_667), .B1(n_694), .B2(n_696), .Y(n_693) );
OAI21xp33_ASAP7_75t_SL g633 ( .A1(n_634), .A2(n_635), .B(n_639), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_634), .B(n_671), .Y(n_670) );
INVx1_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
HB1xp67_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
AOI221xp5_ASAP7_75t_L g681 ( .A1(n_640), .A2(n_682), .B1(n_683), .B2(n_686), .C(n_688), .Y(n_681) );
AOI221xp5_ASAP7_75t_L g641 ( .A1(n_642), .A2(n_644), .B1(n_646), .B2(n_648), .C(n_649), .Y(n_641) );
INVx1_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_L g678 ( .A(n_644), .Y(n_678) );
INVx1_ASAP7_75t_L g700 ( .A(n_645), .Y(n_700) );
INVx1_ASAP7_75t_SL g698 ( .A(n_646), .Y(n_698) );
AOI31xp33_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_651), .A3(n_653), .B(n_657), .Y(n_649) );
OAI221xp5_ASAP7_75t_L g659 ( .A1(n_650), .A2(n_660), .B1(n_662), .B2(n_663), .C(n_754), .Y(n_659) );
INVx2_ASAP7_75t_L g651 ( .A(n_652), .Y(n_651) );
NAND2xp5_ASAP7_75t_L g653 ( .A(n_654), .B(n_656), .Y(n_653) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g660 ( .A(n_661), .Y(n_660) );
AOI211xp5_ASAP7_75t_L g663 ( .A1(n_664), .A2(n_666), .B(n_669), .C(n_677), .Y(n_663) );
INVx1_ASAP7_75t_L g666 ( .A(n_667), .Y(n_666) );
AND2x2_ASAP7_75t_L g675 ( .A(n_668), .B(n_676), .Y(n_675) );
OAI21xp5_ASAP7_75t_SL g669 ( .A1(n_670), .A2(n_672), .B(n_673), .Y(n_669) );
INVx1_ASAP7_75t_L g704 ( .A(n_676), .Y(n_704) );
BUFx2_ASAP7_75t_SL g713 ( .A(n_676), .Y(n_713) );
NAND3xp33_ASAP7_75t_SL g680 ( .A(n_681), .B(n_692), .C(n_702), .Y(n_680) );
INVx2_ASAP7_75t_L g683 ( .A(n_684), .Y(n_683) );
AOI21xp33_ASAP7_75t_L g688 ( .A1(n_689), .A2(n_690), .B(n_691), .Y(n_688) );
AOI21xp33_ASAP7_75t_L g697 ( .A1(n_698), .A2(n_699), .B(n_701), .Y(n_697) );
HB1xp67_ASAP7_75t_L g703 ( .A(n_704), .Y(n_703) );
INVxp67_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g710 ( .A(n_711), .B(n_712), .Y(n_710) );
INVx1_ASAP7_75t_SL g723 ( .A(n_714), .Y(n_723) );
CKINVDCx11_ASAP7_75t_R g714 ( .A(n_715), .Y(n_714) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
INVx4_ASAP7_75t_SL g720 ( .A(n_721), .Y(n_720) );
INVx3_ASAP7_75t_SL g721 ( .A(n_722), .Y(n_721) );
INVx2_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
INVx3_ASAP7_75t_L g725 ( .A(n_726), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_729), .B(n_733), .Y(n_728) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
CKINVDCx20_ASAP7_75t_R g730 ( .A(n_731), .Y(n_730) );
HB1xp67_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
INVxp67_ASAP7_75t_L g733 ( .A(n_734), .Y(n_733) );
AOI21xp5_ASAP7_75t_L g742 ( .A1(n_734), .A2(n_743), .B(n_747), .Y(n_742) );
NOR2xp33_ASAP7_75t_SL g734 ( .A(n_735), .B(n_738), .Y(n_734) );
HB1xp67_ASAP7_75t_L g735 ( .A(n_736), .Y(n_735) );
BUFx3_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
BUFx2_ASAP7_75t_L g748 ( .A(n_737), .Y(n_748) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_740), .B(n_742), .Y(n_739) );
CKINVDCx5p33_ASAP7_75t_R g740 ( .A(n_741), .Y(n_740) );
HB1xp67_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NOR2xp33_ASAP7_75t_L g749 ( .A(n_750), .B(n_751), .Y(n_749) );
endmodule