module fake_netlist_5_1908_n_3736 (n_137, n_924, n_676, n_294, n_431, n_318, n_380, n_419, n_977, n_653, n_611, n_444, n_642, n_469, n_615, n_851, n_82, n_194, n_316, n_785, n_389, n_843, n_855, n_549, n_684, n_850, n_418, n_248, n_124, n_86, n_136, n_146, n_315, n_268, n_523, n_451, n_532, n_705, n_619, n_408, n_865, n_61, n_913, n_678, n_664, n_376, n_697, n_503, n_967, n_127, n_75, n_235, n_226, n_605, n_74, n_776, n_928, n_667, n_515, n_790, n_57, n_353, n_351, n_367, n_620, n_643, n_1055, n_916, n_452, n_885, n_397, n_493, n_111, n_525, n_880, n_703, n_698, n_980, n_483, n_544, n_683, n_1007, n_155, n_780, n_649, n_552, n_1057, n_1051, n_547, n_43, n_721, n_998, n_116, n_841, n_1050, n_956, n_22, n_467, n_564, n_802, n_423, n_840, n_284, n_46, n_245, n_21, n_501, n_823, n_725, n_983, n_139, n_38, n_105, n_280, n_744, n_1021, n_590, n_629, n_672, n_4, n_873, n_378, n_551, n_762, n_17, n_581, n_688, n_382, n_554, n_800, n_898, n_254, n_690, n_33, n_1013, n_23, n_583, n_671, n_718, n_819, n_302, n_265, n_1022, n_526, n_915, n_719, n_293, n_372, n_443, n_244, n_677, n_47, n_173, n_859, n_864, n_951, n_821, n_198, n_714, n_447, n_247, n_314, n_368, n_433, n_604, n_8, n_321, n_292, n_909, n_625, n_854, n_949, n_621, n_753, n_997, n_100, n_455, n_674, n_1008, n_932, n_417, n_946, n_1048, n_612, n_1001, n_212, n_385, n_498, n_516, n_933, n_788, n_507, n_119, n_497, n_689, n_738, n_912, n_606, n_559, n_275, n_640, n_968, n_252, n_624, n_825, n_26, n_295, n_133, n_1010, n_330, n_877, n_508, n_739, n_506, n_2, n_737, n_610, n_972, n_692, n_986, n_755, n_6, n_509, n_568, n_936, n_39, n_147, n_373, n_820, n_757, n_947, n_67, n_307, n_633, n_439, n_87, n_150, n_530, n_1024, n_556, n_106, n_209, n_259, n_448, n_758, n_999, n_668, n_733, n_991, n_375, n_301, n_828, n_779, n_576, n_941, n_929, n_981, n_1032, n_68, n_804, n_93, n_867, n_186, n_537, n_134, n_902, n_191, n_587, n_945, n_659, n_51, n_63, n_492, n_792, n_563, n_171, n_153, n_756, n_878, n_524, n_943, n_399, n_341, n_204, n_394, n_250, n_579, n_992, n_1049, n_938, n_741, n_548, n_543, n_260, n_812, n_842, n_298, n_650, n_984, n_320, n_694, n_518, n_505, n_286, n_883, n_122, n_282, n_752, n_331, n_10, n_905, n_906, n_24, n_406, n_519, n_470, n_908, n_782, n_919, n_325, n_449, n_132, n_862, n_90, n_900, n_724, n_856, n_546, n_1016, n_101, n_760, n_658, n_281, n_918, n_240, n_942, n_381, n_189, n_220, n_291, n_231, n_257, n_390, n_731, n_31, n_456, n_13, n_371, n_959, n_481, n_535, n_709, n_152, n_540, n_317, n_618, n_940, n_896, n_9, n_323, n_569, n_769, n_195, n_42, n_356, n_227, n_592, n_45, n_920, n_894, n_1046, n_271, n_934, n_1017, n_94, n_831, n_826, n_335, n_123, n_886, n_978, n_964, n_1054, n_654, n_370, n_167, n_976, n_234, n_343, n_308, n_379, n_428, n_267, n_514, n_457, n_570, n_833, n_297, n_1045, n_156, n_5, n_853, n_603, n_225, n_377, n_751, n_484, n_775, n_219, n_1033, n_988, n_442, n_157, n_814, n_131, n_192, n_636, n_786, n_600, n_660, n_223, n_392, n_158, n_655, n_704, n_787, n_1009, n_138, n_264, n_109, n_669, n_472, n_742, n_750, n_454, n_961, n_995, n_955, n_387, n_771, n_374, n_163, n_276, n_339, n_95, n_882, n_183, n_185, n_243, n_398, n_396, n_1036, n_635, n_347, n_763, n_169, n_59, n_522, n_550, n_255, n_696, n_897, n_215, n_350, n_196, n_798, n_662, n_459, n_1020, n_646, n_211, n_218, n_400, n_930, n_181, n_436, n_962, n_3, n_290, n_580, n_221, n_178, n_622, n_1040, n_723, n_1035, n_386, n_578, n_994, n_926, n_287, n_344, n_848, n_555, n_783, n_473, n_422, n_475, n_777, n_1030, n_72, n_661, n_104, n_41, n_682, n_415, n_56, n_141, n_485, n_1043, n_496, n_355, n_958, n_849, n_1034, n_486, n_670, n_15, n_816, n_336, n_584, n_681, n_591, n_922, n_145, n_48, n_521, n_614, n_663, n_845, n_50, n_337, n_430, n_313, n_631, n_673, n_837, n_88, n_479, n_528, n_510, n_216, n_680, n_168, n_974, n_395, n_164, n_432, n_553, n_727, n_839, n_901, n_311, n_813, n_957, n_830, n_773, n_208, n_142, n_743, n_214, n_328, n_140, n_801, n_299, n_303, n_369, n_675, n_888, n_296, n_613, n_871, n_241, n_637, n_357, n_875, n_598, n_685, n_608, n_184, n_446, n_445, n_65, n_78, n_749, n_829, n_144, n_858, n_114, n_96, n_923, n_772, n_691, n_881, n_717, n_165, n_468, n_499, n_939, n_213, n_129, n_342, n_482, n_517, n_98, n_588, n_361, n_464, n_789, n_363, n_402, n_413, n_734, n_638, n_700, n_197, n_796, n_107, n_573, n_69, n_866, n_969, n_236, n_388, n_761, n_1012, n_1, n_1019, n_249, n_903, n_1006, n_740, n_304, n_329, n_203, n_274, n_577, n_384, n_582, n_460, n_889, n_80, n_973, n_35, n_73, n_277, n_92, n_19, n_338, n_149, n_477, n_461, n_333, n_571, n_693, n_309, n_30, n_512, n_14, n_836, n_990, n_84, n_462, n_975, n_130, n_322, n_567, n_258, n_652, n_778, n_29, n_79, n_151, n_25, n_306, n_907, n_722, n_458, n_288, n_770, n_188, n_190, n_844, n_201, n_1031, n_263, n_471, n_609, n_852, n_989, n_1041, n_1039, n_44, n_224, n_40, n_34, n_228, n_283, n_1028, n_383, n_711, n_781, n_834, n_474, n_112, n_765, n_542, n_85, n_463, n_488, n_595, n_736, n_502, n_892, n_893, n_1015, n_1000, n_891, n_239, n_466, n_420, n_630, n_489, n_632, n_699, n_55, n_979, n_1002, n_617, n_49, n_310, n_54, n_593, n_504, n_511, n_12, n_748, n_586, n_846, n_874, n_465, n_838, n_76, n_358, n_1058, n_362, n_876, n_170, n_332, n_27, n_1053, n_77, n_102, n_161, n_273, n_349, n_585, n_270, n_616, n_230, n_81, n_118, n_953, n_601, n_279, n_917, n_1014, n_966, n_70, n_987, n_253, n_261, n_174, n_289, n_745, n_963, n_1052, n_954, n_627, n_767, n_172, n_206, n_217, n_993, n_440, n_726, n_478, n_793, n_545, n_982, n_441, n_860, n_450, n_648, n_312, n_476, n_818, n_429, n_861, n_534, n_948, n_884, n_899, n_345, n_210, n_944, n_494, n_641, n_628, n_365, n_774, n_91, n_729, n_730, n_1059, n_176, n_970, n_911, n_557, n_182, n_143, n_83, n_1005, n_354, n_575, n_607, n_480, n_647, n_237, n_425, n_513, n_407, n_527, n_679, n_707, n_710, n_795, n_695, n_832, n_180, n_857, n_560, n_656, n_340, n_207, n_561, n_1044, n_37, n_346, n_937, n_393, n_229, n_108, n_487, n_495, n_602, n_665, n_574, n_437, n_66, n_177, n_60, n_403, n_453, n_421, n_879, n_16, n_720, n_0, n_58, n_623, n_405, n_824, n_18, n_359, n_863, n_910, n_971, n_490, n_805, n_1027, n_117, n_326, n_794, n_768, n_921, n_996, n_233, n_404, n_686, n_205, n_366, n_572, n_113, n_712, n_754, n_847, n_815, n_246, n_596, n_179, n_125, n_410, n_1042, n_558, n_708, n_269, n_529, n_128, n_735, n_702, n_285, n_822, n_412, n_120, n_232, n_327, n_135, n_657, n_126, n_644, n_728, n_895, n_1037, n_202, n_266, n_272, n_491, n_427, n_791, n_732, n_193, n_251, n_352, n_53, n_160, n_565, n_426, n_520, n_566, n_808, n_409, n_797, n_1038, n_1025, n_887, n_589, n_716, n_597, n_500, n_562, n_154, n_62, n_148, n_71, n_300, n_651, n_435, n_809, n_870, n_931, n_159, n_334, n_599, n_766, n_811, n_952, n_541, n_807, n_391, n_701, n_434, n_1023, n_645, n_539, n_835, n_175, n_538, n_666, n_262, n_803, n_868, n_238, n_639, n_799, n_914, n_99, n_687, n_715, n_411, n_414, n_1026, n_319, n_364, n_965, n_927, n_20, n_536, n_531, n_935, n_1004, n_121, n_242, n_817, n_872, n_360, n_36, n_594, n_764, n_200, n_890, n_1056, n_162, n_960, n_64, n_759, n_1018, n_222, n_28, n_89, n_438, n_806, n_115, n_713, n_1011, n_904, n_985, n_1047, n_869, n_324, n_810, n_634, n_416, n_199, n_827, n_187, n_32, n_401, n_103, n_348, n_97, n_1029, n_166, n_626, n_11, n_925, n_424, n_1003, n_7, n_706, n_746, n_256, n_305, n_533, n_950, n_747, n_52, n_278, n_784, n_110, n_3736);

input n_137;
input n_924;
input n_676;
input n_294;
input n_431;
input n_318;
input n_380;
input n_419;
input n_977;
input n_653;
input n_611;
input n_444;
input n_642;
input n_469;
input n_615;
input n_851;
input n_82;
input n_194;
input n_316;
input n_785;
input n_389;
input n_843;
input n_855;
input n_549;
input n_684;
input n_850;
input n_418;
input n_248;
input n_124;
input n_86;
input n_136;
input n_146;
input n_315;
input n_268;
input n_523;
input n_451;
input n_532;
input n_705;
input n_619;
input n_408;
input n_865;
input n_61;
input n_913;
input n_678;
input n_664;
input n_376;
input n_697;
input n_503;
input n_967;
input n_127;
input n_75;
input n_235;
input n_226;
input n_605;
input n_74;
input n_776;
input n_928;
input n_667;
input n_515;
input n_790;
input n_57;
input n_353;
input n_351;
input n_367;
input n_620;
input n_643;
input n_1055;
input n_916;
input n_452;
input n_885;
input n_397;
input n_493;
input n_111;
input n_525;
input n_880;
input n_703;
input n_698;
input n_980;
input n_483;
input n_544;
input n_683;
input n_1007;
input n_155;
input n_780;
input n_649;
input n_552;
input n_1057;
input n_1051;
input n_547;
input n_43;
input n_721;
input n_998;
input n_116;
input n_841;
input n_1050;
input n_956;
input n_22;
input n_467;
input n_564;
input n_802;
input n_423;
input n_840;
input n_284;
input n_46;
input n_245;
input n_21;
input n_501;
input n_823;
input n_725;
input n_983;
input n_139;
input n_38;
input n_105;
input n_280;
input n_744;
input n_1021;
input n_590;
input n_629;
input n_672;
input n_4;
input n_873;
input n_378;
input n_551;
input n_762;
input n_17;
input n_581;
input n_688;
input n_382;
input n_554;
input n_800;
input n_898;
input n_254;
input n_690;
input n_33;
input n_1013;
input n_23;
input n_583;
input n_671;
input n_718;
input n_819;
input n_302;
input n_265;
input n_1022;
input n_526;
input n_915;
input n_719;
input n_293;
input n_372;
input n_443;
input n_244;
input n_677;
input n_47;
input n_173;
input n_859;
input n_864;
input n_951;
input n_821;
input n_198;
input n_714;
input n_447;
input n_247;
input n_314;
input n_368;
input n_433;
input n_604;
input n_8;
input n_321;
input n_292;
input n_909;
input n_625;
input n_854;
input n_949;
input n_621;
input n_753;
input n_997;
input n_100;
input n_455;
input n_674;
input n_1008;
input n_932;
input n_417;
input n_946;
input n_1048;
input n_612;
input n_1001;
input n_212;
input n_385;
input n_498;
input n_516;
input n_933;
input n_788;
input n_507;
input n_119;
input n_497;
input n_689;
input n_738;
input n_912;
input n_606;
input n_559;
input n_275;
input n_640;
input n_968;
input n_252;
input n_624;
input n_825;
input n_26;
input n_295;
input n_133;
input n_1010;
input n_330;
input n_877;
input n_508;
input n_739;
input n_506;
input n_2;
input n_737;
input n_610;
input n_972;
input n_692;
input n_986;
input n_755;
input n_6;
input n_509;
input n_568;
input n_936;
input n_39;
input n_147;
input n_373;
input n_820;
input n_757;
input n_947;
input n_67;
input n_307;
input n_633;
input n_439;
input n_87;
input n_150;
input n_530;
input n_1024;
input n_556;
input n_106;
input n_209;
input n_259;
input n_448;
input n_758;
input n_999;
input n_668;
input n_733;
input n_991;
input n_375;
input n_301;
input n_828;
input n_779;
input n_576;
input n_941;
input n_929;
input n_981;
input n_1032;
input n_68;
input n_804;
input n_93;
input n_867;
input n_186;
input n_537;
input n_134;
input n_902;
input n_191;
input n_587;
input n_945;
input n_659;
input n_51;
input n_63;
input n_492;
input n_792;
input n_563;
input n_171;
input n_153;
input n_756;
input n_878;
input n_524;
input n_943;
input n_399;
input n_341;
input n_204;
input n_394;
input n_250;
input n_579;
input n_992;
input n_1049;
input n_938;
input n_741;
input n_548;
input n_543;
input n_260;
input n_812;
input n_842;
input n_298;
input n_650;
input n_984;
input n_320;
input n_694;
input n_518;
input n_505;
input n_286;
input n_883;
input n_122;
input n_282;
input n_752;
input n_331;
input n_10;
input n_905;
input n_906;
input n_24;
input n_406;
input n_519;
input n_470;
input n_908;
input n_782;
input n_919;
input n_325;
input n_449;
input n_132;
input n_862;
input n_90;
input n_900;
input n_724;
input n_856;
input n_546;
input n_1016;
input n_101;
input n_760;
input n_658;
input n_281;
input n_918;
input n_240;
input n_942;
input n_381;
input n_189;
input n_220;
input n_291;
input n_231;
input n_257;
input n_390;
input n_731;
input n_31;
input n_456;
input n_13;
input n_371;
input n_959;
input n_481;
input n_535;
input n_709;
input n_152;
input n_540;
input n_317;
input n_618;
input n_940;
input n_896;
input n_9;
input n_323;
input n_569;
input n_769;
input n_195;
input n_42;
input n_356;
input n_227;
input n_592;
input n_45;
input n_920;
input n_894;
input n_1046;
input n_271;
input n_934;
input n_1017;
input n_94;
input n_831;
input n_826;
input n_335;
input n_123;
input n_886;
input n_978;
input n_964;
input n_1054;
input n_654;
input n_370;
input n_167;
input n_976;
input n_234;
input n_343;
input n_308;
input n_379;
input n_428;
input n_267;
input n_514;
input n_457;
input n_570;
input n_833;
input n_297;
input n_1045;
input n_156;
input n_5;
input n_853;
input n_603;
input n_225;
input n_377;
input n_751;
input n_484;
input n_775;
input n_219;
input n_1033;
input n_988;
input n_442;
input n_157;
input n_814;
input n_131;
input n_192;
input n_636;
input n_786;
input n_600;
input n_660;
input n_223;
input n_392;
input n_158;
input n_655;
input n_704;
input n_787;
input n_1009;
input n_138;
input n_264;
input n_109;
input n_669;
input n_472;
input n_742;
input n_750;
input n_454;
input n_961;
input n_995;
input n_955;
input n_387;
input n_771;
input n_374;
input n_163;
input n_276;
input n_339;
input n_95;
input n_882;
input n_183;
input n_185;
input n_243;
input n_398;
input n_396;
input n_1036;
input n_635;
input n_347;
input n_763;
input n_169;
input n_59;
input n_522;
input n_550;
input n_255;
input n_696;
input n_897;
input n_215;
input n_350;
input n_196;
input n_798;
input n_662;
input n_459;
input n_1020;
input n_646;
input n_211;
input n_218;
input n_400;
input n_930;
input n_181;
input n_436;
input n_962;
input n_3;
input n_290;
input n_580;
input n_221;
input n_178;
input n_622;
input n_1040;
input n_723;
input n_1035;
input n_386;
input n_578;
input n_994;
input n_926;
input n_287;
input n_344;
input n_848;
input n_555;
input n_783;
input n_473;
input n_422;
input n_475;
input n_777;
input n_1030;
input n_72;
input n_661;
input n_104;
input n_41;
input n_682;
input n_415;
input n_56;
input n_141;
input n_485;
input n_1043;
input n_496;
input n_355;
input n_958;
input n_849;
input n_1034;
input n_486;
input n_670;
input n_15;
input n_816;
input n_336;
input n_584;
input n_681;
input n_591;
input n_922;
input n_145;
input n_48;
input n_521;
input n_614;
input n_663;
input n_845;
input n_50;
input n_337;
input n_430;
input n_313;
input n_631;
input n_673;
input n_837;
input n_88;
input n_479;
input n_528;
input n_510;
input n_216;
input n_680;
input n_168;
input n_974;
input n_395;
input n_164;
input n_432;
input n_553;
input n_727;
input n_839;
input n_901;
input n_311;
input n_813;
input n_957;
input n_830;
input n_773;
input n_208;
input n_142;
input n_743;
input n_214;
input n_328;
input n_140;
input n_801;
input n_299;
input n_303;
input n_369;
input n_675;
input n_888;
input n_296;
input n_613;
input n_871;
input n_241;
input n_637;
input n_357;
input n_875;
input n_598;
input n_685;
input n_608;
input n_184;
input n_446;
input n_445;
input n_65;
input n_78;
input n_749;
input n_829;
input n_144;
input n_858;
input n_114;
input n_96;
input n_923;
input n_772;
input n_691;
input n_881;
input n_717;
input n_165;
input n_468;
input n_499;
input n_939;
input n_213;
input n_129;
input n_342;
input n_482;
input n_517;
input n_98;
input n_588;
input n_361;
input n_464;
input n_789;
input n_363;
input n_402;
input n_413;
input n_734;
input n_638;
input n_700;
input n_197;
input n_796;
input n_107;
input n_573;
input n_69;
input n_866;
input n_969;
input n_236;
input n_388;
input n_761;
input n_1012;
input n_1;
input n_1019;
input n_249;
input n_903;
input n_1006;
input n_740;
input n_304;
input n_329;
input n_203;
input n_274;
input n_577;
input n_384;
input n_582;
input n_460;
input n_889;
input n_80;
input n_973;
input n_35;
input n_73;
input n_277;
input n_92;
input n_19;
input n_338;
input n_149;
input n_477;
input n_461;
input n_333;
input n_571;
input n_693;
input n_309;
input n_30;
input n_512;
input n_14;
input n_836;
input n_990;
input n_84;
input n_462;
input n_975;
input n_130;
input n_322;
input n_567;
input n_258;
input n_652;
input n_778;
input n_29;
input n_79;
input n_151;
input n_25;
input n_306;
input n_907;
input n_722;
input n_458;
input n_288;
input n_770;
input n_188;
input n_190;
input n_844;
input n_201;
input n_1031;
input n_263;
input n_471;
input n_609;
input n_852;
input n_989;
input n_1041;
input n_1039;
input n_44;
input n_224;
input n_40;
input n_34;
input n_228;
input n_283;
input n_1028;
input n_383;
input n_711;
input n_781;
input n_834;
input n_474;
input n_112;
input n_765;
input n_542;
input n_85;
input n_463;
input n_488;
input n_595;
input n_736;
input n_502;
input n_892;
input n_893;
input n_1015;
input n_1000;
input n_891;
input n_239;
input n_466;
input n_420;
input n_630;
input n_489;
input n_632;
input n_699;
input n_55;
input n_979;
input n_1002;
input n_617;
input n_49;
input n_310;
input n_54;
input n_593;
input n_504;
input n_511;
input n_12;
input n_748;
input n_586;
input n_846;
input n_874;
input n_465;
input n_838;
input n_76;
input n_358;
input n_1058;
input n_362;
input n_876;
input n_170;
input n_332;
input n_27;
input n_1053;
input n_77;
input n_102;
input n_161;
input n_273;
input n_349;
input n_585;
input n_270;
input n_616;
input n_230;
input n_81;
input n_118;
input n_953;
input n_601;
input n_279;
input n_917;
input n_1014;
input n_966;
input n_70;
input n_987;
input n_253;
input n_261;
input n_174;
input n_289;
input n_745;
input n_963;
input n_1052;
input n_954;
input n_627;
input n_767;
input n_172;
input n_206;
input n_217;
input n_993;
input n_440;
input n_726;
input n_478;
input n_793;
input n_545;
input n_982;
input n_441;
input n_860;
input n_450;
input n_648;
input n_312;
input n_476;
input n_818;
input n_429;
input n_861;
input n_534;
input n_948;
input n_884;
input n_899;
input n_345;
input n_210;
input n_944;
input n_494;
input n_641;
input n_628;
input n_365;
input n_774;
input n_91;
input n_729;
input n_730;
input n_1059;
input n_176;
input n_970;
input n_911;
input n_557;
input n_182;
input n_143;
input n_83;
input n_1005;
input n_354;
input n_575;
input n_607;
input n_480;
input n_647;
input n_237;
input n_425;
input n_513;
input n_407;
input n_527;
input n_679;
input n_707;
input n_710;
input n_795;
input n_695;
input n_832;
input n_180;
input n_857;
input n_560;
input n_656;
input n_340;
input n_207;
input n_561;
input n_1044;
input n_37;
input n_346;
input n_937;
input n_393;
input n_229;
input n_108;
input n_487;
input n_495;
input n_602;
input n_665;
input n_574;
input n_437;
input n_66;
input n_177;
input n_60;
input n_403;
input n_453;
input n_421;
input n_879;
input n_16;
input n_720;
input n_0;
input n_58;
input n_623;
input n_405;
input n_824;
input n_18;
input n_359;
input n_863;
input n_910;
input n_971;
input n_490;
input n_805;
input n_1027;
input n_117;
input n_326;
input n_794;
input n_768;
input n_921;
input n_996;
input n_233;
input n_404;
input n_686;
input n_205;
input n_366;
input n_572;
input n_113;
input n_712;
input n_754;
input n_847;
input n_815;
input n_246;
input n_596;
input n_179;
input n_125;
input n_410;
input n_1042;
input n_558;
input n_708;
input n_269;
input n_529;
input n_128;
input n_735;
input n_702;
input n_285;
input n_822;
input n_412;
input n_120;
input n_232;
input n_327;
input n_135;
input n_657;
input n_126;
input n_644;
input n_728;
input n_895;
input n_1037;
input n_202;
input n_266;
input n_272;
input n_491;
input n_427;
input n_791;
input n_732;
input n_193;
input n_251;
input n_352;
input n_53;
input n_160;
input n_565;
input n_426;
input n_520;
input n_566;
input n_808;
input n_409;
input n_797;
input n_1038;
input n_1025;
input n_887;
input n_589;
input n_716;
input n_597;
input n_500;
input n_562;
input n_154;
input n_62;
input n_148;
input n_71;
input n_300;
input n_651;
input n_435;
input n_809;
input n_870;
input n_931;
input n_159;
input n_334;
input n_599;
input n_766;
input n_811;
input n_952;
input n_541;
input n_807;
input n_391;
input n_701;
input n_434;
input n_1023;
input n_645;
input n_539;
input n_835;
input n_175;
input n_538;
input n_666;
input n_262;
input n_803;
input n_868;
input n_238;
input n_639;
input n_799;
input n_914;
input n_99;
input n_687;
input n_715;
input n_411;
input n_414;
input n_1026;
input n_319;
input n_364;
input n_965;
input n_927;
input n_20;
input n_536;
input n_531;
input n_935;
input n_1004;
input n_121;
input n_242;
input n_817;
input n_872;
input n_360;
input n_36;
input n_594;
input n_764;
input n_200;
input n_890;
input n_1056;
input n_162;
input n_960;
input n_64;
input n_759;
input n_1018;
input n_222;
input n_28;
input n_89;
input n_438;
input n_806;
input n_115;
input n_713;
input n_1011;
input n_904;
input n_985;
input n_1047;
input n_869;
input n_324;
input n_810;
input n_634;
input n_416;
input n_199;
input n_827;
input n_187;
input n_32;
input n_401;
input n_103;
input n_348;
input n_97;
input n_1029;
input n_166;
input n_626;
input n_11;
input n_925;
input n_424;
input n_1003;
input n_7;
input n_706;
input n_746;
input n_256;
input n_305;
input n_533;
input n_950;
input n_747;
input n_52;
input n_278;
input n_784;
input n_110;

output n_3736;

wire n_1263;
wire n_3304;
wire n_1378;
wire n_2253;
wire n_2417;
wire n_2756;
wire n_1126;
wire n_1423;
wire n_1729;
wire n_2739;
wire n_1166;
wire n_2380;
wire n_1751;
wire n_1508;
wire n_2771;
wire n_3241;
wire n_2617;
wire n_2200;
wire n_3261;
wire n_3006;
wire n_1161;
wire n_3027;
wire n_1859;
wire n_2746;
wire n_1677;
wire n_1150;
wire n_2327;
wire n_3179;
wire n_3127;
wire n_1780;
wire n_3256;
wire n_3732;
wire n_1488;
wire n_2899;
wire n_2955;
wire n_3619;
wire n_3541;
wire n_3622;
wire n_2386;
wire n_3596;
wire n_1501;
wire n_2395;
wire n_3086;
wire n_3297;
wire n_2369;
wire n_2927;
wire n_1528;
wire n_2683;
wire n_1370;
wire n_1292;
wire n_2520;
wire n_2347;
wire n_2821;
wire n_1360;
wire n_1198;
wire n_2388;
wire n_1099;
wire n_2568;
wire n_3641;
wire n_1738;
wire n_2021;
wire n_3728;
wire n_2134;
wire n_3064;
wire n_2391;
wire n_3088;
wire n_1960;
wire n_2843;
wire n_2185;
wire n_3270;
wire n_2143;
wire n_3713;
wire n_2853;
wire n_3615;
wire n_2059;
wire n_1323;
wire n_3663;
wire n_1466;
wire n_1695;
wire n_2487;
wire n_1353;
wire n_3595;
wire n_3246;
wire n_3202;
wire n_1347;
wire n_2495;
wire n_2880;
wire n_1535;
wire n_1789;
wire n_1666;
wire n_3350;
wire n_2389;
wire n_1451;
wire n_2302;
wire n_1545;
wire n_2374;
wire n_3341;
wire n_1947;
wire n_1264;
wire n_3587;
wire n_2114;
wire n_3445;
wire n_2001;
wire n_1494;
wire n_3407;
wire n_3571;
wire n_3599;
wire n_1462;
wire n_1799;
wire n_2069;
wire n_2396;
wire n_3621;
wire n_1580;
wire n_1939;
wire n_2486;
wire n_3434;
wire n_1806;
wire n_2244;
wire n_2257;
wire n_1152;
wire n_3501;
wire n_3448;
wire n_1869;
wire n_1607;
wire n_1563;
wire n_3019;
wire n_3039;
wire n_2011;
wire n_2096;
wire n_2105;
wire n_2538;
wire n_2024;
wire n_2530;
wire n_1696;
wire n_2483;
wire n_3163;
wire n_1118;
wire n_1686;
wire n_1285;
wire n_3710;
wire n_1860;
wire n_2543;
wire n_1359;
wire n_1728;
wire n_1107;
wire n_2031;
wire n_2076;
wire n_2482;
wire n_3036;
wire n_2677;
wire n_1230;
wire n_2165;
wire n_1896;
wire n_2147;
wire n_3010;
wire n_3180;
wire n_3379;
wire n_3532;
wire n_2770;
wire n_1124;
wire n_1818;
wire n_2127;
wire n_1576;
wire n_1104;
wire n_1705;
wire n_1294;
wire n_2584;
wire n_1257;
wire n_2639;
wire n_1182;
wire n_3188;
wire n_3325;
wire n_3107;
wire n_3531;
wire n_3403;
wire n_1698;
wire n_1261;
wire n_2329;
wire n_1098;
wire n_2963;
wire n_3624;
wire n_2142;
wire n_3186;
wire n_3461;
wire n_3082;
wire n_1154;
wire n_2189;
wire n_3332;
wire n_1242;
wire n_3283;
wire n_1135;
wire n_3048;
wire n_3258;
wire n_3696;
wire n_2323;
wire n_2203;
wire n_2597;
wire n_1243;
wire n_2959;
wire n_3340;
wire n_2047;
wire n_1280;
wire n_3277;
wire n_1845;
wire n_2052;
wire n_2193;
wire n_2978;
wire n_2058;
wire n_2458;
wire n_2478;
wire n_3650;
wire n_2761;
wire n_1483;
wire n_2888;
wire n_3638;
wire n_1314;
wire n_1512;
wire n_3157;
wire n_1490;
wire n_1236;
wire n_1633;
wire n_2537;
wire n_2983;
wire n_2669;
wire n_2144;
wire n_1778;
wire n_3214;
wire n_2306;
wire n_2515;
wire n_3022;
wire n_1289;
wire n_1517;
wire n_2091;
wire n_2466;
wire n_2652;
wire n_2635;
wire n_3631;
wire n_2715;
wire n_3087;
wire n_2085;
wire n_3489;
wire n_1669;
wire n_2566;
wire n_1949;
wire n_1449;
wire n_1946;
wire n_2936;
wire n_1566;
wire n_2032;
wire n_2587;
wire n_2149;
wire n_1078;
wire n_2782;
wire n_1670;
wire n_2672;
wire n_3060;
wire n_2651;
wire n_3490;
wire n_3656;
wire n_2071;
wire n_1484;
wire n_2561;
wire n_1374;
wire n_1328;
wire n_2643;
wire n_2141;
wire n_1948;
wire n_3013;
wire n_3183;
wire n_1984;
wire n_3437;
wire n_2099;
wire n_2408;
wire n_3446;
wire n_3353;
wire n_1877;
wire n_3687;
wire n_1831;
wire n_1598;
wire n_3049;
wire n_1723;
wire n_1850;
wire n_3028;
wire n_1146;
wire n_2384;
wire n_1097;
wire n_1749;
wire n_3156;
wire n_3101;
wire n_3669;
wire n_3376;
wire n_1428;
wire n_2663;
wire n_1394;
wire n_2659;
wire n_3653;
wire n_1414;
wire n_1216;
wire n_2693;
wire n_3702;
wire n_2202;
wire n_2648;
wire n_1872;
wire n_3389;
wire n_1852;
wire n_2159;
wire n_2976;
wire n_2249;
wire n_2180;
wire n_2353;
wire n_1218;
wire n_1931;
wire n_2439;
wire n_2632;
wire n_2276;
wire n_3089;
wire n_1070;
wire n_1547;
wire n_2089;
wire n_3420;
wire n_2470;
wire n_1755;
wire n_3222;
wire n_1561;
wire n_1071;
wire n_1165;
wire n_1267;
wire n_1801;
wire n_1391;
wire n_1513;
wire n_2908;
wire n_2970;
wire n_3361;
wire n_1600;
wire n_2235;
wire n_1862;
wire n_1239;
wire n_2915;
wire n_2300;
wire n_2791;
wire n_1796;
wire n_2551;
wire n_3291;
wire n_1587;
wire n_1473;
wire n_2682;
wire n_2432;
wire n_3668;
wire n_1521;
wire n_1284;
wire n_1590;
wire n_3440;
wire n_3405;
wire n_2174;
wire n_2714;
wire n_1748;
wire n_3563;
wire n_2934;
wire n_1672;
wire n_2506;
wire n_2699;
wire n_1880;
wire n_2769;
wire n_3550;
wire n_2337;
wire n_3436;
wire n_1167;
wire n_1626;
wire n_3542;
wire n_2615;
wire n_1384;
wire n_1556;
wire n_1863;
wire n_1064;
wire n_2079;
wire n_2238;
wire n_2118;
wire n_1151;
wire n_2985;
wire n_2944;
wire n_1405;
wire n_2407;
wire n_1706;
wire n_3418;
wire n_2932;
wire n_2753;
wire n_2980;
wire n_1582;
wire n_3637;
wire n_1069;
wire n_3306;
wire n_1784;
wire n_2859;
wire n_2842;
wire n_1075;
wire n_3262;
wire n_3136;
wire n_1836;
wire n_2868;
wire n_3395;
wire n_1450;
wire n_3141;
wire n_1322;
wire n_2101;
wire n_1471;
wire n_1986;
wire n_2863;
wire n_2072;
wire n_3164;
wire n_2738;
wire n_1750;
wire n_3570;
wire n_3690;
wire n_1459;
wire n_2358;
wire n_3716;
wire n_2968;
wire n_1700;
wire n_2833;
wire n_3191;
wire n_1585;
wire n_2712;
wire n_2684;
wire n_3593;
wire n_3193;
wire n_1971;
wire n_1599;
wire n_3252;
wire n_2275;
wire n_2855;
wire n_3507;
wire n_3273;
wire n_2713;
wire n_3544;
wire n_2644;
wire n_2700;
wire n_1211;
wire n_1197;
wire n_3367;
wire n_2951;
wire n_1523;
wire n_2730;
wire n_1950;
wire n_3008;
wire n_3709;
wire n_1447;
wire n_2251;
wire n_3096;
wire n_1377;
wire n_2370;
wire n_3496;
wire n_2544;
wire n_2214;
wire n_3339;
wire n_2055;
wire n_3427;
wire n_3025;
wire n_3349;
wire n_1403;
wire n_3735;
wire n_2248;
wire n_2356;
wire n_3320;
wire n_3007;
wire n_2688;
wire n_1202;
wire n_2750;
wire n_2620;
wire n_1278;
wire n_2622;
wire n_2062;
wire n_2668;
wire n_3714;
wire n_1463;
wire n_1581;
wire n_2100;
wire n_3071;
wire n_3651;
wire n_3310;
wire n_3487;
wire n_2258;
wire n_1667;
wire n_3359;
wire n_2784;
wire n_3718;
wire n_2919;
wire n_3092;
wire n_3470;
wire n_1224;
wire n_2865;
wire n_2557;
wire n_1926;
wire n_2706;
wire n_1248;
wire n_1331;
wire n_1241;
wire n_3676;
wire n_2150;
wire n_3146;
wire n_2241;
wire n_2757;
wire n_2152;
wire n_3598;
wire n_1385;
wire n_2590;
wire n_2776;
wire n_2140;
wire n_2385;
wire n_3580;
wire n_1819;
wire n_2330;
wire n_2139;
wire n_2942;
wire n_2987;
wire n_1527;
wire n_2042;
wire n_3106;
wire n_1882;
wire n_3328;
wire n_1754;
wire n_3611;
wire n_1623;
wire n_2862;
wire n_2175;
wire n_2921;
wire n_2720;
wire n_2324;
wire n_1854;
wire n_2606;
wire n_2674;
wire n_3187;
wire n_1565;
wire n_3508;
wire n_2828;
wire n_3682;
wire n_3371;
wire n_1809;
wire n_1856;
wire n_3433;
wire n_1072;
wire n_2218;
wire n_2267;
wire n_2305;
wire n_3430;
wire n_3392;
wire n_2636;
wire n_2450;
wire n_3208;
wire n_1319;
wire n_2379;
wire n_3331;
wire n_3447;
wire n_2616;
wire n_2911;
wire n_3305;
wire n_2154;
wire n_1825;
wire n_1951;
wire n_1906;
wire n_1883;
wire n_2759;
wire n_1712;
wire n_1387;
wire n_3528;
wire n_3649;
wire n_2262;
wire n_2462;
wire n_2514;
wire n_1532;
wire n_2322;
wire n_2271;
wire n_2625;
wire n_3257;
wire n_3625;
wire n_1156;
wire n_2798;
wire n_2945;
wire n_2331;
wire n_2293;
wire n_2837;
wire n_1393;
wire n_2319;
wire n_1775;
wire n_2979;
wire n_3296;
wire n_2028;
wire n_1368;
wire n_3481;
wire n_2762;
wire n_3655;
wire n_2808;
wire n_1276;
wire n_3009;
wire n_2548;
wire n_1412;
wire n_2676;
wire n_1709;
wire n_2679;
wire n_2108;
wire n_3640;
wire n_1538;
wire n_1162;
wire n_2930;
wire n_1838;
wire n_1199;
wire n_1847;
wire n_1779;
wire n_2767;
wire n_2777;
wire n_2603;
wire n_3514;
wire n_3116;
wire n_1884;
wire n_2434;
wire n_2660;
wire n_3602;
wire n_2967;
wire n_1369;
wire n_2611;
wire n_1841;
wire n_1660;
wire n_1905;
wire n_2553;
wire n_3706;
wire n_3207;
wire n_2581;
wire n_2195;
wire n_2529;
wire n_3224;
wire n_2698;
wire n_1711;
wire n_1891;
wire n_1662;
wire n_1481;
wire n_2626;
wire n_3441;
wire n_3042;
wire n_1942;
wire n_1978;
wire n_1544;
wire n_2510;
wire n_3047;
wire n_3526;
wire n_2454;
wire n_2804;
wire n_3659;
wire n_2120;
wire n_2546;
wire n_1629;
wire n_1293;
wire n_2801;
wire n_3120;
wire n_1876;
wire n_1743;
wire n_3491;
wire n_1175;
wire n_2763;
wire n_1479;
wire n_1810;
wire n_2350;
wire n_2813;
wire n_2825;
wire n_1888;
wire n_2009;
wire n_3643;
wire n_2222;
wire n_1892;
wire n_3510;
wire n_2990;
wire n_1997;
wire n_2667;
wire n_1766;
wire n_3218;
wire n_1477;
wire n_3142;
wire n_1635;
wire n_1963;
wire n_2226;
wire n_1571;
wire n_2891;
wire n_3119;
wire n_1189;
wire n_2690;
wire n_3370;
wire n_2215;
wire n_3479;
wire n_1259;
wire n_1690;
wire n_1649;
wire n_3150;
wire n_2064;
wire n_2449;
wire n_1733;
wire n_1244;
wire n_3500;
wire n_2413;
wire n_1194;
wire n_1925;
wire n_3660;
wire n_2297;
wire n_1815;
wire n_3279;
wire n_2621;
wire n_1759;
wire n_1788;
wire n_2177;
wire n_2491;
wire n_1537;
wire n_2227;
wire n_2671;
wire n_1222;
wire n_1679;
wire n_2190;
wire n_3346;
wire n_1798;
wire n_2022;
wire n_1790;
wire n_2518;
wire n_2876;
wire n_1415;
wire n_2629;
wire n_2592;
wire n_3416;
wire n_3484;
wire n_3620;
wire n_1260;
wire n_1746;
wire n_1647;
wire n_2181;
wire n_2479;
wire n_2838;
wire n_1829;
wire n_1464;
wire n_3133;
wire n_3513;
wire n_2563;
wire n_1444;
wire n_1191;
wire n_2387;
wire n_2992;
wire n_1674;
wire n_3725;
wire n_1833;
wire n_3138;
wire n_1830;
wire n_2517;
wire n_2073;
wire n_1710;
wire n_1128;
wire n_2928;
wire n_3128;
wire n_1734;
wire n_3038;
wire n_2631;
wire n_1308;
wire n_2871;
wire n_2178;
wire n_3068;
wire n_1767;
wire n_3144;
wire n_2943;
wire n_2913;
wire n_2336;
wire n_3143;
wire n_3168;
wire n_1680;
wire n_1233;
wire n_3469;
wire n_2607;
wire n_1615;
wire n_1529;
wire n_2005;
wire n_1916;
wire n_3317;
wire n_1333;
wire n_2469;
wire n_1121;
wire n_2723;
wire n_3355;
wire n_2007;
wire n_3220;
wire n_2539;
wire n_3263;
wire n_2582;
wire n_1443;
wire n_1539;
wire n_2736;
wire n_2054;
wire n_1503;
wire n_1468;
wire n_1559;
wire n_1765;
wire n_3455;
wire n_1866;
wire n_3158;
wire n_1624;
wire n_3000;
wire n_3452;
wire n_1510;
wire n_1380;
wire n_1744;
wire n_2623;
wire n_1617;
wire n_1994;
wire n_1231;
wire n_1279;
wire n_1406;
wire n_3113;
wire n_3108;
wire n_3111;
wire n_2718;
wire n_1195;
wire n_1839;
wire n_1837;
wire n_2577;
wire n_1760;
wire n_2875;
wire n_1500;
wire n_2960;
wire n_1090;
wire n_2796;
wire n_3280;
wire n_2342;
wire n_2856;
wire n_3471;
wire n_1832;
wire n_1851;
wire n_3205;
wire n_2046;
wire n_2848;
wire n_2741;
wire n_2937;
wire n_3666;
wire n_3003;
wire n_3610;
wire n_1933;
wire n_2290;
wire n_1656;
wire n_3564;
wire n_3288;
wire n_1158;
wire n_3095;
wire n_2045;
wire n_3369;
wire n_1509;
wire n_1874;
wire n_2040;
wire n_2060;
wire n_3199;
wire n_2613;
wire n_1987;
wire n_2805;
wire n_3667;
wire n_1145;
wire n_3457;
wire n_1678;
wire n_1153;
wire n_2145;
wire n_1639;
wire n_1306;
wire n_3703;
wire n_1068;
wire n_3030;
wire n_3558;
wire n_1871;
wire n_2580;
wire n_3630;
wire n_2545;
wire n_2787;
wire n_3685;
wire n_2914;
wire n_1964;
wire n_2869;
wire n_1163;
wire n_3271;
wire n_2039;
wire n_1207;
wire n_2412;
wire n_2406;
wire n_3623;
wire n_2846;
wire n_1781;
wire n_2084;
wire n_2925;
wire n_3648;
wire n_2035;
wire n_2061;
wire n_3555;
wire n_3579;
wire n_3075;
wire n_3173;
wire n_2378;
wire n_2509;
wire n_1740;
wire n_3236;
wire n_2398;
wire n_1362;
wire n_2857;
wire n_1586;
wire n_2459;
wire n_3031;
wire n_3396;
wire n_3701;
wire n_1445;
wire n_3516;
wire n_1492;
wire n_2155;
wire n_2516;
wire n_1923;
wire n_1773;
wire n_3243;
wire n_1169;
wire n_1596;
wire n_1692;
wire n_2666;
wire n_2982;
wire n_3385;
wire n_2481;
wire n_2947;
wire n_3545;
wire n_2171;
wire n_2768;
wire n_2116;
wire n_2314;
wire n_1434;
wire n_2507;
wire n_1474;
wire n_1665;
wire n_1269;
wire n_2420;
wire n_2900;
wire n_1095;
wire n_3343;
wire n_3515;
wire n_1828;
wire n_1614;
wire n_2886;
wire n_2093;
wire n_1079;
wire n_2473;
wire n_1208;
wire n_2320;
wire n_2038;
wire n_2339;
wire n_3287;
wire n_2137;
wire n_3378;
wire n_1431;
wire n_2583;
wire n_1593;
wire n_3426;
wire n_3454;
wire n_2299;
wire n_2540;
wire n_2873;
wire n_3410;
wire n_2087;
wire n_1640;
wire n_2162;
wire n_1732;
wire n_2847;
wire n_1148;
wire n_2051;
wire n_2029;
wire n_3221;
wire n_2168;
wire n_2790;
wire n_1609;
wire n_3629;
wire n_3021;
wire n_1989;
wire n_2359;
wire n_2941;
wire n_3674;
wire n_1887;
wire n_3502;
wire n_2523;
wire n_1383;
wire n_3098;
wire n_1073;
wire n_2346;
wire n_2457;
wire n_2312;
wire n_3475;
wire n_1215;
wire n_3015;
wire n_1171;
wire n_1578;
wire n_1920;
wire n_1065;
wire n_1592;
wire n_2536;
wire n_1336;
wire n_2882;
wire n_3719;
wire n_1721;
wire n_1959;
wire n_1758;
wire n_2338;
wire n_3681;
wire n_2952;
wire n_2737;
wire n_1574;
wire n_3672;
wire n_2399;
wire n_3058;
wire n_2812;
wire n_2048;
wire n_3197;
wire n_3109;
wire n_3607;
wire n_2355;
wire n_2133;
wire n_1921;
wire n_2721;
wire n_1309;
wire n_1878;
wire n_1426;
wire n_2585;
wire n_3505;
wire n_3002;
wire n_1800;
wire n_1548;
wire n_2725;
wire n_1421;
wire n_2571;
wire n_1286;
wire n_3730;
wire n_1177;
wire n_3276;
wire n_1355;
wire n_2565;
wire n_1159;
wire n_2124;
wire n_3001;
wire n_2081;
wire n_3149;
wire n_1119;
wire n_2261;
wire n_1240;
wire n_2156;
wire n_1820;
wire n_2729;
wire n_3268;
wire n_3597;
wire n_2418;
wire n_2519;
wire n_3354;
wire n_2724;
wire n_1612;
wire n_2179;
wire n_1416;
wire n_2077;
wire n_2897;
wire n_3614;
wire n_2909;
wire n_1724;
wire n_2111;
wire n_2521;
wire n_3301;
wire n_3466;
wire n_3458;
wire n_1237;
wire n_1420;
wire n_3185;
wire n_1132;
wire n_3330;
wire n_1366;
wire n_1300;
wire n_2595;
wire n_1127;
wire n_3248;
wire n_2277;
wire n_2477;
wire n_3523;
wire n_1785;
wire n_1568;
wire n_2829;
wire n_3411;
wire n_2110;
wire n_1270;
wire n_1664;
wire n_3200;
wire n_1486;
wire n_3586;
wire n_1332;
wire n_3519;
wire n_2231;
wire n_1390;
wire n_2017;
wire n_2474;
wire n_2879;
wire n_2604;
wire n_2090;
wire n_3374;
wire n_3153;
wire n_3045;
wire n_1870;
wire n_2367;
wire n_1591;
wire n_2033;
wire n_3453;
wire n_1682;
wire n_1980;
wire n_2390;
wire n_2628;
wire n_1249;
wire n_3399;
wire n_2896;
wire n_1111;
wire n_3213;
wire n_1365;
wire n_1927;
wire n_3065;
wire n_2132;
wire n_1349;
wire n_1093;
wire n_2400;
wire n_3645;
wire n_1265;
wire n_3223;
wire n_1909;
wire n_3077;
wire n_2681;
wire n_1562;
wire n_3103;
wire n_3474;
wire n_3675;
wire n_2255;
wire n_2424;
wire n_2272;
wire n_1140;
wire n_1651;
wire n_1965;
wire n_3387;
wire n_1902;
wire n_2151;
wire n_1941;
wire n_2106;
wire n_2775;
wire n_2716;
wire n_1913;
wire n_2878;
wire n_1823;
wire n_3679;
wire n_2464;
wire n_3422;
wire n_1101;
wire n_2831;
wire n_1106;
wire n_1456;
wire n_3557;
wire n_2230;
wire n_3498;
wire n_2015;
wire n_2365;
wire n_1875;
wire n_1982;
wire n_1304;
wire n_2803;
wire n_1324;
wire n_2851;
wire n_3707;
wire n_3189;
wire n_1846;
wire n_3037;
wire n_2066;
wire n_1885;
wire n_1455;
wire n_3429;
wire n_1903;
wire n_2490;
wire n_1407;
wire n_2452;
wire n_1551;
wire n_3154;
wire n_3229;
wire n_2849;
wire n_1805;
wire n_2176;
wire n_2204;
wire n_2905;
wire n_1816;
wire n_3692;
wire n_3566;
wire n_1217;
wire n_2220;
wire n_2455;
wire n_1849;
wire n_2410;
wire n_1131;
wire n_1084;
wire n_1961;
wire n_1935;
wire n_2922;
wire n_1430;
wire n_3275;
wire n_3499;
wire n_2645;
wire n_2467;
wire n_3366;
wire n_2727;
wire n_1094;
wire n_1354;
wire n_1534;
wire n_2288;
wire n_3421;
wire n_1351;
wire n_2240;
wire n_2696;
wire n_1205;
wire n_2436;
wire n_1209;
wire n_3029;
wire n_1552;
wire n_2508;
wire n_3242;
wire n_3592;
wire n_3618;
wire n_3525;
wire n_2593;
wire n_3486;
wire n_1435;
wire n_3394;
wire n_3683;
wire n_2416;
wire n_2405;
wire n_3642;
wire n_3286;
wire n_2088;
wire n_2953;
wire n_1645;
wire n_2461;
wire n_1327;
wire n_2858;
wire n_2243;
wire n_1684;
wire n_2658;
wire n_3590;
wire n_1717;
wire n_2895;
wire n_1795;
wire n_2128;
wire n_2578;
wire n_3097;
wire n_3483;
wire n_1821;
wire n_2929;
wire n_3424;
wire n_3478;
wire n_1381;
wire n_2555;
wire n_2662;
wire n_2740;
wire n_1611;
wire n_2368;
wire n_3388;
wire n_2656;
wire n_1080;
wire n_2301;
wire n_1274;
wire n_3583;
wire n_2890;
wire n_3560;
wire n_3059;
wire n_3524;
wire n_2554;
wire n_3465;
wire n_1316;
wire n_1708;
wire n_2419;
wire n_3215;
wire n_1438;
wire n_3698;
wire n_1082;
wire n_1840;
wire n_1630;
wire n_2122;
wire n_2512;
wire n_3589;
wire n_1436;
wire n_3549;
wire n_1691;
wire n_2786;
wire n_2534;
wire n_2092;
wire n_3171;
wire n_1229;
wire n_1437;
wire n_2075;
wire n_3658;
wire n_3449;
wire n_1092;
wire n_2694;
wire n_1776;
wire n_3559;
wire n_2198;
wire n_2610;
wire n_2661;
wire n_2572;
wire n_2989;
wire n_2281;
wire n_2131;
wire n_2789;
wire n_3026;
wire n_2216;
wire n_3020;
wire n_3677;
wire n_1757;
wire n_1897;
wire n_1919;
wire n_1424;
wire n_3462;
wire n_3588;
wire n_2933;
wire n_2308;
wire n_3468;
wire n_1893;
wire n_2910;
wire n_3419;
wire n_1290;
wire n_1123;
wire n_1467;
wire n_2053;
wire n_2163;
wire n_2328;
wire n_1958;
wire n_2254;
wire n_1252;
wire n_1382;
wire n_3546;
wire n_1206;
wire n_2647;
wire n_3160;
wire n_1311;
wire n_2191;
wire n_2864;
wire n_2969;
wire n_3195;
wire n_1519;
wire n_3190;
wire n_2428;
wire n_1553;
wire n_3678;
wire n_2664;
wire n_1811;
wire n_2443;
wire n_2624;
wire n_3012;
wire n_3456;
wire n_1346;
wire n_3053;
wire n_1299;
wire n_3244;
wire n_2158;
wire n_1808;
wire n_3290;
wire n_1060;
wire n_1141;
wire n_2266;
wire n_3130;
wire n_2465;
wire n_2824;
wire n_3033;
wire n_2650;
wire n_3298;
wire n_3548;
wire n_2440;
wire n_1699;
wire n_1386;
wire n_3334;
wire n_1442;
wire n_2923;
wire n_3665;
wire n_3494;
wire n_2541;
wire n_1139;
wire n_2731;
wire n_3264;
wire n_2333;
wire n_2916;
wire n_3166;
wire n_1432;
wire n_1357;
wire n_2125;
wire n_1632;
wire n_3110;
wire n_2998;
wire n_1085;
wire n_1066;
wire n_2402;
wire n_1157;
wire n_3073;
wire n_2403;
wire n_1954;
wire n_2265;
wire n_3162;
wire n_1608;
wire n_1844;
wire n_2760;
wire n_2792;
wire n_3554;
wire n_3377;
wire n_2870;
wire n_1305;
wire n_3178;
wire n_1826;
wire n_1112;
wire n_3134;
wire n_2304;
wire n_2999;
wire n_1283;
wire n_1644;
wire n_2334;
wire n_2637;
wire n_3695;
wire n_1974;
wire n_2463;
wire n_2086;
wire n_3537;
wire n_2289;
wire n_3080;
wire n_3051;
wire n_1343;
wire n_2701;
wire n_2783;
wire n_2263;
wire n_3362;
wire n_2881;
wire n_1631;
wire n_1203;
wire n_3282;
wire n_2472;
wire n_1763;
wire n_2341;
wire n_3105;
wire n_3231;
wire n_1966;
wire n_3632;
wire n_1768;
wire n_2294;
wire n_1179;
wire n_2475;
wire n_2733;
wire n_1719;
wire n_2993;
wire n_1288;
wire n_2785;
wire n_2556;
wire n_2269;
wire n_2732;
wire n_3569;
wire n_2309;
wire n_2415;
wire n_2948;
wire n_3299;
wire n_3041;
wire n_3274;
wire n_2646;
wire n_1560;
wire n_3715;
wire n_1605;
wire n_2236;
wire n_1228;
wire n_2816;
wire n_2123;
wire n_3209;
wire n_3504;
wire n_2037;
wire n_2685;
wire n_3040;
wire n_1953;
wire n_1938;
wire n_1200;
wire n_2499;
wire n_1911;
wire n_3616;
wire n_2460;
wire n_3568;
wire n_3664;
wire n_2589;
wire n_3203;
wire n_1363;
wire n_1668;
wire n_1301;
wire n_1185;
wire n_2903;
wire n_3417;
wire n_3482;
wire n_1967;
wire n_1143;
wire n_1579;
wire n_2233;
wire n_3717;
wire n_1329;
wire n_2743;
wire n_2675;
wire n_3255;
wire n_1312;
wire n_1439;
wire n_2827;
wire n_1688;
wire n_3052;
wire n_2997;
wire n_3327;
wire n_1504;
wire n_3326;
wire n_3572;
wire n_3067;
wire n_1932;
wire n_3375;
wire n_2755;
wire n_3734;
wire n_3237;
wire n_2082;
wire n_1992;
wire n_2429;
wire n_1643;
wire n_1983;
wire n_3167;
wire n_3400;
wire n_1594;
wire n_1400;
wire n_1342;
wire n_1214;
wire n_3423;
wire n_2362;
wire n_2609;
wire n_1793;
wire n_3382;
wire n_1976;
wire n_2223;
wire n_3044;
wire n_3574;
wire n_3529;
wire n_2169;
wire n_1804;
wire n_1147;
wire n_1977;
wire n_1557;
wire n_2153;
wire n_2468;
wire n_1610;
wire n_1077;
wire n_1422;
wire n_3196;
wire n_3078;
wire n_2533;
wire n_2364;
wire n_3492;
wire n_3094;
wire n_2310;
wire n_2780;
wire n_2287;
wire n_2860;
wire n_3316;
wire n_2291;
wire n_3099;
wire n_3704;
wire n_2596;
wire n_1636;
wire n_2056;
wire n_3253;
wire n_1730;
wire n_3601;
wire n_3603;
wire n_2280;
wire n_2192;
wire n_3633;
wire n_3363;
wire n_1373;
wire n_1350;
wire n_1511;
wire n_1865;
wire n_2973;
wire n_1470;
wire n_1096;
wire n_2094;
wire n_2670;
wire n_1575;
wire n_1697;
wire n_1735;
wire n_2318;
wire n_2393;
wire n_3689;
wire n_2020;
wire n_1646;
wire n_2502;
wire n_2504;
wire n_1307;
wire n_1881;
wire n_2974;
wire n_2749;
wire n_2043;
wire n_2901;
wire n_1940;
wire n_2707;
wire n_2793;
wire n_2751;
wire n_3372;
wire n_3451;
wire n_2971;
wire n_3442;
wire n_1549;
wire n_1934;
wire n_2311;
wire n_1201;
wire n_1114;
wire n_3240;
wire n_2025;
wire n_1616;
wire n_1446;
wire n_2285;
wire n_3147;
wire n_2758;
wire n_1458;
wire n_2471;
wire n_1176;
wire n_1472;
wire n_2298;
wire n_1807;
wire n_1149;
wire n_2618;
wire n_1671;
wire n_2559;
wire n_3230;
wire n_1062;
wire n_3342;
wire n_2303;
wire n_1824;
wire n_1917;
wire n_2295;
wire n_1219;
wire n_3386;
wire n_3708;
wire n_1204;
wire n_2840;
wire n_3729;
wire n_2810;
wire n_2325;
wire n_2747;
wire n_2446;
wire n_3488;
wire n_1814;
wire n_2822;
wire n_1848;
wire n_1928;
wire n_2126;
wire n_2893;
wire n_3636;
wire n_1188;
wire n_2588;
wire n_2962;
wire n_1722;
wire n_2441;
wire n_1802;
wire n_3083;
wire n_2600;
wire n_2795;
wire n_1638;
wire n_1786;
wire n_2981;
wire n_2002;
wire n_2282;
wire n_3608;
wire n_2800;
wire n_3712;
wire n_2371;
wire n_2935;
wire n_3233;
wire n_3380;
wire n_3177;
wire n_2098;
wire n_1296;
wire n_2627;
wire n_3409;
wire n_3460;
wire n_2352;
wire n_3538;
wire n_1413;
wire n_2207;
wire n_2080;
wire n_2377;
wire n_2619;
wire n_2340;
wire n_3085;
wire n_2444;
wire n_2068;
wire n_3552;
wire n_1110;
wire n_1655;
wire n_2641;
wire n_3198;
wire n_1895;
wire n_3123;
wire n_3684;
wire n_3137;
wire n_2574;
wire n_1134;
wire n_1358;
wire n_3697;
wire n_2361;
wire n_1088;
wire n_1173;
wire n_3393;
wire n_1603;
wire n_1232;
wire n_2638;
wire n_1401;
wire n_3520;
wire n_2492;
wire n_1998;
wire n_1105;
wire n_1338;
wire n_2016;
wire n_1522;
wire n_2949;
wire n_1687;
wire n_1637;
wire n_2034;
wire n_1419;
wire n_2711;
wire n_1653;
wire n_2270;
wire n_1506;
wire n_3206;
wire n_2653;
wire n_3578;
wire n_2867;
wire n_2496;
wire n_1886;
wire n_1389;
wire n_1894;
wire n_1908;
wire n_1256;
wire n_1702;
wire n_2259;
wire n_2794;
wire n_1465;
wire n_3145;
wire n_3124;
wire n_1122;
wire n_3192;
wire n_2608;
wire n_2657;
wire n_2995;
wire n_1375;
wire n_2494;
wire n_3547;
wire n_2649;
wire n_1102;
wire n_3727;
wire n_2852;
wire n_2392;
wire n_3459;
wire n_3093;
wire n_1843;
wire n_1499;
wire n_3061;
wire n_3155;
wire n_1187;
wire n_3517;
wire n_2633;
wire n_1441;
wire n_3100;
wire n_2522;
wire n_2435;
wire n_1597;
wire n_1392;
wire n_1929;
wire n_2807;
wire n_1164;
wire n_1659;
wire n_1834;
wire n_2097;
wire n_2542;
wire n_2313;
wire n_3324;
wire n_1174;
wire n_2431;
wire n_3356;
wire n_2835;
wire n_2558;
wire n_1371;
wire n_1303;
wire n_2206;
wire n_2063;
wire n_3182;
wire n_1572;
wire n_1968;
wire n_3269;
wire n_2564;
wire n_2252;
wire n_1516;
wire n_1190;
wire n_3506;
wire n_1736;
wire n_3605;
wire n_1685;
wire n_2409;
wire n_3450;
wire n_1714;
wire n_1116;
wire n_2000;
wire n_1661;
wire n_3402;
wire n_1212;
wire n_2074;
wire n_1541;
wire n_2576;
wire n_3565;
wire n_3174;
wire n_2575;
wire n_2988;
wire n_3390;
wire n_1573;
wire n_1731;
wire n_1453;
wire n_2217;
wire n_2373;
wire n_1970;
wire n_1713;
wire n_1183;
wire n_3398;
wire n_2307;
wire n_2766;
wire n_1658;
wire n_1253;
wire n_2722;
wire n_1737;
wire n_2201;
wire n_2745;
wire n_2117;
wire n_3408;
wire n_1904;
wire n_2640;
wire n_1993;
wire n_1628;
wire n_2493;
wire n_2205;
wire n_3432;
wire n_1777;
wire n_1335;
wire n_1514;
wire n_1957;
wire n_1345;
wire n_1133;
wire n_1771;
wire n_1912;
wire n_3401;
wire n_1899;
wire n_3226;
wire n_1410;
wire n_3090;
wire n_2067;
wire n_1168;
wire n_2219;
wire n_2437;
wire n_2885;
wire n_3533;
wire n_2877;
wire n_3318;
wire n_2148;
wire n_2445;
wire n_1427;
wire n_2779;
wire n_3485;
wire n_1584;
wire n_1726;
wire n_1835;
wire n_3035;
wire n_3654;
wire n_1440;
wire n_2164;
wire n_1988;
wire n_3333;
wire n_2115;
wire n_1853;
wire n_1356;
wire n_2845;
wire n_1787;
wire n_2634;
wire n_2232;
wire n_3034;
wire n_2212;
wire n_2602;
wire n_1657;
wire n_1475;
wire n_1302;
wire n_1774;
wire n_1725;
wire n_1136;
wire n_1313;
wire n_1491;
wire n_2811;
wire n_1496;
wire n_3348;
wire n_1125;
wire n_2547;
wire n_3014;
wire n_3639;
wire n_1812;
wire n_2501;
wire n_3079;
wire n_1915;
wire n_1109;
wire n_2532;
wire n_1310;
wire n_2605;
wire n_3358;
wire n_2121;
wire n_1803;
wire n_3308;
wire n_2665;
wire n_1991;
wire n_1399;
wire n_1543;
wire n_1979;
wire n_1533;
wire n_2224;
wire n_3368;
wire n_2924;
wire n_3467;
wire n_2484;
wire n_3530;
wire n_1930;
wire n_1955;
wire n_3731;
wire n_2765;
wire n_3329;
wire n_2994;
wire n_1067;
wire n_2946;
wire n_1720;
wire n_2830;
wire n_2401;
wire n_3135;
wire n_3657;
wire n_2003;
wire n_1457;
wire n_2692;
wire n_3573;
wire n_3148;
wire n_2354;
wire n_2246;
wire n_2008;
wire n_1117;
wire n_2264;
wire n_2754;
wire n_3534;
wire n_1742;
wire n_1480;
wire n_1482;
wire n_1213;
wire n_2489;
wire n_1266;
wire n_3438;
wire n_2012;
wire n_1291;
wire n_3381;
wire n_3503;
wire n_1297;
wire n_1753;
wire n_2283;
wire n_2866;
wire n_3278;
wire n_1782;
wire n_2245;
wire n_3561;
wire n_1155;
wire n_1418;
wire n_1972;
wire n_1689;
wire n_1524;
wire n_1485;
wire n_2806;
wire n_1184;
wire n_2184;
wire n_1855;
wire n_2425;
wire n_2917;
wire n_2965;
wire n_3536;
wire n_3661;
wire n_3635;
wire n_3217;
wire n_3404;
wire n_3425;
wire n_1703;
wire n_3312;
wire n_1352;
wire n_2926;
wire n_2197;
wire n_2199;
wire n_3540;
wire n_1650;
wire n_3670;
wire n_1144;
wire n_1137;
wire n_1570;
wire n_2814;
wire n_3046;
wire n_1170;
wire n_2213;
wire n_2023;
wire n_3249;
wire n_3211;
wire n_3285;
wire n_2351;
wire n_2211;
wire n_2095;
wire n_3121;
wire n_2103;
wire n_2160;
wire n_3337;
wire n_2228;
wire n_2527;
wire n_1602;
wire n_2498;
wire n_1178;
wire n_1461;
wire n_2697;
wire n_3074;
wire n_3204;
wire n_2421;
wire n_2286;
wire n_2902;
wire n_1999;
wire n_2372;
wire n_2065;
wire n_2136;
wire n_3673;
wire n_2480;
wire n_1372;
wire n_2861;
wire n_2630;
wire n_1273;
wire n_1822;
wire n_3397;
wire n_2363;
wire n_2430;
wire n_1081;
wire n_2549;
wire n_2705;
wire n_3005;
wire n_2332;
wire n_1235;
wire n_1115;
wire n_2433;
wire n_3293;
wire n_3129;
wire n_1282;
wire n_1318;
wire n_1783;
wire n_2977;
wire n_3606;
wire n_2601;
wire n_3043;
wire n_2375;
wire n_2550;
wire n_1454;
wire n_3723;
wire n_1227;
wire n_1531;
wire n_1334;
wire n_1907;
wire n_3600;
wire n_2686;
wire n_2528;
wire n_2344;
wire n_1388;
wire n_1417;
wire n_1295;
wire n_2836;
wire n_2316;
wire n_1985;
wire n_3055;
wire n_1898;
wire n_2107;
wire n_3294;
wire n_3219;
wire n_3711;
wire n_3315;
wire n_2906;
wire n_1625;
wire n_2130;
wire n_3415;
wire n_2187;
wire n_2284;
wire n_2817;
wire n_3172;
wire n_3139;
wire n_2773;
wire n_3239;
wire n_3292;
wire n_2598;
wire n_1762;
wire n_3365;
wire n_3476;
wire n_3686;
wire n_1452;
wire n_2687;
wire n_3023;
wire n_3553;
wire n_1120;
wire n_1791;
wire n_1890;
wire n_1747;
wire n_2850;
wire n_1683;
wire n_1817;
wire n_1944;
wire n_1530;
wire n_1497;
wire n_2654;
wire n_3431;
wire n_3104;
wire n_3169;
wire n_3151;
wire n_3131;
wire n_2078;
wire n_1409;
wire n_1326;
wire n_3070;
wire n_3284;
wire n_3647;
wire n_3176;
wire n_2884;
wire n_1268;
wire n_2996;
wire n_2819;
wire n_3126;
wire n_1981;
wire n_2186;
wire n_1320;
wire n_1663;
wire n_1718;
wire n_3700;
wire n_3609;
wire n_2315;
wire n_3228;
wire n_1317;
wire n_1518;
wire n_1715;
wire n_2102;
wire n_3581;
wire n_2562;
wire n_1281;
wire n_1952;
wire n_1192;
wire n_2221;
wire n_3576;
wire n_1063;
wire n_3720;
wire n_1889;
wire n_1792;
wire n_1564;
wire n_1868;
wire n_1613;
wire n_1489;
wire n_1922;
wire n_2966;
wire n_1376;
wire n_2560;
wire n_2326;
wire n_1569;
wire n_2188;
wire n_3495;
wire n_2348;
wire n_2422;
wire n_2239;
wire n_2950;
wire n_1429;
wire n_1238;
wire n_2448;
wire n_3140;
wire n_3170;
wire n_3724;
wire n_2104;
wire n_2748;
wire n_3311;
wire n_2057;
wire n_3272;
wire n_3011;
wire n_1772;
wire n_1476;
wire n_1108;
wire n_2898;
wire n_2717;
wire n_2818;
wire n_1100;
wire n_3646;
wire n_1861;
wire n_2129;
wire n_1395;
wire n_3345;
wire n_3584;
wire n_1425;
wire n_1901;
wire n_3069;
wire n_1900;
wire n_1620;
wire n_3032;
wire n_3628;
wire n_2889;
wire n_3691;
wire n_1867;
wire n_1330;
wire n_1945;
wire n_2772;
wire n_3018;
wire n_1675;
wire n_3072;
wire n_1924;
wire n_2573;
wire n_3084;
wire n_3081;
wire n_3313;
wire n_1727;
wire n_2710;
wire n_1554;
wire n_2939;
wire n_1745;
wire n_2735;
wire n_2497;
wire n_2006;
wire n_3412;
wire n_2844;
wire n_1995;
wire n_2411;
wire n_2138;
wire n_1618;
wire n_2260;
wire n_2343;
wire n_1813;
wire n_2447;
wire n_3439;
wire n_2014;
wire n_3056;
wire n_1221;
wire n_2345;
wire n_2986;
wire n_1172;
wire n_2535;
wire n_1341;
wire n_2726;
wire n_2774;
wire n_3295;
wire n_1641;
wire n_1361;
wire n_3184;
wire n_2382;
wire n_1707;
wire n_3062;
wire n_3161;
wire n_2317;
wire n_3289;
wire n_2799;
wire n_2172;
wire n_1973;
wire n_1083;
wire n_1142;
wire n_2376;
wire n_2488;
wire n_1129;
wire n_2579;
wire n_3477;
wire n_3017;
wire n_3626;
wire n_2476;
wire n_1770;
wire n_2781;
wire n_2456;
wire n_2250;
wire n_2678;
wire n_1756;
wire n_2778;
wire n_1716;
wire n_2788;
wire n_2872;
wire n_1225;
wire n_2984;
wire n_1520;
wire n_2451;
wire n_2887;
wire n_3364;
wire n_1287;
wire n_1262;
wire n_2691;
wire n_1873;
wire n_1411;
wire n_3201;
wire n_3054;
wire n_1962;
wire n_1577;
wire n_2423;
wire n_3671;
wire n_1087;
wire n_3472;
wire n_2526;
wire n_2854;
wire n_1701;
wire n_3344;
wire n_2194;
wire n_1550;
wire n_2874;
wire n_2764;
wire n_2703;
wire n_1498;
wire n_2167;
wire n_3302;
wire n_3235;
wire n_1223;
wire n_1272;
wire n_2680;
wire n_3391;
wire n_1567;
wire n_2567;
wire n_3543;
wire n_1247;
wire n_2709;
wire n_3102;
wire n_3122;
wire n_1648;
wire n_1536;
wire n_3050;
wire n_3265;
wire n_1857;
wire n_1344;
wire n_2041;
wire n_3627;
wire n_1246;
wire n_1478;
wire n_1339;
wire n_1797;
wire n_1769;
wire n_2957;
wire n_3551;
wire n_1210;
wire n_3518;
wire n_2964;
wire n_1364;
wire n_2956;
wire n_2357;
wire n_3733;
wire n_2183;
wire n_2673;
wire n_2742;
wire n_3314;
wire n_2360;
wire n_3254;
wire n_2292;
wire n_1250;
wire n_2173;
wire n_3722;
wire n_1842;
wire n_2442;
wire n_3309;
wire n_1367;
wire n_1943;
wire n_3634;
wire n_1460;
wire n_2018;
wire n_3464;
wire n_3260;
wire n_1555;
wire n_3117;
wire n_2834;
wire n_3245;
wire n_3357;
wire n_2531;
wire n_1589;
wire n_3428;
wire n_2961;
wire n_1086;
wire n_2570;
wire n_2702;
wire n_1858;
wire n_3351;
wire n_1619;
wire n_3527;
wire n_2815;
wire n_2119;
wire n_1502;
wire n_2157;
wire n_2552;
wire n_1469;
wire n_1396;
wire n_2744;
wire n_1348;
wire n_2030;
wire n_2453;
wire n_1752;
wire n_1525;
wire n_2397;
wire n_2883;
wire n_3115;
wire n_3509;
wire n_3352;
wire n_2208;
wire n_3076;
wire n_1404;
wire n_3063;
wire n_3617;
wire n_2912;
wire n_1794;
wire n_3535;
wire n_2182;
wire n_1315;
wire n_2234;
wire n_1061;
wire n_3251;
wire n_1910;
wire n_1298;
wire n_2931;
wire n_1652;
wire n_2209;
wire n_2809;
wire n_2050;
wire n_1193;
wire n_2797;
wire n_1676;
wire n_1255;
wire n_1113;
wire n_3118;
wire n_3227;
wire n_3300;
wire n_2321;
wire n_3511;
wire n_1226;
wire n_1277;
wire n_3680;
wire n_2591;
wire n_3443;
wire n_2146;
wire n_3384;
wire n_3497;
wire n_1487;
wire n_1864;
wire n_3644;
wire n_1601;
wire n_3336;
wire n_2940;
wire n_3435;
wire n_3521;
wire n_3575;
wire n_1546;
wire n_3562;
wire n_2612;
wire n_1337;
wire n_1495;
wire n_1515;
wire n_2841;
wire n_3165;
wire n_1627;
wire n_2918;
wire n_3232;
wire n_3322;
wire n_3652;
wire n_1245;
wire n_2427;
wire n_2438;
wire n_2505;
wire n_1673;
wire n_2832;
wire n_1321;
wire n_1975;
wire n_2296;
wire n_2070;
wire n_1937;
wire n_2112;
wire n_3250;
wire n_1739;
wire n_3181;
wire n_2958;
wire n_2278;
wire n_2594;
wire n_3114;
wire n_3125;
wire n_2394;
wire n_3234;
wire n_1914;
wire n_3612;
wire n_2954;
wire n_2135;
wire n_2335;
wire n_2904;
wire n_3493;
wire n_2381;
wire n_3303;
wire n_1654;
wire n_3004;
wire n_3323;
wire n_2569;
wire n_3112;
wire n_2349;
wire n_1103;
wire n_3132;
wire n_3556;
wire n_1379;
wire n_2734;
wire n_2196;
wire n_3591;
wire n_3024;
wire n_2170;
wire n_1076;
wire n_2823;
wire n_1091;
wire n_1408;
wire n_3512;
wire n_1761;
wire n_3238;
wire n_3210;
wire n_3175;
wire n_3522;
wire n_2036;
wire n_1325;
wire n_3267;
wire n_1595;
wire n_2161;
wire n_2404;
wire n_2083;
wire n_3281;
wire n_3307;
wire n_1606;
wire n_2503;
wire n_1220;
wire n_1694;
wire n_1540;
wire n_3266;
wire n_2485;
wire n_1956;
wire n_1936;
wire n_1642;
wire n_2279;
wire n_3373;
wire n_2655;
wire n_2027;
wire n_2642;
wire n_1130;
wire n_2500;
wire n_2366;
wire n_1918;
wire n_1526;
wire n_3726;
wire n_2210;
wire n_3247;
wire n_1604;
wire n_1275;
wire n_2513;
wire n_2525;
wire n_3091;
wire n_2695;
wire n_1764;
wire n_3480;
wire n_2892;
wire n_3057;
wire n_3194;
wire n_3582;
wire n_3066;
wire n_2414;
wire n_2907;
wire n_1583;
wire n_2426;
wire n_2826;
wire n_3577;
wire n_3539;
wire n_1402;
wire n_2820;
wire n_3662;
wire n_2049;
wire n_2273;
wire n_2719;
wire n_1493;
wire n_1741;
wire n_2229;
wire n_1160;
wire n_1397;
wire n_1258;
wire n_1074;
wire n_3347;
wire n_2004;
wire n_3216;
wire n_1621;
wire n_2708;
wire n_2113;
wire n_2586;
wire n_3694;
wire n_1448;
wire n_2225;
wire n_3567;
wire n_3613;
wire n_1507;
wire n_1398;
wire n_2383;
wire n_1879;
wire n_1996;
wire n_3406;
wire n_3604;
wire n_3444;
wire n_1181;
wire n_1505;
wire n_1634;
wire n_1196;
wire n_2019;
wire n_1340;
wire n_2274;
wire n_2972;
wire n_1558;
wire n_3225;
wire n_3321;
wire n_2166;
wire n_2938;
wire n_3212;
wire n_3319;
wire n_1433;
wire n_3594;
wire n_1704;
wire n_2256;
wire n_3152;
wire n_3721;
wire n_3335;
wire n_1254;
wire n_3413;
wire n_2026;
wire n_1969;
wire n_1234;
wire n_2109;
wire n_2044;
wire n_1138;
wire n_1089;
wire n_2013;
wire n_1990;
wire n_2689;
wire n_2920;
wire n_3259;
wire n_1186;
wire n_2614;
wire n_2511;
wire n_1681;
wire n_2010;
wire n_2991;
wire n_3688;
wire n_3383;
wire n_2242;
wire n_2247;
wire n_2752;
wire n_2894;
wire n_3016;
wire n_1693;
wire n_3585;
wire n_2975;
wire n_3473;
wire n_2599;
wire n_2704;
wire n_2839;
wire n_3338;
wire n_1588;
wire n_1622;
wire n_2237;
wire n_3414;
wire n_3463;
wire n_3699;
wire n_1827;
wire n_1180;
wire n_3360;
wire n_2524;
wire n_1271;
wire n_3705;
wire n_2802;
wire n_1542;
wire n_1251;
wire n_3693;
wire n_3159;
wire n_2728;
wire n_2268;

INVx1_ASAP7_75t_L g1060 ( 
.A(n_894),
.Y(n_1060)
);

BUFx10_ASAP7_75t_L g1061 ( 
.A(n_573),
.Y(n_1061)
);

INVx1_ASAP7_75t_L g1062 ( 
.A(n_479),
.Y(n_1062)
);

CKINVDCx5p33_ASAP7_75t_R g1063 ( 
.A(n_994),
.Y(n_1063)
);

BUFx6f_ASAP7_75t_L g1064 ( 
.A(n_775),
.Y(n_1064)
);

CKINVDCx20_ASAP7_75t_R g1065 ( 
.A(n_890),
.Y(n_1065)
);

INVx1_ASAP7_75t_L g1066 ( 
.A(n_5),
.Y(n_1066)
);

INVx1_ASAP7_75t_L g1067 ( 
.A(n_620),
.Y(n_1067)
);

CKINVDCx5p33_ASAP7_75t_R g1068 ( 
.A(n_1056),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_957),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_804),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_920),
.Y(n_1071)
);

BUFx2_ASAP7_75t_L g1072 ( 
.A(n_1040),
.Y(n_1072)
);

INVx1_ASAP7_75t_L g1073 ( 
.A(n_162),
.Y(n_1073)
);

INVx1_ASAP7_75t_L g1074 ( 
.A(n_664),
.Y(n_1074)
);

INVx2_ASAP7_75t_L g1075 ( 
.A(n_1043),
.Y(n_1075)
);

CKINVDCx5p33_ASAP7_75t_R g1076 ( 
.A(n_735),
.Y(n_1076)
);

CKINVDCx20_ASAP7_75t_R g1077 ( 
.A(n_115),
.Y(n_1077)
);

INVx1_ASAP7_75t_L g1078 ( 
.A(n_654),
.Y(n_1078)
);

INVx1_ASAP7_75t_L g1079 ( 
.A(n_657),
.Y(n_1079)
);

BUFx6f_ASAP7_75t_L g1080 ( 
.A(n_237),
.Y(n_1080)
);

BUFx5_ASAP7_75t_L g1081 ( 
.A(n_649),
.Y(n_1081)
);

INVx1_ASAP7_75t_L g1082 ( 
.A(n_1022),
.Y(n_1082)
);

CKINVDCx5p33_ASAP7_75t_R g1083 ( 
.A(n_252),
.Y(n_1083)
);

INVx1_ASAP7_75t_L g1084 ( 
.A(n_178),
.Y(n_1084)
);

CKINVDCx5p33_ASAP7_75t_R g1085 ( 
.A(n_553),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_549),
.Y(n_1086)
);

CKINVDCx5p33_ASAP7_75t_R g1087 ( 
.A(n_190),
.Y(n_1087)
);

BUFx10_ASAP7_75t_L g1088 ( 
.A(n_309),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_672),
.Y(n_1089)
);

INVx1_ASAP7_75t_L g1090 ( 
.A(n_1049),
.Y(n_1090)
);

INVx2_ASAP7_75t_L g1091 ( 
.A(n_844),
.Y(n_1091)
);

INVx1_ASAP7_75t_L g1092 ( 
.A(n_653),
.Y(n_1092)
);

INVx1_ASAP7_75t_L g1093 ( 
.A(n_154),
.Y(n_1093)
);

INVx1_ASAP7_75t_L g1094 ( 
.A(n_743),
.Y(n_1094)
);

INVx1_ASAP7_75t_L g1095 ( 
.A(n_458),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_432),
.Y(n_1096)
);

INVx1_ASAP7_75t_L g1097 ( 
.A(n_794),
.Y(n_1097)
);

INVx1_ASAP7_75t_L g1098 ( 
.A(n_853),
.Y(n_1098)
);

INVx1_ASAP7_75t_L g1099 ( 
.A(n_689),
.Y(n_1099)
);

BUFx6f_ASAP7_75t_L g1100 ( 
.A(n_459),
.Y(n_1100)
);

BUFx6f_ASAP7_75t_L g1101 ( 
.A(n_556),
.Y(n_1101)
);

INVx1_ASAP7_75t_L g1102 ( 
.A(n_393),
.Y(n_1102)
);

INVx1_ASAP7_75t_L g1103 ( 
.A(n_391),
.Y(n_1103)
);

CKINVDCx5p33_ASAP7_75t_R g1104 ( 
.A(n_1014),
.Y(n_1104)
);

CKINVDCx5p33_ASAP7_75t_R g1105 ( 
.A(n_260),
.Y(n_1105)
);

INVx1_ASAP7_75t_L g1106 ( 
.A(n_108),
.Y(n_1106)
);

INVx1_ASAP7_75t_L g1107 ( 
.A(n_686),
.Y(n_1107)
);

INVx1_ASAP7_75t_L g1108 ( 
.A(n_392),
.Y(n_1108)
);

CKINVDCx5p33_ASAP7_75t_R g1109 ( 
.A(n_209),
.Y(n_1109)
);

CKINVDCx5p33_ASAP7_75t_R g1110 ( 
.A(n_696),
.Y(n_1110)
);

CKINVDCx5p33_ASAP7_75t_R g1111 ( 
.A(n_650),
.Y(n_1111)
);

CKINVDCx5p33_ASAP7_75t_R g1112 ( 
.A(n_749),
.Y(n_1112)
);

CKINVDCx20_ASAP7_75t_R g1113 ( 
.A(n_1051),
.Y(n_1113)
);

INVx1_ASAP7_75t_L g1114 ( 
.A(n_271),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_746),
.Y(n_1115)
);

INVx1_ASAP7_75t_L g1116 ( 
.A(n_15),
.Y(n_1116)
);

INVx1_ASAP7_75t_L g1117 ( 
.A(n_101),
.Y(n_1117)
);

BUFx3_ASAP7_75t_L g1118 ( 
.A(n_647),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_577),
.Y(n_1119)
);

CKINVDCx5p33_ASAP7_75t_R g1120 ( 
.A(n_684),
.Y(n_1120)
);

CKINVDCx5p33_ASAP7_75t_R g1121 ( 
.A(n_75),
.Y(n_1121)
);

CKINVDCx5p33_ASAP7_75t_R g1122 ( 
.A(n_212),
.Y(n_1122)
);

INVx1_ASAP7_75t_L g1123 ( 
.A(n_371),
.Y(n_1123)
);

BUFx2_ASAP7_75t_SL g1124 ( 
.A(n_610),
.Y(n_1124)
);

CKINVDCx20_ASAP7_75t_R g1125 ( 
.A(n_812),
.Y(n_1125)
);

CKINVDCx5p33_ASAP7_75t_R g1126 ( 
.A(n_786),
.Y(n_1126)
);

INVx1_ASAP7_75t_L g1127 ( 
.A(n_1041),
.Y(n_1127)
);

INVx2_ASAP7_75t_L g1128 ( 
.A(n_112),
.Y(n_1128)
);

INVx1_ASAP7_75t_L g1129 ( 
.A(n_1055),
.Y(n_1129)
);

CKINVDCx5p33_ASAP7_75t_R g1130 ( 
.A(n_425),
.Y(n_1130)
);

INVx1_ASAP7_75t_L g1131 ( 
.A(n_1050),
.Y(n_1131)
);

CKINVDCx5p33_ASAP7_75t_R g1132 ( 
.A(n_632),
.Y(n_1132)
);

CKINVDCx20_ASAP7_75t_R g1133 ( 
.A(n_578),
.Y(n_1133)
);

CKINVDCx5p33_ASAP7_75t_R g1134 ( 
.A(n_585),
.Y(n_1134)
);

CKINVDCx5p33_ASAP7_75t_R g1135 ( 
.A(n_1007),
.Y(n_1135)
);

INVx1_ASAP7_75t_L g1136 ( 
.A(n_441),
.Y(n_1136)
);

CKINVDCx5p33_ASAP7_75t_R g1137 ( 
.A(n_194),
.Y(n_1137)
);

INVx1_ASAP7_75t_L g1138 ( 
.A(n_49),
.Y(n_1138)
);

CKINVDCx5p33_ASAP7_75t_R g1139 ( 
.A(n_43),
.Y(n_1139)
);

INVx1_ASAP7_75t_L g1140 ( 
.A(n_607),
.Y(n_1140)
);

CKINVDCx5p33_ASAP7_75t_R g1141 ( 
.A(n_14),
.Y(n_1141)
);

CKINVDCx5p33_ASAP7_75t_R g1142 ( 
.A(n_576),
.Y(n_1142)
);

CKINVDCx5p33_ASAP7_75t_R g1143 ( 
.A(n_654),
.Y(n_1143)
);

INVx1_ASAP7_75t_L g1144 ( 
.A(n_1030),
.Y(n_1144)
);

INVx1_ASAP7_75t_L g1145 ( 
.A(n_502),
.Y(n_1145)
);

INVx1_ASAP7_75t_L g1146 ( 
.A(n_230),
.Y(n_1146)
);

INVx1_ASAP7_75t_L g1147 ( 
.A(n_1032),
.Y(n_1147)
);

CKINVDCx5p33_ASAP7_75t_R g1148 ( 
.A(n_377),
.Y(n_1148)
);

CKINVDCx5p33_ASAP7_75t_R g1149 ( 
.A(n_988),
.Y(n_1149)
);

CKINVDCx5p33_ASAP7_75t_R g1150 ( 
.A(n_638),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_477),
.Y(n_1151)
);

CKINVDCx5p33_ASAP7_75t_R g1152 ( 
.A(n_670),
.Y(n_1152)
);

CKINVDCx5p33_ASAP7_75t_R g1153 ( 
.A(n_924),
.Y(n_1153)
);

INVx2_ASAP7_75t_L g1154 ( 
.A(n_861),
.Y(n_1154)
);

BUFx3_ASAP7_75t_L g1155 ( 
.A(n_966),
.Y(n_1155)
);

CKINVDCx14_ASAP7_75t_R g1156 ( 
.A(n_699),
.Y(n_1156)
);

CKINVDCx5p33_ASAP7_75t_R g1157 ( 
.A(n_138),
.Y(n_1157)
);

INVx2_ASAP7_75t_L g1158 ( 
.A(n_616),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_277),
.Y(n_1159)
);

INVx1_ASAP7_75t_L g1160 ( 
.A(n_663),
.Y(n_1160)
);

CKINVDCx20_ASAP7_75t_R g1161 ( 
.A(n_965),
.Y(n_1161)
);

CKINVDCx5p33_ASAP7_75t_R g1162 ( 
.A(n_435),
.Y(n_1162)
);

CKINVDCx5p33_ASAP7_75t_R g1163 ( 
.A(n_876),
.Y(n_1163)
);

INVx2_ASAP7_75t_SL g1164 ( 
.A(n_1025),
.Y(n_1164)
);

HB1xp67_ASAP7_75t_L g1165 ( 
.A(n_578),
.Y(n_1165)
);

BUFx10_ASAP7_75t_L g1166 ( 
.A(n_729),
.Y(n_1166)
);

BUFx10_ASAP7_75t_L g1167 ( 
.A(n_1039),
.Y(n_1167)
);

CKINVDCx5p33_ASAP7_75t_R g1168 ( 
.A(n_382),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_1031),
.Y(n_1169)
);

CKINVDCx16_ASAP7_75t_R g1170 ( 
.A(n_534),
.Y(n_1170)
);

INVx2_ASAP7_75t_L g1171 ( 
.A(n_49),
.Y(n_1171)
);

INVx1_ASAP7_75t_L g1172 ( 
.A(n_549),
.Y(n_1172)
);

BUFx2_ASAP7_75t_L g1173 ( 
.A(n_146),
.Y(n_1173)
);

INVx1_ASAP7_75t_L g1174 ( 
.A(n_249),
.Y(n_1174)
);

CKINVDCx5p33_ASAP7_75t_R g1175 ( 
.A(n_1058),
.Y(n_1175)
);

CKINVDCx5p33_ASAP7_75t_R g1176 ( 
.A(n_850),
.Y(n_1176)
);

INVx4_ASAP7_75t_R g1177 ( 
.A(n_950),
.Y(n_1177)
);

CKINVDCx5p33_ASAP7_75t_R g1178 ( 
.A(n_198),
.Y(n_1178)
);

BUFx3_ASAP7_75t_L g1179 ( 
.A(n_93),
.Y(n_1179)
);

CKINVDCx5p33_ASAP7_75t_R g1180 ( 
.A(n_169),
.Y(n_1180)
);

BUFx2_ASAP7_75t_L g1181 ( 
.A(n_222),
.Y(n_1181)
);

CKINVDCx5p33_ASAP7_75t_R g1182 ( 
.A(n_1047),
.Y(n_1182)
);

CKINVDCx20_ASAP7_75t_R g1183 ( 
.A(n_126),
.Y(n_1183)
);

CKINVDCx5p33_ASAP7_75t_R g1184 ( 
.A(n_78),
.Y(n_1184)
);

CKINVDCx20_ASAP7_75t_R g1185 ( 
.A(n_641),
.Y(n_1185)
);

INVx1_ASAP7_75t_L g1186 ( 
.A(n_691),
.Y(n_1186)
);

CKINVDCx20_ASAP7_75t_R g1187 ( 
.A(n_579),
.Y(n_1187)
);

CKINVDCx5p33_ASAP7_75t_R g1188 ( 
.A(n_480),
.Y(n_1188)
);

CKINVDCx5p33_ASAP7_75t_R g1189 ( 
.A(n_1011),
.Y(n_1189)
);

CKINVDCx14_ASAP7_75t_R g1190 ( 
.A(n_262),
.Y(n_1190)
);

CKINVDCx5p33_ASAP7_75t_R g1191 ( 
.A(n_564),
.Y(n_1191)
);

CKINVDCx20_ASAP7_75t_R g1192 ( 
.A(n_839),
.Y(n_1192)
);

CKINVDCx20_ASAP7_75t_R g1193 ( 
.A(n_720),
.Y(n_1193)
);

CKINVDCx5p33_ASAP7_75t_R g1194 ( 
.A(n_637),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_673),
.Y(n_1195)
);

CKINVDCx5p33_ASAP7_75t_R g1196 ( 
.A(n_377),
.Y(n_1196)
);

CKINVDCx5p33_ASAP7_75t_R g1197 ( 
.A(n_433),
.Y(n_1197)
);

CKINVDCx5p33_ASAP7_75t_R g1198 ( 
.A(n_53),
.Y(n_1198)
);

CKINVDCx5p33_ASAP7_75t_R g1199 ( 
.A(n_789),
.Y(n_1199)
);

CKINVDCx5p33_ASAP7_75t_R g1200 ( 
.A(n_215),
.Y(n_1200)
);

CKINVDCx5p33_ASAP7_75t_R g1201 ( 
.A(n_177),
.Y(n_1201)
);

BUFx8_ASAP7_75t_SL g1202 ( 
.A(n_287),
.Y(n_1202)
);

CKINVDCx5p33_ASAP7_75t_R g1203 ( 
.A(n_508),
.Y(n_1203)
);

CKINVDCx5p33_ASAP7_75t_R g1204 ( 
.A(n_819),
.Y(n_1204)
);

CKINVDCx5p33_ASAP7_75t_R g1205 ( 
.A(n_1024),
.Y(n_1205)
);

INVx1_ASAP7_75t_L g1206 ( 
.A(n_656),
.Y(n_1206)
);

INVx1_ASAP7_75t_L g1207 ( 
.A(n_646),
.Y(n_1207)
);

INVx1_ASAP7_75t_L g1208 ( 
.A(n_39),
.Y(n_1208)
);

INVx1_ASAP7_75t_L g1209 ( 
.A(n_403),
.Y(n_1209)
);

INVx1_ASAP7_75t_L g1210 ( 
.A(n_657),
.Y(n_1210)
);

INVx1_ASAP7_75t_SL g1211 ( 
.A(n_921),
.Y(n_1211)
);

INVx1_ASAP7_75t_L g1212 ( 
.A(n_223),
.Y(n_1212)
);

INVx1_ASAP7_75t_L g1213 ( 
.A(n_455),
.Y(n_1213)
);

CKINVDCx5p33_ASAP7_75t_R g1214 ( 
.A(n_475),
.Y(n_1214)
);

INVx1_ASAP7_75t_L g1215 ( 
.A(n_754),
.Y(n_1215)
);

CKINVDCx5p33_ASAP7_75t_R g1216 ( 
.A(n_98),
.Y(n_1216)
);

INVx1_ASAP7_75t_L g1217 ( 
.A(n_621),
.Y(n_1217)
);

CKINVDCx5p33_ASAP7_75t_R g1218 ( 
.A(n_182),
.Y(n_1218)
);

INVx1_ASAP7_75t_L g1219 ( 
.A(n_655),
.Y(n_1219)
);

CKINVDCx5p33_ASAP7_75t_R g1220 ( 
.A(n_285),
.Y(n_1220)
);

INVx1_ASAP7_75t_L g1221 ( 
.A(n_1057),
.Y(n_1221)
);

INVx2_ASAP7_75t_L g1222 ( 
.A(n_398),
.Y(n_1222)
);

INVx1_ASAP7_75t_SL g1223 ( 
.A(n_1034),
.Y(n_1223)
);

CKINVDCx5p33_ASAP7_75t_R g1224 ( 
.A(n_1036),
.Y(n_1224)
);

INVx1_ASAP7_75t_L g1225 ( 
.A(n_117),
.Y(n_1225)
);

CKINVDCx20_ASAP7_75t_R g1226 ( 
.A(n_669),
.Y(n_1226)
);

BUFx2_ASAP7_75t_L g1227 ( 
.A(n_1016),
.Y(n_1227)
);

CKINVDCx5p33_ASAP7_75t_R g1228 ( 
.A(n_608),
.Y(n_1228)
);

CKINVDCx5p33_ASAP7_75t_R g1229 ( 
.A(n_721),
.Y(n_1229)
);

CKINVDCx5p33_ASAP7_75t_R g1230 ( 
.A(n_727),
.Y(n_1230)
);

CKINVDCx5p33_ASAP7_75t_R g1231 ( 
.A(n_590),
.Y(n_1231)
);

INVx2_ASAP7_75t_L g1232 ( 
.A(n_256),
.Y(n_1232)
);

CKINVDCx5p33_ASAP7_75t_R g1233 ( 
.A(n_38),
.Y(n_1233)
);

CKINVDCx5p33_ASAP7_75t_R g1234 ( 
.A(n_593),
.Y(n_1234)
);

INVx1_ASAP7_75t_L g1235 ( 
.A(n_608),
.Y(n_1235)
);

CKINVDCx5p33_ASAP7_75t_R g1236 ( 
.A(n_892),
.Y(n_1236)
);

BUFx6f_ASAP7_75t_L g1237 ( 
.A(n_37),
.Y(n_1237)
);

CKINVDCx5p33_ASAP7_75t_R g1238 ( 
.A(n_838),
.Y(n_1238)
);

CKINVDCx5p33_ASAP7_75t_R g1239 ( 
.A(n_931),
.Y(n_1239)
);

CKINVDCx5p33_ASAP7_75t_R g1240 ( 
.A(n_384),
.Y(n_1240)
);

CKINVDCx20_ASAP7_75t_R g1241 ( 
.A(n_177),
.Y(n_1241)
);

INVx1_ASAP7_75t_L g1242 ( 
.A(n_534),
.Y(n_1242)
);

INVx1_ASAP7_75t_L g1243 ( 
.A(n_410),
.Y(n_1243)
);

CKINVDCx5p33_ASAP7_75t_R g1244 ( 
.A(n_849),
.Y(n_1244)
);

CKINVDCx16_ASAP7_75t_R g1245 ( 
.A(n_633),
.Y(n_1245)
);

CKINVDCx5p33_ASAP7_75t_R g1246 ( 
.A(n_494),
.Y(n_1246)
);

CKINVDCx5p33_ASAP7_75t_R g1247 ( 
.A(n_387),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_688),
.Y(n_1248)
);

CKINVDCx5p33_ASAP7_75t_R g1249 ( 
.A(n_687),
.Y(n_1249)
);

CKINVDCx5p33_ASAP7_75t_R g1250 ( 
.A(n_643),
.Y(n_1250)
);

CKINVDCx20_ASAP7_75t_R g1251 ( 
.A(n_569),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_695),
.Y(n_1252)
);

CKINVDCx5p33_ASAP7_75t_R g1253 ( 
.A(n_648),
.Y(n_1253)
);

CKINVDCx5p33_ASAP7_75t_R g1254 ( 
.A(n_694),
.Y(n_1254)
);

CKINVDCx5p33_ASAP7_75t_R g1255 ( 
.A(n_87),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_813),
.Y(n_1256)
);

BUFx5_ASAP7_75t_L g1257 ( 
.A(n_22),
.Y(n_1257)
);

CKINVDCx5p33_ASAP7_75t_R g1258 ( 
.A(n_520),
.Y(n_1258)
);

CKINVDCx5p33_ASAP7_75t_R g1259 ( 
.A(n_705),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_313),
.Y(n_1260)
);

BUFx6f_ASAP7_75t_L g1261 ( 
.A(n_545),
.Y(n_1261)
);

CKINVDCx5p33_ASAP7_75t_R g1262 ( 
.A(n_579),
.Y(n_1262)
);

CKINVDCx5p33_ASAP7_75t_R g1263 ( 
.A(n_673),
.Y(n_1263)
);

INVx1_ASAP7_75t_L g1264 ( 
.A(n_1048),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_640),
.Y(n_1265)
);

INVx1_ASAP7_75t_L g1266 ( 
.A(n_1037),
.Y(n_1266)
);

CKINVDCx5p33_ASAP7_75t_R g1267 ( 
.A(n_708),
.Y(n_1267)
);

BUFx6f_ASAP7_75t_L g1268 ( 
.A(n_607),
.Y(n_1268)
);

CKINVDCx5p33_ASAP7_75t_R g1269 ( 
.A(n_575),
.Y(n_1269)
);

CKINVDCx5p33_ASAP7_75t_R g1270 ( 
.A(n_122),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_930),
.Y(n_1271)
);

INVx1_ASAP7_75t_L g1272 ( 
.A(n_830),
.Y(n_1272)
);

INVx1_ASAP7_75t_L g1273 ( 
.A(n_485),
.Y(n_1273)
);

BUFx10_ASAP7_75t_L g1274 ( 
.A(n_495),
.Y(n_1274)
);

INVx1_ASAP7_75t_L g1275 ( 
.A(n_61),
.Y(n_1275)
);

BUFx8_ASAP7_75t_SL g1276 ( 
.A(n_145),
.Y(n_1276)
);

CKINVDCx5p33_ASAP7_75t_R g1277 ( 
.A(n_327),
.Y(n_1277)
);

CKINVDCx5p33_ASAP7_75t_R g1278 ( 
.A(n_638),
.Y(n_1278)
);

BUFx3_ASAP7_75t_L g1279 ( 
.A(n_1023),
.Y(n_1279)
);

CKINVDCx20_ASAP7_75t_R g1280 ( 
.A(n_250),
.Y(n_1280)
);

INVx1_ASAP7_75t_L g1281 ( 
.A(n_702),
.Y(n_1281)
);

CKINVDCx5p33_ASAP7_75t_R g1282 ( 
.A(n_599),
.Y(n_1282)
);

CKINVDCx5p33_ASAP7_75t_R g1283 ( 
.A(n_769),
.Y(n_1283)
);

CKINVDCx5p33_ASAP7_75t_R g1284 ( 
.A(n_365),
.Y(n_1284)
);

CKINVDCx20_ASAP7_75t_R g1285 ( 
.A(n_784),
.Y(n_1285)
);

CKINVDCx5p33_ASAP7_75t_R g1286 ( 
.A(n_260),
.Y(n_1286)
);

CKINVDCx5p33_ASAP7_75t_R g1287 ( 
.A(n_493),
.Y(n_1287)
);

CKINVDCx5p33_ASAP7_75t_R g1288 ( 
.A(n_473),
.Y(n_1288)
);

CKINVDCx5p33_ASAP7_75t_R g1289 ( 
.A(n_259),
.Y(n_1289)
);

INVx2_ASAP7_75t_SL g1290 ( 
.A(n_1054),
.Y(n_1290)
);

INVx2_ASAP7_75t_L g1291 ( 
.A(n_96),
.Y(n_1291)
);

CKINVDCx5p33_ASAP7_75t_R g1292 ( 
.A(n_100),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_874),
.Y(n_1293)
);

CKINVDCx5p33_ASAP7_75t_R g1294 ( 
.A(n_741),
.Y(n_1294)
);

BUFx6f_ASAP7_75t_L g1295 ( 
.A(n_353),
.Y(n_1295)
);

INVx2_ASAP7_75t_L g1296 ( 
.A(n_170),
.Y(n_1296)
);

INVx2_ASAP7_75t_SL g1297 ( 
.A(n_392),
.Y(n_1297)
);

CKINVDCx5p33_ASAP7_75t_R g1298 ( 
.A(n_742),
.Y(n_1298)
);

INVx4_ASAP7_75t_R g1299 ( 
.A(n_541),
.Y(n_1299)
);

CKINVDCx5p33_ASAP7_75t_R g1300 ( 
.A(n_461),
.Y(n_1300)
);

CKINVDCx5p33_ASAP7_75t_R g1301 ( 
.A(n_601),
.Y(n_1301)
);

CKINVDCx5p33_ASAP7_75t_R g1302 ( 
.A(n_875),
.Y(n_1302)
);

CKINVDCx20_ASAP7_75t_R g1303 ( 
.A(n_548),
.Y(n_1303)
);

CKINVDCx5p33_ASAP7_75t_R g1304 ( 
.A(n_451),
.Y(n_1304)
);

CKINVDCx5p33_ASAP7_75t_R g1305 ( 
.A(n_83),
.Y(n_1305)
);

CKINVDCx5p33_ASAP7_75t_R g1306 ( 
.A(n_668),
.Y(n_1306)
);

CKINVDCx5p33_ASAP7_75t_R g1307 ( 
.A(n_181),
.Y(n_1307)
);

INVx2_ASAP7_75t_L g1308 ( 
.A(n_1020),
.Y(n_1308)
);

CKINVDCx5p33_ASAP7_75t_R g1309 ( 
.A(n_1038),
.Y(n_1309)
);

CKINVDCx5p33_ASAP7_75t_R g1310 ( 
.A(n_528),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_384),
.Y(n_1311)
);

CKINVDCx5p33_ASAP7_75t_R g1312 ( 
.A(n_935),
.Y(n_1312)
);

BUFx10_ASAP7_75t_L g1313 ( 
.A(n_67),
.Y(n_1313)
);

INVx1_ASAP7_75t_L g1314 ( 
.A(n_414),
.Y(n_1314)
);

INVx1_ASAP7_75t_L g1315 ( 
.A(n_700),
.Y(n_1315)
);

INVx1_ASAP7_75t_L g1316 ( 
.A(n_34),
.Y(n_1316)
);

INVx1_ASAP7_75t_SL g1317 ( 
.A(n_680),
.Y(n_1317)
);

INVx1_ASAP7_75t_L g1318 ( 
.A(n_310),
.Y(n_1318)
);

CKINVDCx5p33_ASAP7_75t_R g1319 ( 
.A(n_778),
.Y(n_1319)
);

CKINVDCx5p33_ASAP7_75t_R g1320 ( 
.A(n_440),
.Y(n_1320)
);

CKINVDCx5p33_ASAP7_75t_R g1321 ( 
.A(n_693),
.Y(n_1321)
);

BUFx3_ASAP7_75t_L g1322 ( 
.A(n_617),
.Y(n_1322)
);

INVx1_ASAP7_75t_L g1323 ( 
.A(n_83),
.Y(n_1323)
);

CKINVDCx5p33_ASAP7_75t_R g1324 ( 
.A(n_761),
.Y(n_1324)
);

INVx1_ASAP7_75t_L g1325 ( 
.A(n_1033),
.Y(n_1325)
);

INVx1_ASAP7_75t_L g1326 ( 
.A(n_855),
.Y(n_1326)
);

CKINVDCx5p33_ASAP7_75t_R g1327 ( 
.A(n_681),
.Y(n_1327)
);

CKINVDCx5p33_ASAP7_75t_R g1328 ( 
.A(n_790),
.Y(n_1328)
);

INVx1_ASAP7_75t_L g1329 ( 
.A(n_1027),
.Y(n_1329)
);

CKINVDCx5p33_ASAP7_75t_R g1330 ( 
.A(n_565),
.Y(n_1330)
);

BUFx10_ASAP7_75t_L g1331 ( 
.A(n_973),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_369),
.Y(n_1332)
);

CKINVDCx5p33_ASAP7_75t_R g1333 ( 
.A(n_206),
.Y(n_1333)
);

INVx1_ASAP7_75t_L g1334 ( 
.A(n_234),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_485),
.Y(n_1335)
);

CKINVDCx5p33_ASAP7_75t_R g1336 ( 
.A(n_58),
.Y(n_1336)
);

INVx1_ASAP7_75t_L g1337 ( 
.A(n_677),
.Y(n_1337)
);

CKINVDCx5p33_ASAP7_75t_R g1338 ( 
.A(n_107),
.Y(n_1338)
);

CKINVDCx5p33_ASAP7_75t_R g1339 ( 
.A(n_585),
.Y(n_1339)
);

CKINVDCx5p33_ASAP7_75t_R g1340 ( 
.A(n_880),
.Y(n_1340)
);

INVx1_ASAP7_75t_SL g1341 ( 
.A(n_731),
.Y(n_1341)
);

HB1xp67_ASAP7_75t_L g1342 ( 
.A(n_1008),
.Y(n_1342)
);

INVx2_ASAP7_75t_SL g1343 ( 
.A(n_511),
.Y(n_1343)
);

INVx1_ASAP7_75t_L g1344 ( 
.A(n_1026),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_631),
.Y(n_1345)
);

BUFx5_ASAP7_75t_L g1346 ( 
.A(n_954),
.Y(n_1346)
);

CKINVDCx5p33_ASAP7_75t_R g1347 ( 
.A(n_715),
.Y(n_1347)
);

CKINVDCx5p33_ASAP7_75t_R g1348 ( 
.A(n_528),
.Y(n_1348)
);

BUFx3_ASAP7_75t_L g1349 ( 
.A(n_531),
.Y(n_1349)
);

CKINVDCx20_ASAP7_75t_R g1350 ( 
.A(n_542),
.Y(n_1350)
);

CKINVDCx5p33_ASAP7_75t_R g1351 ( 
.A(n_863),
.Y(n_1351)
);

CKINVDCx5p33_ASAP7_75t_R g1352 ( 
.A(n_675),
.Y(n_1352)
);

CKINVDCx5p33_ASAP7_75t_R g1353 ( 
.A(n_652),
.Y(n_1353)
);

INVx2_ASAP7_75t_SL g1354 ( 
.A(n_893),
.Y(n_1354)
);

CKINVDCx5p33_ASAP7_75t_R g1355 ( 
.A(n_983),
.Y(n_1355)
);

INVx1_ASAP7_75t_SL g1356 ( 
.A(n_770),
.Y(n_1356)
);

BUFx3_ASAP7_75t_L g1357 ( 
.A(n_685),
.Y(n_1357)
);

INVx1_ASAP7_75t_L g1358 ( 
.A(n_480),
.Y(n_1358)
);

INVx1_ASAP7_75t_L g1359 ( 
.A(n_678),
.Y(n_1359)
);

INVx1_ASAP7_75t_L g1360 ( 
.A(n_351),
.Y(n_1360)
);

BUFx10_ASAP7_75t_L g1361 ( 
.A(n_1044),
.Y(n_1361)
);

CKINVDCx5p33_ASAP7_75t_R g1362 ( 
.A(n_281),
.Y(n_1362)
);

CKINVDCx5p33_ASAP7_75t_R g1363 ( 
.A(n_828),
.Y(n_1363)
);

CKINVDCx5p33_ASAP7_75t_R g1364 ( 
.A(n_597),
.Y(n_1364)
);

CKINVDCx5p33_ASAP7_75t_R g1365 ( 
.A(n_550),
.Y(n_1365)
);

CKINVDCx5p33_ASAP7_75t_R g1366 ( 
.A(n_1053),
.Y(n_1366)
);

CKINVDCx5p33_ASAP7_75t_R g1367 ( 
.A(n_929),
.Y(n_1367)
);

INVx1_ASAP7_75t_L g1368 ( 
.A(n_477),
.Y(n_1368)
);

INVx1_ASAP7_75t_L g1369 ( 
.A(n_367),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_905),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_717),
.Y(n_1371)
);

HB1xp67_ASAP7_75t_L g1372 ( 
.A(n_42),
.Y(n_1372)
);

INVx1_ASAP7_75t_L g1373 ( 
.A(n_3),
.Y(n_1373)
);

CKINVDCx5p33_ASAP7_75t_R g1374 ( 
.A(n_79),
.Y(n_1374)
);

INVx1_ASAP7_75t_L g1375 ( 
.A(n_523),
.Y(n_1375)
);

INVx1_ASAP7_75t_SL g1376 ( 
.A(n_219),
.Y(n_1376)
);

INVx1_ASAP7_75t_L g1377 ( 
.A(n_560),
.Y(n_1377)
);

INVx1_ASAP7_75t_L g1378 ( 
.A(n_149),
.Y(n_1378)
);

CKINVDCx20_ASAP7_75t_R g1379 ( 
.A(n_615),
.Y(n_1379)
);

INVx2_ASAP7_75t_SL g1380 ( 
.A(n_293),
.Y(n_1380)
);

CKINVDCx5p33_ASAP7_75t_R g1381 ( 
.A(n_101),
.Y(n_1381)
);

BUFx3_ASAP7_75t_L g1382 ( 
.A(n_659),
.Y(n_1382)
);

CKINVDCx5p33_ASAP7_75t_R g1383 ( 
.A(n_133),
.Y(n_1383)
);

CKINVDCx5p33_ASAP7_75t_R g1384 ( 
.A(n_26),
.Y(n_1384)
);

CKINVDCx5p33_ASAP7_75t_R g1385 ( 
.A(n_679),
.Y(n_1385)
);

CKINVDCx5p33_ASAP7_75t_R g1386 ( 
.A(n_580),
.Y(n_1386)
);

INVx1_ASAP7_75t_L g1387 ( 
.A(n_980),
.Y(n_1387)
);

CKINVDCx5p33_ASAP7_75t_R g1388 ( 
.A(n_676),
.Y(n_1388)
);

CKINVDCx5p33_ASAP7_75t_R g1389 ( 
.A(n_533),
.Y(n_1389)
);

INVx1_ASAP7_75t_L g1390 ( 
.A(n_856),
.Y(n_1390)
);

CKINVDCx14_ASAP7_75t_R g1391 ( 
.A(n_644),
.Y(n_1391)
);

CKINVDCx5p33_ASAP7_75t_R g1392 ( 
.A(n_1028),
.Y(n_1392)
);

INVx1_ASAP7_75t_L g1393 ( 
.A(n_1046),
.Y(n_1393)
);

INVx1_ASAP7_75t_L g1394 ( 
.A(n_1010),
.Y(n_1394)
);

CKINVDCx5p33_ASAP7_75t_R g1395 ( 
.A(n_648),
.Y(n_1395)
);

INVx1_ASAP7_75t_L g1396 ( 
.A(n_205),
.Y(n_1396)
);

CKINVDCx5p33_ASAP7_75t_R g1397 ( 
.A(n_194),
.Y(n_1397)
);

BUFx5_ASAP7_75t_L g1398 ( 
.A(n_645),
.Y(n_1398)
);

CKINVDCx5p33_ASAP7_75t_R g1399 ( 
.A(n_389),
.Y(n_1399)
);

CKINVDCx5p33_ASAP7_75t_R g1400 ( 
.A(n_1052),
.Y(n_1400)
);

INVx1_ASAP7_75t_L g1401 ( 
.A(n_486),
.Y(n_1401)
);

CKINVDCx5p33_ASAP7_75t_R g1402 ( 
.A(n_926),
.Y(n_1402)
);

CKINVDCx20_ASAP7_75t_R g1403 ( 
.A(n_613),
.Y(n_1403)
);

CKINVDCx5p33_ASAP7_75t_R g1404 ( 
.A(n_690),
.Y(n_1404)
);

HB1xp67_ASAP7_75t_L g1405 ( 
.A(n_617),
.Y(n_1405)
);

CKINVDCx5p33_ASAP7_75t_R g1406 ( 
.A(n_12),
.Y(n_1406)
);

CKINVDCx5p33_ASAP7_75t_R g1407 ( 
.A(n_755),
.Y(n_1407)
);

INVx1_ASAP7_75t_L g1408 ( 
.A(n_172),
.Y(n_1408)
);

CKINVDCx5p33_ASAP7_75t_R g1409 ( 
.A(n_886),
.Y(n_1409)
);

CKINVDCx5p33_ASAP7_75t_R g1410 ( 
.A(n_514),
.Y(n_1410)
);

CKINVDCx20_ASAP7_75t_R g1411 ( 
.A(n_189),
.Y(n_1411)
);

CKINVDCx20_ASAP7_75t_R g1412 ( 
.A(n_993),
.Y(n_1412)
);

INVx1_ASAP7_75t_L g1413 ( 
.A(n_563),
.Y(n_1413)
);

CKINVDCx5p33_ASAP7_75t_R g1414 ( 
.A(n_692),
.Y(n_1414)
);

CKINVDCx5p33_ASAP7_75t_R g1415 ( 
.A(n_366),
.Y(n_1415)
);

CKINVDCx5p33_ASAP7_75t_R g1416 ( 
.A(n_236),
.Y(n_1416)
);

CKINVDCx5p33_ASAP7_75t_R g1417 ( 
.A(n_270),
.Y(n_1417)
);

BUFx3_ASAP7_75t_L g1418 ( 
.A(n_1029),
.Y(n_1418)
);

CKINVDCx5p33_ASAP7_75t_R g1419 ( 
.A(n_128),
.Y(n_1419)
);

CKINVDCx20_ASAP7_75t_R g1420 ( 
.A(n_171),
.Y(n_1420)
);

INVx1_ASAP7_75t_L g1421 ( 
.A(n_214),
.Y(n_1421)
);

INVx1_ASAP7_75t_L g1422 ( 
.A(n_156),
.Y(n_1422)
);

CKINVDCx5p33_ASAP7_75t_R g1423 ( 
.A(n_559),
.Y(n_1423)
);

INVx1_ASAP7_75t_L g1424 ( 
.A(n_991),
.Y(n_1424)
);

INVxp67_ASAP7_75t_L g1425 ( 
.A(n_667),
.Y(n_1425)
);

INVx1_ASAP7_75t_L g1426 ( 
.A(n_810),
.Y(n_1426)
);

INVx1_ASAP7_75t_L g1427 ( 
.A(n_703),
.Y(n_1427)
);

INVx1_ASAP7_75t_SL g1428 ( 
.A(n_511),
.Y(n_1428)
);

INVx1_ASAP7_75t_L g1429 ( 
.A(n_728),
.Y(n_1429)
);

CKINVDCx5p33_ASAP7_75t_R g1430 ( 
.A(n_111),
.Y(n_1430)
);

CKINVDCx5p33_ASAP7_75t_R g1431 ( 
.A(n_1035),
.Y(n_1431)
);

CKINVDCx5p33_ASAP7_75t_R g1432 ( 
.A(n_252),
.Y(n_1432)
);

CKINVDCx16_ASAP7_75t_R g1433 ( 
.A(n_1005),
.Y(n_1433)
);

CKINVDCx20_ASAP7_75t_R g1434 ( 
.A(n_406),
.Y(n_1434)
);

INVx2_ASAP7_75t_L g1435 ( 
.A(n_548),
.Y(n_1435)
);

INVx1_ASAP7_75t_L g1436 ( 
.A(n_1045),
.Y(n_1436)
);

BUFx5_ASAP7_75t_L g1437 ( 
.A(n_701),
.Y(n_1437)
);

CKINVDCx14_ASAP7_75t_R g1438 ( 
.A(n_556),
.Y(n_1438)
);

CKINVDCx5p33_ASAP7_75t_R g1439 ( 
.A(n_47),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_91),
.Y(n_1440)
);

INVx2_ASAP7_75t_SL g1441 ( 
.A(n_908),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_674),
.Y(n_1442)
);

CKINVDCx5p33_ASAP7_75t_R g1443 ( 
.A(n_599),
.Y(n_1443)
);

CKINVDCx5p33_ASAP7_75t_R g1444 ( 
.A(n_372),
.Y(n_1444)
);

INVx1_ASAP7_75t_L g1445 ( 
.A(n_842),
.Y(n_1445)
);

INVx1_ASAP7_75t_L g1446 ( 
.A(n_304),
.Y(n_1446)
);

CKINVDCx5p33_ASAP7_75t_R g1447 ( 
.A(n_577),
.Y(n_1447)
);

CKINVDCx5p33_ASAP7_75t_R g1448 ( 
.A(n_665),
.Y(n_1448)
);

CKINVDCx5p33_ASAP7_75t_R g1449 ( 
.A(n_958),
.Y(n_1449)
);

CKINVDCx5p33_ASAP7_75t_R g1450 ( 
.A(n_158),
.Y(n_1450)
);

CKINVDCx5p33_ASAP7_75t_R g1451 ( 
.A(n_323),
.Y(n_1451)
);

BUFx3_ASAP7_75t_L g1452 ( 
.A(n_643),
.Y(n_1452)
);

CKINVDCx5p33_ASAP7_75t_R g1453 ( 
.A(n_427),
.Y(n_1453)
);

CKINVDCx5p33_ASAP7_75t_R g1454 ( 
.A(n_119),
.Y(n_1454)
);

BUFx2_ASAP7_75t_L g1455 ( 
.A(n_1042),
.Y(n_1455)
);

CKINVDCx20_ASAP7_75t_R g1456 ( 
.A(n_945),
.Y(n_1456)
);

CKINVDCx5p33_ASAP7_75t_R g1457 ( 
.A(n_48),
.Y(n_1457)
);

CKINVDCx5p33_ASAP7_75t_R g1458 ( 
.A(n_642),
.Y(n_1458)
);

CKINVDCx5p33_ASAP7_75t_R g1459 ( 
.A(n_666),
.Y(n_1459)
);

INVx2_ASAP7_75t_SL g1460 ( 
.A(n_788),
.Y(n_1460)
);

CKINVDCx5p33_ASAP7_75t_R g1461 ( 
.A(n_967),
.Y(n_1461)
);

CKINVDCx5p33_ASAP7_75t_R g1462 ( 
.A(n_989),
.Y(n_1462)
);

INVx1_ASAP7_75t_L g1463 ( 
.A(n_998),
.Y(n_1463)
);

CKINVDCx5p33_ASAP7_75t_R g1464 ( 
.A(n_67),
.Y(n_1464)
);

CKINVDCx5p33_ASAP7_75t_R g1465 ( 
.A(n_313),
.Y(n_1465)
);

CKINVDCx20_ASAP7_75t_R g1466 ( 
.A(n_698),
.Y(n_1466)
);

CKINVDCx5p33_ASAP7_75t_R g1467 ( 
.A(n_59),
.Y(n_1467)
);

CKINVDCx5p33_ASAP7_75t_R g1468 ( 
.A(n_464),
.Y(n_1468)
);

CKINVDCx5p33_ASAP7_75t_R g1469 ( 
.A(n_661),
.Y(n_1469)
);

CKINVDCx5p33_ASAP7_75t_R g1470 ( 
.A(n_639),
.Y(n_1470)
);

BUFx5_ASAP7_75t_L g1471 ( 
.A(n_249),
.Y(n_1471)
);

INVx1_ASAP7_75t_SL g1472 ( 
.A(n_625),
.Y(n_1472)
);

INVx1_ASAP7_75t_L g1473 ( 
.A(n_716),
.Y(n_1473)
);

CKINVDCx5p33_ASAP7_75t_R g1474 ( 
.A(n_806),
.Y(n_1474)
);

BUFx6f_ASAP7_75t_L g1475 ( 
.A(n_171),
.Y(n_1475)
);

INVx1_ASAP7_75t_L g1476 ( 
.A(n_531),
.Y(n_1476)
);

CKINVDCx5p33_ASAP7_75t_R g1477 ( 
.A(n_495),
.Y(n_1477)
);

BUFx10_ASAP7_75t_L g1478 ( 
.A(n_299),
.Y(n_1478)
);

CKINVDCx5p33_ASAP7_75t_R g1479 ( 
.A(n_723),
.Y(n_1479)
);

CKINVDCx5p33_ASAP7_75t_R g1480 ( 
.A(n_799),
.Y(n_1480)
);

CKINVDCx5p33_ASAP7_75t_R g1481 ( 
.A(n_136),
.Y(n_1481)
);

INVx1_ASAP7_75t_L g1482 ( 
.A(n_697),
.Y(n_1482)
);

INVx2_ASAP7_75t_SL g1483 ( 
.A(n_25),
.Y(n_1483)
);

CKINVDCx5p33_ASAP7_75t_R g1484 ( 
.A(n_665),
.Y(n_1484)
);

INVx1_ASAP7_75t_L g1485 ( 
.A(n_624),
.Y(n_1485)
);

CKINVDCx5p33_ASAP7_75t_R g1486 ( 
.A(n_662),
.Y(n_1486)
);

INVx1_ASAP7_75t_L g1487 ( 
.A(n_747),
.Y(n_1487)
);

INVx1_ASAP7_75t_L g1488 ( 
.A(n_431),
.Y(n_1488)
);

CKINVDCx5p33_ASAP7_75t_R g1489 ( 
.A(n_547),
.Y(n_1489)
);

BUFx6f_ASAP7_75t_L g1490 ( 
.A(n_332),
.Y(n_1490)
);

CKINVDCx5p33_ASAP7_75t_R g1491 ( 
.A(n_269),
.Y(n_1491)
);

BUFx8_ASAP7_75t_SL g1492 ( 
.A(n_199),
.Y(n_1492)
);

CKINVDCx5p33_ASAP7_75t_R g1493 ( 
.A(n_111),
.Y(n_1493)
);

CKINVDCx5p33_ASAP7_75t_R g1494 ( 
.A(n_773),
.Y(n_1494)
);

CKINVDCx5p33_ASAP7_75t_R g1495 ( 
.A(n_79),
.Y(n_1495)
);

CKINVDCx5p33_ASAP7_75t_R g1496 ( 
.A(n_581),
.Y(n_1496)
);

INVx1_ASAP7_75t_L g1497 ( 
.A(n_271),
.Y(n_1497)
);

CKINVDCx5p33_ASAP7_75t_R g1498 ( 
.A(n_837),
.Y(n_1498)
);

CKINVDCx5p33_ASAP7_75t_R g1499 ( 
.A(n_138),
.Y(n_1499)
);

INVx1_ASAP7_75t_L g1500 ( 
.A(n_658),
.Y(n_1500)
);

CKINVDCx5p33_ASAP7_75t_R g1501 ( 
.A(n_230),
.Y(n_1501)
);

INVx1_ASAP7_75t_L g1502 ( 
.A(n_1000),
.Y(n_1502)
);

CKINVDCx5p33_ASAP7_75t_R g1503 ( 
.A(n_592),
.Y(n_1503)
);

CKINVDCx5p33_ASAP7_75t_R g1504 ( 
.A(n_768),
.Y(n_1504)
);

INVx1_ASAP7_75t_L g1505 ( 
.A(n_1017),
.Y(n_1505)
);

INVx2_ASAP7_75t_L g1506 ( 
.A(n_933),
.Y(n_1506)
);

INVx1_ASAP7_75t_SL g1507 ( 
.A(n_925),
.Y(n_1507)
);

INVx1_ASAP7_75t_L g1508 ( 
.A(n_671),
.Y(n_1508)
);

BUFx5_ASAP7_75t_L g1509 ( 
.A(n_437),
.Y(n_1509)
);

INVx1_ASAP7_75t_L g1510 ( 
.A(n_625),
.Y(n_1510)
);

INVx1_ASAP7_75t_L g1511 ( 
.A(n_80),
.Y(n_1511)
);

INVx1_ASAP7_75t_L g1512 ( 
.A(n_144),
.Y(n_1512)
);

CKINVDCx5p33_ASAP7_75t_R g1513 ( 
.A(n_157),
.Y(n_1513)
);

CKINVDCx5p33_ASAP7_75t_R g1514 ( 
.A(n_354),
.Y(n_1514)
);

CKINVDCx5p33_ASAP7_75t_R g1515 ( 
.A(n_636),
.Y(n_1515)
);

CKINVDCx5p33_ASAP7_75t_R g1516 ( 
.A(n_475),
.Y(n_1516)
);

CKINVDCx5p33_ASAP7_75t_R g1517 ( 
.A(n_750),
.Y(n_1517)
);

HB1xp67_ASAP7_75t_L g1518 ( 
.A(n_297),
.Y(n_1518)
);

BUFx8_ASAP7_75t_SL g1519 ( 
.A(n_411),
.Y(n_1519)
);

CKINVDCx20_ASAP7_75t_R g1520 ( 
.A(n_192),
.Y(n_1520)
);

INVx2_ASAP7_75t_L g1521 ( 
.A(n_902),
.Y(n_1521)
);

CKINVDCx5p33_ASAP7_75t_R g1522 ( 
.A(n_557),
.Y(n_1522)
);

CKINVDCx5p33_ASAP7_75t_R g1523 ( 
.A(n_947),
.Y(n_1523)
);

CKINVDCx5p33_ASAP7_75t_R g1524 ( 
.A(n_575),
.Y(n_1524)
);

CKINVDCx20_ASAP7_75t_R g1525 ( 
.A(n_463),
.Y(n_1525)
);

CKINVDCx5p33_ASAP7_75t_R g1526 ( 
.A(n_391),
.Y(n_1526)
);

CKINVDCx5p33_ASAP7_75t_R g1527 ( 
.A(n_982),
.Y(n_1527)
);

CKINVDCx5p33_ASAP7_75t_R g1528 ( 
.A(n_52),
.Y(n_1528)
);

CKINVDCx5p33_ASAP7_75t_R g1529 ( 
.A(n_21),
.Y(n_1529)
);

INVx1_ASAP7_75t_L g1530 ( 
.A(n_1059),
.Y(n_1530)
);

CKINVDCx20_ASAP7_75t_R g1531 ( 
.A(n_634),
.Y(n_1531)
);

CKINVDCx5p33_ASAP7_75t_R g1532 ( 
.A(n_724),
.Y(n_1532)
);

CKINVDCx20_ASAP7_75t_R g1533 ( 
.A(n_263),
.Y(n_1533)
);

CKINVDCx5p33_ASAP7_75t_R g1534 ( 
.A(n_626),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_859),
.Y(n_1535)
);

INVx1_ASAP7_75t_L g1536 ( 
.A(n_943),
.Y(n_1536)
);

INVx2_ASAP7_75t_L g1537 ( 
.A(n_757),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_241),
.Y(n_1538)
);

CKINVDCx20_ASAP7_75t_R g1539 ( 
.A(n_683),
.Y(n_1539)
);

BUFx10_ASAP7_75t_L g1540 ( 
.A(n_686),
.Y(n_1540)
);

CKINVDCx5p33_ASAP7_75t_R g1541 ( 
.A(n_539),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_405),
.Y(n_1542)
);

CKINVDCx5p33_ASAP7_75t_R g1543 ( 
.A(n_682),
.Y(n_1543)
);

INVx1_ASAP7_75t_L g1544 ( 
.A(n_910),
.Y(n_1544)
);

CKINVDCx5p33_ASAP7_75t_R g1545 ( 
.A(n_394),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_257),
.Y(n_1546)
);

CKINVDCx5p33_ASAP7_75t_R g1547 ( 
.A(n_651),
.Y(n_1547)
);

BUFx5_ASAP7_75t_L g1548 ( 
.A(n_166),
.Y(n_1548)
);

INVx1_ASAP7_75t_L g1549 ( 
.A(n_130),
.Y(n_1549)
);

INVx1_ASAP7_75t_L g1550 ( 
.A(n_722),
.Y(n_1550)
);

CKINVDCx5p33_ASAP7_75t_R g1551 ( 
.A(n_92),
.Y(n_1551)
);

INVx1_ASAP7_75t_SL g1552 ( 
.A(n_202),
.Y(n_1552)
);

CKINVDCx5p33_ASAP7_75t_R g1553 ( 
.A(n_331),
.Y(n_1553)
);

CKINVDCx5p33_ASAP7_75t_R g1554 ( 
.A(n_439),
.Y(n_1554)
);

INVx2_ASAP7_75t_SL g1555 ( 
.A(n_660),
.Y(n_1555)
);

CKINVDCx5p33_ASAP7_75t_R g1556 ( 
.A(n_300),
.Y(n_1556)
);

CKINVDCx5p33_ASAP7_75t_R g1557 ( 
.A(n_250),
.Y(n_1557)
);

CKINVDCx5p33_ASAP7_75t_R g1558 ( 
.A(n_383),
.Y(n_1558)
);

CKINVDCx5p33_ASAP7_75t_R g1559 ( 
.A(n_292),
.Y(n_1559)
);

BUFx2_ASAP7_75t_L g1560 ( 
.A(n_627),
.Y(n_1560)
);

INVx1_ASAP7_75t_SL g1561 ( 
.A(n_766),
.Y(n_1561)
);

INVx1_ASAP7_75t_L g1562 ( 
.A(n_635),
.Y(n_1562)
);

CKINVDCx5p33_ASAP7_75t_R g1563 ( 
.A(n_669),
.Y(n_1563)
);

CKINVDCx5p33_ASAP7_75t_R g1564 ( 
.A(n_734),
.Y(n_1564)
);

BUFx6f_ASAP7_75t_L g1565 ( 
.A(n_563),
.Y(n_1565)
);

INVx1_ASAP7_75t_L g1566 ( 
.A(n_1081),
.Y(n_1566)
);

CKINVDCx20_ASAP7_75t_R g1567 ( 
.A(n_1065),
.Y(n_1567)
);

INVx1_ASAP7_75t_L g1568 ( 
.A(n_1081),
.Y(n_1568)
);

INVxp67_ASAP7_75t_L g1569 ( 
.A(n_1173),
.Y(n_1569)
);

CKINVDCx20_ASAP7_75t_R g1570 ( 
.A(n_1113),
.Y(n_1570)
);

INVx1_ASAP7_75t_L g1571 ( 
.A(n_1081),
.Y(n_1571)
);

INVx1_ASAP7_75t_L g1572 ( 
.A(n_1081),
.Y(n_1572)
);

CKINVDCx5p33_ASAP7_75t_R g1573 ( 
.A(n_1202),
.Y(n_1573)
);

INVx1_ASAP7_75t_L g1574 ( 
.A(n_1081),
.Y(n_1574)
);

INVx1_ASAP7_75t_L g1575 ( 
.A(n_1257),
.Y(n_1575)
);

CKINVDCx16_ASAP7_75t_R g1576 ( 
.A(n_1170),
.Y(n_1576)
);

INVxp67_ASAP7_75t_SL g1577 ( 
.A(n_1342),
.Y(n_1577)
);

CKINVDCx20_ASAP7_75t_R g1578 ( 
.A(n_1125),
.Y(n_1578)
);

CKINVDCx5p33_ASAP7_75t_R g1579 ( 
.A(n_1276),
.Y(n_1579)
);

INVx1_ASAP7_75t_L g1580 ( 
.A(n_1257),
.Y(n_1580)
);

INVx1_ASAP7_75t_L g1581 ( 
.A(n_1257),
.Y(n_1581)
);

INVxp67_ASAP7_75t_L g1582 ( 
.A(n_1165),
.Y(n_1582)
);

INVx1_ASAP7_75t_L g1583 ( 
.A(n_1257),
.Y(n_1583)
);

CKINVDCx16_ASAP7_75t_R g1584 ( 
.A(n_1245),
.Y(n_1584)
);

CKINVDCx20_ASAP7_75t_R g1585 ( 
.A(n_1161),
.Y(n_1585)
);

INVx1_ASAP7_75t_L g1586 ( 
.A(n_1257),
.Y(n_1586)
);

CKINVDCx20_ASAP7_75t_R g1587 ( 
.A(n_1192),
.Y(n_1587)
);

NOR2xp67_ASAP7_75t_L g1588 ( 
.A(n_1425),
.B(n_0),
.Y(n_1588)
);

CKINVDCx5p33_ASAP7_75t_R g1589 ( 
.A(n_1492),
.Y(n_1589)
);

INVxp67_ASAP7_75t_SL g1590 ( 
.A(n_1072),
.Y(n_1590)
);

CKINVDCx20_ASAP7_75t_R g1591 ( 
.A(n_1193),
.Y(n_1591)
);

CKINVDCx20_ASAP7_75t_R g1592 ( 
.A(n_1285),
.Y(n_1592)
);

INVx1_ASAP7_75t_L g1593 ( 
.A(n_1398),
.Y(n_1593)
);

INVxp67_ASAP7_75t_SL g1594 ( 
.A(n_1227),
.Y(n_1594)
);

INVx1_ASAP7_75t_L g1595 ( 
.A(n_1398),
.Y(n_1595)
);

CKINVDCx5p33_ASAP7_75t_R g1596 ( 
.A(n_1519),
.Y(n_1596)
);

INVx1_ASAP7_75t_L g1597 ( 
.A(n_1398),
.Y(n_1597)
);

CKINVDCx5p33_ASAP7_75t_R g1598 ( 
.A(n_1063),
.Y(n_1598)
);

CKINVDCx5p33_ASAP7_75t_R g1599 ( 
.A(n_1068),
.Y(n_1599)
);

HB1xp67_ASAP7_75t_L g1600 ( 
.A(n_1372),
.Y(n_1600)
);

INVxp67_ASAP7_75t_L g1601 ( 
.A(n_1181),
.Y(n_1601)
);

CKINVDCx5p33_ASAP7_75t_R g1602 ( 
.A(n_1069),
.Y(n_1602)
);

INVxp67_ASAP7_75t_SL g1603 ( 
.A(n_1455),
.Y(n_1603)
);

NOR2xp33_ASAP7_75t_L g1604 ( 
.A(n_1156),
.B(n_1),
.Y(n_1604)
);

NOR2xp33_ASAP7_75t_L g1605 ( 
.A(n_1190),
.B(n_1),
.Y(n_1605)
);

BUFx2_ASAP7_75t_L g1606 ( 
.A(n_1560),
.Y(n_1606)
);

INVx1_ASAP7_75t_L g1607 ( 
.A(n_1398),
.Y(n_1607)
);

CKINVDCx5p33_ASAP7_75t_R g1608 ( 
.A(n_1070),
.Y(n_1608)
);

BUFx3_ASAP7_75t_L g1609 ( 
.A(n_1166),
.Y(n_1609)
);

INVx1_ASAP7_75t_L g1610 ( 
.A(n_1398),
.Y(n_1610)
);

NOR2xp33_ASAP7_75t_L g1611 ( 
.A(n_1391),
.B(n_2),
.Y(n_1611)
);

INVx1_ASAP7_75t_L g1612 ( 
.A(n_1437),
.Y(n_1612)
);

CKINVDCx5p33_ASAP7_75t_R g1613 ( 
.A(n_1071),
.Y(n_1613)
);

INVx1_ASAP7_75t_L g1614 ( 
.A(n_1437),
.Y(n_1614)
);

HB1xp67_ASAP7_75t_L g1615 ( 
.A(n_1405),
.Y(n_1615)
);

CKINVDCx20_ASAP7_75t_R g1616 ( 
.A(n_1412),
.Y(n_1616)
);

CKINVDCx5p33_ASAP7_75t_R g1617 ( 
.A(n_1076),
.Y(n_1617)
);

INVx1_ASAP7_75t_L g1618 ( 
.A(n_1437),
.Y(n_1618)
);

INVxp33_ASAP7_75t_SL g1619 ( 
.A(n_1518),
.Y(n_1619)
);

CKINVDCx20_ASAP7_75t_R g1620 ( 
.A(n_1456),
.Y(n_1620)
);

CKINVDCx5p33_ASAP7_75t_R g1621 ( 
.A(n_1104),
.Y(n_1621)
);

INVx1_ASAP7_75t_L g1622 ( 
.A(n_1437),
.Y(n_1622)
);

CKINVDCx5p33_ASAP7_75t_R g1623 ( 
.A(n_1112),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1437),
.Y(n_1624)
);

NOR2xp33_ASAP7_75t_L g1625 ( 
.A(n_1438),
.B(n_2),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1164),
.B(n_0),
.Y(n_1626)
);

CKINVDCx16_ASAP7_75t_R g1627 ( 
.A(n_1433),
.Y(n_1627)
);

CKINVDCx20_ASAP7_75t_R g1628 ( 
.A(n_1126),
.Y(n_1628)
);

CKINVDCx5p33_ASAP7_75t_R g1629 ( 
.A(n_1135),
.Y(n_1629)
);

BUFx3_ASAP7_75t_L g1630 ( 
.A(n_1166),
.Y(n_1630)
);

INVx2_ASAP7_75t_L g1631 ( 
.A(n_1471),
.Y(n_1631)
);

INVx1_ASAP7_75t_L g1632 ( 
.A(n_1471),
.Y(n_1632)
);

INVx1_ASAP7_75t_L g1633 ( 
.A(n_1471),
.Y(n_1633)
);

INVx1_ASAP7_75t_L g1634 ( 
.A(n_1471),
.Y(n_1634)
);

CKINVDCx20_ASAP7_75t_R g1635 ( 
.A(n_1149),
.Y(n_1635)
);

INVx1_ASAP7_75t_L g1636 ( 
.A(n_1471),
.Y(n_1636)
);

CKINVDCx5p33_ASAP7_75t_R g1637 ( 
.A(n_1153),
.Y(n_1637)
);

INVx1_ASAP7_75t_L g1638 ( 
.A(n_1509),
.Y(n_1638)
);

CKINVDCx5p33_ASAP7_75t_R g1639 ( 
.A(n_1163),
.Y(n_1639)
);

INVx1_ASAP7_75t_L g1640 ( 
.A(n_1509),
.Y(n_1640)
);

INVxp67_ASAP7_75t_SL g1641 ( 
.A(n_1155),
.Y(n_1641)
);

INVx1_ASAP7_75t_L g1642 ( 
.A(n_1566),
.Y(n_1642)
);

INVx1_ASAP7_75t_L g1643 ( 
.A(n_1568),
.Y(n_1643)
);

INVx4_ASAP7_75t_L g1644 ( 
.A(n_1598),
.Y(n_1644)
);

INVx3_ASAP7_75t_L g1645 ( 
.A(n_1631),
.Y(n_1645)
);

INVx2_ASAP7_75t_L g1646 ( 
.A(n_1571),
.Y(n_1646)
);

INVx1_ASAP7_75t_L g1647 ( 
.A(n_1572),
.Y(n_1647)
);

INVx3_ASAP7_75t_L g1648 ( 
.A(n_1609),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_L g1649 ( 
.A(n_1599),
.B(n_1290),
.Y(n_1649)
);

INVx2_ASAP7_75t_L g1650 ( 
.A(n_1574),
.Y(n_1650)
);

NAND2xp5_ASAP7_75t_L g1651 ( 
.A(n_1602),
.B(n_1354),
.Y(n_1651)
);

CKINVDCx5p33_ASAP7_75t_R g1652 ( 
.A(n_1608),
.Y(n_1652)
);

BUFx6f_ASAP7_75t_L g1653 ( 
.A(n_1575),
.Y(n_1653)
);

INVx1_ASAP7_75t_L g1654 ( 
.A(n_1580),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1581),
.Y(n_1655)
);

INVxp67_ASAP7_75t_L g1656 ( 
.A(n_1630),
.Y(n_1656)
);

INVx1_ASAP7_75t_L g1657 ( 
.A(n_1583),
.Y(n_1657)
);

HB1xp67_ASAP7_75t_L g1658 ( 
.A(n_1576),
.Y(n_1658)
);

INVx1_ASAP7_75t_L g1659 ( 
.A(n_1586),
.Y(n_1659)
);

INVxp67_ASAP7_75t_L g1660 ( 
.A(n_1606),
.Y(n_1660)
);

INVx1_ASAP7_75t_L g1661 ( 
.A(n_1593),
.Y(n_1661)
);

NAND2xp5_ASAP7_75t_L g1662 ( 
.A(n_1613),
.B(n_1441),
.Y(n_1662)
);

INVx1_ASAP7_75t_L g1663 ( 
.A(n_1595),
.Y(n_1663)
);

INVx1_ASAP7_75t_L g1664 ( 
.A(n_1597),
.Y(n_1664)
);

INVx2_ASAP7_75t_L g1665 ( 
.A(n_1607),
.Y(n_1665)
);

INVx2_ASAP7_75t_L g1666 ( 
.A(n_1610),
.Y(n_1666)
);

INVx1_ASAP7_75t_L g1667 ( 
.A(n_1612),
.Y(n_1667)
);

NAND2xp5_ASAP7_75t_L g1668 ( 
.A(n_1617),
.B(n_1460),
.Y(n_1668)
);

INVx1_ASAP7_75t_L g1669 ( 
.A(n_1614),
.Y(n_1669)
);

NAND2xp5_ASAP7_75t_L g1670 ( 
.A(n_1621),
.B(n_1279),
.Y(n_1670)
);

CKINVDCx8_ASAP7_75t_R g1671 ( 
.A(n_1584),
.Y(n_1671)
);

AND2x2_ASAP7_75t_L g1672 ( 
.A(n_1641),
.B(n_1118),
.Y(n_1672)
);

BUFx6f_ASAP7_75t_L g1673 ( 
.A(n_1618),
.Y(n_1673)
);

INVx1_ASAP7_75t_L g1674 ( 
.A(n_1622),
.Y(n_1674)
);

NOR2xp33_ASAP7_75t_L g1675 ( 
.A(n_1623),
.B(n_1211),
.Y(n_1675)
);

BUFx6f_ASAP7_75t_L g1676 ( 
.A(n_1624),
.Y(n_1676)
);

AND2x2_ASAP7_75t_L g1677 ( 
.A(n_1590),
.B(n_1179),
.Y(n_1677)
);

NAND3xp33_ASAP7_75t_L g1678 ( 
.A(n_1604),
.B(n_1085),
.C(n_1083),
.Y(n_1678)
);

INVx2_ASAP7_75t_L g1679 ( 
.A(n_1640),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1629),
.B(n_1418),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1632),
.Y(n_1681)
);

NAND2xp5_ASAP7_75t_SL g1682 ( 
.A(n_1627),
.B(n_1167),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1637),
.B(n_1075),
.Y(n_1683)
);

INVx1_ASAP7_75t_L g1684 ( 
.A(n_1633),
.Y(n_1684)
);

CKINVDCx5p33_ASAP7_75t_R g1685 ( 
.A(n_1639),
.Y(n_1685)
);

INVx1_ASAP7_75t_L g1686 ( 
.A(n_1634),
.Y(n_1686)
);

NAND2xp5_ASAP7_75t_L g1687 ( 
.A(n_1577),
.B(n_1091),
.Y(n_1687)
);

HB1xp67_ASAP7_75t_L g1688 ( 
.A(n_1569),
.Y(n_1688)
);

INVx1_ASAP7_75t_L g1689 ( 
.A(n_1636),
.Y(n_1689)
);

INVx1_ASAP7_75t_L g1690 ( 
.A(n_1638),
.Y(n_1690)
);

NAND2xp5_ASAP7_75t_L g1691 ( 
.A(n_1594),
.B(n_1154),
.Y(n_1691)
);

INVx2_ASAP7_75t_L g1692 ( 
.A(n_1626),
.Y(n_1692)
);

NAND2xp5_ASAP7_75t_L g1693 ( 
.A(n_1603),
.B(n_1308),
.Y(n_1693)
);

INVx1_ASAP7_75t_L g1694 ( 
.A(n_1588),
.Y(n_1694)
);

INVx2_ASAP7_75t_L g1695 ( 
.A(n_1582),
.Y(n_1695)
);

BUFx6f_ASAP7_75t_L g1696 ( 
.A(n_1605),
.Y(n_1696)
);

HB1xp67_ASAP7_75t_L g1697 ( 
.A(n_1601),
.Y(n_1697)
);

AND2x2_ASAP7_75t_L g1698 ( 
.A(n_1582),
.B(n_1322),
.Y(n_1698)
);

AND2x2_ASAP7_75t_L g1699 ( 
.A(n_1600),
.B(n_1349),
.Y(n_1699)
);

INVx1_ASAP7_75t_L g1700 ( 
.A(n_1615),
.Y(n_1700)
);

BUFx3_ASAP7_75t_L g1701 ( 
.A(n_1628),
.Y(n_1701)
);

INVxp33_ASAP7_75t_L g1702 ( 
.A(n_1611),
.Y(n_1702)
);

NAND2xp5_ASAP7_75t_L g1703 ( 
.A(n_1625),
.B(n_1506),
.Y(n_1703)
);

BUFx6f_ASAP7_75t_L g1704 ( 
.A(n_1573),
.Y(n_1704)
);

INVx4_ASAP7_75t_L g1705 ( 
.A(n_1704),
.Y(n_1705)
);

INVx1_ASAP7_75t_L g1706 ( 
.A(n_1653),
.Y(n_1706)
);

AND2x4_ASAP7_75t_L g1707 ( 
.A(n_1672),
.B(n_1635),
.Y(n_1707)
);

INVx1_ASAP7_75t_L g1708 ( 
.A(n_1653),
.Y(n_1708)
);

NAND2xp5_ASAP7_75t_L g1709 ( 
.A(n_1675),
.B(n_1223),
.Y(n_1709)
);

AO21x2_ASAP7_75t_L g1710 ( 
.A1(n_1683),
.A2(n_1082),
.B(n_1060),
.Y(n_1710)
);

INVx2_ASAP7_75t_L g1711 ( 
.A(n_1673),
.Y(n_1711)
);

INVx1_ASAP7_75t_L g1712 ( 
.A(n_1673),
.Y(n_1712)
);

INVx1_ASAP7_75t_L g1713 ( 
.A(n_1676),
.Y(n_1713)
);

INVx1_ASAP7_75t_L g1714 ( 
.A(n_1676),
.Y(n_1714)
);

INVx5_ASAP7_75t_L g1715 ( 
.A(n_1648),
.Y(n_1715)
);

AND2x6_ASAP7_75t_L g1716 ( 
.A(n_1692),
.B(n_1064),
.Y(n_1716)
);

NOR2xp33_ASAP7_75t_L g1717 ( 
.A(n_1702),
.B(n_1619),
.Y(n_1717)
);

NAND2xp5_ASAP7_75t_L g1718 ( 
.A(n_1703),
.B(n_1670),
.Y(n_1718)
);

INVx3_ASAP7_75t_L g1719 ( 
.A(n_1645),
.Y(n_1719)
);

OR2x2_ASAP7_75t_L g1720 ( 
.A(n_1660),
.B(n_1579),
.Y(n_1720)
);

NAND2xp5_ASAP7_75t_L g1721 ( 
.A(n_1680),
.B(n_1341),
.Y(n_1721)
);

NOR2xp33_ASAP7_75t_L g1722 ( 
.A(n_1649),
.B(n_1589),
.Y(n_1722)
);

BUFx2_ASAP7_75t_L g1723 ( 
.A(n_1658),
.Y(n_1723)
);

NAND2xp5_ASAP7_75t_SL g1724 ( 
.A(n_1696),
.B(n_1596),
.Y(n_1724)
);

AND2x2_ASAP7_75t_SL g1725 ( 
.A(n_1696),
.B(n_1688),
.Y(n_1725)
);

BUFx3_ASAP7_75t_L g1726 ( 
.A(n_1704),
.Y(n_1726)
);

NOR2xp33_ASAP7_75t_SL g1727 ( 
.A(n_1671),
.B(n_1567),
.Y(n_1727)
);

INVx2_ASAP7_75t_L g1728 ( 
.A(n_1646),
.Y(n_1728)
);

CKINVDCx5p33_ASAP7_75t_R g1729 ( 
.A(n_1652),
.Y(n_1729)
);

NAND2xp5_ASAP7_75t_SL g1730 ( 
.A(n_1685),
.B(n_1695),
.Y(n_1730)
);

INVxp67_ASAP7_75t_L g1731 ( 
.A(n_1697),
.Y(n_1731)
);

NAND2xp5_ASAP7_75t_L g1732 ( 
.A(n_1651),
.B(n_1356),
.Y(n_1732)
);

INVx1_ASAP7_75t_L g1733 ( 
.A(n_1642),
.Y(n_1733)
);

OR2x6_ASAP7_75t_L g1734 ( 
.A(n_1701),
.B(n_1124),
.Y(n_1734)
);

INVx5_ASAP7_75t_L g1735 ( 
.A(n_1698),
.Y(n_1735)
);

INVx1_ASAP7_75t_L g1736 ( 
.A(n_1643),
.Y(n_1736)
);

AND2x2_ASAP7_75t_SL g1737 ( 
.A(n_1700),
.B(n_1080),
.Y(n_1737)
);

NAND2xp5_ASAP7_75t_SL g1738 ( 
.A(n_1662),
.B(n_1167),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_SL g1739 ( 
.A(n_1668),
.B(n_1331),
.Y(n_1739)
);

NAND2xp5_ASAP7_75t_L g1740 ( 
.A(n_1647),
.B(n_1507),
.Y(n_1740)
);

AND2x2_ASAP7_75t_SL g1741 ( 
.A(n_1644),
.B(n_1080),
.Y(n_1741)
);

INVx1_ASAP7_75t_L g1742 ( 
.A(n_1654),
.Y(n_1742)
);

AND2x2_ASAP7_75t_L g1743 ( 
.A(n_1677),
.B(n_1061),
.Y(n_1743)
);

BUFx3_ASAP7_75t_L g1744 ( 
.A(n_1655),
.Y(n_1744)
);

INVx1_ASAP7_75t_L g1745 ( 
.A(n_1657),
.Y(n_1745)
);

INVx2_ASAP7_75t_L g1746 ( 
.A(n_1650),
.Y(n_1746)
);

INVx1_ASAP7_75t_L g1747 ( 
.A(n_1659),
.Y(n_1747)
);

AOI22xp5_ASAP7_75t_L g1748 ( 
.A1(n_1678),
.A2(n_1570),
.B1(n_1585),
.B2(n_1578),
.Y(n_1748)
);

INVx2_ASAP7_75t_SL g1749 ( 
.A(n_1699),
.Y(n_1749)
);

NAND2xp5_ASAP7_75t_SL g1750 ( 
.A(n_1656),
.B(n_1331),
.Y(n_1750)
);

AND2x2_ASAP7_75t_L g1751 ( 
.A(n_1694),
.B(n_1061),
.Y(n_1751)
);

INVx1_ASAP7_75t_L g1752 ( 
.A(n_1661),
.Y(n_1752)
);

OR2x2_ASAP7_75t_L g1753 ( 
.A(n_1691),
.B(n_1317),
.Y(n_1753)
);

AND2x2_ASAP7_75t_L g1754 ( 
.A(n_1693),
.B(n_1687),
.Y(n_1754)
);

NOR2xp33_ASAP7_75t_L g1755 ( 
.A(n_1663),
.B(n_1587),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1664),
.Y(n_1756)
);

NAND2xp5_ASAP7_75t_L g1757 ( 
.A(n_1667),
.B(n_1561),
.Y(n_1757)
);

BUFx6f_ASAP7_75t_L g1758 ( 
.A(n_1665),
.Y(n_1758)
);

AND3x4_ASAP7_75t_L g1759 ( 
.A(n_1682),
.B(n_1382),
.C(n_1357),
.Y(n_1759)
);

INVx4_ASAP7_75t_L g1760 ( 
.A(n_1666),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1679),
.Y(n_1761)
);

INVx1_ASAP7_75t_L g1762 ( 
.A(n_1669),
.Y(n_1762)
);

INVx1_ASAP7_75t_L g1763 ( 
.A(n_1674),
.Y(n_1763)
);

NAND2xp5_ASAP7_75t_L g1764 ( 
.A(n_1681),
.B(n_1175),
.Y(n_1764)
);

NAND2xp5_ASAP7_75t_SL g1765 ( 
.A(n_1684),
.B(n_1361),
.Y(n_1765)
);

BUFx6f_ASAP7_75t_L g1766 ( 
.A(n_1686),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1689),
.Y(n_1767)
);

NAND2xp5_ASAP7_75t_L g1768 ( 
.A(n_1690),
.B(n_1176),
.Y(n_1768)
);

INVx2_ASAP7_75t_L g1769 ( 
.A(n_1653),
.Y(n_1769)
);

NAND2xp5_ASAP7_75t_SL g1770 ( 
.A(n_1696),
.B(n_1361),
.Y(n_1770)
);

INVx1_ASAP7_75t_L g1771 ( 
.A(n_1653),
.Y(n_1771)
);

OR2x2_ASAP7_75t_L g1772 ( 
.A(n_1660),
.B(n_1376),
.Y(n_1772)
);

AND2x4_ASAP7_75t_L g1773 ( 
.A(n_1672),
.B(n_1452),
.Y(n_1773)
);

INVx2_ASAP7_75t_L g1774 ( 
.A(n_1653),
.Y(n_1774)
);

NAND2xp5_ASAP7_75t_SL g1775 ( 
.A(n_1696),
.B(n_1182),
.Y(n_1775)
);

INVxp33_ASAP7_75t_L g1776 ( 
.A(n_1688),
.Y(n_1776)
);

OAI22xp33_ASAP7_75t_SL g1777 ( 
.A1(n_1703),
.A2(n_1343),
.B1(n_1380),
.B2(n_1297),
.Y(n_1777)
);

NAND3xp33_ASAP7_75t_L g1778 ( 
.A(n_1703),
.B(n_1087),
.C(n_1086),
.Y(n_1778)
);

BUFx3_ASAP7_75t_L g1779 ( 
.A(n_1648),
.Y(n_1779)
);

BUFx6f_ASAP7_75t_L g1780 ( 
.A(n_1653),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1733),
.Y(n_1781)
);

CKINVDCx5p33_ASAP7_75t_R g1782 ( 
.A(n_1729),
.Y(n_1782)
);

BUFx2_ASAP7_75t_L g1783 ( 
.A(n_1723),
.Y(n_1783)
);

INVx2_ASAP7_75t_L g1784 ( 
.A(n_1728),
.Y(n_1784)
);

INVx1_ASAP7_75t_SL g1785 ( 
.A(n_1725),
.Y(n_1785)
);

INVx2_ASAP7_75t_L g1786 ( 
.A(n_1746),
.Y(n_1786)
);

AO22x2_ASAP7_75t_L g1787 ( 
.A1(n_1759),
.A2(n_1472),
.B1(n_1552),
.B2(n_1428),
.Y(n_1787)
);

AOI22xp5_ASAP7_75t_L g1788 ( 
.A1(n_1754),
.A2(n_1592),
.B1(n_1616),
.B2(n_1591),
.Y(n_1788)
);

NAND2xp5_ASAP7_75t_L g1789 ( 
.A(n_1718),
.B(n_1090),
.Y(n_1789)
);

INVx1_ASAP7_75t_L g1790 ( 
.A(n_1736),
.Y(n_1790)
);

AO22x2_ASAP7_75t_L g1791 ( 
.A1(n_1772),
.A2(n_1555),
.B1(n_1483),
.B2(n_1066),
.Y(n_1791)
);

INVx1_ASAP7_75t_L g1792 ( 
.A(n_1742),
.Y(n_1792)
);

AO22x2_ASAP7_75t_L g1793 ( 
.A1(n_1770),
.A2(n_1067),
.B1(n_1073),
.B2(n_1062),
.Y(n_1793)
);

NAND2xp5_ASAP7_75t_L g1794 ( 
.A(n_1709),
.B(n_1721),
.Y(n_1794)
);

INVx1_ASAP7_75t_L g1795 ( 
.A(n_1745),
.Y(n_1795)
);

NAND2xp5_ASAP7_75t_L g1796 ( 
.A(n_1732),
.B(n_1094),
.Y(n_1796)
);

AO22x2_ASAP7_75t_L g1797 ( 
.A1(n_1753),
.A2(n_1078),
.B1(n_1079),
.B2(n_1074),
.Y(n_1797)
);

OAI221xp5_ASAP7_75t_L g1798 ( 
.A1(n_1778),
.A2(n_1092),
.B1(n_1095),
.B2(n_1093),
.C(n_1084),
.Y(n_1798)
);

NAND2xp5_ASAP7_75t_L g1799 ( 
.A(n_1747),
.B(n_1097),
.Y(n_1799)
);

INVx1_ASAP7_75t_L g1800 ( 
.A(n_1752),
.Y(n_1800)
);

INVx2_ASAP7_75t_L g1801 ( 
.A(n_1761),
.Y(n_1801)
);

INVx1_ASAP7_75t_L g1802 ( 
.A(n_1756),
.Y(n_1802)
);

INVx1_ASAP7_75t_L g1803 ( 
.A(n_1762),
.Y(n_1803)
);

BUFx6f_ASAP7_75t_SL g1804 ( 
.A(n_1726),
.Y(n_1804)
);

INVx1_ASAP7_75t_L g1805 ( 
.A(n_1763),
.Y(n_1805)
);

INVx3_ASAP7_75t_L g1806 ( 
.A(n_1780),
.Y(n_1806)
);

INVx1_ASAP7_75t_L g1807 ( 
.A(n_1767),
.Y(n_1807)
);

NOR2xp33_ASAP7_75t_L g1808 ( 
.A(n_1717),
.B(n_1620),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1735),
.B(n_1098),
.Y(n_1809)
);

OAI221xp5_ASAP7_75t_L g1810 ( 
.A1(n_1740),
.A2(n_1099),
.B1(n_1106),
.B2(n_1103),
.C(n_1102),
.Y(n_1810)
);

OR2x2_ASAP7_75t_L g1811 ( 
.A(n_1749),
.B(n_1089),
.Y(n_1811)
);

OAI221xp5_ASAP7_75t_L g1812 ( 
.A1(n_1757),
.A2(n_1107),
.B1(n_1116),
.B2(n_1114),
.C(n_1108),
.Y(n_1812)
);

INVx1_ASAP7_75t_L g1813 ( 
.A(n_1744),
.Y(n_1813)
);

BUFx12f_ASAP7_75t_L g1814 ( 
.A(n_1705),
.Y(n_1814)
);

AO22x2_ASAP7_75t_L g1815 ( 
.A1(n_1743),
.A2(n_1119),
.B1(n_1123),
.B2(n_1117),
.Y(n_1815)
);

OAI221xp5_ASAP7_75t_L g1816 ( 
.A1(n_1777),
.A2(n_1140),
.B1(n_1145),
.B2(n_1138),
.C(n_1136),
.Y(n_1816)
);

INVx2_ASAP7_75t_L g1817 ( 
.A(n_1758),
.Y(n_1817)
);

XNOR2xp5_ASAP7_75t_L g1818 ( 
.A(n_1748),
.B(n_1077),
.Y(n_1818)
);

NOR2xp33_ASAP7_75t_L g1819 ( 
.A(n_1776),
.B(n_1096),
.Y(n_1819)
);

AO22x2_ASAP7_75t_L g1820 ( 
.A1(n_1731),
.A2(n_1146),
.B1(n_1172),
.B2(n_1160),
.Y(n_1820)
);

NAND2xp5_ASAP7_75t_SL g1821 ( 
.A(n_1735),
.B(n_1189),
.Y(n_1821)
);

INVx1_ASAP7_75t_L g1822 ( 
.A(n_1719),
.Y(n_1822)
);

AO22x1_ASAP7_75t_L g1823 ( 
.A1(n_1773),
.A2(n_1186),
.B1(n_1206),
.B2(n_1174),
.Y(n_1823)
);

INVx1_ASAP7_75t_L g1824 ( 
.A(n_1711),
.Y(n_1824)
);

AND2x2_ASAP7_75t_L g1825 ( 
.A(n_1751),
.B(n_1088),
.Y(n_1825)
);

AOI22xp5_ASAP7_75t_L g1826 ( 
.A1(n_1741),
.A2(n_1204),
.B1(n_1205),
.B2(n_1199),
.Y(n_1826)
);

INVx1_ASAP7_75t_L g1827 ( 
.A(n_1769),
.Y(n_1827)
);

AO22x2_ASAP7_75t_L g1828 ( 
.A1(n_1707),
.A2(n_1208),
.B1(n_1235),
.B2(n_1217),
.Y(n_1828)
);

NAND2x1p5_ASAP7_75t_L g1829 ( 
.A(n_1715),
.B(n_1115),
.Y(n_1829)
);

AND2x6_ASAP7_75t_L g1830 ( 
.A(n_1722),
.B(n_1755),
.Y(n_1830)
);

NAND2xp5_ASAP7_75t_L g1831 ( 
.A(n_1710),
.B(n_1127),
.Y(n_1831)
);

INVx1_ASAP7_75t_L g1832 ( 
.A(n_1774),
.Y(n_1832)
);

AO22x2_ASAP7_75t_L g1833 ( 
.A1(n_1738),
.A2(n_1401),
.B1(n_1442),
.B2(n_1212),
.Y(n_1833)
);

NOR2xp33_ASAP7_75t_L g1834 ( 
.A(n_1775),
.B(n_1105),
.Y(n_1834)
);

HB1xp67_ASAP7_75t_L g1835 ( 
.A(n_1734),
.Y(n_1835)
);

INVx1_ASAP7_75t_L g1836 ( 
.A(n_1766),
.Y(n_1836)
);

OR2x6_ASAP7_75t_L g1837 ( 
.A(n_1734),
.B(n_1128),
.Y(n_1837)
);

INVx1_ASAP7_75t_L g1838 ( 
.A(n_1766),
.Y(n_1838)
);

AND2x4_ASAP7_75t_L g1839 ( 
.A(n_1779),
.B(n_1207),
.Y(n_1839)
);

AO22x2_ASAP7_75t_L g1840 ( 
.A1(n_1739),
.A2(n_1335),
.B1(n_1358),
.B2(n_1316),
.Y(n_1840)
);

AO22x2_ASAP7_75t_L g1841 ( 
.A1(n_1750),
.A2(n_1337),
.B1(n_1562),
.B2(n_1318),
.Y(n_1841)
);

INVx2_ASAP7_75t_L g1842 ( 
.A(n_1758),
.Y(n_1842)
);

NAND2xp5_ASAP7_75t_L g1843 ( 
.A(n_1764),
.B(n_1129),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1706),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1708),
.Y(n_1845)
);

INVx1_ASAP7_75t_L g1846 ( 
.A(n_1712),
.Y(n_1846)
);

NAND2x1p5_ASAP7_75t_L g1847 ( 
.A(n_1715),
.B(n_1131),
.Y(n_1847)
);

BUFx8_ASAP7_75t_L g1848 ( 
.A(n_1720),
.Y(n_1848)
);

BUFx6f_ASAP7_75t_L g1849 ( 
.A(n_1780),
.Y(n_1849)
);

NOR2xp33_ASAP7_75t_L g1850 ( 
.A(n_1730),
.B(n_1109),
.Y(n_1850)
);

AO22x2_ASAP7_75t_L g1851 ( 
.A1(n_1765),
.A2(n_1248),
.B1(n_1273),
.B2(n_1209),
.Y(n_1851)
);

INVx1_ASAP7_75t_L g1852 ( 
.A(n_1713),
.Y(n_1852)
);

INVx2_ASAP7_75t_L g1853 ( 
.A(n_1714),
.Y(n_1853)
);

AO22x2_ASAP7_75t_L g1854 ( 
.A1(n_1724),
.A2(n_1314),
.B1(n_1210),
.B2(n_1219),
.Y(n_1854)
);

NAND2xp5_ASAP7_75t_L g1855 ( 
.A(n_1768),
.B(n_1144),
.Y(n_1855)
);

INVx1_ASAP7_75t_L g1856 ( 
.A(n_1771),
.Y(n_1856)
);

AO22x2_ASAP7_75t_L g1857 ( 
.A1(n_1737),
.A2(n_1225),
.B1(n_1281),
.B2(n_1243),
.Y(n_1857)
);

OR2x6_ASAP7_75t_L g1858 ( 
.A(n_1760),
.B(n_1158),
.Y(n_1858)
);

INVx1_ASAP7_75t_L g1859 ( 
.A(n_1716),
.Y(n_1859)
);

INVxp67_ASAP7_75t_L g1860 ( 
.A(n_1727),
.Y(n_1860)
);

HB1xp67_ASAP7_75t_L g1861 ( 
.A(n_1716),
.Y(n_1861)
);

INVx1_ASAP7_75t_L g1862 ( 
.A(n_1716),
.Y(n_1862)
);

INVxp67_ASAP7_75t_L g1863 ( 
.A(n_1717),
.Y(n_1863)
);

AO22x2_ASAP7_75t_L g1864 ( 
.A1(n_1759),
.A2(n_1213),
.B1(n_1252),
.B2(n_1242),
.Y(n_1864)
);

AND2x2_ASAP7_75t_L g1865 ( 
.A(n_1743),
.B(n_1088),
.Y(n_1865)
);

BUFx8_ASAP7_75t_L g1866 ( 
.A(n_1723),
.Y(n_1866)
);

INVx2_ASAP7_75t_L g1867 ( 
.A(n_1728),
.Y(n_1867)
);

AO22x2_ASAP7_75t_L g1868 ( 
.A1(n_1759),
.A2(n_1375),
.B1(n_1275),
.B2(n_1315),
.Y(n_1868)
);

NAND2xp5_ASAP7_75t_L g1869 ( 
.A(n_1718),
.B(n_1147),
.Y(n_1869)
);

INVx1_ASAP7_75t_L g1870 ( 
.A(n_1733),
.Y(n_1870)
);

AND2x2_ASAP7_75t_SL g1871 ( 
.A(n_1741),
.B(n_1080),
.Y(n_1871)
);

BUFx6f_ASAP7_75t_SL g1872 ( 
.A(n_1726),
.Y(n_1872)
);

INVx1_ASAP7_75t_L g1873 ( 
.A(n_1733),
.Y(n_1873)
);

INVx1_ASAP7_75t_L g1874 ( 
.A(n_1733),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1733),
.Y(n_1875)
);

NAND2xp5_ASAP7_75t_L g1876 ( 
.A(n_1718),
.B(n_1169),
.Y(n_1876)
);

AO22x2_ASAP7_75t_L g1877 ( 
.A1(n_1759),
.A2(n_1422),
.B1(n_1511),
.B2(n_1413),
.Y(n_1877)
);

BUFx8_ASAP7_75t_L g1878 ( 
.A(n_1723),
.Y(n_1878)
);

AOI22xp5_ASAP7_75t_L g1879 ( 
.A1(n_1754),
.A2(n_1229),
.B1(n_1230),
.B2(n_1224),
.Y(n_1879)
);

AO22x2_ASAP7_75t_L g1880 ( 
.A1(n_1759),
.A2(n_1396),
.B1(n_1440),
.B2(n_1377),
.Y(n_1880)
);

INVx1_ASAP7_75t_L g1881 ( 
.A(n_1733),
.Y(n_1881)
);

AOI22xp5_ASAP7_75t_L g1882 ( 
.A1(n_1754),
.A2(n_1238),
.B1(n_1239),
.B2(n_1236),
.Y(n_1882)
);

INVx1_ASAP7_75t_L g1883 ( 
.A(n_1733),
.Y(n_1883)
);

INVxp67_ASAP7_75t_L g1884 ( 
.A(n_1717),
.Y(n_1884)
);

AO22x2_ASAP7_75t_L g1885 ( 
.A1(n_1759),
.A2(n_1360),
.B1(n_1369),
.B2(n_1334),
.Y(n_1885)
);

INVx1_ASAP7_75t_L g1886 ( 
.A(n_1733),
.Y(n_1886)
);

AND2x2_ASAP7_75t_L g1887 ( 
.A(n_1743),
.B(n_1274),
.Y(n_1887)
);

INVx1_ASAP7_75t_L g1888 ( 
.A(n_1733),
.Y(n_1888)
);

BUFx8_ASAP7_75t_L g1889 ( 
.A(n_1723),
.Y(n_1889)
);

NAND2x1p5_ASAP7_75t_L g1890 ( 
.A(n_1705),
.B(n_1215),
.Y(n_1890)
);

AO22x2_ASAP7_75t_L g1891 ( 
.A1(n_1759),
.A2(n_1482),
.B1(n_1500),
.B2(n_1408),
.Y(n_1891)
);

INVx1_ASAP7_75t_L g1892 ( 
.A(n_1733),
.Y(n_1892)
);

INVx2_ASAP7_75t_L g1893 ( 
.A(n_1728),
.Y(n_1893)
);

NAND2xp5_ASAP7_75t_L g1894 ( 
.A(n_1718),
.B(n_1221),
.Y(n_1894)
);

OA22x2_ASAP7_75t_L g1895 ( 
.A1(n_1759),
.A2(n_1111),
.B1(n_1120),
.B2(n_1110),
.Y(n_1895)
);

INVx1_ASAP7_75t_L g1896 ( 
.A(n_1733),
.Y(n_1896)
);

NAND2x1p5_ASAP7_75t_L g1897 ( 
.A(n_1705),
.B(n_1256),
.Y(n_1897)
);

INVx1_ASAP7_75t_L g1898 ( 
.A(n_1733),
.Y(n_1898)
);

INVx1_ASAP7_75t_L g1899 ( 
.A(n_1733),
.Y(n_1899)
);

NAND2x1p5_ASAP7_75t_L g1900 ( 
.A(n_1705),
.B(n_1264),
.Y(n_1900)
);

AO22x2_ASAP7_75t_L g1901 ( 
.A1(n_1759),
.A2(n_1512),
.B1(n_1538),
.B2(n_1260),
.Y(n_1901)
);

NOR2xp33_ASAP7_75t_L g1902 ( 
.A(n_1709),
.B(n_1121),
.Y(n_1902)
);

INVx2_ASAP7_75t_L g1903 ( 
.A(n_1728),
.Y(n_1903)
);

AO22x2_ASAP7_75t_L g1904 ( 
.A1(n_1759),
.A2(n_1542),
.B1(n_1485),
.B2(n_1345),
.Y(n_1904)
);

CKINVDCx20_ASAP7_75t_R g1905 ( 
.A(n_1729),
.Y(n_1905)
);

AO22x2_ASAP7_75t_L g1906 ( 
.A1(n_1759),
.A2(n_1421),
.B1(n_1446),
.B2(n_1378),
.Y(n_1906)
);

NAND2x1p5_ASAP7_75t_L g1907 ( 
.A(n_1705),
.B(n_1266),
.Y(n_1907)
);

NAND2x1p5_ASAP7_75t_L g1908 ( 
.A(n_1705),
.B(n_1271),
.Y(n_1908)
);

INVx2_ASAP7_75t_SL g1909 ( 
.A(n_1773),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1735),
.B(n_1564),
.Y(n_1910)
);

INVx2_ASAP7_75t_SL g1911 ( 
.A(n_1773),
.Y(n_1911)
);

CKINVDCx5p33_ASAP7_75t_R g1912 ( 
.A(n_1729),
.Y(n_1912)
);

INVxp67_ASAP7_75t_L g1913 ( 
.A(n_1717),
.Y(n_1913)
);

NOR2xp33_ASAP7_75t_L g1914 ( 
.A(n_1709),
.B(n_1122),
.Y(n_1914)
);

NAND3xp33_ASAP7_75t_L g1915 ( 
.A(n_1709),
.B(n_1132),
.C(n_1130),
.Y(n_1915)
);

AO22x2_ASAP7_75t_L g1916 ( 
.A1(n_1759),
.A2(n_1476),
.B1(n_1323),
.B2(n_1368),
.Y(n_1916)
);

INVx1_ASAP7_75t_L g1917 ( 
.A(n_1733),
.Y(n_1917)
);

AND2x2_ASAP7_75t_SL g1918 ( 
.A(n_1741),
.B(n_1100),
.Y(n_1918)
);

INVx1_ASAP7_75t_L g1919 ( 
.A(n_1733),
.Y(n_1919)
);

INVx1_ASAP7_75t_L g1920 ( 
.A(n_1733),
.Y(n_1920)
);

CKINVDCx5p33_ASAP7_75t_R g1921 ( 
.A(n_1729),
.Y(n_1921)
);

AND2x6_ASAP7_75t_SL g1922 ( 
.A(n_1717),
.B(n_1359),
.Y(n_1922)
);

NAND2xp5_ASAP7_75t_SL g1923 ( 
.A(n_1871),
.B(n_1244),
.Y(n_1923)
);

NAND2xp33_ASAP7_75t_SL g1924 ( 
.A(n_1782),
.B(n_1133),
.Y(n_1924)
);

NAND2xp5_ASAP7_75t_L g1925 ( 
.A(n_1794),
.B(n_1272),
.Y(n_1925)
);

NAND2xp5_ASAP7_75t_SL g1926 ( 
.A(n_1918),
.B(n_1259),
.Y(n_1926)
);

NAND2xp33_ASAP7_75t_SL g1927 ( 
.A(n_1912),
.B(n_1183),
.Y(n_1927)
);

NAND2xp5_ASAP7_75t_SL g1928 ( 
.A(n_1863),
.B(n_1267),
.Y(n_1928)
);

NAND2xp33_ASAP7_75t_SL g1929 ( 
.A(n_1921),
.B(n_1185),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_L g1930 ( 
.A(n_1902),
.B(n_1293),
.Y(n_1930)
);

NAND2xp5_ASAP7_75t_SL g1931 ( 
.A(n_1884),
.B(n_1913),
.Y(n_1931)
);

NAND2xp5_ASAP7_75t_L g1932 ( 
.A(n_1914),
.B(n_1325),
.Y(n_1932)
);

NAND2xp5_ASAP7_75t_SL g1933 ( 
.A(n_1785),
.B(n_1283),
.Y(n_1933)
);

NAND2xp33_ASAP7_75t_SL g1934 ( 
.A(n_1804),
.B(n_1187),
.Y(n_1934)
);

NAND2xp33_ASAP7_75t_SL g1935 ( 
.A(n_1872),
.B(n_1226),
.Y(n_1935)
);

NAND2xp5_ASAP7_75t_SL g1936 ( 
.A(n_1860),
.B(n_1294),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_SL g1937 ( 
.A(n_1789),
.B(n_1869),
.Y(n_1937)
);

AND2x2_ASAP7_75t_L g1938 ( 
.A(n_1865),
.B(n_1274),
.Y(n_1938)
);

NAND2xp33_ASAP7_75t_SL g1939 ( 
.A(n_1887),
.B(n_1241),
.Y(n_1939)
);

NAND2xp33_ASAP7_75t_SL g1940 ( 
.A(n_1849),
.B(n_1251),
.Y(n_1940)
);

NAND2xp5_ASAP7_75t_SL g1941 ( 
.A(n_1876),
.B(n_1298),
.Y(n_1941)
);

NAND2xp5_ASAP7_75t_SL g1942 ( 
.A(n_1894),
.B(n_1302),
.Y(n_1942)
);

NAND2xp33_ASAP7_75t_SL g1943 ( 
.A(n_1849),
.B(n_1280),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1879),
.B(n_1309),
.Y(n_1944)
);

NAND2xp5_ASAP7_75t_SL g1945 ( 
.A(n_1882),
.B(n_1312),
.Y(n_1945)
);

NAND2xp5_ASAP7_75t_SL g1946 ( 
.A(n_1850),
.B(n_1319),
.Y(n_1946)
);

NAND2xp5_ASAP7_75t_SL g1947 ( 
.A(n_1788),
.B(n_1324),
.Y(n_1947)
);

AND2x2_ASAP7_75t_L g1948 ( 
.A(n_1825),
.B(n_1313),
.Y(n_1948)
);

NAND2xp5_ASAP7_75t_L g1949 ( 
.A(n_1796),
.B(n_1781),
.Y(n_1949)
);

NAND2xp5_ASAP7_75t_SL g1950 ( 
.A(n_1834),
.B(n_1328),
.Y(n_1950)
);

NAND2xp5_ASAP7_75t_SL g1951 ( 
.A(n_1915),
.B(n_1340),
.Y(n_1951)
);

NAND2xp33_ASAP7_75t_SL g1952 ( 
.A(n_1905),
.B(n_1303),
.Y(n_1952)
);

NAND2xp5_ASAP7_75t_SL g1953 ( 
.A(n_1790),
.B(n_1792),
.Y(n_1953)
);

NAND2xp5_ASAP7_75t_SL g1954 ( 
.A(n_1795),
.B(n_1347),
.Y(n_1954)
);

NAND2xp33_ASAP7_75t_SL g1955 ( 
.A(n_1861),
.B(n_1350),
.Y(n_1955)
);

NAND2xp5_ASAP7_75t_SL g1956 ( 
.A(n_1800),
.B(n_1351),
.Y(n_1956)
);

NAND2xp5_ASAP7_75t_L g1957 ( 
.A(n_1802),
.B(n_1326),
.Y(n_1957)
);

NOR2xp33_ASAP7_75t_L g1958 ( 
.A(n_1808),
.B(n_1379),
.Y(n_1958)
);

NAND2xp33_ASAP7_75t_SL g1959 ( 
.A(n_1909),
.B(n_1403),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_SL g1960 ( 
.A(n_1803),
.B(n_1355),
.Y(n_1960)
);

NAND2xp5_ASAP7_75t_SL g1961 ( 
.A(n_1805),
.B(n_1363),
.Y(n_1961)
);

NAND2xp33_ASAP7_75t_SL g1962 ( 
.A(n_1911),
.B(n_1411),
.Y(n_1962)
);

NAND2xp5_ASAP7_75t_SL g1963 ( 
.A(n_1807),
.B(n_1366),
.Y(n_1963)
);

NAND2xp5_ASAP7_75t_SL g1964 ( 
.A(n_1870),
.B(n_1367),
.Y(n_1964)
);

NAND2xp5_ASAP7_75t_L g1965 ( 
.A(n_1873),
.B(n_1329),
.Y(n_1965)
);

NAND2xp33_ASAP7_75t_SL g1966 ( 
.A(n_1783),
.B(n_1420),
.Y(n_1966)
);

NAND2xp5_ASAP7_75t_L g1967 ( 
.A(n_1874),
.B(n_1344),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_SL g1968 ( 
.A(n_1875),
.B(n_1371),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_L g1969 ( 
.A(n_1881),
.B(n_1370),
.Y(n_1969)
);

AND2x4_ASAP7_75t_L g1970 ( 
.A(n_1817),
.B(n_1373),
.Y(n_1970)
);

NAND2xp5_ASAP7_75t_SL g1971 ( 
.A(n_1883),
.B(n_1392),
.Y(n_1971)
);

NAND2xp5_ASAP7_75t_SL g1972 ( 
.A(n_1886),
.B(n_1400),
.Y(n_1972)
);

NAND2xp5_ASAP7_75t_SL g1973 ( 
.A(n_1888),
.B(n_1402),
.Y(n_1973)
);

NAND2xp33_ASAP7_75t_SL g1974 ( 
.A(n_1835),
.B(n_1434),
.Y(n_1974)
);

NAND2xp5_ASAP7_75t_SL g1975 ( 
.A(n_1892),
.B(n_1407),
.Y(n_1975)
);

NAND2xp5_ASAP7_75t_SL g1976 ( 
.A(n_1896),
.B(n_1409),
.Y(n_1976)
);

NAND2xp5_ASAP7_75t_SL g1977 ( 
.A(n_1898),
.B(n_1431),
.Y(n_1977)
);

NAND2xp5_ASAP7_75t_SL g1978 ( 
.A(n_1899),
.B(n_1449),
.Y(n_1978)
);

NAND2xp5_ASAP7_75t_SL g1979 ( 
.A(n_1917),
.B(n_1919),
.Y(n_1979)
);

NOR2xp33_ASAP7_75t_L g1980 ( 
.A(n_1819),
.B(n_1466),
.Y(n_1980)
);

AND2x2_ASAP7_75t_L g1981 ( 
.A(n_1811),
.B(n_1313),
.Y(n_1981)
);

NAND2xp5_ASAP7_75t_SL g1982 ( 
.A(n_1920),
.B(n_1461),
.Y(n_1982)
);

NAND2xp33_ASAP7_75t_SL g1983 ( 
.A(n_1813),
.B(n_1520),
.Y(n_1983)
);

NAND2xp5_ASAP7_75t_SL g1984 ( 
.A(n_1826),
.B(n_1462),
.Y(n_1984)
);

NAND2xp5_ASAP7_75t_SL g1985 ( 
.A(n_1836),
.B(n_1474),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_SL g1986 ( 
.A(n_1838),
.B(n_1479),
.Y(n_1986)
);

NAND2xp5_ASAP7_75t_SL g1987 ( 
.A(n_1809),
.B(n_1843),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1855),
.B(n_1387),
.Y(n_1988)
);

NAND2xp5_ASAP7_75t_L g1989 ( 
.A(n_1830),
.B(n_1390),
.Y(n_1989)
);

NAND2xp5_ASAP7_75t_L g1990 ( 
.A(n_1830),
.B(n_1393),
.Y(n_1990)
);

NAND2xp5_ASAP7_75t_SL g1991 ( 
.A(n_1842),
.B(n_1480),
.Y(n_1991)
);

NAND2xp5_ASAP7_75t_SL g1992 ( 
.A(n_1784),
.B(n_1494),
.Y(n_1992)
);

NAND2xp5_ASAP7_75t_SL g1993 ( 
.A(n_1786),
.B(n_1498),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_SL g1994 ( 
.A(n_1801),
.B(n_1504),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1830),
.B(n_1394),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_SL g1996 ( 
.A(n_1867),
.B(n_1517),
.Y(n_1996)
);

NAND2xp5_ASAP7_75t_SL g1997 ( 
.A(n_1893),
.B(n_1523),
.Y(n_1997)
);

NAND2xp5_ASAP7_75t_SL g1998 ( 
.A(n_1903),
.B(n_1527),
.Y(n_1998)
);

NAND2xp33_ASAP7_75t_SL g1999 ( 
.A(n_1859),
.B(n_1525),
.Y(n_1999)
);

AND2x4_ASAP7_75t_L g2000 ( 
.A(n_1822),
.B(n_1427),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1799),
.B(n_1831),
.Y(n_2001)
);

NAND2xp33_ASAP7_75t_SL g2002 ( 
.A(n_1862),
.B(n_1531),
.Y(n_2002)
);

NAND2xp5_ASAP7_75t_SL g2003 ( 
.A(n_1853),
.B(n_1532),
.Y(n_2003)
);

NAND2xp5_ASAP7_75t_SL g2004 ( 
.A(n_1844),
.B(n_1064),
.Y(n_2004)
);

NAND2xp5_ASAP7_75t_SL g2005 ( 
.A(n_1845),
.B(n_1064),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1846),
.B(n_1488),
.Y(n_2006)
);

NAND2xp5_ASAP7_75t_SL g2007 ( 
.A(n_1852),
.B(n_1424),
.Y(n_2007)
);

NAND2xp5_ASAP7_75t_SL g2008 ( 
.A(n_1856),
.B(n_1426),
.Y(n_2008)
);

NAND2xp5_ASAP7_75t_SL g2009 ( 
.A(n_1824),
.B(n_1429),
.Y(n_2009)
);

NAND2xp33_ASAP7_75t_SL g2010 ( 
.A(n_1806),
.B(n_1821),
.Y(n_2010)
);

NAND2xp5_ASAP7_75t_SL g2011 ( 
.A(n_1827),
.B(n_1832),
.Y(n_2011)
);

NAND2xp5_ASAP7_75t_SL g2012 ( 
.A(n_1839),
.B(n_1436),
.Y(n_2012)
);

NAND2xp5_ASAP7_75t_L g2013 ( 
.A(n_1854),
.B(n_1445),
.Y(n_2013)
);

AND2x4_ASAP7_75t_L g2014 ( 
.A(n_1858),
.B(n_1837),
.Y(n_2014)
);

NAND2xp33_ASAP7_75t_SL g2015 ( 
.A(n_1910),
.B(n_1533),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_SL g2016 ( 
.A(n_1890),
.B(n_1897),
.Y(n_2016)
);

NAND2xp5_ASAP7_75t_SL g2017 ( 
.A(n_1900),
.B(n_1463),
.Y(n_2017)
);

NAND2xp5_ASAP7_75t_SL g2018 ( 
.A(n_1907),
.B(n_1473),
.Y(n_2018)
);

AND2x2_ASAP7_75t_L g2019 ( 
.A(n_1797),
.B(n_1478),
.Y(n_2019)
);

NAND2xp5_ASAP7_75t_SL g2020 ( 
.A(n_1908),
.B(n_1487),
.Y(n_2020)
);

NAND2xp5_ASAP7_75t_SL g2021 ( 
.A(n_1814),
.B(n_1502),
.Y(n_2021)
);

NAND2xp5_ASAP7_75t_SL g2022 ( 
.A(n_1895),
.B(n_1505),
.Y(n_2022)
);

NAND2xp33_ASAP7_75t_SL g2023 ( 
.A(n_1818),
.B(n_1539),
.Y(n_2023)
);

NAND2xp5_ASAP7_75t_SL g2024 ( 
.A(n_1829),
.B(n_1530),
.Y(n_2024)
);

AND2x4_ASAP7_75t_L g2025 ( 
.A(n_1793),
.B(n_1497),
.Y(n_2025)
);

NAND2xp33_ASAP7_75t_SL g2026 ( 
.A(n_1833),
.B(n_1134),
.Y(n_2026)
);

NAND2xp5_ASAP7_75t_L g2027 ( 
.A(n_1823),
.B(n_1840),
.Y(n_2027)
);

NAND2xp5_ASAP7_75t_SL g2028 ( 
.A(n_1847),
.B(n_1535),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1866),
.B(n_1536),
.Y(n_2029)
);

NAND2xp33_ASAP7_75t_SL g2030 ( 
.A(n_1857),
.B(n_1137),
.Y(n_2030)
);

NAND2xp5_ASAP7_75t_SL g2031 ( 
.A(n_1878),
.B(n_1544),
.Y(n_2031)
);

NAND2xp5_ASAP7_75t_SL g2032 ( 
.A(n_1889),
.B(n_1550),
.Y(n_2032)
);

NAND2xp33_ASAP7_75t_SL g2033 ( 
.A(n_1841),
.B(n_1139),
.Y(n_2033)
);

NAND2xp5_ASAP7_75t_SL g2034 ( 
.A(n_1848),
.B(n_1346),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1815),
.B(n_1346),
.Y(n_2035)
);

NAND2xp5_ASAP7_75t_L g2036 ( 
.A(n_1851),
.B(n_1521),
.Y(n_2036)
);

NAND2xp33_ASAP7_75t_SL g2037 ( 
.A(n_1864),
.B(n_1141),
.Y(n_2037)
);

NAND2xp5_ASAP7_75t_SL g2038 ( 
.A(n_1868),
.B(n_1346),
.Y(n_2038)
);

NAND2xp33_ASAP7_75t_SL g2039 ( 
.A(n_1877),
.B(n_1142),
.Y(n_2039)
);

NAND2xp5_ASAP7_75t_L g2040 ( 
.A(n_1820),
.B(n_1537),
.Y(n_2040)
);

NAND2xp5_ASAP7_75t_SL g2041 ( 
.A(n_1880),
.B(n_1346),
.Y(n_2041)
);

NAND2xp5_ASAP7_75t_SL g2042 ( 
.A(n_1885),
.B(n_1346),
.Y(n_2042)
);

NAND2xp5_ASAP7_75t_L g2043 ( 
.A(n_1828),
.B(n_1509),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_SL g2044 ( 
.A(n_1891),
.B(n_1100),
.Y(n_2044)
);

NAND2xp33_ASAP7_75t_SL g2045 ( 
.A(n_1901),
.B(n_1143),
.Y(n_2045)
);

AND2x4_ASAP7_75t_L g2046 ( 
.A(n_1798),
.B(n_1508),
.Y(n_2046)
);

NAND2xp5_ASAP7_75t_SL g2047 ( 
.A(n_1904),
.B(n_1100),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_SL g2048 ( 
.A(n_1906),
.B(n_1101),
.Y(n_2048)
);

NAND2xp5_ASAP7_75t_SL g2049 ( 
.A(n_1916),
.B(n_1101),
.Y(n_2049)
);

AND3x1_ASAP7_75t_L g2050 ( 
.A(n_1787),
.B(n_1549),
.C(n_1546),
.Y(n_2050)
);

NAND2xp5_ASAP7_75t_SL g2051 ( 
.A(n_1922),
.B(n_1101),
.Y(n_2051)
);

NAND2xp5_ASAP7_75t_SL g2052 ( 
.A(n_1791),
.B(n_1237),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_SL g2053 ( 
.A(n_1816),
.B(n_1237),
.Y(n_2053)
);

NAND2xp5_ASAP7_75t_L g2054 ( 
.A(n_1810),
.B(n_1509),
.Y(n_2054)
);

NAND2xp5_ASAP7_75t_SL g2055 ( 
.A(n_1812),
.B(n_1237),
.Y(n_2055)
);

NAND2xp5_ASAP7_75t_SL g2056 ( 
.A(n_1871),
.B(n_1261),
.Y(n_2056)
);

NAND2xp5_ASAP7_75t_L g2057 ( 
.A(n_1794),
.B(n_1509),
.Y(n_2057)
);

NAND2xp5_ASAP7_75t_SL g2058 ( 
.A(n_1871),
.B(n_1261),
.Y(n_2058)
);

NAND2xp5_ASAP7_75t_SL g2059 ( 
.A(n_1871),
.B(n_1261),
.Y(n_2059)
);

NAND2xp5_ASAP7_75t_L g2060 ( 
.A(n_1794),
.B(n_1548),
.Y(n_2060)
);

NAND2xp5_ASAP7_75t_SL g2061 ( 
.A(n_1871),
.B(n_1265),
.Y(n_2061)
);

NAND2xp5_ASAP7_75t_L g2062 ( 
.A(n_1794),
.B(n_1548),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_SL g2063 ( 
.A(n_1871),
.B(n_1265),
.Y(n_2063)
);

NAND2xp5_ASAP7_75t_SL g2064 ( 
.A(n_1871),
.B(n_1265),
.Y(n_2064)
);

NAND2xp5_ASAP7_75t_SL g2065 ( 
.A(n_1871),
.B(n_1268),
.Y(n_2065)
);

NAND2xp5_ASAP7_75t_SL g2066 ( 
.A(n_1871),
.B(n_1268),
.Y(n_2066)
);

NAND2xp33_ASAP7_75t_SL g2067 ( 
.A(n_1782),
.B(n_1148),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_SL g2068 ( 
.A(n_1871),
.B(n_1268),
.Y(n_2068)
);

NAND2xp5_ASAP7_75t_SL g2069 ( 
.A(n_1871),
.B(n_1295),
.Y(n_2069)
);

NAND2xp5_ASAP7_75t_SL g2070 ( 
.A(n_1871),
.B(n_1295),
.Y(n_2070)
);

NAND2xp33_ASAP7_75t_SL g2071 ( 
.A(n_1782),
.B(n_1150),
.Y(n_2071)
);

NAND2xp5_ASAP7_75t_SL g2072 ( 
.A(n_1871),
.B(n_1295),
.Y(n_2072)
);

NAND2xp33_ASAP7_75t_SL g2073 ( 
.A(n_1782),
.B(n_1151),
.Y(n_2073)
);

NAND2xp5_ASAP7_75t_L g2074 ( 
.A(n_1794),
.B(n_1548),
.Y(n_2074)
);

NAND2xp5_ASAP7_75t_SL g2075 ( 
.A(n_1871),
.B(n_1475),
.Y(n_2075)
);

NAND2xp33_ASAP7_75t_SL g2076 ( 
.A(n_1782),
.B(n_1152),
.Y(n_2076)
);

NAND2xp5_ASAP7_75t_L g2077 ( 
.A(n_1794),
.B(n_1548),
.Y(n_2077)
);

NAND2xp5_ASAP7_75t_SL g2078 ( 
.A(n_1871),
.B(n_1475),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_SL g2079 ( 
.A(n_1871),
.B(n_1475),
.Y(n_2079)
);

NAND2xp5_ASAP7_75t_L g2080 ( 
.A(n_1794),
.B(n_1490),
.Y(n_2080)
);

NAND2xp5_ASAP7_75t_SL g2081 ( 
.A(n_1871),
.B(n_1490),
.Y(n_2081)
);

NAND2xp5_ASAP7_75t_SL g2082 ( 
.A(n_1871),
.B(n_1490),
.Y(n_2082)
);

NOR2xp33_ASAP7_75t_L g2083 ( 
.A(n_1863),
.B(n_1157),
.Y(n_2083)
);

NAND2xp5_ASAP7_75t_SL g2084 ( 
.A(n_1871),
.B(n_1565),
.Y(n_2084)
);

NAND2xp5_ASAP7_75t_L g2085 ( 
.A(n_1794),
.B(n_1565),
.Y(n_2085)
);

NAND2xp33_ASAP7_75t_SL g2086 ( 
.A(n_1782),
.B(n_1162),
.Y(n_2086)
);

NAND2xp5_ASAP7_75t_SL g2087 ( 
.A(n_1871),
.B(n_1565),
.Y(n_2087)
);

NAND2xp33_ASAP7_75t_R g2088 ( 
.A(n_1783),
.B(n_1168),
.Y(n_2088)
);

NAND2xp33_ASAP7_75t_SL g2089 ( 
.A(n_1782),
.B(n_1178),
.Y(n_2089)
);

NAND2xp5_ASAP7_75t_SL g2090 ( 
.A(n_1871),
.B(n_1180),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_SL g2091 ( 
.A(n_1871),
.B(n_1184),
.Y(n_2091)
);

NAND2xp5_ASAP7_75t_SL g2092 ( 
.A(n_1871),
.B(n_1188),
.Y(n_2092)
);

NAND2xp5_ASAP7_75t_SL g2093 ( 
.A(n_1871),
.B(n_1191),
.Y(n_2093)
);

NAND2xp33_ASAP7_75t_SL g2094 ( 
.A(n_1782),
.B(n_1194),
.Y(n_2094)
);

AND2x2_ASAP7_75t_L g2095 ( 
.A(n_1863),
.B(n_1478),
.Y(n_2095)
);

NAND2xp5_ASAP7_75t_SL g2096 ( 
.A(n_1871),
.B(n_1195),
.Y(n_2096)
);

NAND2xp33_ASAP7_75t_SL g2097 ( 
.A(n_1782),
.B(n_1196),
.Y(n_2097)
);

NAND2xp5_ASAP7_75t_SL g2098 ( 
.A(n_1871),
.B(n_1197),
.Y(n_2098)
);

NAND2xp33_ASAP7_75t_SL g2099 ( 
.A(n_1782),
.B(n_1198),
.Y(n_2099)
);

NAND2xp5_ASAP7_75t_SL g2100 ( 
.A(n_1871),
.B(n_1200),
.Y(n_2100)
);

NAND2xp5_ASAP7_75t_SL g2101 ( 
.A(n_1871),
.B(n_1201),
.Y(n_2101)
);

NAND2xp5_ASAP7_75t_L g2102 ( 
.A(n_1794),
.B(n_1203),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_SL g2103 ( 
.A(n_1871),
.B(n_1214),
.Y(n_2103)
);

NAND2xp33_ASAP7_75t_SL g2104 ( 
.A(n_1782),
.B(n_1216),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_SL g2105 ( 
.A(n_1871),
.B(n_1218),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_SL g2106 ( 
.A(n_1871),
.B(n_1220),
.Y(n_2106)
);

NAND2xp5_ASAP7_75t_SL g2107 ( 
.A(n_1871),
.B(n_1228),
.Y(n_2107)
);

NAND2xp5_ASAP7_75t_SL g2108 ( 
.A(n_1871),
.B(n_1231),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_SL g2109 ( 
.A(n_1871),
.B(n_1233),
.Y(n_2109)
);

NAND2xp5_ASAP7_75t_SL g2110 ( 
.A(n_1871),
.B(n_1234),
.Y(n_2110)
);

NAND2xp5_ASAP7_75t_SL g2111 ( 
.A(n_1871),
.B(n_1240),
.Y(n_2111)
);

AND2x4_ASAP7_75t_L g2112 ( 
.A(n_1817),
.B(n_1510),
.Y(n_2112)
);

NAND2xp5_ASAP7_75t_SL g2113 ( 
.A(n_1871),
.B(n_1246),
.Y(n_2113)
);

NAND2xp5_ASAP7_75t_L g2114 ( 
.A(n_1794),
.B(n_1247),
.Y(n_2114)
);

NAND2xp33_ASAP7_75t_SL g2115 ( 
.A(n_1782),
.B(n_1249),
.Y(n_2115)
);

NAND2xp5_ASAP7_75t_SL g2116 ( 
.A(n_1871),
.B(n_1250),
.Y(n_2116)
);

NAND2xp5_ASAP7_75t_SL g2117 ( 
.A(n_1871),
.B(n_1253),
.Y(n_2117)
);

NAND2xp5_ASAP7_75t_SL g2118 ( 
.A(n_1871),
.B(n_1254),
.Y(n_2118)
);

NAND2xp5_ASAP7_75t_SL g2119 ( 
.A(n_1871),
.B(n_1255),
.Y(n_2119)
);

NAND2xp33_ASAP7_75t_SL g2120 ( 
.A(n_1782),
.B(n_1258),
.Y(n_2120)
);

NAND2xp5_ASAP7_75t_SL g2121 ( 
.A(n_1871),
.B(n_1262),
.Y(n_2121)
);

NAND2xp33_ASAP7_75t_SL g2122 ( 
.A(n_1782),
.B(n_1263),
.Y(n_2122)
);

INVx1_ASAP7_75t_L g2123 ( 
.A(n_1970),
.Y(n_2123)
);

AND2x2_ASAP7_75t_L g2124 ( 
.A(n_1980),
.B(n_1540),
.Y(n_2124)
);

INVx2_ASAP7_75t_L g2125 ( 
.A(n_2000),
.Y(n_2125)
);

OAI21x1_ASAP7_75t_L g2126 ( 
.A1(n_2011),
.A2(n_1171),
.B(n_1159),
.Y(n_2126)
);

AO21x1_ASAP7_75t_L g2127 ( 
.A1(n_1930),
.A2(n_1232),
.B(n_1222),
.Y(n_2127)
);

NOR4xp25_ASAP7_75t_L g2128 ( 
.A(n_1958),
.B(n_1932),
.C(n_2035),
.D(n_2038),
.Y(n_2128)
);

OAI21x1_ASAP7_75t_L g2129 ( 
.A1(n_2057),
.A2(n_1296),
.B(n_1291),
.Y(n_2129)
);

NAND2xp5_ASAP7_75t_L g2130 ( 
.A(n_2102),
.B(n_1269),
.Y(n_2130)
);

INVx1_ASAP7_75t_L g2131 ( 
.A(n_1970),
.Y(n_2131)
);

INVx8_ASAP7_75t_L g2132 ( 
.A(n_2014),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_2095),
.B(n_1540),
.Y(n_2133)
);

AOI221xp5_ASAP7_75t_L g2134 ( 
.A1(n_2050),
.A2(n_1277),
.B1(n_1282),
.B2(n_1278),
.C(n_1270),
.Y(n_2134)
);

BUFx2_ASAP7_75t_SL g2135 ( 
.A(n_2014),
.Y(n_2135)
);

AOI21xp5_ASAP7_75t_L g2136 ( 
.A1(n_2001),
.A2(n_1937),
.B(n_1987),
.Y(n_2136)
);

HB1xp67_ASAP7_75t_L g2137 ( 
.A(n_2112),
.Y(n_2137)
);

AOI21xp5_ASAP7_75t_L g2138 ( 
.A1(n_1949),
.A2(n_1925),
.B(n_2060),
.Y(n_2138)
);

OAI21x1_ASAP7_75t_L g2139 ( 
.A1(n_2062),
.A2(n_1435),
.B(n_1311),
.Y(n_2139)
);

NAND2xp5_ASAP7_75t_L g2140 ( 
.A(n_2114),
.B(n_2080),
.Y(n_2140)
);

AOI21xp33_ASAP7_75t_L g2141 ( 
.A1(n_2083),
.A2(n_1286),
.B(n_1284),
.Y(n_2141)
);

NAND2xp5_ASAP7_75t_L g2142 ( 
.A(n_2085),
.B(n_1287),
.Y(n_2142)
);

NAND2xp5_ASAP7_75t_L g2143 ( 
.A(n_2074),
.B(n_1288),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_2077),
.B(n_1289),
.Y(n_2144)
);

AOI21xp5_ASAP7_75t_L g2145 ( 
.A1(n_1953),
.A2(n_1979),
.B(n_1950),
.Y(n_2145)
);

NOR3xp33_ASAP7_75t_SL g2146 ( 
.A(n_2088),
.B(n_1300),
.C(n_1292),
.Y(n_2146)
);

OAI21x1_ASAP7_75t_L g2147 ( 
.A1(n_1989),
.A2(n_706),
.B(n_704),
.Y(n_2147)
);

INVx1_ASAP7_75t_L g2148 ( 
.A(n_2112),
.Y(n_2148)
);

AOI21x1_ASAP7_75t_SL g2149 ( 
.A1(n_1990),
.A2(n_1177),
.B(n_1299),
.Y(n_2149)
);

A2O1A1Ixp33_ASAP7_75t_L g2150 ( 
.A1(n_1995),
.A2(n_1304),
.B(n_1305),
.C(n_1301),
.Y(n_2150)
);

INVxp67_ASAP7_75t_SL g2151 ( 
.A(n_1931),
.Y(n_2151)
);

AOI21xp5_ASAP7_75t_L g2152 ( 
.A1(n_1946),
.A2(n_709),
.B(n_707),
.Y(n_2152)
);

AOI211x1_ASAP7_75t_L g2153 ( 
.A1(n_2022),
.A2(n_1307),
.B(n_1310),
.C(n_1306),
.Y(n_2153)
);

INVx3_ASAP7_75t_L g2154 ( 
.A(n_2000),
.Y(n_2154)
);

NAND2xp5_ASAP7_75t_L g2155 ( 
.A(n_1988),
.B(n_1320),
.Y(n_2155)
);

OA21x2_ASAP7_75t_L g2156 ( 
.A1(n_1957),
.A2(n_1327),
.B(n_1321),
.Y(n_2156)
);

AO31x2_ASAP7_75t_L g2157 ( 
.A1(n_2013),
.A2(n_711),
.A3(n_712),
.B(n_710),
.Y(n_2157)
);

OAI21x1_ASAP7_75t_L g2158 ( 
.A1(n_1965),
.A2(n_714),
.B(n_713),
.Y(n_2158)
);

AO21x2_ASAP7_75t_L g2159 ( 
.A1(n_1941),
.A2(n_719),
.B(n_718),
.Y(n_2159)
);

NAND3x1_ASAP7_75t_L g2160 ( 
.A(n_2027),
.B(n_1332),
.C(n_1330),
.Y(n_2160)
);

OAI22xp5_ASAP7_75t_L g2161 ( 
.A1(n_1923),
.A2(n_1336),
.B1(n_1338),
.B2(n_1333),
.Y(n_2161)
);

OAI22xp5_ASAP7_75t_L g2162 ( 
.A1(n_1926),
.A2(n_2058),
.B1(n_2059),
.B2(n_2056),
.Y(n_2162)
);

INVx1_ASAP7_75t_L g2163 ( 
.A(n_2006),
.Y(n_2163)
);

OAI21x1_ASAP7_75t_L g2164 ( 
.A1(n_1967),
.A2(n_726),
.B(n_725),
.Y(n_2164)
);

AOI21xp5_ASAP7_75t_L g2165 ( 
.A1(n_1942),
.A2(n_732),
.B(n_730),
.Y(n_2165)
);

NOR2x1p5_ASAP7_75t_L g2166 ( 
.A(n_2040),
.B(n_1339),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_SL g2167 ( 
.A(n_1939),
.B(n_1348),
.Y(n_2167)
);

OAI21x1_ASAP7_75t_L g2168 ( 
.A1(n_1969),
.A2(n_736),
.B(n_733),
.Y(n_2168)
);

AO21x2_ASAP7_75t_L g2169 ( 
.A1(n_1951),
.A2(n_738),
.B(n_737),
.Y(n_2169)
);

INVx1_ASAP7_75t_SL g2170 ( 
.A(n_1966),
.Y(n_2170)
);

AOI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_1954),
.A2(n_740),
.B(n_739),
.Y(n_2171)
);

OAI21x1_ASAP7_75t_L g2172 ( 
.A1(n_1992),
.A2(n_745),
.B(n_744),
.Y(n_2172)
);

OA21x2_ASAP7_75t_L g2173 ( 
.A1(n_1993),
.A2(n_1353),
.B(n_1352),
.Y(n_2173)
);

AOI21xp5_ASAP7_75t_L g2174 ( 
.A1(n_1956),
.A2(n_751),
.B(n_748),
.Y(n_2174)
);

OAI21x1_ASAP7_75t_L g2175 ( 
.A1(n_1994),
.A2(n_1997),
.B(n_1996),
.Y(n_2175)
);

AOI21xp5_ASAP7_75t_L g2176 ( 
.A1(n_1960),
.A2(n_753),
.B(n_752),
.Y(n_2176)
);

AOI211x1_ASAP7_75t_L g2177 ( 
.A1(n_2041),
.A2(n_1364),
.B(n_1365),
.C(n_1362),
.Y(n_2177)
);

NAND3xp33_ASAP7_75t_L g2178 ( 
.A(n_2023),
.B(n_1381),
.C(n_1374),
.Y(n_2178)
);

NAND2xp5_ASAP7_75t_L g2179 ( 
.A(n_1938),
.B(n_1383),
.Y(n_2179)
);

NAND2x1p5_ASAP7_75t_L g2180 ( 
.A(n_2016),
.B(n_756),
.Y(n_2180)
);

OAI21x1_ASAP7_75t_SL g2181 ( 
.A1(n_2036),
.A2(n_759),
.B(n_758),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_2006),
.Y(n_2182)
);

NAND2xp5_ASAP7_75t_L g2183 ( 
.A(n_1948),
.B(n_1384),
.Y(n_2183)
);

INVx2_ASAP7_75t_SL g2184 ( 
.A(n_1981),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_2061),
.B(n_1385),
.Y(n_2185)
);

OR2x6_ASAP7_75t_L g2186 ( 
.A(n_2044),
.B(n_3),
.Y(n_2186)
);

OAI21x1_ASAP7_75t_L g2187 ( 
.A1(n_1998),
.A2(n_762),
.B(n_760),
.Y(n_2187)
);

AOI21xp5_ASAP7_75t_L g2188 ( 
.A1(n_1961),
.A2(n_764),
.B(n_763),
.Y(n_2188)
);

OAI21x1_ASAP7_75t_L g2189 ( 
.A1(n_1991),
.A2(n_767),
.B(n_765),
.Y(n_2189)
);

AOI21xp5_ASAP7_75t_L g2190 ( 
.A1(n_1963),
.A2(n_772),
.B(n_771),
.Y(n_2190)
);

OAI21x1_ASAP7_75t_L g2191 ( 
.A1(n_2009),
.A2(n_776),
.B(n_774),
.Y(n_2191)
);

NAND2xp5_ASAP7_75t_L g2192 ( 
.A(n_2063),
.B(n_1386),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_2064),
.B(n_1388),
.Y(n_2193)
);

OA21x2_ASAP7_75t_L g2194 ( 
.A1(n_2007),
.A2(n_1395),
.B(n_1389),
.Y(n_2194)
);

OR2x2_ASAP7_75t_L g2195 ( 
.A(n_1924),
.B(n_1397),
.Y(n_2195)
);

BUFx2_ASAP7_75t_L g2196 ( 
.A(n_1940),
.Y(n_2196)
);

OAI21x1_ASAP7_75t_L g2197 ( 
.A1(n_2003),
.A2(n_1986),
.B(n_1985),
.Y(n_2197)
);

OR2x2_ASAP7_75t_L g2198 ( 
.A(n_1927),
.B(n_1929),
.Y(n_2198)
);

BUFx6f_ASAP7_75t_L g2199 ( 
.A(n_2025),
.Y(n_2199)
);

INVx1_ASAP7_75t_L g2200 ( 
.A(n_2043),
.Y(n_2200)
);

AOI21xp5_ASAP7_75t_L g2201 ( 
.A1(n_1964),
.A2(n_779),
.B(n_777),
.Y(n_2201)
);

NAND3x1_ASAP7_75t_L g2202 ( 
.A(n_2019),
.B(n_1404),
.C(n_1399),
.Y(n_2202)
);

NAND2xp5_ASAP7_75t_L g2203 ( 
.A(n_2065),
.B(n_1406),
.Y(n_2203)
);

OR2x2_ASAP7_75t_L g2204 ( 
.A(n_1952),
.B(n_1410),
.Y(n_2204)
);

INVx1_ASAP7_75t_L g2205 ( 
.A(n_2054),
.Y(n_2205)
);

CKINVDCx5p33_ASAP7_75t_R g2206 ( 
.A(n_1934),
.Y(n_2206)
);

OAI22xp5_ASAP7_75t_L g2207 ( 
.A1(n_2066),
.A2(n_1415),
.B1(n_1416),
.B2(n_1414),
.Y(n_2207)
);

BUFx3_ASAP7_75t_L g2208 ( 
.A(n_2046),
.Y(n_2208)
);

INVx1_ASAP7_75t_L g2209 ( 
.A(n_2008),
.Y(n_2209)
);

OAI21x1_ASAP7_75t_L g2210 ( 
.A1(n_1968),
.A2(n_781),
.B(n_780),
.Y(n_2210)
);

NAND2xp5_ASAP7_75t_L g2211 ( 
.A(n_2068),
.B(n_1417),
.Y(n_2211)
);

INVx1_ASAP7_75t_L g2212 ( 
.A(n_2046),
.Y(n_2212)
);

INVx2_ASAP7_75t_L g2213 ( 
.A(n_2004),
.Y(n_2213)
);

AND2x2_ASAP7_75t_SL g2214 ( 
.A(n_2015),
.B(n_4),
.Y(n_2214)
);

NAND2xp5_ASAP7_75t_L g2215 ( 
.A(n_2069),
.B(n_1419),
.Y(n_2215)
);

INVx3_ASAP7_75t_SL g2216 ( 
.A(n_2029),
.Y(n_2216)
);

NAND2xp5_ASAP7_75t_L g2217 ( 
.A(n_2070),
.B(n_1423),
.Y(n_2217)
);

CKINVDCx8_ASAP7_75t_R g2218 ( 
.A(n_1935),
.Y(n_2218)
);

AOI221xp5_ASAP7_75t_SL g2219 ( 
.A1(n_2072),
.A2(n_1439),
.B1(n_1443),
.B2(n_1432),
.C(n_1430),
.Y(n_2219)
);

INVx2_ASAP7_75t_L g2220 ( 
.A(n_2005),
.Y(n_2220)
);

AOI21xp5_ASAP7_75t_L g2221 ( 
.A1(n_1971),
.A2(n_783),
.B(n_782),
.Y(n_2221)
);

NOR2xp67_ASAP7_75t_L g2222 ( 
.A(n_1933),
.B(n_785),
.Y(n_2222)
);

NOR2xp33_ASAP7_75t_L g2223 ( 
.A(n_2090),
.B(n_1444),
.Y(n_2223)
);

BUFx4f_ASAP7_75t_SL g2224 ( 
.A(n_2021),
.Y(n_2224)
);

OAI21x1_ASAP7_75t_L g2225 ( 
.A1(n_1972),
.A2(n_1975),
.B(n_1973),
.Y(n_2225)
);

NAND2xp5_ASAP7_75t_SL g2226 ( 
.A(n_1999),
.B(n_2002),
.Y(n_2226)
);

NAND2xp5_ASAP7_75t_L g2227 ( 
.A(n_2075),
.B(n_1447),
.Y(n_2227)
);

INVxp67_ASAP7_75t_SL g2228 ( 
.A(n_2047),
.Y(n_2228)
);

INVx1_ASAP7_75t_L g2229 ( 
.A(n_2042),
.Y(n_2229)
);

BUFx2_ASAP7_75t_L g2230 ( 
.A(n_1943),
.Y(n_2230)
);

A2O1A1Ixp33_ASAP7_75t_L g2231 ( 
.A1(n_2091),
.A2(n_1450),
.B(n_1451),
.C(n_1448),
.Y(n_2231)
);

NAND2xp5_ASAP7_75t_L g2232 ( 
.A(n_2078),
.B(n_1453),
.Y(n_2232)
);

NAND2xp5_ASAP7_75t_L g2233 ( 
.A(n_2079),
.B(n_1454),
.Y(n_2233)
);

OAI21x1_ASAP7_75t_L g2234 ( 
.A1(n_1976),
.A2(n_791),
.B(n_787),
.Y(n_2234)
);

AND2x4_ASAP7_75t_L g2235 ( 
.A(n_2012),
.B(n_792),
.Y(n_2235)
);

O2A1O1Ixp5_ASAP7_75t_L g2236 ( 
.A1(n_1984),
.A2(n_795),
.B(n_796),
.C(n_793),
.Y(n_2236)
);

AO21x1_ASAP7_75t_L g2237 ( 
.A1(n_2026),
.A2(n_4),
.B(n_5),
.Y(n_2237)
);

NAND2xp5_ASAP7_75t_L g2238 ( 
.A(n_2081),
.B(n_1457),
.Y(n_2238)
);

AOI31xp67_ASAP7_75t_L g2239 ( 
.A1(n_1944),
.A2(n_798),
.A3(n_800),
.B(n_797),
.Y(n_2239)
);

AOI21xp5_ASAP7_75t_L g2240 ( 
.A1(n_1977),
.A2(n_1982),
.B(n_1978),
.Y(n_2240)
);

NAND2xp5_ASAP7_75t_SL g2241 ( 
.A(n_1983),
.B(n_1458),
.Y(n_2241)
);

OAI21x1_ASAP7_75t_L g2242 ( 
.A1(n_1936),
.A2(n_802),
.B(n_801),
.Y(n_2242)
);

AOI21xp5_ASAP7_75t_L g2243 ( 
.A1(n_1945),
.A2(n_805),
.B(n_803),
.Y(n_2243)
);

NOR2xp67_ASAP7_75t_L g2244 ( 
.A(n_1928),
.B(n_807),
.Y(n_2244)
);

CKINVDCx5p33_ASAP7_75t_R g2245 ( 
.A(n_2067),
.Y(n_2245)
);

NAND2xp5_ASAP7_75t_L g2246 ( 
.A(n_2082),
.B(n_1459),
.Y(n_2246)
);

OAI22xp5_ASAP7_75t_L g2247 ( 
.A1(n_2084),
.A2(n_1465),
.B1(n_1467),
.B2(n_1464),
.Y(n_2247)
);

AOI21xp5_ASAP7_75t_L g2248 ( 
.A1(n_2010),
.A2(n_809),
.B(n_808),
.Y(n_2248)
);

INVx6_ASAP7_75t_L g2249 ( 
.A(n_2071),
.Y(n_2249)
);

INVx2_ASAP7_75t_SL g2250 ( 
.A(n_2052),
.Y(n_2250)
);

OAI21x1_ASAP7_75t_L g2251 ( 
.A1(n_2087),
.A2(n_814),
.B(n_811),
.Y(n_2251)
);

NAND2xp5_ASAP7_75t_L g2252 ( 
.A(n_2092),
.B(n_1468),
.Y(n_2252)
);

INVx1_ASAP7_75t_L g2253 ( 
.A(n_2053),
.Y(n_2253)
);

NOR2xp33_ASAP7_75t_L g2254 ( 
.A(n_2093),
.B(n_1469),
.Y(n_2254)
);

AOI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2017),
.A2(n_816),
.B(n_815),
.Y(n_2255)
);

INVxp67_ASAP7_75t_L g2256 ( 
.A(n_2048),
.Y(n_2256)
);

NOR2x1_ASAP7_75t_R g2257 ( 
.A(n_2031),
.B(n_1470),
.Y(n_2257)
);

OAI21xp5_ASAP7_75t_L g2258 ( 
.A1(n_2096),
.A2(n_1481),
.B(n_1477),
.Y(n_2258)
);

NOR2xp67_ASAP7_75t_L g2259 ( 
.A(n_2098),
.B(n_817),
.Y(n_2259)
);

OR2x2_ASAP7_75t_L g2260 ( 
.A(n_1947),
.B(n_1484),
.Y(n_2260)
);

CKINVDCx20_ASAP7_75t_R g2261 ( 
.A(n_2073),
.Y(n_2261)
);

NAND2xp33_ASAP7_75t_L g2262 ( 
.A(n_2100),
.B(n_1554),
.Y(n_2262)
);

NAND2xp5_ASAP7_75t_L g2263 ( 
.A(n_2101),
.B(n_1486),
.Y(n_2263)
);

OA21x2_ASAP7_75t_L g2264 ( 
.A1(n_2103),
.A2(n_1491),
.B(n_1489),
.Y(n_2264)
);

NAND2xp5_ASAP7_75t_L g2265 ( 
.A(n_2105),
.B(n_1493),
.Y(n_2265)
);

OAI21x1_ASAP7_75t_L g2266 ( 
.A1(n_2018),
.A2(n_820),
.B(n_818),
.Y(n_2266)
);

INVx3_ASAP7_75t_L g2267 ( 
.A(n_2076),
.Y(n_2267)
);

CKINVDCx16_ASAP7_75t_R g2268 ( 
.A(n_1974),
.Y(n_2268)
);

BUFx6f_ASAP7_75t_L g2269 ( 
.A(n_2034),
.Y(n_2269)
);

OAI21x1_ASAP7_75t_L g2270 ( 
.A1(n_2020),
.A2(n_822),
.B(n_821),
.Y(n_2270)
);

OAI21x1_ASAP7_75t_SL g2271 ( 
.A1(n_2033),
.A2(n_824),
.B(n_823),
.Y(n_2271)
);

A2O1A1Ixp33_ASAP7_75t_L g2272 ( 
.A1(n_2106),
.A2(n_1496),
.B(n_1499),
.C(n_1495),
.Y(n_2272)
);

OAI21x1_ASAP7_75t_L g2273 ( 
.A1(n_2107),
.A2(n_826),
.B(n_825),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_2055),
.Y(n_2274)
);

OAI21xp5_ASAP7_75t_L g2275 ( 
.A1(n_2138),
.A2(n_2109),
.B(n_2108),
.Y(n_2275)
);

AND2x4_ASAP7_75t_L g2276 ( 
.A(n_2208),
.B(n_2049),
.Y(n_2276)
);

NAND2xp5_ASAP7_75t_L g2277 ( 
.A(n_2140),
.B(n_2110),
.Y(n_2277)
);

INVxp67_ASAP7_75t_SL g2278 ( 
.A(n_2137),
.Y(n_2278)
);

INVx2_ASAP7_75t_L g2279 ( 
.A(n_2212),
.Y(n_2279)
);

INVxp67_ASAP7_75t_L g2280 ( 
.A(n_2135),
.Y(n_2280)
);

INVx1_ASAP7_75t_L g2281 ( 
.A(n_2163),
.Y(n_2281)
);

INVx1_ASAP7_75t_L g2282 ( 
.A(n_2182),
.Y(n_2282)
);

INVx2_ASAP7_75t_L g2283 ( 
.A(n_2126),
.Y(n_2283)
);

INVx2_ASAP7_75t_L g2284 ( 
.A(n_2205),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2200),
.Y(n_2285)
);

OAI21xp5_ASAP7_75t_L g2286 ( 
.A1(n_2136),
.A2(n_2113),
.B(n_2111),
.Y(n_2286)
);

INVx1_ASAP7_75t_L g2287 ( 
.A(n_2123),
.Y(n_2287)
);

AO21x2_ASAP7_75t_L g2288 ( 
.A1(n_2128),
.A2(n_2117),
.B(n_2116),
.Y(n_2288)
);

AO21x2_ASAP7_75t_L g2289 ( 
.A1(n_2129),
.A2(n_2119),
.B(n_2118),
.Y(n_2289)
);

INVxp67_ASAP7_75t_L g2290 ( 
.A(n_2151),
.Y(n_2290)
);

INVx4_ASAP7_75t_L g2291 ( 
.A(n_2132),
.Y(n_2291)
);

AND2x4_ASAP7_75t_L g2292 ( 
.A(n_2154),
.B(n_2121),
.Y(n_2292)
);

OAI22xp5_ASAP7_75t_L g2293 ( 
.A1(n_2229),
.A2(n_2051),
.B1(n_2028),
.B2(n_2024),
.Y(n_2293)
);

OAI21x1_ASAP7_75t_SL g2294 ( 
.A1(n_2271),
.A2(n_2030),
.B(n_1962),
.Y(n_2294)
);

AND2x2_ASAP7_75t_L g2295 ( 
.A(n_2124),
.B(n_2032),
.Y(n_2295)
);

OAI21xp5_ASAP7_75t_L g2296 ( 
.A1(n_2145),
.A2(n_1955),
.B(n_2037),
.Y(n_2296)
);

AND2x2_ASAP7_75t_L g2297 ( 
.A(n_2133),
.B(n_1501),
.Y(n_2297)
);

NAND2xp5_ASAP7_75t_L g2298 ( 
.A(n_2130),
.B(n_1959),
.Y(n_2298)
);

NOR2xp33_ASAP7_75t_SL g2299 ( 
.A(n_2218),
.B(n_1503),
.Y(n_2299)
);

OAI21x1_ASAP7_75t_L g2300 ( 
.A1(n_2139),
.A2(n_829),
.B(n_827),
.Y(n_2300)
);

INVx3_ASAP7_75t_L g2301 ( 
.A(n_2132),
.Y(n_2301)
);

BUFx10_ASAP7_75t_L g2302 ( 
.A(n_2166),
.Y(n_2302)
);

INVx1_ASAP7_75t_L g2303 ( 
.A(n_2131),
.Y(n_2303)
);

INVx1_ASAP7_75t_L g2304 ( 
.A(n_2148),
.Y(n_2304)
);

AO21x2_ASAP7_75t_L g2305 ( 
.A1(n_2181),
.A2(n_2045),
.B(n_2039),
.Y(n_2305)
);

OAI22xp5_ASAP7_75t_L g2306 ( 
.A1(n_2228),
.A2(n_1514),
.B1(n_1515),
.B2(n_1513),
.Y(n_2306)
);

AND2x4_ASAP7_75t_L g2307 ( 
.A(n_2125),
.B(n_2086),
.Y(n_2307)
);

INVx2_ASAP7_75t_L g2308 ( 
.A(n_2274),
.Y(n_2308)
);

INVx2_ASAP7_75t_SL g2309 ( 
.A(n_2269),
.Y(n_2309)
);

AO32x2_ASAP7_75t_L g2310 ( 
.A1(n_2162),
.A2(n_2097),
.A3(n_2099),
.B1(n_2094),
.B2(n_2089),
.Y(n_2310)
);

INVx2_ASAP7_75t_L g2311 ( 
.A(n_2253),
.Y(n_2311)
);

AOI21xp5_ASAP7_75t_SL g2312 ( 
.A1(n_2226),
.A2(n_832),
.B(n_831),
.Y(n_2312)
);

AO31x2_ASAP7_75t_L g2313 ( 
.A1(n_2127),
.A2(n_834),
.A3(n_835),
.B(n_833),
.Y(n_2313)
);

OAI21x1_ASAP7_75t_L g2314 ( 
.A1(n_2149),
.A2(n_840),
.B(n_836),
.Y(n_2314)
);

INVx1_ASAP7_75t_L g2315 ( 
.A(n_2209),
.Y(n_2315)
);

AO31x2_ASAP7_75t_L g2316 ( 
.A1(n_2237),
.A2(n_843),
.A3(n_845),
.B(n_841),
.Y(n_2316)
);

AOI21xp5_ASAP7_75t_L g2317 ( 
.A1(n_2240),
.A2(n_2115),
.B(n_2104),
.Y(n_2317)
);

AND2x2_ASAP7_75t_L g2318 ( 
.A(n_2214),
.B(n_1516),
.Y(n_2318)
);

NAND2xp5_ASAP7_75t_L g2319 ( 
.A(n_2155),
.B(n_2120),
.Y(n_2319)
);

A2O1A1Ixp33_ASAP7_75t_L g2320 ( 
.A1(n_2223),
.A2(n_2122),
.B(n_1524),
.C(n_1526),
.Y(n_2320)
);

NAND2x1p5_ASAP7_75t_L g2321 ( 
.A(n_2199),
.B(n_846),
.Y(n_2321)
);

AOI22xp33_ASAP7_75t_L g2322 ( 
.A1(n_2141),
.A2(n_1528),
.B1(n_1529),
.B2(n_1522),
.Y(n_2322)
);

OA21x2_ASAP7_75t_L g2323 ( 
.A1(n_2175),
.A2(n_1541),
.B(n_1534),
.Y(n_2323)
);

A2O1A1Ixp33_ASAP7_75t_L g2324 ( 
.A1(n_2254),
.A2(n_1545),
.B(n_1551),
.C(n_1547),
.Y(n_2324)
);

AO32x2_ASAP7_75t_L g2325 ( 
.A1(n_2161),
.A2(n_8),
.A3(n_6),
.B1(n_7),
.B2(n_9),
.Y(n_2325)
);

AOI222xp33_ASAP7_75t_L g2326 ( 
.A1(n_2134),
.A2(n_1557),
.B1(n_1553),
.B2(n_1558),
.C1(n_1556),
.C2(n_1543),
.Y(n_2326)
);

AND2x4_ASAP7_75t_L g2327 ( 
.A(n_2199),
.B(n_847),
.Y(n_2327)
);

AOI22xp33_ASAP7_75t_L g2328 ( 
.A1(n_2196),
.A2(n_1563),
.B1(n_1559),
.B2(n_8),
.Y(n_2328)
);

NOR2xp33_ASAP7_75t_L g2329 ( 
.A(n_2170),
.B(n_6),
.Y(n_2329)
);

AOI21x1_ASAP7_75t_L g2330 ( 
.A1(n_2142),
.A2(n_851),
.B(n_848),
.Y(n_2330)
);

INVx4_ASAP7_75t_L g2331 ( 
.A(n_2269),
.Y(n_2331)
);

INVx2_ASAP7_75t_SL g2332 ( 
.A(n_2249),
.Y(n_2332)
);

INVx1_ASAP7_75t_SL g2333 ( 
.A(n_2216),
.Y(n_2333)
);

OAI21xp5_ASAP7_75t_L g2334 ( 
.A1(n_2143),
.A2(n_854),
.B(n_852),
.Y(n_2334)
);

INVx1_ASAP7_75t_L g2335 ( 
.A(n_2256),
.Y(n_2335)
);

OAI21x1_ASAP7_75t_L g2336 ( 
.A1(n_2172),
.A2(n_858),
.B(n_857),
.Y(n_2336)
);

INVx2_ASAP7_75t_L g2337 ( 
.A(n_2213),
.Y(n_2337)
);

INVxp67_ASAP7_75t_L g2338 ( 
.A(n_2184),
.Y(n_2338)
);

O2A1O1Ixp33_ASAP7_75t_SL g2339 ( 
.A1(n_2150),
.A2(n_862),
.B(n_864),
.C(n_860),
.Y(n_2339)
);

AO21x2_ASAP7_75t_L g2340 ( 
.A1(n_2144),
.A2(n_866),
.B(n_865),
.Y(n_2340)
);

NOR2xp33_ASAP7_75t_L g2341 ( 
.A(n_2230),
.B(n_7),
.Y(n_2341)
);

OAI21x1_ASAP7_75t_L g2342 ( 
.A1(n_2187),
.A2(n_2234),
.B(n_2210),
.Y(n_2342)
);

OAI21xp5_ASAP7_75t_L g2343 ( 
.A1(n_2225),
.A2(n_868),
.B(n_867),
.Y(n_2343)
);

BUFx2_ASAP7_75t_L g2344 ( 
.A(n_2186),
.Y(n_2344)
);

INVx1_ASAP7_75t_L g2345 ( 
.A(n_2220),
.Y(n_2345)
);

AND2x2_ASAP7_75t_L g2346 ( 
.A(n_2268),
.B(n_9),
.Y(n_2346)
);

AO21x2_ASAP7_75t_L g2347 ( 
.A1(n_2248),
.A2(n_870),
.B(n_869),
.Y(n_2347)
);

OAI21xp5_ASAP7_75t_L g2348 ( 
.A1(n_2236),
.A2(n_872),
.B(n_871),
.Y(n_2348)
);

INVx1_ASAP7_75t_L g2349 ( 
.A(n_2250),
.Y(n_2349)
);

OAI21xp5_ASAP7_75t_L g2350 ( 
.A1(n_2197),
.A2(n_877),
.B(n_873),
.Y(n_2350)
);

NOR2x1_ASAP7_75t_SL g2351 ( 
.A(n_2159),
.B(n_878),
.Y(n_2351)
);

INVx1_ASAP7_75t_L g2352 ( 
.A(n_2273),
.Y(n_2352)
);

OAI21x1_ASAP7_75t_L g2353 ( 
.A1(n_2189),
.A2(n_2242),
.B(n_2191),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_2194),
.Y(n_2354)
);

A2O1A1Ixp33_ASAP7_75t_L g2355 ( 
.A1(n_2259),
.A2(n_12),
.B(n_10),
.C(n_11),
.Y(n_2355)
);

OAI21x1_ASAP7_75t_L g2356 ( 
.A1(n_2158),
.A2(n_881),
.B(n_879),
.Y(n_2356)
);

OR2x2_ASAP7_75t_L g2357 ( 
.A(n_2179),
.B(n_10),
.Y(n_2357)
);

OAI21x1_ASAP7_75t_L g2358 ( 
.A1(n_2164),
.A2(n_883),
.B(n_882),
.Y(n_2358)
);

OR2x2_ASAP7_75t_L g2359 ( 
.A(n_2183),
.B(n_11),
.Y(n_2359)
);

A2O1A1Ixp33_ASAP7_75t_L g2360 ( 
.A1(n_2260),
.A2(n_15),
.B(n_13),
.C(n_14),
.Y(n_2360)
);

NAND3xp33_ASAP7_75t_L g2361 ( 
.A(n_2153),
.B(n_13),
.C(n_16),
.Y(n_2361)
);

OAI21x1_ASAP7_75t_L g2362 ( 
.A1(n_2168),
.A2(n_885),
.B(n_884),
.Y(n_2362)
);

NAND3xp33_ASAP7_75t_L g2363 ( 
.A(n_2177),
.B(n_16),
.C(n_17),
.Y(n_2363)
);

OAI21x1_ASAP7_75t_L g2364 ( 
.A1(n_2266),
.A2(n_888),
.B(n_887),
.Y(n_2364)
);

AOI21xp5_ASAP7_75t_L g2365 ( 
.A1(n_2243),
.A2(n_891),
.B(n_889),
.Y(n_2365)
);

OAI21xp5_ASAP7_75t_L g2366 ( 
.A1(n_2252),
.A2(n_2265),
.B(n_2263),
.Y(n_2366)
);

AO21x2_ASAP7_75t_L g2367 ( 
.A1(n_2147),
.A2(n_896),
.B(n_895),
.Y(n_2367)
);

AOI22xp5_ASAP7_75t_L g2368 ( 
.A1(n_2261),
.A2(n_19),
.B1(n_17),
.B2(n_18),
.Y(n_2368)
);

OAI21x1_ASAP7_75t_L g2369 ( 
.A1(n_2270),
.A2(n_898),
.B(n_897),
.Y(n_2369)
);

OAI21x1_ASAP7_75t_L g2370 ( 
.A1(n_2251),
.A2(n_900),
.B(n_899),
.Y(n_2370)
);

AOI21xp5_ASAP7_75t_L g2371 ( 
.A1(n_2152),
.A2(n_903),
.B(n_901),
.Y(n_2371)
);

AND2x4_ASAP7_75t_L g2372 ( 
.A(n_2267),
.B(n_904),
.Y(n_2372)
);

CKINVDCx20_ASAP7_75t_R g2373 ( 
.A(n_2245),
.Y(n_2373)
);

OAI22xp5_ASAP7_75t_L g2374 ( 
.A1(n_2198),
.A2(n_20),
.B1(n_18),
.B2(n_19),
.Y(n_2374)
);

NOR2xp33_ASAP7_75t_L g2375 ( 
.A(n_2204),
.B(n_20),
.Y(n_2375)
);

BUFx10_ASAP7_75t_L g2376 ( 
.A(n_2206),
.Y(n_2376)
);

OR2x2_ASAP7_75t_L g2377 ( 
.A(n_2195),
.B(n_2185),
.Y(n_2377)
);

OA21x2_ASAP7_75t_L g2378 ( 
.A1(n_2219),
.A2(n_907),
.B(n_906),
.Y(n_2378)
);

OAI22xp33_ASAP7_75t_L g2379 ( 
.A1(n_2186),
.A2(n_23),
.B1(n_21),
.B2(n_22),
.Y(n_2379)
);

OAI21xp5_ASAP7_75t_L g2380 ( 
.A1(n_2272),
.A2(n_911),
.B(n_909),
.Y(n_2380)
);

OAI21x1_ASAP7_75t_L g2381 ( 
.A1(n_2165),
.A2(n_913),
.B(n_912),
.Y(n_2381)
);

OAI21x1_ASAP7_75t_L g2382 ( 
.A1(n_2171),
.A2(n_2176),
.B(n_2174),
.Y(n_2382)
);

AND2x2_ASAP7_75t_L g2383 ( 
.A(n_2146),
.B(n_23),
.Y(n_2383)
);

OAI21xp5_ASAP7_75t_L g2384 ( 
.A1(n_2231),
.A2(n_915),
.B(n_914),
.Y(n_2384)
);

INVx1_ASAP7_75t_L g2385 ( 
.A(n_2180),
.Y(n_2385)
);

OR2x2_ASAP7_75t_L g2386 ( 
.A(n_2192),
.B(n_24),
.Y(n_2386)
);

NOR2x1_ASAP7_75t_R g2387 ( 
.A(n_2249),
.B(n_916),
.Y(n_2387)
);

AOI22xp33_ASAP7_75t_L g2388 ( 
.A1(n_2178),
.A2(n_26),
.B1(n_24),
.B2(n_25),
.Y(n_2388)
);

OAI22xp33_ASAP7_75t_L g2389 ( 
.A1(n_2224),
.A2(n_29),
.B1(n_27),
.B2(n_28),
.Y(n_2389)
);

OAI21x1_ASAP7_75t_L g2390 ( 
.A1(n_2188),
.A2(n_918),
.B(n_917),
.Y(n_2390)
);

AO31x2_ASAP7_75t_L g2391 ( 
.A1(n_2190),
.A2(n_922),
.A3(n_923),
.B(n_919),
.Y(n_2391)
);

OAI21x1_ASAP7_75t_L g2392 ( 
.A1(n_2201),
.A2(n_2221),
.B(n_2255),
.Y(n_2392)
);

INVx2_ASAP7_75t_L g2393 ( 
.A(n_2169),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_2156),
.Y(n_2394)
);

INVx2_ASAP7_75t_L g2395 ( 
.A(n_2239),
.Y(n_2395)
);

OAI21x1_ASAP7_75t_L g2396 ( 
.A1(n_2173),
.A2(n_928),
.B(n_927),
.Y(n_2396)
);

AO21x2_ASAP7_75t_L g2397 ( 
.A1(n_2244),
.A2(n_934),
.B(n_932),
.Y(n_2397)
);

INVx2_ASAP7_75t_L g2398 ( 
.A(n_2157),
.Y(n_2398)
);

OAI21x1_ASAP7_75t_L g2399 ( 
.A1(n_2264),
.A2(n_937),
.B(n_936),
.Y(n_2399)
);

NAND2xp5_ASAP7_75t_L g2400 ( 
.A(n_2235),
.B(n_27),
.Y(n_2400)
);

OAI21x1_ASAP7_75t_L g2401 ( 
.A1(n_2160),
.A2(n_939),
.B(n_938),
.Y(n_2401)
);

AOI21xp5_ASAP7_75t_L g2402 ( 
.A1(n_2222),
.A2(n_941),
.B(n_940),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_2157),
.Y(n_2403)
);

AOI22xp5_ASAP7_75t_L g2404 ( 
.A1(n_2262),
.A2(n_2167),
.B1(n_2241),
.B2(n_2202),
.Y(n_2404)
);

AO21x2_ASAP7_75t_L g2405 ( 
.A1(n_2258),
.A2(n_944),
.B(n_942),
.Y(n_2405)
);

OAI21xp5_ASAP7_75t_L g2406 ( 
.A1(n_2193),
.A2(n_948),
.B(n_946),
.Y(n_2406)
);

NAND2xp5_ASAP7_75t_L g2407 ( 
.A(n_2203),
.B(n_28),
.Y(n_2407)
);

AND2x4_ASAP7_75t_L g2408 ( 
.A(n_2211),
.B(n_949),
.Y(n_2408)
);

INVx1_ASAP7_75t_L g2409 ( 
.A(n_2215),
.Y(n_2409)
);

INVx2_ASAP7_75t_L g2410 ( 
.A(n_2217),
.Y(n_2410)
);

AO31x2_ASAP7_75t_L g2411 ( 
.A1(n_2227),
.A2(n_952),
.A3(n_953),
.B(n_951),
.Y(n_2411)
);

OAI22xp5_ASAP7_75t_L g2412 ( 
.A1(n_2232),
.A2(n_31),
.B1(n_29),
.B2(n_30),
.Y(n_2412)
);

CKINVDCx20_ASAP7_75t_R g2413 ( 
.A(n_2233),
.Y(n_2413)
);

OAI21x1_ASAP7_75t_L g2414 ( 
.A1(n_2238),
.A2(n_956),
.B(n_955),
.Y(n_2414)
);

NOR2xp67_ASAP7_75t_L g2415 ( 
.A(n_2246),
.B(n_959),
.Y(n_2415)
);

OAI21x1_ASAP7_75t_L g2416 ( 
.A1(n_2207),
.A2(n_961),
.B(n_960),
.Y(n_2416)
);

BUFx3_ASAP7_75t_L g2417 ( 
.A(n_2247),
.Y(n_2417)
);

CKINVDCx5p33_ASAP7_75t_R g2418 ( 
.A(n_2257),
.Y(n_2418)
);

OA21x2_ASAP7_75t_L g2419 ( 
.A1(n_2129),
.A2(n_963),
.B(n_962),
.Y(n_2419)
);

OAI21x1_ASAP7_75t_L g2420 ( 
.A1(n_2126),
.A2(n_968),
.B(n_964),
.Y(n_2420)
);

OAI21x1_ASAP7_75t_SL g2421 ( 
.A1(n_2271),
.A2(n_970),
.B(n_969),
.Y(n_2421)
);

INVx1_ASAP7_75t_L g2422 ( 
.A(n_2212),
.Y(n_2422)
);

NAND2xp5_ASAP7_75t_L g2423 ( 
.A(n_2140),
.B(n_30),
.Y(n_2423)
);

INVx2_ASAP7_75t_SL g2424 ( 
.A(n_2132),
.Y(n_2424)
);

OAI21x1_ASAP7_75t_L g2425 ( 
.A1(n_2126),
.A2(n_972),
.B(n_971),
.Y(n_2425)
);

INVxp67_ASAP7_75t_SL g2426 ( 
.A(n_2137),
.Y(n_2426)
);

OAI21xp5_ASAP7_75t_L g2427 ( 
.A1(n_2138),
.A2(n_975),
.B(n_974),
.Y(n_2427)
);

INVx2_ASAP7_75t_L g2428 ( 
.A(n_2212),
.Y(n_2428)
);

AOI22xp33_ASAP7_75t_SL g2429 ( 
.A1(n_2124),
.A2(n_33),
.B1(n_31),
.B2(n_32),
.Y(n_2429)
);

OAI21x1_ASAP7_75t_L g2430 ( 
.A1(n_2126),
.A2(n_977),
.B(n_976),
.Y(n_2430)
);

OA21x2_ASAP7_75t_L g2431 ( 
.A1(n_2350),
.A2(n_2343),
.B(n_2427),
.Y(n_2431)
);

INVx1_ASAP7_75t_L g2432 ( 
.A(n_2315),
.Y(n_2432)
);

BUFx2_ASAP7_75t_L g2433 ( 
.A(n_2338),
.Y(n_2433)
);

BUFx2_ASAP7_75t_L g2434 ( 
.A(n_2278),
.Y(n_2434)
);

BUFx2_ASAP7_75t_L g2435 ( 
.A(n_2426),
.Y(n_2435)
);

INVx2_ASAP7_75t_L g2436 ( 
.A(n_2337),
.Y(n_2436)
);

AO21x2_ASAP7_75t_L g2437 ( 
.A1(n_2403),
.A2(n_979),
.B(n_978),
.Y(n_2437)
);

INVx2_ASAP7_75t_L g2438 ( 
.A(n_2308),
.Y(n_2438)
);

OAI21x1_ASAP7_75t_L g2439 ( 
.A1(n_2342),
.A2(n_984),
.B(n_981),
.Y(n_2439)
);

NOR2xp33_ASAP7_75t_L g2440 ( 
.A(n_2298),
.B(n_985),
.Y(n_2440)
);

OR2x2_ASAP7_75t_L g2441 ( 
.A(n_2423),
.B(n_32),
.Y(n_2441)
);

OR2x2_ASAP7_75t_L g2442 ( 
.A(n_2377),
.B(n_33),
.Y(n_2442)
);

INVx1_ASAP7_75t_L g2443 ( 
.A(n_2284),
.Y(n_2443)
);

INVx4_ASAP7_75t_L g2444 ( 
.A(n_2291),
.Y(n_2444)
);

INVx1_ASAP7_75t_L g2445 ( 
.A(n_2285),
.Y(n_2445)
);

INVx1_ASAP7_75t_L g2446 ( 
.A(n_2287),
.Y(n_2446)
);

INVx1_ASAP7_75t_L g2447 ( 
.A(n_2303),
.Y(n_2447)
);

AND2x4_ASAP7_75t_L g2448 ( 
.A(n_2332),
.B(n_2331),
.Y(n_2448)
);

NOR2xp33_ASAP7_75t_L g2449 ( 
.A(n_2319),
.B(n_2277),
.Y(n_2449)
);

AO21x2_ASAP7_75t_L g2450 ( 
.A1(n_2398),
.A2(n_987),
.B(n_986),
.Y(n_2450)
);

AND2x2_ASAP7_75t_L g2451 ( 
.A(n_2318),
.B(n_34),
.Y(n_2451)
);

AOI21x1_ASAP7_75t_L g2452 ( 
.A1(n_2394),
.A2(n_992),
.B(n_990),
.Y(n_2452)
);

INVx2_ASAP7_75t_L g2453 ( 
.A(n_2311),
.Y(n_2453)
);

AND2x2_ASAP7_75t_L g2454 ( 
.A(n_2295),
.B(n_35),
.Y(n_2454)
);

OR2x2_ASAP7_75t_L g2455 ( 
.A(n_2279),
.B(n_35),
.Y(n_2455)
);

INVx3_ASAP7_75t_L g2456 ( 
.A(n_2376),
.Y(n_2456)
);

INVx2_ASAP7_75t_L g2457 ( 
.A(n_2345),
.Y(n_2457)
);

INVx1_ASAP7_75t_L g2458 ( 
.A(n_2304),
.Y(n_2458)
);

HB1xp67_ASAP7_75t_L g2459 ( 
.A(n_2290),
.Y(n_2459)
);

INVx2_ASAP7_75t_L g2460 ( 
.A(n_2428),
.Y(n_2460)
);

BUFx6f_ASAP7_75t_L g2461 ( 
.A(n_2309),
.Y(n_2461)
);

NOR2xp33_ASAP7_75t_L g2462 ( 
.A(n_2333),
.B(n_995),
.Y(n_2462)
);

INVx2_ASAP7_75t_L g2463 ( 
.A(n_2281),
.Y(n_2463)
);

HB1xp67_ASAP7_75t_L g2464 ( 
.A(n_2335),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_2282),
.Y(n_2465)
);

INVx1_ASAP7_75t_L g2466 ( 
.A(n_2422),
.Y(n_2466)
);

INVx2_ASAP7_75t_L g2467 ( 
.A(n_2349),
.Y(n_2467)
);

NAND2xp5_ASAP7_75t_L g2468 ( 
.A(n_2410),
.B(n_36),
.Y(n_2468)
);

OR2x2_ASAP7_75t_L g2469 ( 
.A(n_2357),
.B(n_36),
.Y(n_2469)
);

INVx1_ASAP7_75t_L g2470 ( 
.A(n_2354),
.Y(n_2470)
);

INVx1_ASAP7_75t_L g2471 ( 
.A(n_2407),
.Y(n_2471)
);

HB1xp67_ASAP7_75t_L g2472 ( 
.A(n_2280),
.Y(n_2472)
);

INVx1_ASAP7_75t_L g2473 ( 
.A(n_2409),
.Y(n_2473)
);

INVx1_ASAP7_75t_L g2474 ( 
.A(n_2325),
.Y(n_2474)
);

OAI21x1_ASAP7_75t_L g2475 ( 
.A1(n_2353),
.A2(n_997),
.B(n_996),
.Y(n_2475)
);

INVx2_ASAP7_75t_L g2476 ( 
.A(n_2385),
.Y(n_2476)
);

OAI22xp5_ASAP7_75t_L g2477 ( 
.A1(n_2417),
.A2(n_39),
.B1(n_37),
.B2(n_38),
.Y(n_2477)
);

AND2x2_ASAP7_75t_L g2478 ( 
.A(n_2297),
.B(n_40),
.Y(n_2478)
);

AOI22xp33_ASAP7_75t_L g2479 ( 
.A1(n_2375),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_2479)
);

AO21x2_ASAP7_75t_L g2480 ( 
.A1(n_2296),
.A2(n_1001),
.B(n_999),
.Y(n_2480)
);

INVx2_ASAP7_75t_SL g2481 ( 
.A(n_2302),
.Y(n_2481)
);

INVx2_ASAP7_75t_L g2482 ( 
.A(n_2288),
.Y(n_2482)
);

INVx1_ASAP7_75t_L g2483 ( 
.A(n_2325),
.Y(n_2483)
);

INVx1_ASAP7_75t_L g2484 ( 
.A(n_2386),
.Y(n_2484)
);

INVx1_ASAP7_75t_L g2485 ( 
.A(n_2361),
.Y(n_2485)
);

AND2x2_ASAP7_75t_L g2486 ( 
.A(n_2346),
.B(n_41),
.Y(n_2486)
);

INVx1_ASAP7_75t_L g2487 ( 
.A(n_2359),
.Y(n_2487)
);

OR2x2_ASAP7_75t_L g2488 ( 
.A(n_2344),
.B(n_44),
.Y(n_2488)
);

OR2x2_ASAP7_75t_L g2489 ( 
.A(n_2400),
.B(n_44),
.Y(n_2489)
);

INVx2_ASAP7_75t_L g2490 ( 
.A(n_2307),
.Y(n_2490)
);

BUFx6f_ASAP7_75t_L g2491 ( 
.A(n_2424),
.Y(n_2491)
);

INVx1_ASAP7_75t_L g2492 ( 
.A(n_2363),
.Y(n_2492)
);

INVx2_ASAP7_75t_L g2493 ( 
.A(n_2399),
.Y(n_2493)
);

INVx3_ASAP7_75t_L g2494 ( 
.A(n_2301),
.Y(n_2494)
);

INVx1_ASAP7_75t_L g2495 ( 
.A(n_2292),
.Y(n_2495)
);

AO31x2_ASAP7_75t_L g2496 ( 
.A1(n_2395),
.A2(n_1003),
.A3(n_1004),
.B(n_1002),
.Y(n_2496)
);

INVx2_ASAP7_75t_L g2497 ( 
.A(n_2396),
.Y(n_2497)
);

INVx2_ASAP7_75t_L g2498 ( 
.A(n_2330),
.Y(n_2498)
);

HB1xp67_ASAP7_75t_L g2499 ( 
.A(n_2276),
.Y(n_2499)
);

INVx1_ASAP7_75t_L g2500 ( 
.A(n_2411),
.Y(n_2500)
);

NAND2xp5_ASAP7_75t_SL g2501 ( 
.A(n_2366),
.B(n_45),
.Y(n_2501)
);

BUFx2_ASAP7_75t_SL g2502 ( 
.A(n_2373),
.Y(n_2502)
);

AND2x2_ASAP7_75t_L g2503 ( 
.A(n_2383),
.B(n_45),
.Y(n_2503)
);

CKINVDCx6p67_ASAP7_75t_R g2504 ( 
.A(n_2413),
.Y(n_2504)
);

INVx1_ASAP7_75t_L g2505 ( 
.A(n_2411),
.Y(n_2505)
);

INVx4_ASAP7_75t_L g2506 ( 
.A(n_2327),
.Y(n_2506)
);

INVx2_ASAP7_75t_L g2507 ( 
.A(n_2352),
.Y(n_2507)
);

INVx1_ASAP7_75t_L g2508 ( 
.A(n_2372),
.Y(n_2508)
);

BUFx6f_ASAP7_75t_L g2509 ( 
.A(n_2418),
.Y(n_2509)
);

INVx1_ASAP7_75t_L g2510 ( 
.A(n_2391),
.Y(n_2510)
);

AOI22xp33_ASAP7_75t_L g2511 ( 
.A1(n_2380),
.A2(n_48),
.B1(n_46),
.B2(n_47),
.Y(n_2511)
);

OAI21xp5_ASAP7_75t_L g2512 ( 
.A1(n_2275),
.A2(n_46),
.B(n_50),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_2391),
.Y(n_2513)
);

INVx1_ASAP7_75t_L g2514 ( 
.A(n_2412),
.Y(n_2514)
);

AOI22xp33_ASAP7_75t_SL g2515 ( 
.A1(n_2384),
.A2(n_58),
.B1(n_66),
.B2(n_50),
.Y(n_2515)
);

INVx2_ASAP7_75t_L g2516 ( 
.A(n_2289),
.Y(n_2516)
);

O2A1O1Ixp33_ASAP7_75t_L g2517 ( 
.A1(n_2360),
.A2(n_53),
.B(n_51),
.C(n_52),
.Y(n_2517)
);

BUFx2_ASAP7_75t_L g2518 ( 
.A(n_2310),
.Y(n_2518)
);

AND2x2_ASAP7_75t_L g2519 ( 
.A(n_2429),
.B(n_51),
.Y(n_2519)
);

INVx2_ASAP7_75t_L g2520 ( 
.A(n_2381),
.Y(n_2520)
);

BUFx2_ASAP7_75t_L g2521 ( 
.A(n_2310),
.Y(n_2521)
);

AND2x2_ASAP7_75t_L g2522 ( 
.A(n_2329),
.B(n_54),
.Y(n_2522)
);

INVx1_ASAP7_75t_L g2523 ( 
.A(n_2414),
.Y(n_2523)
);

OAI21x1_ASAP7_75t_L g2524 ( 
.A1(n_2420),
.A2(n_1009),
.B(n_1006),
.Y(n_2524)
);

AO31x2_ASAP7_75t_L g2525 ( 
.A1(n_2393),
.A2(n_2351),
.A3(n_2283),
.B(n_2317),
.Y(n_2525)
);

AND2x2_ASAP7_75t_L g2526 ( 
.A(n_2341),
.B(n_54),
.Y(n_2526)
);

AND2x2_ASAP7_75t_L g2527 ( 
.A(n_2328),
.B(n_55),
.Y(n_2527)
);

BUFx2_ASAP7_75t_L g2528 ( 
.A(n_2408),
.Y(n_2528)
);

INVx2_ASAP7_75t_L g2529 ( 
.A(n_2390),
.Y(n_2529)
);

BUFx6f_ASAP7_75t_L g2530 ( 
.A(n_2321),
.Y(n_2530)
);

INVx1_ASAP7_75t_L g2531 ( 
.A(n_2355),
.Y(n_2531)
);

AOI22xp33_ASAP7_75t_L g2532 ( 
.A1(n_2388),
.A2(n_57),
.B1(n_55),
.B2(n_56),
.Y(n_2532)
);

INVx1_ASAP7_75t_L g2533 ( 
.A(n_2316),
.Y(n_2533)
);

NAND2xp5_ASAP7_75t_L g2534 ( 
.A(n_2449),
.B(n_2404),
.Y(n_2534)
);

BUFx3_ASAP7_75t_L g2535 ( 
.A(n_2461),
.Y(n_2535)
);

NAND2xp33_ASAP7_75t_R g2536 ( 
.A(n_2456),
.B(n_2378),
.Y(n_2536)
);

BUFx3_ASAP7_75t_L g2537 ( 
.A(n_2461),
.Y(n_2537)
);

AND2x2_ASAP7_75t_L g2538 ( 
.A(n_2454),
.B(n_2368),
.Y(n_2538)
);

INVx2_ASAP7_75t_SL g2539 ( 
.A(n_2448),
.Y(n_2539)
);

NAND2xp33_ASAP7_75t_R g2540 ( 
.A(n_2528),
.B(n_2323),
.Y(n_2540)
);

AND2x4_ASAP7_75t_L g2541 ( 
.A(n_2506),
.B(n_2415),
.Y(n_2541)
);

INVx1_ASAP7_75t_L g2542 ( 
.A(n_2470),
.Y(n_2542)
);

NOR2xp33_ASAP7_75t_R g2543 ( 
.A(n_2504),
.B(n_2299),
.Y(n_2543)
);

BUFx10_ASAP7_75t_L g2544 ( 
.A(n_2509),
.Y(n_2544)
);

CKINVDCx11_ASAP7_75t_R g2545 ( 
.A(n_2509),
.Y(n_2545)
);

NOR2x1_ASAP7_75t_L g2546 ( 
.A(n_2471),
.B(n_2473),
.Y(n_2546)
);

INVx1_ASAP7_75t_L g2547 ( 
.A(n_2432),
.Y(n_2547)
);

XNOR2xp5_ASAP7_75t_L g2548 ( 
.A(n_2502),
.B(n_2306),
.Y(n_2548)
);

AND2x2_ASAP7_75t_L g2549 ( 
.A(n_2503),
.B(n_2286),
.Y(n_2549)
);

NOR2xp33_ASAP7_75t_R g2550 ( 
.A(n_2508),
.B(n_2481),
.Y(n_2550)
);

AND2x4_ASAP7_75t_L g2551 ( 
.A(n_2490),
.B(n_2305),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2446),
.Y(n_2552)
);

BUFx10_ASAP7_75t_L g2553 ( 
.A(n_2491),
.Y(n_2553)
);

NOR2xp33_ASAP7_75t_R g2554 ( 
.A(n_2530),
.B(n_2387),
.Y(n_2554)
);

AND2x2_ASAP7_75t_L g2555 ( 
.A(n_2451),
.B(n_2487),
.Y(n_2555)
);

NOR2xp33_ASAP7_75t_R g2556 ( 
.A(n_2530),
.B(n_1012),
.Y(n_2556)
);

AND2x4_ASAP7_75t_L g2557 ( 
.A(n_2495),
.B(n_2397),
.Y(n_2557)
);

AND2x2_ASAP7_75t_L g2558 ( 
.A(n_2484),
.B(n_2316),
.Y(n_2558)
);

XNOR2xp5_ASAP7_75t_SL g2559 ( 
.A(n_2499),
.B(n_2374),
.Y(n_2559)
);

NOR2xp33_ASAP7_75t_R g2560 ( 
.A(n_2494),
.B(n_2433),
.Y(n_2560)
);

XNOR2xp5_ASAP7_75t_L g2561 ( 
.A(n_2486),
.B(n_2389),
.Y(n_2561)
);

NOR2xp33_ASAP7_75t_R g2562 ( 
.A(n_2491),
.B(n_1013),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2447),
.Y(n_2563)
);

INVxp67_ASAP7_75t_L g2564 ( 
.A(n_2464),
.Y(n_2564)
);

NAND2xp33_ASAP7_75t_R g2565 ( 
.A(n_2442),
.B(n_2440),
.Y(n_2565)
);

XNOR2xp5_ASAP7_75t_L g2566 ( 
.A(n_2478),
.B(n_2522),
.Y(n_2566)
);

NAND2xp5_ASAP7_75t_L g2567 ( 
.A(n_2459),
.B(n_2379),
.Y(n_2567)
);

INVx1_ASAP7_75t_L g2568 ( 
.A(n_2458),
.Y(n_2568)
);

NOR2xp33_ASAP7_75t_R g2569 ( 
.A(n_2444),
.B(n_1015),
.Y(n_2569)
);

AND2x2_ASAP7_75t_L g2570 ( 
.A(n_2519),
.B(n_2406),
.Y(n_2570)
);

NAND2xp33_ASAP7_75t_R g2571 ( 
.A(n_2434),
.B(n_2419),
.Y(n_2571)
);

NAND2xp33_ASAP7_75t_R g2572 ( 
.A(n_2435),
.B(n_2401),
.Y(n_2572)
);

OR2x6_ASAP7_75t_L g2573 ( 
.A(n_2517),
.B(n_2312),
.Y(n_2573)
);

NAND2xp5_ASAP7_75t_L g2574 ( 
.A(n_2438),
.B(n_2324),
.Y(n_2574)
);

AND2x2_ASAP7_75t_L g2575 ( 
.A(n_2467),
.B(n_2320),
.Y(n_2575)
);

INVx1_ASAP7_75t_L g2576 ( 
.A(n_2465),
.Y(n_2576)
);

AND2x2_ASAP7_75t_L g2577 ( 
.A(n_2460),
.B(n_2340),
.Y(n_2577)
);

AND2x2_ASAP7_75t_L g2578 ( 
.A(n_2526),
.B(n_2405),
.Y(n_2578)
);

INVx1_ASAP7_75t_L g2579 ( 
.A(n_2466),
.Y(n_2579)
);

INVxp67_ASAP7_75t_L g2580 ( 
.A(n_2472),
.Y(n_2580)
);

NAND2xp5_ASAP7_75t_L g2581 ( 
.A(n_2453),
.B(n_2322),
.Y(n_2581)
);

NOR2xp33_ASAP7_75t_R g2582 ( 
.A(n_2489),
.B(n_1018),
.Y(n_2582)
);

INVxp67_ASAP7_75t_L g2583 ( 
.A(n_2488),
.Y(n_2583)
);

AND2x4_ASAP7_75t_L g2584 ( 
.A(n_2436),
.B(n_2402),
.Y(n_2584)
);

NOR2xp33_ASAP7_75t_R g2585 ( 
.A(n_2441),
.B(n_1019),
.Y(n_2585)
);

INVxp67_ASAP7_75t_L g2586 ( 
.A(n_2443),
.Y(n_2586)
);

NAND2xp33_ASAP7_75t_R g2587 ( 
.A(n_2527),
.B(n_2334),
.Y(n_2587)
);

NAND2xp5_ASAP7_75t_L g2588 ( 
.A(n_2445),
.B(n_2293),
.Y(n_2588)
);

NOR2xp33_ASAP7_75t_R g2589 ( 
.A(n_2468),
.B(n_1021),
.Y(n_2589)
);

XNOR2xp5_ASAP7_75t_L g2590 ( 
.A(n_2469),
.B(n_2314),
.Y(n_2590)
);

INVx1_ASAP7_75t_L g2591 ( 
.A(n_2463),
.Y(n_2591)
);

AND2x4_ASAP7_75t_L g2592 ( 
.A(n_2476),
.B(n_2416),
.Y(n_2592)
);

CKINVDCx5p33_ASAP7_75t_R g2593 ( 
.A(n_2545),
.Y(n_2593)
);

HB1xp67_ASAP7_75t_L g2594 ( 
.A(n_2546),
.Y(n_2594)
);

INVx1_ASAP7_75t_L g2595 ( 
.A(n_2542),
.Y(n_2595)
);

OAI22xp5_ASAP7_75t_L g2596 ( 
.A1(n_2534),
.A2(n_2511),
.B1(n_2515),
.B2(n_2479),
.Y(n_2596)
);

INVx1_ASAP7_75t_L g2597 ( 
.A(n_2547),
.Y(n_2597)
);

INVx1_ASAP7_75t_L g2598 ( 
.A(n_2552),
.Y(n_2598)
);

INVx2_ASAP7_75t_L g2599 ( 
.A(n_2591),
.Y(n_2599)
);

OR2x2_ASAP7_75t_L g2600 ( 
.A(n_2564),
.B(n_2518),
.Y(n_2600)
);

AND2x2_ASAP7_75t_L g2601 ( 
.A(n_2578),
.B(n_2521),
.Y(n_2601)
);

INVx2_ASAP7_75t_SL g2602 ( 
.A(n_2553),
.Y(n_2602)
);

INVx2_ASAP7_75t_SL g2603 ( 
.A(n_2560),
.Y(n_2603)
);

NAND2xp5_ASAP7_75t_L g2604 ( 
.A(n_2549),
.B(n_2457),
.Y(n_2604)
);

NOR2xp33_ASAP7_75t_L g2605 ( 
.A(n_2548),
.B(n_2462),
.Y(n_2605)
);

OR2x2_ASAP7_75t_L g2606 ( 
.A(n_2563),
.B(n_2507),
.Y(n_2606)
);

AND2x2_ASAP7_75t_L g2607 ( 
.A(n_2555),
.B(n_2510),
.Y(n_2607)
);

INVx1_ASAP7_75t_L g2608 ( 
.A(n_2568),
.Y(n_2608)
);

NAND2xp5_ASAP7_75t_L g2609 ( 
.A(n_2586),
.B(n_2514),
.Y(n_2609)
);

INVxp67_ASAP7_75t_SL g2610 ( 
.A(n_2588),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2558),
.B(n_2576),
.Y(n_2611)
);

AND2x2_ASAP7_75t_L g2612 ( 
.A(n_2579),
.B(n_2513),
.Y(n_2612)
);

HB1xp67_ASAP7_75t_L g2613 ( 
.A(n_2577),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2551),
.Y(n_2614)
);

INVx2_ASAP7_75t_L g2615 ( 
.A(n_2557),
.Y(n_2615)
);

INVxp67_ASAP7_75t_L g2616 ( 
.A(n_2580),
.Y(n_2616)
);

INVx1_ASAP7_75t_L g2617 ( 
.A(n_2592),
.Y(n_2617)
);

AND2x2_ASAP7_75t_L g2618 ( 
.A(n_2590),
.B(n_2485),
.Y(n_2618)
);

AND2x2_ASAP7_75t_L g2619 ( 
.A(n_2570),
.B(n_2492),
.Y(n_2619)
);

AND2x2_ASAP7_75t_L g2620 ( 
.A(n_2575),
.B(n_2538),
.Y(n_2620)
);

INVx3_ASAP7_75t_L g2621 ( 
.A(n_2535),
.Y(n_2621)
);

NAND3xp33_ASAP7_75t_L g2622 ( 
.A(n_2587),
.B(n_2512),
.C(n_2501),
.Y(n_2622)
);

INVx2_ASAP7_75t_L g2623 ( 
.A(n_2584),
.Y(n_2623)
);

AND2x2_ASAP7_75t_L g2624 ( 
.A(n_2583),
.B(n_2500),
.Y(n_2624)
);

INVx3_ASAP7_75t_L g2625 ( 
.A(n_2537),
.Y(n_2625)
);

INVxp67_ASAP7_75t_L g2626 ( 
.A(n_2539),
.Y(n_2626)
);

INVx1_ASAP7_75t_L g2627 ( 
.A(n_2567),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2574),
.Y(n_2628)
);

BUFx2_ASAP7_75t_L g2629 ( 
.A(n_2550),
.Y(n_2629)
);

INVx2_ASAP7_75t_L g2630 ( 
.A(n_2581),
.Y(n_2630)
);

INVx1_ASAP7_75t_L g2631 ( 
.A(n_2559),
.Y(n_2631)
);

INVx1_ASAP7_75t_L g2632 ( 
.A(n_2573),
.Y(n_2632)
);

OR2x6_ASAP7_75t_L g2633 ( 
.A(n_2573),
.B(n_2439),
.Y(n_2633)
);

AND2x4_ASAP7_75t_SL g2634 ( 
.A(n_2544),
.B(n_2482),
.Y(n_2634)
);

INVx1_ASAP7_75t_L g2635 ( 
.A(n_2541),
.Y(n_2635)
);

AND2x2_ASAP7_75t_L g2636 ( 
.A(n_2566),
.B(n_2505),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2561),
.Y(n_2637)
);

NAND2xp5_ASAP7_75t_L g2638 ( 
.A(n_2585),
.B(n_2455),
.Y(n_2638)
);

AOI22xp33_ASAP7_75t_L g2639 ( 
.A1(n_2582),
.A2(n_2532),
.B1(n_2531),
.B2(n_2431),
.Y(n_2639)
);

INVx1_ASAP7_75t_L g2640 ( 
.A(n_2589),
.Y(n_2640)
);

NAND2xp5_ASAP7_75t_L g2641 ( 
.A(n_2554),
.B(n_2474),
.Y(n_2641)
);

INVx3_ASAP7_75t_SL g2642 ( 
.A(n_2543),
.Y(n_2642)
);

INVx2_ASAP7_75t_L g2643 ( 
.A(n_2571),
.Y(n_2643)
);

AND2x4_ASAP7_75t_L g2644 ( 
.A(n_2572),
.B(n_2523),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2569),
.Y(n_2645)
);

INVx1_ASAP7_75t_L g2646 ( 
.A(n_2556),
.Y(n_2646)
);

INVx1_ASAP7_75t_L g2647 ( 
.A(n_2562),
.Y(n_2647)
);

AND2x2_ASAP7_75t_L g2648 ( 
.A(n_2565),
.B(n_2533),
.Y(n_2648)
);

NAND2xp5_ASAP7_75t_L g2649 ( 
.A(n_2540),
.B(n_2483),
.Y(n_2649)
);

AOI22xp33_ASAP7_75t_L g2650 ( 
.A1(n_2536),
.A2(n_2477),
.B1(n_2294),
.B2(n_2480),
.Y(n_2650)
);

INVx1_ASAP7_75t_L g2651 ( 
.A(n_2542),
.Y(n_2651)
);

NAND2xp5_ASAP7_75t_L g2652 ( 
.A(n_2564),
.B(n_2498),
.Y(n_2652)
);

OAI31xp33_ASAP7_75t_L g2653 ( 
.A1(n_2622),
.A2(n_2339),
.A3(n_2371),
.B(n_2365),
.Y(n_2653)
);

INVx1_ASAP7_75t_L g2654 ( 
.A(n_2595),
.Y(n_2654)
);

OAI22xp5_ASAP7_75t_L g2655 ( 
.A1(n_2639),
.A2(n_2348),
.B1(n_2529),
.B2(n_2520),
.Y(n_2655)
);

AND2x2_ASAP7_75t_SL g2656 ( 
.A(n_2644),
.B(n_2516),
.Y(n_2656)
);

INVx1_ASAP7_75t_L g2657 ( 
.A(n_2597),
.Y(n_2657)
);

AND2x2_ASAP7_75t_L g2658 ( 
.A(n_2601),
.B(n_2437),
.Y(n_2658)
);

BUFx2_ASAP7_75t_L g2659 ( 
.A(n_2613),
.Y(n_2659)
);

INVx2_ASAP7_75t_L g2660 ( 
.A(n_2599),
.Y(n_2660)
);

OAI22xp5_ASAP7_75t_L g2661 ( 
.A1(n_2596),
.A2(n_2629),
.B1(n_2640),
.B2(n_2638),
.Y(n_2661)
);

NAND2xp5_ASAP7_75t_L g2662 ( 
.A(n_2610),
.B(n_2525),
.Y(n_2662)
);

AND2x4_ASAP7_75t_L g2663 ( 
.A(n_2615),
.B(n_2525),
.Y(n_2663)
);

AND2x2_ASAP7_75t_L g2664 ( 
.A(n_2620),
.B(n_2450),
.Y(n_2664)
);

INVx1_ASAP7_75t_L g2665 ( 
.A(n_2598),
.Y(n_2665)
);

INVx1_ASAP7_75t_L g2666 ( 
.A(n_2608),
.Y(n_2666)
);

OR2x2_ASAP7_75t_L g2667 ( 
.A(n_2600),
.B(n_2313),
.Y(n_2667)
);

INVx2_ASAP7_75t_L g2668 ( 
.A(n_2651),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2594),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2612),
.Y(n_2670)
);

INVx1_ASAP7_75t_L g2671 ( 
.A(n_2606),
.Y(n_2671)
);

INVxp67_ASAP7_75t_SL g2672 ( 
.A(n_2643),
.Y(n_2672)
);

AND2x2_ASAP7_75t_L g2673 ( 
.A(n_2636),
.B(n_2496),
.Y(n_2673)
);

AND2x2_ASAP7_75t_L g2674 ( 
.A(n_2648),
.B(n_2496),
.Y(n_2674)
);

NAND2xp5_ASAP7_75t_L g2675 ( 
.A(n_2630),
.B(n_2313),
.Y(n_2675)
);

HB1xp67_ASAP7_75t_L g2676 ( 
.A(n_2611),
.Y(n_2676)
);

OR2x2_ASAP7_75t_L g2677 ( 
.A(n_2649),
.B(n_2493),
.Y(n_2677)
);

BUFx2_ASAP7_75t_L g2678 ( 
.A(n_2644),
.Y(n_2678)
);

INVx1_ASAP7_75t_SL g2679 ( 
.A(n_2629),
.Y(n_2679)
);

AND2x2_ASAP7_75t_L g2680 ( 
.A(n_2618),
.B(n_2497),
.Y(n_2680)
);

INVx2_ASAP7_75t_L g2681 ( 
.A(n_2624),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2652),
.Y(n_2682)
);

OR2x2_ASAP7_75t_L g2683 ( 
.A(n_2604),
.B(n_2367),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2607),
.Y(n_2684)
);

AND2x2_ASAP7_75t_L g2685 ( 
.A(n_2619),
.B(n_2475),
.Y(n_2685)
);

OR2x6_ASAP7_75t_L g2686 ( 
.A(n_2632),
.B(n_2452),
.Y(n_2686)
);

INVx1_ASAP7_75t_L g2687 ( 
.A(n_2609),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2617),
.Y(n_2688)
);

INVx2_ASAP7_75t_L g2689 ( 
.A(n_2614),
.Y(n_2689)
);

NAND2xp5_ASAP7_75t_L g2690 ( 
.A(n_2628),
.B(n_2627),
.Y(n_2690)
);

AOI31xp33_ASAP7_75t_L g2691 ( 
.A1(n_2631),
.A2(n_2326),
.A3(n_2421),
.B(n_59),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2616),
.B(n_2524),
.Y(n_2692)
);

INVx2_ASAP7_75t_L g2693 ( 
.A(n_2623),
.Y(n_2693)
);

AND2x4_ASAP7_75t_L g2694 ( 
.A(n_2634),
.B(n_2356),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2641),
.Y(n_2695)
);

AND2x2_ASAP7_75t_L g2696 ( 
.A(n_2603),
.B(n_2358),
.Y(n_2696)
);

INVx2_ASAP7_75t_SL g2697 ( 
.A(n_2621),
.Y(n_2697)
);

AND2x2_ASAP7_75t_L g2698 ( 
.A(n_2635),
.B(n_2362),
.Y(n_2698)
);

AND2x2_ASAP7_75t_L g2699 ( 
.A(n_2625),
.B(n_2347),
.Y(n_2699)
);

AOI222xp33_ASAP7_75t_L g2700 ( 
.A1(n_2605),
.A2(n_85),
.B1(n_66),
.B2(n_93),
.C1(n_75),
.C2(n_56),
.Y(n_2700)
);

INVx2_ASAP7_75t_L g2701 ( 
.A(n_2626),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2633),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2633),
.Y(n_2703)
);

INVx2_ASAP7_75t_L g2704 ( 
.A(n_2602),
.Y(n_2704)
);

INVx2_ASAP7_75t_L g2705 ( 
.A(n_2645),
.Y(n_2705)
);

NAND2x1_ASAP7_75t_L g2706 ( 
.A(n_2650),
.B(n_2382),
.Y(n_2706)
);

AND2x2_ASAP7_75t_L g2707 ( 
.A(n_2647),
.B(n_2336),
.Y(n_2707)
);

AND2x2_ASAP7_75t_L g2708 ( 
.A(n_2646),
.B(n_2364),
.Y(n_2708)
);

INVx2_ASAP7_75t_L g2709 ( 
.A(n_2637),
.Y(n_2709)
);

OR2x2_ASAP7_75t_L g2710 ( 
.A(n_2642),
.B(n_2300),
.Y(n_2710)
);

AND2x2_ASAP7_75t_L g2711 ( 
.A(n_2593),
.B(n_2369),
.Y(n_2711)
);

INVx2_ASAP7_75t_L g2712 ( 
.A(n_2599),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2595),
.Y(n_2713)
);

AO21x2_ASAP7_75t_L g2714 ( 
.A1(n_2643),
.A2(n_2392),
.B(n_2425),
.Y(n_2714)
);

OAI221xp5_ASAP7_75t_L g2715 ( 
.A1(n_2622),
.A2(n_61),
.B1(n_57),
.B2(n_60),
.C(n_62),
.Y(n_2715)
);

OR2x2_ASAP7_75t_L g2716 ( 
.A(n_2613),
.B(n_2370),
.Y(n_2716)
);

INVx2_ASAP7_75t_SL g2717 ( 
.A(n_2621),
.Y(n_2717)
);

AOI221xp5_ASAP7_75t_L g2718 ( 
.A1(n_2622),
.A2(n_63),
.B1(n_60),
.B2(n_62),
.C(n_64),
.Y(n_2718)
);

AND2x2_ASAP7_75t_L g2719 ( 
.A(n_2601),
.B(n_2430),
.Y(n_2719)
);

AND2x2_ASAP7_75t_L g2720 ( 
.A(n_2601),
.B(n_63),
.Y(n_2720)
);

AOI22xp33_ASAP7_75t_L g2721 ( 
.A1(n_2622),
.A2(n_68),
.B1(n_64),
.B2(n_65),
.Y(n_2721)
);

NAND2xp5_ASAP7_75t_L g2722 ( 
.A(n_2610),
.B(n_65),
.Y(n_2722)
);

INVx2_ASAP7_75t_L g2723 ( 
.A(n_2599),
.Y(n_2723)
);

INVx2_ASAP7_75t_L g2724 ( 
.A(n_2599),
.Y(n_2724)
);

NAND4xp25_ASAP7_75t_L g2725 ( 
.A(n_2622),
.B(n_70),
.C(n_68),
.D(n_69),
.Y(n_2725)
);

INVx1_ASAP7_75t_L g2726 ( 
.A(n_2595),
.Y(n_2726)
);

BUFx2_ASAP7_75t_SL g2727 ( 
.A(n_2603),
.Y(n_2727)
);

OAI21xp33_ASAP7_75t_L g2728 ( 
.A1(n_2622),
.A2(n_69),
.B(n_70),
.Y(n_2728)
);

INVx1_ASAP7_75t_L g2729 ( 
.A(n_2595),
.Y(n_2729)
);

AND2x2_ASAP7_75t_L g2730 ( 
.A(n_2601),
.B(n_71),
.Y(n_2730)
);

INVx5_ASAP7_75t_L g2731 ( 
.A(n_2633),
.Y(n_2731)
);

NAND2xp5_ASAP7_75t_L g2732 ( 
.A(n_2610),
.B(n_71),
.Y(n_2732)
);

AOI22xp33_ASAP7_75t_L g2733 ( 
.A1(n_2622),
.A2(n_74),
.B1(n_72),
.B2(n_73),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2695),
.B(n_72),
.Y(n_2734)
);

NAND2xp5_ASAP7_75t_L g2735 ( 
.A(n_2687),
.B(n_73),
.Y(n_2735)
);

AND2x2_ASAP7_75t_L g2736 ( 
.A(n_2659),
.B(n_74),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2654),
.Y(n_2737)
);

AND2x2_ASAP7_75t_L g2738 ( 
.A(n_2678),
.B(n_76),
.Y(n_2738)
);

AND2x4_ASAP7_75t_L g2739 ( 
.A(n_2702),
.B(n_76),
.Y(n_2739)
);

AND2x2_ASAP7_75t_L g2740 ( 
.A(n_2678),
.B(n_77),
.Y(n_2740)
);

INVx2_ASAP7_75t_L g2741 ( 
.A(n_2669),
.Y(n_2741)
);

INVx1_ASAP7_75t_L g2742 ( 
.A(n_2657),
.Y(n_2742)
);

AOI22xp5_ASAP7_75t_L g2743 ( 
.A1(n_2728),
.A2(n_80),
.B1(n_77),
.B2(n_78),
.Y(n_2743)
);

AND2x2_ASAP7_75t_L g2744 ( 
.A(n_2676),
.B(n_81),
.Y(n_2744)
);

NAND2xp5_ASAP7_75t_L g2745 ( 
.A(n_2682),
.B(n_81),
.Y(n_2745)
);

BUFx2_ASAP7_75t_L g2746 ( 
.A(n_2703),
.Y(n_2746)
);

OR2x2_ASAP7_75t_L g2747 ( 
.A(n_2671),
.B(n_82),
.Y(n_2747)
);

AND2x4_ASAP7_75t_L g2748 ( 
.A(n_2705),
.B(n_82),
.Y(n_2748)
);

INVx2_ASAP7_75t_L g2749 ( 
.A(n_2668),
.Y(n_2749)
);

NAND2xp5_ASAP7_75t_L g2750 ( 
.A(n_2672),
.B(n_84),
.Y(n_2750)
);

NAND2xp5_ASAP7_75t_L g2751 ( 
.A(n_2690),
.B(n_84),
.Y(n_2751)
);

NAND2xp5_ASAP7_75t_L g2752 ( 
.A(n_2680),
.B(n_85),
.Y(n_2752)
);

NOR2xp33_ASAP7_75t_L g2753 ( 
.A(n_2661),
.B(n_86),
.Y(n_2753)
);

INVx3_ASAP7_75t_L g2754 ( 
.A(n_2704),
.Y(n_2754)
);

NAND2xp5_ASAP7_75t_L g2755 ( 
.A(n_2677),
.B(n_86),
.Y(n_2755)
);

AND2x4_ASAP7_75t_L g2756 ( 
.A(n_2681),
.B(n_2693),
.Y(n_2756)
);

INVx1_ASAP7_75t_L g2757 ( 
.A(n_2665),
.Y(n_2757)
);

INVx2_ASAP7_75t_L g2758 ( 
.A(n_2666),
.Y(n_2758)
);

INVx1_ASAP7_75t_L g2759 ( 
.A(n_2713),
.Y(n_2759)
);

AND2x2_ASAP7_75t_L g2760 ( 
.A(n_2679),
.B(n_87),
.Y(n_2760)
);

NAND2xp5_ASAP7_75t_L g2761 ( 
.A(n_2660),
.B(n_88),
.Y(n_2761)
);

INVx1_ASAP7_75t_L g2762 ( 
.A(n_2726),
.Y(n_2762)
);

NAND2xp5_ASAP7_75t_L g2763 ( 
.A(n_2712),
.B(n_88),
.Y(n_2763)
);

INVxp67_ASAP7_75t_SL g2764 ( 
.A(n_2662),
.Y(n_2764)
);

NAND2xp5_ASAP7_75t_L g2765 ( 
.A(n_2723),
.B(n_89),
.Y(n_2765)
);

INVx1_ASAP7_75t_L g2766 ( 
.A(n_2729),
.Y(n_2766)
);

INVx1_ASAP7_75t_L g2767 ( 
.A(n_2724),
.Y(n_2767)
);

INVx3_ASAP7_75t_SL g2768 ( 
.A(n_2697),
.Y(n_2768)
);

INVx1_ASAP7_75t_L g2769 ( 
.A(n_2670),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2684),
.Y(n_2770)
);

AND2x2_ASAP7_75t_L g2771 ( 
.A(n_2656),
.B(n_89),
.Y(n_2771)
);

AND2x2_ASAP7_75t_L g2772 ( 
.A(n_2658),
.B(n_90),
.Y(n_2772)
);

OR2x2_ASAP7_75t_L g2773 ( 
.A(n_2667),
.B(n_90),
.Y(n_2773)
);

INVx2_ASAP7_75t_L g2774 ( 
.A(n_2688),
.Y(n_2774)
);

AND2x2_ASAP7_75t_L g2775 ( 
.A(n_2689),
.B(n_91),
.Y(n_2775)
);

INVx1_ASAP7_75t_L g2776 ( 
.A(n_2692),
.Y(n_2776)
);

AND2x2_ASAP7_75t_L g2777 ( 
.A(n_2717),
.B(n_92),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2675),
.Y(n_2778)
);

INVx1_ASAP7_75t_L g2779 ( 
.A(n_2674),
.Y(n_2779)
);

AND2x2_ASAP7_75t_L g2780 ( 
.A(n_2727),
.B(n_94),
.Y(n_2780)
);

OR2x2_ASAP7_75t_L g2781 ( 
.A(n_2683),
.B(n_94),
.Y(n_2781)
);

INVx2_ASAP7_75t_L g2782 ( 
.A(n_2701),
.Y(n_2782)
);

INVx1_ASAP7_75t_L g2783 ( 
.A(n_2716),
.Y(n_2783)
);

AND2x2_ASAP7_75t_L g2784 ( 
.A(n_2673),
.B(n_2731),
.Y(n_2784)
);

INVxp67_ASAP7_75t_L g2785 ( 
.A(n_2722),
.Y(n_2785)
);

INVx1_ASAP7_75t_L g2786 ( 
.A(n_2663),
.Y(n_2786)
);

AND2x2_ASAP7_75t_L g2787 ( 
.A(n_2731),
.B(n_95),
.Y(n_2787)
);

AND2x2_ASAP7_75t_L g2788 ( 
.A(n_2731),
.B(n_95),
.Y(n_2788)
);

HB1xp67_ASAP7_75t_L g2789 ( 
.A(n_2685),
.Y(n_2789)
);

INVx1_ASAP7_75t_L g2790 ( 
.A(n_2732),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2664),
.B(n_96),
.Y(n_2791)
);

INVx3_ASAP7_75t_L g2792 ( 
.A(n_2709),
.Y(n_2792)
);

NAND2xp5_ASAP7_75t_L g2793 ( 
.A(n_2720),
.B(n_97),
.Y(n_2793)
);

AND2x2_ASAP7_75t_L g2794 ( 
.A(n_2719),
.B(n_97),
.Y(n_2794)
);

AND2x2_ASAP7_75t_L g2795 ( 
.A(n_2711),
.B(n_98),
.Y(n_2795)
);

INVx2_ASAP7_75t_L g2796 ( 
.A(n_2698),
.Y(n_2796)
);

AND2x2_ASAP7_75t_L g2797 ( 
.A(n_2730),
.B(n_99),
.Y(n_2797)
);

INVx1_ASAP7_75t_L g2798 ( 
.A(n_2699),
.Y(n_2798)
);

OR2x2_ASAP7_75t_L g2799 ( 
.A(n_2706),
.B(n_99),
.Y(n_2799)
);

OR2x2_ASAP7_75t_L g2800 ( 
.A(n_2710),
.B(n_100),
.Y(n_2800)
);

AND2x2_ASAP7_75t_L g2801 ( 
.A(n_2696),
.B(n_102),
.Y(n_2801)
);

AND2x2_ASAP7_75t_L g2802 ( 
.A(n_2707),
.B(n_103),
.Y(n_2802)
);

OR2x2_ASAP7_75t_L g2803 ( 
.A(n_2686),
.B(n_103),
.Y(n_2803)
);

AND2x2_ASAP7_75t_L g2804 ( 
.A(n_2708),
.B(n_104),
.Y(n_2804)
);

AND2x2_ASAP7_75t_L g2805 ( 
.A(n_2686),
.B(n_2714),
.Y(n_2805)
);

INVx1_ASAP7_75t_L g2806 ( 
.A(n_2655),
.Y(n_2806)
);

INVx1_ASAP7_75t_L g2807 ( 
.A(n_2694),
.Y(n_2807)
);

AND2x2_ASAP7_75t_L g2808 ( 
.A(n_2653),
.B(n_104),
.Y(n_2808)
);

INVx4_ASAP7_75t_L g2809 ( 
.A(n_2691),
.Y(n_2809)
);

AND2x4_ASAP7_75t_L g2810 ( 
.A(n_2721),
.B(n_105),
.Y(n_2810)
);

INVx3_ASAP7_75t_L g2811 ( 
.A(n_2725),
.Y(n_2811)
);

OR2x2_ASAP7_75t_L g2812 ( 
.A(n_2715),
.B(n_105),
.Y(n_2812)
);

NAND2xp5_ASAP7_75t_L g2813 ( 
.A(n_2700),
.B(n_106),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2733),
.B(n_106),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2718),
.Y(n_2815)
);

AND2x2_ASAP7_75t_L g2816 ( 
.A(n_2659),
.B(n_107),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2654),
.Y(n_2817)
);

AND2x2_ASAP7_75t_L g2818 ( 
.A(n_2659),
.B(n_108),
.Y(n_2818)
);

NAND2x1_ASAP7_75t_L g2819 ( 
.A(n_2678),
.B(n_109),
.Y(n_2819)
);

OR2x2_ASAP7_75t_L g2820 ( 
.A(n_2659),
.B(n_109),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2654),
.Y(n_2821)
);

NAND2xp5_ASAP7_75t_L g2822 ( 
.A(n_2695),
.B(n_110),
.Y(n_2822)
);

AND2x2_ASAP7_75t_L g2823 ( 
.A(n_2659),
.B(n_110),
.Y(n_2823)
);

NOR2x1_ASAP7_75t_L g2824 ( 
.A(n_2669),
.B(n_112),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2659),
.B(n_113),
.Y(n_2825)
);

INVx1_ASAP7_75t_L g2826 ( 
.A(n_2654),
.Y(n_2826)
);

AND2x2_ASAP7_75t_L g2827 ( 
.A(n_2659),
.B(n_113),
.Y(n_2827)
);

INVx1_ASAP7_75t_L g2828 ( 
.A(n_2654),
.Y(n_2828)
);

OR2x2_ASAP7_75t_L g2829 ( 
.A(n_2659),
.B(n_114),
.Y(n_2829)
);

AND2x4_ASAP7_75t_L g2830 ( 
.A(n_2702),
.B(n_114),
.Y(n_2830)
);

AND2x2_ASAP7_75t_L g2831 ( 
.A(n_2659),
.B(n_115),
.Y(n_2831)
);

INVx1_ASAP7_75t_L g2832 ( 
.A(n_2654),
.Y(n_2832)
);

AND2x2_ASAP7_75t_L g2833 ( 
.A(n_2659),
.B(n_116),
.Y(n_2833)
);

AND2x2_ASAP7_75t_L g2834 ( 
.A(n_2659),
.B(n_116),
.Y(n_2834)
);

INVx2_ASAP7_75t_SL g2835 ( 
.A(n_2697),
.Y(n_2835)
);

AND2x2_ASAP7_75t_L g2836 ( 
.A(n_2659),
.B(n_117),
.Y(n_2836)
);

INVx2_ASAP7_75t_L g2837 ( 
.A(n_2669),
.Y(n_2837)
);

AND2x4_ASAP7_75t_L g2838 ( 
.A(n_2702),
.B(n_118),
.Y(n_2838)
);

AND2x2_ASAP7_75t_L g2839 ( 
.A(n_2659),
.B(n_118),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2654),
.Y(n_2840)
);

AND2x4_ASAP7_75t_L g2841 ( 
.A(n_2702),
.B(n_119),
.Y(n_2841)
);

AND2x2_ASAP7_75t_L g2842 ( 
.A(n_2659),
.B(n_120),
.Y(n_2842)
);

NAND2xp5_ASAP7_75t_L g2843 ( 
.A(n_2695),
.B(n_120),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2659),
.B(n_121),
.Y(n_2844)
);

NOR2xp33_ASAP7_75t_L g2845 ( 
.A(n_2661),
.B(n_122),
.Y(n_2845)
);

INVx1_ASAP7_75t_L g2846 ( 
.A(n_2654),
.Y(n_2846)
);

AND3x2_ASAP7_75t_L g2847 ( 
.A(n_2718),
.B(n_123),
.C(n_124),
.Y(n_2847)
);

NAND2xp5_ASAP7_75t_L g2848 ( 
.A(n_2695),
.B(n_123),
.Y(n_2848)
);

OR2x2_ASAP7_75t_L g2849 ( 
.A(n_2659),
.B(n_124),
.Y(n_2849)
);

INVx1_ASAP7_75t_L g2850 ( 
.A(n_2737),
.Y(n_2850)
);

OAI22xp33_ASAP7_75t_L g2851 ( 
.A1(n_2809),
.A2(n_127),
.B1(n_125),
.B2(n_126),
.Y(n_2851)
);

CKINVDCx5p33_ASAP7_75t_R g2852 ( 
.A(n_2768),
.Y(n_2852)
);

NOR2x1_ASAP7_75t_L g2853 ( 
.A(n_2819),
.B(n_125),
.Y(n_2853)
);

INVx1_ASAP7_75t_L g2854 ( 
.A(n_2742),
.Y(n_2854)
);

OAI22xp33_ASAP7_75t_L g2855 ( 
.A1(n_2799),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_2855)
);

BUFx3_ASAP7_75t_L g2856 ( 
.A(n_2754),
.Y(n_2856)
);

AOI22xp5_ASAP7_75t_L g2857 ( 
.A1(n_2815),
.A2(n_131),
.B1(n_129),
.B2(n_130),
.Y(n_2857)
);

NAND2xp5_ASAP7_75t_L g2858 ( 
.A(n_2790),
.B(n_131),
.Y(n_2858)
);

NAND2xp33_ASAP7_75t_L g2859 ( 
.A(n_2808),
.B(n_132),
.Y(n_2859)
);

OAI22xp33_ASAP7_75t_L g2860 ( 
.A1(n_2806),
.A2(n_134),
.B1(n_132),
.B2(n_133),
.Y(n_2860)
);

INVxp33_ASAP7_75t_SL g2861 ( 
.A(n_2780),
.Y(n_2861)
);

NAND2xp5_ASAP7_75t_L g2862 ( 
.A(n_2764),
.B(n_134),
.Y(n_2862)
);

INVx3_ASAP7_75t_L g2863 ( 
.A(n_2756),
.Y(n_2863)
);

INVx1_ASAP7_75t_L g2864 ( 
.A(n_2757),
.Y(n_2864)
);

INVx2_ASAP7_75t_L g2865 ( 
.A(n_2746),
.Y(n_2865)
);

INVx1_ASAP7_75t_L g2866 ( 
.A(n_2759),
.Y(n_2866)
);

NAND2xp33_ASAP7_75t_SL g2867 ( 
.A(n_2819),
.B(n_135),
.Y(n_2867)
);

XNOR2xp5_ASAP7_75t_L g2868 ( 
.A(n_2797),
.B(n_135),
.Y(n_2868)
);

AOI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2753),
.A2(n_139),
.B1(n_136),
.B2(n_137),
.Y(n_2869)
);

CKINVDCx5p33_ASAP7_75t_R g2870 ( 
.A(n_2835),
.Y(n_2870)
);

AOI22xp5_ASAP7_75t_L g2871 ( 
.A1(n_2845),
.A2(n_140),
.B1(n_137),
.B2(n_139),
.Y(n_2871)
);

BUFx2_ASAP7_75t_L g2872 ( 
.A(n_2746),
.Y(n_2872)
);

NAND2xp5_ASAP7_75t_L g2873 ( 
.A(n_2785),
.B(n_140),
.Y(n_2873)
);

AO221x2_ASAP7_75t_L g2874 ( 
.A1(n_2813),
.A2(n_143),
.B1(n_141),
.B2(n_142),
.C(n_144),
.Y(n_2874)
);

CKINVDCx5p33_ASAP7_75t_R g2875 ( 
.A(n_2739),
.Y(n_2875)
);

NAND2xp33_ASAP7_75t_SL g2876 ( 
.A(n_2771),
.B(n_141),
.Y(n_2876)
);

CKINVDCx5p33_ASAP7_75t_R g2877 ( 
.A(n_2830),
.Y(n_2877)
);

OAI22xp33_ASAP7_75t_L g2878 ( 
.A1(n_2743),
.A2(n_145),
.B1(n_142),
.B2(n_143),
.Y(n_2878)
);

NAND2xp33_ASAP7_75t_SL g2879 ( 
.A(n_2787),
.B(n_146),
.Y(n_2879)
);

NOR2x1_ASAP7_75t_L g2880 ( 
.A(n_2824),
.B(n_147),
.Y(n_2880)
);

CKINVDCx20_ASAP7_75t_R g2881 ( 
.A(n_2793),
.Y(n_2881)
);

NAND2xp5_ASAP7_75t_L g2882 ( 
.A(n_2778),
.B(n_147),
.Y(n_2882)
);

INVxp67_ASAP7_75t_SL g2883 ( 
.A(n_2750),
.Y(n_2883)
);

NAND2xp5_ASAP7_75t_L g2884 ( 
.A(n_2782),
.B(n_148),
.Y(n_2884)
);

NAND2xp5_ASAP7_75t_L g2885 ( 
.A(n_2781),
.B(n_2783),
.Y(n_2885)
);

AO221x2_ASAP7_75t_L g2886 ( 
.A1(n_2734),
.A2(n_150),
.B1(n_148),
.B2(n_149),
.C(n_151),
.Y(n_2886)
);

NAND2xp5_ASAP7_75t_L g2887 ( 
.A(n_2741),
.B(n_150),
.Y(n_2887)
);

CKINVDCx5p33_ASAP7_75t_R g2888 ( 
.A(n_2838),
.Y(n_2888)
);

INVxp67_ASAP7_75t_L g2889 ( 
.A(n_2800),
.Y(n_2889)
);

NOR2xp33_ASAP7_75t_SL g2890 ( 
.A(n_2788),
.B(n_151),
.Y(n_2890)
);

NAND2xp5_ASAP7_75t_L g2891 ( 
.A(n_2837),
.B(n_152),
.Y(n_2891)
);

NAND2xp5_ASAP7_75t_L g2892 ( 
.A(n_2773),
.B(n_152),
.Y(n_2892)
);

OAI22xp33_ASAP7_75t_L g2893 ( 
.A1(n_2812),
.A2(n_155),
.B1(n_153),
.B2(n_154),
.Y(n_2893)
);

OAI22xp33_ASAP7_75t_L g2894 ( 
.A1(n_2803),
.A2(n_156),
.B1(n_153),
.B2(n_155),
.Y(n_2894)
);

INVx1_ASAP7_75t_L g2895 ( 
.A(n_2762),
.Y(n_2895)
);

NAND2xp5_ASAP7_75t_L g2896 ( 
.A(n_2776),
.B(n_2792),
.Y(n_2896)
);

INVx3_ASAP7_75t_L g2897 ( 
.A(n_2796),
.Y(n_2897)
);

NAND2xp5_ASAP7_75t_L g2898 ( 
.A(n_2798),
.B(n_2766),
.Y(n_2898)
);

NAND2xp33_ASAP7_75t_SL g2899 ( 
.A(n_2738),
.B(n_157),
.Y(n_2899)
);

AO221x2_ASAP7_75t_L g2900 ( 
.A1(n_2822),
.A2(n_160),
.B1(n_158),
.B2(n_159),
.C(n_161),
.Y(n_2900)
);

AO221x2_ASAP7_75t_L g2901 ( 
.A1(n_2843),
.A2(n_161),
.B1(n_159),
.B2(n_160),
.C(n_162),
.Y(n_2901)
);

NAND2xp5_ASAP7_75t_L g2902 ( 
.A(n_2817),
.B(n_163),
.Y(n_2902)
);

INVx2_ASAP7_75t_SL g2903 ( 
.A(n_2769),
.Y(n_2903)
);

NAND2xp5_ASAP7_75t_L g2904 ( 
.A(n_2821),
.B(n_163),
.Y(n_2904)
);

OAI22xp33_ASAP7_75t_L g2905 ( 
.A1(n_2811),
.A2(n_166),
.B1(n_164),
.B2(n_165),
.Y(n_2905)
);

NAND2xp5_ASAP7_75t_L g2906 ( 
.A(n_2826),
.B(n_164),
.Y(n_2906)
);

OAI22xp5_ASAP7_75t_SL g2907 ( 
.A1(n_2810),
.A2(n_168),
.B1(n_165),
.B2(n_167),
.Y(n_2907)
);

OAI22xp33_ASAP7_75t_L g2908 ( 
.A1(n_2820),
.A2(n_169),
.B1(n_167),
.B2(n_168),
.Y(n_2908)
);

NOR2xp33_ASAP7_75t_L g2909 ( 
.A(n_2751),
.B(n_170),
.Y(n_2909)
);

BUFx2_ASAP7_75t_L g2910 ( 
.A(n_2784),
.Y(n_2910)
);

NOR2xp33_ASAP7_75t_SL g2911 ( 
.A(n_2740),
.B(n_2760),
.Y(n_2911)
);

NAND2xp5_ASAP7_75t_L g2912 ( 
.A(n_2828),
.B(n_2832),
.Y(n_2912)
);

AO221x2_ASAP7_75t_L g2913 ( 
.A1(n_2848),
.A2(n_174),
.B1(n_172),
.B2(n_173),
.C(n_175),
.Y(n_2913)
);

AOI22xp5_ASAP7_75t_L g2914 ( 
.A1(n_2810),
.A2(n_2847),
.B1(n_2814),
.B2(n_2772),
.Y(n_2914)
);

NAND2xp5_ASAP7_75t_L g2915 ( 
.A(n_2840),
.B(n_173),
.Y(n_2915)
);

OAI22xp33_ASAP7_75t_L g2916 ( 
.A1(n_2829),
.A2(n_176),
.B1(n_174),
.B2(n_175),
.Y(n_2916)
);

NAND3xp33_ASAP7_75t_L g2917 ( 
.A(n_2805),
.B(n_178),
.C(n_179),
.Y(n_2917)
);

NAND2xp5_ASAP7_75t_L g2918 ( 
.A(n_2846),
.B(n_179),
.Y(n_2918)
);

OAI22xp33_ASAP7_75t_L g2919 ( 
.A1(n_2849),
.A2(n_182),
.B1(n_180),
.B2(n_181),
.Y(n_2919)
);

NOR2x1_ASAP7_75t_L g2920 ( 
.A(n_2735),
.B(n_180),
.Y(n_2920)
);

NAND2xp5_ASAP7_75t_L g2921 ( 
.A(n_2779),
.B(n_183),
.Y(n_2921)
);

NAND2xp5_ASAP7_75t_L g2922 ( 
.A(n_2767),
.B(n_183),
.Y(n_2922)
);

NOR2xp33_ASAP7_75t_L g2923 ( 
.A(n_2745),
.B(n_184),
.Y(n_2923)
);

AND2x4_ASAP7_75t_L g2924 ( 
.A(n_2807),
.B(n_184),
.Y(n_2924)
);

NAND2xp5_ASAP7_75t_L g2925 ( 
.A(n_2758),
.B(n_185),
.Y(n_2925)
);

BUFx2_ASAP7_75t_L g2926 ( 
.A(n_2786),
.Y(n_2926)
);

CKINVDCx5p33_ASAP7_75t_R g2927 ( 
.A(n_2841),
.Y(n_2927)
);

OAI221xp5_ASAP7_75t_L g2928 ( 
.A1(n_2755),
.A2(n_187),
.B1(n_185),
.B2(n_186),
.C(n_188),
.Y(n_2928)
);

NOR2x1_ASAP7_75t_L g2929 ( 
.A(n_2736),
.B(n_186),
.Y(n_2929)
);

AND2x2_ASAP7_75t_L g2930 ( 
.A(n_2789),
.B(n_2770),
.Y(n_2930)
);

NAND2xp5_ASAP7_75t_L g2931 ( 
.A(n_2774),
.B(n_187),
.Y(n_2931)
);

NAND2xp33_ASAP7_75t_SL g2932 ( 
.A(n_2816),
.B(n_188),
.Y(n_2932)
);

NAND2xp5_ASAP7_75t_SL g2933 ( 
.A(n_2748),
.B(n_189),
.Y(n_2933)
);

OAI22xp33_ASAP7_75t_L g2934 ( 
.A1(n_2747),
.A2(n_192),
.B1(n_190),
.B2(n_191),
.Y(n_2934)
);

AOI22xp5_ASAP7_75t_L g2935 ( 
.A1(n_2795),
.A2(n_195),
.B1(n_191),
.B2(n_193),
.Y(n_2935)
);

NOR2xp33_ASAP7_75t_SL g2936 ( 
.A(n_2818),
.B(n_193),
.Y(n_2936)
);

OAI22xp33_ASAP7_75t_L g2937 ( 
.A1(n_2752),
.A2(n_197),
.B1(n_195),
.B2(n_196),
.Y(n_2937)
);

AND2x2_ASAP7_75t_L g2938 ( 
.A(n_2749),
.B(n_196),
.Y(n_2938)
);

NAND2xp5_ASAP7_75t_L g2939 ( 
.A(n_2791),
.B(n_197),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2794),
.B(n_198),
.Y(n_2940)
);

AOI22xp5_ASAP7_75t_L g2941 ( 
.A1(n_2802),
.A2(n_202),
.B1(n_200),
.B2(n_201),
.Y(n_2941)
);

NAND2xp5_ASAP7_75t_L g2942 ( 
.A(n_2801),
.B(n_200),
.Y(n_2942)
);

NAND2xp5_ASAP7_75t_L g2943 ( 
.A(n_2823),
.B(n_201),
.Y(n_2943)
);

NAND2xp5_ASAP7_75t_L g2944 ( 
.A(n_2825),
.B(n_203),
.Y(n_2944)
);

AO221x2_ASAP7_75t_L g2945 ( 
.A1(n_2761),
.A2(n_205),
.B1(n_203),
.B2(n_204),
.C(n_206),
.Y(n_2945)
);

AO221x2_ASAP7_75t_L g2946 ( 
.A1(n_2763),
.A2(n_208),
.B1(n_204),
.B2(n_207),
.C(n_209),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2765),
.Y(n_2947)
);

OAI22xp33_ASAP7_75t_L g2948 ( 
.A1(n_2804),
.A2(n_210),
.B1(n_207),
.B2(n_208),
.Y(n_2948)
);

AOI22xp5_ASAP7_75t_L g2949 ( 
.A1(n_2744),
.A2(n_212),
.B1(n_210),
.B2(n_211),
.Y(n_2949)
);

NAND2xp5_ASAP7_75t_L g2950 ( 
.A(n_2827),
.B(n_211),
.Y(n_2950)
);

AOI22xp5_ASAP7_75t_L g2951 ( 
.A1(n_2831),
.A2(n_215),
.B1(n_213),
.B2(n_214),
.Y(n_2951)
);

INVxp33_ASAP7_75t_SL g2952 ( 
.A(n_2833),
.Y(n_2952)
);

INVx1_ASAP7_75t_L g2953 ( 
.A(n_2775),
.Y(n_2953)
);

NAND2xp5_ASAP7_75t_L g2954 ( 
.A(n_2834),
.B(n_213),
.Y(n_2954)
);

AOI221xp5_ASAP7_75t_L g2955 ( 
.A1(n_2836),
.A2(n_218),
.B1(n_216),
.B2(n_217),
.C(n_219),
.Y(n_2955)
);

NAND2xp33_ASAP7_75t_SL g2956 ( 
.A(n_2839),
.B(n_216),
.Y(n_2956)
);

CKINVDCx5p33_ASAP7_75t_R g2957 ( 
.A(n_2777),
.Y(n_2957)
);

NAND2xp5_ASAP7_75t_L g2958 ( 
.A(n_2842),
.B(n_217),
.Y(n_2958)
);

NOR2xp67_ASAP7_75t_L g2959 ( 
.A(n_2844),
.B(n_218),
.Y(n_2959)
);

BUFx2_ASAP7_75t_L g2960 ( 
.A(n_2768),
.Y(n_2960)
);

OAI22xp33_ASAP7_75t_L g2961 ( 
.A1(n_2809),
.A2(n_222),
.B1(n_220),
.B2(n_221),
.Y(n_2961)
);

NOR2x1_ASAP7_75t_L g2962 ( 
.A(n_2819),
.B(n_220),
.Y(n_2962)
);

CKINVDCx5p33_ASAP7_75t_R g2963 ( 
.A(n_2768),
.Y(n_2963)
);

NAND2xp5_ASAP7_75t_L g2964 ( 
.A(n_2790),
.B(n_221),
.Y(n_2964)
);

NOR2x1_ASAP7_75t_L g2965 ( 
.A(n_2819),
.B(n_223),
.Y(n_2965)
);

OR2x2_ASAP7_75t_L g2966 ( 
.A(n_2783),
.B(n_224),
.Y(n_2966)
);

NAND2xp33_ASAP7_75t_SL g2967 ( 
.A(n_2809),
.B(n_224),
.Y(n_2967)
);

NAND2xp5_ASAP7_75t_L g2968 ( 
.A(n_2790),
.B(n_225),
.Y(n_2968)
);

NAND2xp5_ASAP7_75t_L g2969 ( 
.A(n_2790),
.B(n_225),
.Y(n_2969)
);

AO221x2_ASAP7_75t_L g2970 ( 
.A1(n_2815),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.C(n_229),
.Y(n_2970)
);

OAI221xp5_ASAP7_75t_L g2971 ( 
.A1(n_2809),
.A2(n_228),
.B1(n_226),
.B2(n_227),
.C(n_229),
.Y(n_2971)
);

INVx4_ASAP7_75t_L g2972 ( 
.A(n_2768),
.Y(n_2972)
);

A2O1A1Ixp33_ASAP7_75t_L g2973 ( 
.A1(n_2753),
.A2(n_239),
.B(n_247),
.C(n_231),
.Y(n_2973)
);

NAND2xp5_ASAP7_75t_L g2974 ( 
.A(n_2790),
.B(n_231),
.Y(n_2974)
);

NAND2xp5_ASAP7_75t_L g2975 ( 
.A(n_2790),
.B(n_232),
.Y(n_2975)
);

INVx1_ASAP7_75t_L g2976 ( 
.A(n_2737),
.Y(n_2976)
);

NAND2xp5_ASAP7_75t_L g2977 ( 
.A(n_2790),
.B(n_233),
.Y(n_2977)
);

AOI22xp5_ASAP7_75t_L g2978 ( 
.A1(n_2809),
.A2(n_237),
.B1(n_235),
.B2(n_236),
.Y(n_2978)
);

NOR2xp33_ASAP7_75t_L g2979 ( 
.A(n_2809),
.B(n_235),
.Y(n_2979)
);

NAND2xp5_ASAP7_75t_L g2980 ( 
.A(n_2790),
.B(n_238),
.Y(n_2980)
);

NAND2xp5_ASAP7_75t_L g2981 ( 
.A(n_2790),
.B(n_238),
.Y(n_2981)
);

OAI22xp33_ASAP7_75t_L g2982 ( 
.A1(n_2809),
.A2(n_241),
.B1(n_239),
.B2(n_240),
.Y(n_2982)
);

AO221x1_ASAP7_75t_L g2983 ( 
.A1(n_2806),
.A2(n_243),
.B1(n_240),
.B2(n_242),
.C(n_244),
.Y(n_2983)
);

AND2x4_ASAP7_75t_L g2984 ( 
.A(n_2807),
.B(n_242),
.Y(n_2984)
);

CKINVDCx5p33_ASAP7_75t_R g2985 ( 
.A(n_2768),
.Y(n_2985)
);

OAI22xp33_ASAP7_75t_L g2986 ( 
.A1(n_2809),
.A2(n_245),
.B1(n_243),
.B2(n_244),
.Y(n_2986)
);

NAND2xp5_ASAP7_75t_L g2987 ( 
.A(n_2790),
.B(n_245),
.Y(n_2987)
);

AOI22xp5_ASAP7_75t_L g2988 ( 
.A1(n_2809),
.A2(n_248),
.B1(n_246),
.B2(n_247),
.Y(n_2988)
);

AOI22xp5_ASAP7_75t_L g2989 ( 
.A1(n_2809),
.A2(n_251),
.B1(n_246),
.B2(n_248),
.Y(n_2989)
);

AO221x2_ASAP7_75t_L g2990 ( 
.A1(n_2815),
.A2(n_254),
.B1(n_251),
.B2(n_253),
.C(n_255),
.Y(n_2990)
);

OR2x2_ASAP7_75t_L g2991 ( 
.A(n_2783),
.B(n_253),
.Y(n_2991)
);

NAND2xp5_ASAP7_75t_L g2992 ( 
.A(n_2790),
.B(n_254),
.Y(n_2992)
);

NAND2xp33_ASAP7_75t_R g2993 ( 
.A(n_2787),
.B(n_255),
.Y(n_2993)
);

NOR2x1_ASAP7_75t_L g2994 ( 
.A(n_2819),
.B(n_256),
.Y(n_2994)
);

INVx3_ASAP7_75t_SL g2995 ( 
.A(n_2852),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2850),
.Y(n_2996)
);

AND2x2_ASAP7_75t_L g2997 ( 
.A(n_2910),
.B(n_257),
.Y(n_2997)
);

AOI22xp33_ASAP7_75t_L g2998 ( 
.A1(n_2874),
.A2(n_261),
.B1(n_258),
.B2(n_259),
.Y(n_2998)
);

INVx1_ASAP7_75t_SL g2999 ( 
.A(n_2963),
.Y(n_2999)
);

NAND2xp33_ASAP7_75t_L g3000 ( 
.A(n_2880),
.B(n_258),
.Y(n_3000)
);

AND2x4_ASAP7_75t_L g3001 ( 
.A(n_2960),
.B(n_261),
.Y(n_3001)
);

AO21x2_ASAP7_75t_L g3002 ( 
.A1(n_2983),
.A2(n_262),
.B(n_263),
.Y(n_3002)
);

INVx1_ASAP7_75t_L g3003 ( 
.A(n_2854),
.Y(n_3003)
);

NAND2xp5_ASAP7_75t_L g3004 ( 
.A(n_2883),
.B(n_264),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2864),
.Y(n_3005)
);

NAND2xp5_ASAP7_75t_L g3006 ( 
.A(n_2947),
.B(n_2889),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2866),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2863),
.B(n_264),
.Y(n_3008)
);

INVx2_ASAP7_75t_L g3009 ( 
.A(n_2872),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2862),
.B(n_265),
.Y(n_3010)
);

INVx2_ASAP7_75t_L g3011 ( 
.A(n_2865),
.Y(n_3011)
);

INVxp67_ASAP7_75t_L g3012 ( 
.A(n_2993),
.Y(n_3012)
);

INVx1_ASAP7_75t_SL g3013 ( 
.A(n_2985),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2895),
.Y(n_3014)
);

BUFx3_ASAP7_75t_L g3015 ( 
.A(n_2870),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2976),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2882),
.B(n_265),
.Y(n_3017)
);

INVx1_ASAP7_75t_L g3018 ( 
.A(n_2912),
.Y(n_3018)
);

OR2x2_ASAP7_75t_L g3019 ( 
.A(n_2885),
.B(n_266),
.Y(n_3019)
);

CKINVDCx16_ASAP7_75t_R g3020 ( 
.A(n_2911),
.Y(n_3020)
);

OR2x2_ASAP7_75t_L g3021 ( 
.A(n_2953),
.B(n_266),
.Y(n_3021)
);

INVx1_ASAP7_75t_SL g3022 ( 
.A(n_2861),
.Y(n_3022)
);

NAND2xp5_ASAP7_75t_L g3023 ( 
.A(n_2922),
.B(n_267),
.Y(n_3023)
);

BUFx3_ASAP7_75t_L g3024 ( 
.A(n_2875),
.Y(n_3024)
);

INVx1_ASAP7_75t_SL g3025 ( 
.A(n_2952),
.Y(n_3025)
);

INVx1_ASAP7_75t_L g3026 ( 
.A(n_2898),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2903),
.Y(n_3027)
);

INVx2_ASAP7_75t_L g3028 ( 
.A(n_2926),
.Y(n_3028)
);

AOI22xp5_ASAP7_75t_L g3029 ( 
.A1(n_2874),
.A2(n_269),
.B1(n_267),
.B2(n_268),
.Y(n_3029)
);

OR2x2_ASAP7_75t_L g3030 ( 
.A(n_2966),
.B(n_2991),
.Y(n_3030)
);

OAI22xp5_ASAP7_75t_L g3031 ( 
.A1(n_2917),
.A2(n_272),
.B1(n_268),
.B2(n_270),
.Y(n_3031)
);

OR2x2_ASAP7_75t_L g3032 ( 
.A(n_2896),
.B(n_272),
.Y(n_3032)
);

INVx1_ASAP7_75t_SL g3033 ( 
.A(n_2929),
.Y(n_3033)
);

INVx2_ASAP7_75t_SL g3034 ( 
.A(n_2856),
.Y(n_3034)
);

INVx1_ASAP7_75t_SL g3035 ( 
.A(n_2879),
.Y(n_3035)
);

NOR2xp33_ASAP7_75t_L g3036 ( 
.A(n_2979),
.B(n_2858),
.Y(n_3036)
);

NOR2xp33_ASAP7_75t_L g3037 ( 
.A(n_2964),
.B(n_273),
.Y(n_3037)
);

INVx1_ASAP7_75t_L g3038 ( 
.A(n_2930),
.Y(n_3038)
);

NOR2xp33_ASAP7_75t_L g3039 ( 
.A(n_2968),
.B(n_273),
.Y(n_3039)
);

NAND2xp5_ASAP7_75t_L g3040 ( 
.A(n_2938),
.B(n_274),
.Y(n_3040)
);

AOI22xp33_ASAP7_75t_L g3041 ( 
.A1(n_2859),
.A2(n_276),
.B1(n_274),
.B2(n_275),
.Y(n_3041)
);

INVx1_ASAP7_75t_L g3042 ( 
.A(n_2925),
.Y(n_3042)
);

INVx1_ASAP7_75t_L g3043 ( 
.A(n_2931),
.Y(n_3043)
);

INVx2_ASAP7_75t_L g3044 ( 
.A(n_2897),
.Y(n_3044)
);

AOI22xp33_ASAP7_75t_L g3045 ( 
.A1(n_2970),
.A2(n_277),
.B1(n_275),
.B2(n_276),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2884),
.Y(n_3046)
);

AND2x2_ASAP7_75t_L g3047 ( 
.A(n_2921),
.B(n_278),
.Y(n_3047)
);

INVx2_ASAP7_75t_L g3048 ( 
.A(n_2924),
.Y(n_3048)
);

INVx1_ASAP7_75t_SL g3049 ( 
.A(n_2876),
.Y(n_3049)
);

INVx1_ASAP7_75t_L g3050 ( 
.A(n_2887),
.Y(n_3050)
);

INVx3_ASAP7_75t_L g3051 ( 
.A(n_2984),
.Y(n_3051)
);

OR2x2_ASAP7_75t_L g3052 ( 
.A(n_2891),
.B(n_278),
.Y(n_3052)
);

INVx2_ASAP7_75t_L g3053 ( 
.A(n_2853),
.Y(n_3053)
);

INVx1_ASAP7_75t_L g3054 ( 
.A(n_2902),
.Y(n_3054)
);

OR2x2_ASAP7_75t_L g3055 ( 
.A(n_2904),
.B(n_2906),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2915),
.Y(n_3056)
);

OR2x2_ASAP7_75t_L g3057 ( 
.A(n_2918),
.B(n_2969),
.Y(n_3057)
);

INVx2_ASAP7_75t_L g3058 ( 
.A(n_2962),
.Y(n_3058)
);

INVxp67_ASAP7_75t_SL g3059 ( 
.A(n_2959),
.Y(n_3059)
);

INVx1_ASAP7_75t_L g3060 ( 
.A(n_2974),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2975),
.Y(n_3061)
);

INVx2_ASAP7_75t_SL g3062 ( 
.A(n_2877),
.Y(n_3062)
);

INVx1_ASAP7_75t_L g3063 ( 
.A(n_2977),
.Y(n_3063)
);

AND2x2_ASAP7_75t_L g3064 ( 
.A(n_2957),
.B(n_2888),
.Y(n_3064)
);

INVx2_ASAP7_75t_L g3065 ( 
.A(n_2965),
.Y(n_3065)
);

OAI21xp5_ASAP7_75t_SL g3066 ( 
.A1(n_2914),
.A2(n_279),
.B(n_280),
.Y(n_3066)
);

INVx1_ASAP7_75t_L g3067 ( 
.A(n_2980),
.Y(n_3067)
);

NAND2xp5_ASAP7_75t_L g3068 ( 
.A(n_2981),
.B(n_279),
.Y(n_3068)
);

INVx1_ASAP7_75t_L g3069 ( 
.A(n_2987),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2992),
.Y(n_3070)
);

INVx1_ASAP7_75t_SL g3071 ( 
.A(n_2932),
.Y(n_3071)
);

INVx1_ASAP7_75t_L g3072 ( 
.A(n_2892),
.Y(n_3072)
);

INVx2_ASAP7_75t_L g3073 ( 
.A(n_2994),
.Y(n_3073)
);

AND2x2_ASAP7_75t_SL g3074 ( 
.A(n_2890),
.B(n_280),
.Y(n_3074)
);

AND2x2_ASAP7_75t_L g3075 ( 
.A(n_2927),
.B(n_281),
.Y(n_3075)
);

INVx1_ASAP7_75t_L g3076 ( 
.A(n_2873),
.Y(n_3076)
);

AND2x2_ASAP7_75t_L g3077 ( 
.A(n_2920),
.B(n_282),
.Y(n_3077)
);

NAND2xp5_ASAP7_75t_L g3078 ( 
.A(n_2923),
.B(n_2909),
.Y(n_3078)
);

INVx1_ASAP7_75t_SL g3079 ( 
.A(n_2956),
.Y(n_3079)
);

AOI222xp33_ASAP7_75t_L g3080 ( 
.A1(n_2907),
.A2(n_284),
.B1(n_286),
.B2(n_282),
.C1(n_283),
.C2(n_285),
.Y(n_3080)
);

NAND2xp5_ASAP7_75t_L g3081 ( 
.A(n_2886),
.B(n_283),
.Y(n_3081)
);

CKINVDCx16_ASAP7_75t_R g3082 ( 
.A(n_2967),
.Y(n_3082)
);

OR2x2_ASAP7_75t_L g3083 ( 
.A(n_2943),
.B(n_284),
.Y(n_3083)
);

NAND2xp5_ASAP7_75t_L g3084 ( 
.A(n_2886),
.B(n_286),
.Y(n_3084)
);

INVxp33_ASAP7_75t_L g3085 ( 
.A(n_2868),
.Y(n_3085)
);

INVxp67_ASAP7_75t_L g3086 ( 
.A(n_2936),
.Y(n_3086)
);

AND2x4_ASAP7_75t_L g3087 ( 
.A(n_2933),
.B(n_288),
.Y(n_3087)
);

CKINVDCx16_ASAP7_75t_R g3088 ( 
.A(n_2899),
.Y(n_3088)
);

AND2x2_ASAP7_75t_L g3089 ( 
.A(n_2942),
.B(n_287),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_2939),
.B(n_288),
.Y(n_3090)
);

INVx2_ASAP7_75t_L g3091 ( 
.A(n_2881),
.Y(n_3091)
);

OAI21x1_ASAP7_75t_L g3092 ( 
.A1(n_2940),
.A2(n_289),
.B(n_290),
.Y(n_3092)
);

INVx2_ASAP7_75t_SL g3093 ( 
.A(n_2970),
.Y(n_3093)
);

INVx2_ASAP7_75t_SL g3094 ( 
.A(n_2990),
.Y(n_3094)
);

NAND2xp5_ASAP7_75t_L g3095 ( 
.A(n_2900),
.B(n_289),
.Y(n_3095)
);

INVxp67_ASAP7_75t_SL g3096 ( 
.A(n_2944),
.Y(n_3096)
);

HB1xp67_ASAP7_75t_L g3097 ( 
.A(n_2900),
.Y(n_3097)
);

INVx1_ASAP7_75t_L g3098 ( 
.A(n_2950),
.Y(n_3098)
);

INVx4_ASAP7_75t_L g3099 ( 
.A(n_2990),
.Y(n_3099)
);

NAND2xp5_ASAP7_75t_L g3100 ( 
.A(n_2901),
.B(n_290),
.Y(n_3100)
);

INVx1_ASAP7_75t_L g3101 ( 
.A(n_2954),
.Y(n_3101)
);

INVx1_ASAP7_75t_SL g3102 ( 
.A(n_2867),
.Y(n_3102)
);

NOR2xp33_ASAP7_75t_L g3103 ( 
.A(n_2958),
.B(n_291),
.Y(n_3103)
);

AND2x2_ASAP7_75t_L g3104 ( 
.A(n_2945),
.B(n_2946),
.Y(n_3104)
);

HB1xp67_ASAP7_75t_L g3105 ( 
.A(n_2901),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2941),
.B(n_291),
.Y(n_3106)
);

INVx4_ASAP7_75t_L g3107 ( 
.A(n_2913),
.Y(n_3107)
);

AND2x2_ASAP7_75t_L g3108 ( 
.A(n_2945),
.B(n_292),
.Y(n_3108)
);

NAND2xp5_ASAP7_75t_L g3109 ( 
.A(n_2913),
.B(n_293),
.Y(n_3109)
);

AND2x2_ASAP7_75t_L g3110 ( 
.A(n_2946),
.B(n_2935),
.Y(n_3110)
);

INVx1_ASAP7_75t_L g3111 ( 
.A(n_2855),
.Y(n_3111)
);

CKINVDCx16_ASAP7_75t_R g3112 ( 
.A(n_2978),
.Y(n_3112)
);

INVx1_ASAP7_75t_SL g3113 ( 
.A(n_2988),
.Y(n_3113)
);

INVxp67_ASAP7_75t_L g3114 ( 
.A(n_2928),
.Y(n_3114)
);

NOR2x1_ASAP7_75t_L g3115 ( 
.A(n_2908),
.B(n_294),
.Y(n_3115)
);

INVx1_ASAP7_75t_SL g3116 ( 
.A(n_2989),
.Y(n_3116)
);

AND2x2_ASAP7_75t_L g3117 ( 
.A(n_2951),
.B(n_294),
.Y(n_3117)
);

BUFx2_ASAP7_75t_L g3118 ( 
.A(n_2949),
.Y(n_3118)
);

INVxp67_ASAP7_75t_L g3119 ( 
.A(n_2971),
.Y(n_3119)
);

AND2x4_ASAP7_75t_L g3120 ( 
.A(n_2973),
.B(n_295),
.Y(n_3120)
);

NOR2xp33_ASAP7_75t_L g3121 ( 
.A(n_2893),
.B(n_295),
.Y(n_3121)
);

OR2x2_ASAP7_75t_L g3122 ( 
.A(n_2894),
.B(n_296),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2934),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2869),
.B(n_296),
.Y(n_3124)
);

AOI22x1_ASAP7_75t_L g3125 ( 
.A1(n_2851),
.A2(n_299),
.B1(n_297),
.B2(n_298),
.Y(n_3125)
);

INVx1_ASAP7_75t_L g3126 ( 
.A(n_2937),
.Y(n_3126)
);

INVx2_ASAP7_75t_L g3127 ( 
.A(n_2871),
.Y(n_3127)
);

HB1xp67_ASAP7_75t_L g3128 ( 
.A(n_2916),
.Y(n_3128)
);

INVx2_ASAP7_75t_L g3129 ( 
.A(n_2857),
.Y(n_3129)
);

AND2x2_ASAP7_75t_L g3130 ( 
.A(n_2955),
.B(n_298),
.Y(n_3130)
);

AND2x2_ASAP7_75t_L g3131 ( 
.A(n_2919),
.B(n_300),
.Y(n_3131)
);

AOI22xp33_ASAP7_75t_SL g3132 ( 
.A1(n_2878),
.A2(n_303),
.B1(n_301),
.B2(n_302),
.Y(n_3132)
);

INVx2_ASAP7_75t_L g3133 ( 
.A(n_2948),
.Y(n_3133)
);

CKINVDCx16_ASAP7_75t_R g3134 ( 
.A(n_2961),
.Y(n_3134)
);

INVx1_ASAP7_75t_L g3135 ( 
.A(n_2860),
.Y(n_3135)
);

BUFx2_ASAP7_75t_L g3136 ( 
.A(n_2982),
.Y(n_3136)
);

NAND2xp5_ASAP7_75t_L g3137 ( 
.A(n_2986),
.B(n_301),
.Y(n_3137)
);

BUFx2_ASAP7_75t_L g3138 ( 
.A(n_2905),
.Y(n_3138)
);

OR2x2_ASAP7_75t_L g3139 ( 
.A(n_2885),
.B(n_302),
.Y(n_3139)
);

BUFx3_ASAP7_75t_L g3140 ( 
.A(n_2960),
.Y(n_3140)
);

INVx1_ASAP7_75t_L g3141 ( 
.A(n_2850),
.Y(n_3141)
);

AND2x2_ASAP7_75t_L g3142 ( 
.A(n_2910),
.B(n_303),
.Y(n_3142)
);

INVx1_ASAP7_75t_L g3143 ( 
.A(n_2850),
.Y(n_3143)
);

INVx1_ASAP7_75t_SL g3144 ( 
.A(n_2852),
.Y(n_3144)
);

INVx1_ASAP7_75t_L g3145 ( 
.A(n_2850),
.Y(n_3145)
);

CKINVDCx16_ASAP7_75t_R g3146 ( 
.A(n_2993),
.Y(n_3146)
);

OR2x2_ASAP7_75t_L g3147 ( 
.A(n_2885),
.B(n_304),
.Y(n_3147)
);

AND2x2_ASAP7_75t_L g3148 ( 
.A(n_2910),
.B(n_305),
.Y(n_3148)
);

AND2x4_ASAP7_75t_L g3149 ( 
.A(n_2960),
.B(n_306),
.Y(n_3149)
);

INVx1_ASAP7_75t_L g3150 ( 
.A(n_2850),
.Y(n_3150)
);

INVx1_ASAP7_75t_L g3151 ( 
.A(n_2850),
.Y(n_3151)
);

OAI221xp5_ASAP7_75t_L g3152 ( 
.A1(n_2967),
.A2(n_307),
.B1(n_305),
.B2(n_306),
.C(n_308),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2910),
.B(n_307),
.Y(n_3153)
);

INVx1_ASAP7_75t_L g3154 ( 
.A(n_2850),
.Y(n_3154)
);

OR2x2_ASAP7_75t_L g3155 ( 
.A(n_2885),
.B(n_308),
.Y(n_3155)
);

INVx1_ASAP7_75t_L g3156 ( 
.A(n_2850),
.Y(n_3156)
);

NOR3xp33_ASAP7_75t_L g3157 ( 
.A(n_2928),
.B(n_309),
.C(n_310),
.Y(n_3157)
);

INVx1_ASAP7_75t_SL g3158 ( 
.A(n_2852),
.Y(n_3158)
);

AND2x2_ASAP7_75t_L g3159 ( 
.A(n_2910),
.B(n_311),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_2850),
.Y(n_3160)
);

INVx2_ASAP7_75t_L g3161 ( 
.A(n_2910),
.Y(n_3161)
);

NAND2xp5_ASAP7_75t_L g3162 ( 
.A(n_2883),
.B(n_312),
.Y(n_3162)
);

AO21x2_ASAP7_75t_L g3163 ( 
.A1(n_2983),
.A2(n_312),
.B(n_314),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_2910),
.B(n_314),
.Y(n_3164)
);

OR2x2_ASAP7_75t_L g3165 ( 
.A(n_2885),
.B(n_315),
.Y(n_3165)
);

INVx1_ASAP7_75t_L g3166 ( 
.A(n_2850),
.Y(n_3166)
);

INVx1_ASAP7_75t_L g3167 ( 
.A(n_2850),
.Y(n_3167)
);

INVx1_ASAP7_75t_L g3168 ( 
.A(n_2850),
.Y(n_3168)
);

NAND2xp5_ASAP7_75t_L g3169 ( 
.A(n_2883),
.B(n_315),
.Y(n_3169)
);

NOR2x1_ASAP7_75t_L g3170 ( 
.A(n_2972),
.B(n_316),
.Y(n_3170)
);

INVx2_ASAP7_75t_SL g3171 ( 
.A(n_2852),
.Y(n_3171)
);

INVx3_ASAP7_75t_SL g3172 ( 
.A(n_2852),
.Y(n_3172)
);

INVx1_ASAP7_75t_L g3173 ( 
.A(n_2850),
.Y(n_3173)
);

INVx2_ASAP7_75t_L g3174 ( 
.A(n_2910),
.Y(n_3174)
);

INVx1_ASAP7_75t_L g3175 ( 
.A(n_2850),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_2850),
.Y(n_3176)
);

NAND2xp5_ASAP7_75t_L g3177 ( 
.A(n_2883),
.B(n_316),
.Y(n_3177)
);

AND2x2_ASAP7_75t_L g3178 ( 
.A(n_2910),
.B(n_317),
.Y(n_3178)
);

INVx2_ASAP7_75t_L g3179 ( 
.A(n_2910),
.Y(n_3179)
);

AND2x2_ASAP7_75t_L g3180 ( 
.A(n_2910),
.B(n_317),
.Y(n_3180)
);

INVx1_ASAP7_75t_L g3181 ( 
.A(n_2850),
.Y(n_3181)
);

CKINVDCx16_ASAP7_75t_R g3182 ( 
.A(n_2993),
.Y(n_3182)
);

HB1xp67_ASAP7_75t_L g3183 ( 
.A(n_2872),
.Y(n_3183)
);

OR2x2_ASAP7_75t_L g3184 ( 
.A(n_2885),
.B(n_318),
.Y(n_3184)
);

INVx1_ASAP7_75t_L g3185 ( 
.A(n_2850),
.Y(n_3185)
);

AO21x2_ASAP7_75t_L g3186 ( 
.A1(n_2983),
.A2(n_318),
.B(n_319),
.Y(n_3186)
);

NAND2xp5_ASAP7_75t_L g3187 ( 
.A(n_2883),
.B(n_319),
.Y(n_3187)
);

INVx1_ASAP7_75t_L g3188 ( 
.A(n_2850),
.Y(n_3188)
);

AOI21xp5_ASAP7_75t_L g3189 ( 
.A1(n_2859),
.A2(n_320),
.B(n_321),
.Y(n_3189)
);

OR2x2_ASAP7_75t_L g3190 ( 
.A(n_2885),
.B(n_321),
.Y(n_3190)
);

INVx1_ASAP7_75t_L g3191 ( 
.A(n_2850),
.Y(n_3191)
);

INVx2_ASAP7_75t_L g3192 ( 
.A(n_2910),
.Y(n_3192)
);

AND2x2_ASAP7_75t_L g3193 ( 
.A(n_2910),
.B(n_322),
.Y(n_3193)
);

NAND2xp5_ASAP7_75t_L g3194 ( 
.A(n_2883),
.B(n_322),
.Y(n_3194)
);

INVxp67_ASAP7_75t_SL g3195 ( 
.A(n_2872),
.Y(n_3195)
);

INVx1_ASAP7_75t_L g3196 ( 
.A(n_2996),
.Y(n_3196)
);

INVx1_ASAP7_75t_L g3197 ( 
.A(n_3003),
.Y(n_3197)
);

INVx1_ASAP7_75t_L g3198 ( 
.A(n_3005),
.Y(n_3198)
);

NAND2xp5_ASAP7_75t_L g3199 ( 
.A(n_3053),
.B(n_324),
.Y(n_3199)
);

AND2x2_ASAP7_75t_L g3200 ( 
.A(n_3140),
.B(n_324),
.Y(n_3200)
);

AOI222xp33_ASAP7_75t_L g3201 ( 
.A1(n_3114),
.A2(n_327),
.B1(n_329),
.B2(n_325),
.C1(n_326),
.C2(n_328),
.Y(n_3201)
);

INVxp67_ASAP7_75t_SL g3202 ( 
.A(n_3012),
.Y(n_3202)
);

O2A1O1Ixp5_ASAP7_75t_SL g3203 ( 
.A1(n_3119),
.A2(n_3128),
.B(n_3031),
.C(n_3105),
.Y(n_3203)
);

NAND2xp5_ASAP7_75t_L g3204 ( 
.A(n_3058),
.B(n_325),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3007),
.Y(n_3205)
);

AOI22xp5_ASAP7_75t_L g3206 ( 
.A1(n_3134),
.A2(n_329),
.B1(n_326),
.B2(n_328),
.Y(n_3206)
);

INVxp67_ASAP7_75t_SL g3207 ( 
.A(n_3059),
.Y(n_3207)
);

INVx1_ASAP7_75t_L g3208 ( 
.A(n_3014),
.Y(n_3208)
);

NAND2xp5_ASAP7_75t_L g3209 ( 
.A(n_3065),
.B(n_330),
.Y(n_3209)
);

AOI21xp5_ASAP7_75t_L g3210 ( 
.A1(n_3000),
.A2(n_330),
.B(n_331),
.Y(n_3210)
);

AOI21xp5_ASAP7_75t_L g3211 ( 
.A1(n_3146),
.A2(n_332),
.B(n_333),
.Y(n_3211)
);

NAND2xp5_ASAP7_75t_SL g3212 ( 
.A(n_3020),
.B(n_333),
.Y(n_3212)
);

OAI22xp5_ASAP7_75t_L g3213 ( 
.A1(n_3182),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3213)
);

OAI22xp5_ASAP7_75t_L g3214 ( 
.A1(n_3107),
.A2(n_336),
.B1(n_334),
.B2(n_335),
.Y(n_3214)
);

INVx3_ASAP7_75t_L g3215 ( 
.A(n_3015),
.Y(n_3215)
);

INVx2_ASAP7_75t_L g3216 ( 
.A(n_3034),
.Y(n_3216)
);

AOI221xp5_ASAP7_75t_L g3217 ( 
.A1(n_3099),
.A2(n_339),
.B1(n_337),
.B2(n_338),
.C(n_340),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3006),
.B(n_339),
.Y(n_3218)
);

OAI22xp5_ASAP7_75t_L g3219 ( 
.A1(n_3097),
.A2(n_342),
.B1(n_340),
.B2(n_341),
.Y(n_3219)
);

AND2x2_ASAP7_75t_L g3220 ( 
.A(n_3096),
.B(n_341),
.Y(n_3220)
);

OAI22xp33_ASAP7_75t_L g3221 ( 
.A1(n_3082),
.A2(n_344),
.B1(n_342),
.B2(n_343),
.Y(n_3221)
);

INVx1_ASAP7_75t_L g3222 ( 
.A(n_3016),
.Y(n_3222)
);

INVxp67_ASAP7_75t_L g3223 ( 
.A(n_3033),
.Y(n_3223)
);

AOI21xp5_ASAP7_75t_L g3224 ( 
.A1(n_3066),
.A2(n_343),
.B(n_344),
.Y(n_3224)
);

INVx1_ASAP7_75t_L g3225 ( 
.A(n_3141),
.Y(n_3225)
);

NAND2xp5_ASAP7_75t_L g3226 ( 
.A(n_3073),
.B(n_3093),
.Y(n_3226)
);

NAND2xp33_ASAP7_75t_L g3227 ( 
.A(n_3157),
.B(n_345),
.Y(n_3227)
);

OAI21xp5_ASAP7_75t_L g3228 ( 
.A1(n_3115),
.A2(n_345),
.B(n_346),
.Y(n_3228)
);

AOI22x1_ASAP7_75t_L g3229 ( 
.A1(n_3112),
.A2(n_3088),
.B1(n_3136),
.B2(n_3138),
.Y(n_3229)
);

OR2x2_ASAP7_75t_L g3230 ( 
.A(n_3038),
.B(n_346),
.Y(n_3230)
);

NAND4xp25_ASAP7_75t_L g3231 ( 
.A(n_2998),
.B(n_349),
.C(n_350),
.D(n_348),
.Y(n_3231)
);

INVx1_ASAP7_75t_L g3232 ( 
.A(n_3143),
.Y(n_3232)
);

INVx2_ASAP7_75t_L g3233 ( 
.A(n_3161),
.Y(n_3233)
);

AND2x2_ASAP7_75t_L g3234 ( 
.A(n_3174),
.B(n_347),
.Y(n_3234)
);

INVx1_ASAP7_75t_SL g3235 ( 
.A(n_2995),
.Y(n_3235)
);

NAND2xp5_ASAP7_75t_L g3236 ( 
.A(n_3094),
.B(n_347),
.Y(n_3236)
);

NAND2x1_ASAP7_75t_L g3237 ( 
.A(n_3028),
.B(n_348),
.Y(n_3237)
);

NAND2xp5_ASAP7_75t_L g3238 ( 
.A(n_3110),
.B(n_349),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3145),
.Y(n_3239)
);

OA21x2_ASAP7_75t_L g3240 ( 
.A1(n_3118),
.A2(n_350),
.B(n_351),
.Y(n_3240)
);

AOI321xp33_ASAP7_75t_L g3241 ( 
.A1(n_3104),
.A2(n_354),
.A3(n_356),
.B1(n_352),
.B2(n_353),
.C(n_355),
.Y(n_3241)
);

NOR3xp33_ASAP7_75t_SL g3242 ( 
.A(n_3152),
.B(n_352),
.C(n_355),
.Y(n_3242)
);

OAI221xp5_ASAP7_75t_L g3243 ( 
.A1(n_3029),
.A2(n_358),
.B1(n_356),
.B2(n_357),
.C(n_359),
.Y(n_3243)
);

AOI21xp5_ASAP7_75t_L g3244 ( 
.A1(n_3189),
.A2(n_3074),
.B(n_3078),
.Y(n_3244)
);

AOI22xp5_ASAP7_75t_L g3245 ( 
.A1(n_3120),
.A2(n_359),
.B1(n_357),
.B2(n_358),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3150),
.Y(n_3246)
);

NAND2xp5_ASAP7_75t_L g3247 ( 
.A(n_3129),
.B(n_360),
.Y(n_3247)
);

INVx2_ASAP7_75t_SL g3248 ( 
.A(n_3172),
.Y(n_3248)
);

AOI22xp33_ASAP7_75t_SL g3249 ( 
.A1(n_3126),
.A2(n_362),
.B1(n_360),
.B2(n_361),
.Y(n_3249)
);

NAND2xp5_ASAP7_75t_L g3250 ( 
.A(n_3072),
.B(n_361),
.Y(n_3250)
);

NAND2xp5_ASAP7_75t_L g3251 ( 
.A(n_3113),
.B(n_362),
.Y(n_3251)
);

INVx2_ASAP7_75t_L g3252 ( 
.A(n_3179),
.Y(n_3252)
);

NAND4xp25_ASAP7_75t_SL g3253 ( 
.A(n_3080),
.B(n_365),
.C(n_363),
.D(n_364),
.Y(n_3253)
);

AOI21xp33_ASAP7_75t_L g3254 ( 
.A1(n_3002),
.A2(n_363),
.B(n_364),
.Y(n_3254)
);

AOI21xp5_ASAP7_75t_L g3255 ( 
.A1(n_3163),
.A2(n_366),
.B(n_367),
.Y(n_3255)
);

NAND2xp5_ASAP7_75t_SL g3256 ( 
.A(n_3022),
.B(n_368),
.Y(n_3256)
);

NAND2xp5_ASAP7_75t_L g3257 ( 
.A(n_3116),
.B(n_368),
.Y(n_3257)
);

NAND2xp5_ASAP7_75t_L g3258 ( 
.A(n_3098),
.B(n_369),
.Y(n_3258)
);

NOR2xp33_ASAP7_75t_L g3259 ( 
.A(n_3025),
.B(n_370),
.Y(n_3259)
);

AOI221xp5_ASAP7_75t_L g3260 ( 
.A1(n_3135),
.A2(n_372),
.B1(n_370),
.B2(n_371),
.C(n_373),
.Y(n_3260)
);

NAND2xp5_ASAP7_75t_L g3261 ( 
.A(n_3101),
.B(n_373),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3151),
.Y(n_3262)
);

OAI322xp33_ASAP7_75t_L g3263 ( 
.A1(n_3081),
.A2(n_380),
.A3(n_379),
.B1(n_376),
.B2(n_374),
.C1(n_375),
.C2(n_378),
.Y(n_3263)
);

OAI211xp5_ASAP7_75t_L g3264 ( 
.A1(n_3045),
.A2(n_376),
.B(n_374),
.C(n_375),
.Y(n_3264)
);

AOI32xp33_ASAP7_75t_L g3265 ( 
.A1(n_3108),
.A2(n_380),
.A3(n_378),
.B1(n_379),
.B2(n_381),
.Y(n_3265)
);

AOI222xp33_ASAP7_75t_L g3266 ( 
.A1(n_3130),
.A2(n_383),
.B1(n_386),
.B2(n_381),
.C1(n_382),
.C2(n_385),
.Y(n_3266)
);

NAND2xp5_ASAP7_75t_L g3267 ( 
.A(n_3127),
.B(n_385),
.Y(n_3267)
);

HB1xp67_ASAP7_75t_L g3268 ( 
.A(n_3183),
.Y(n_3268)
);

OAI22xp33_ASAP7_75t_L g3269 ( 
.A1(n_3049),
.A2(n_388),
.B1(n_386),
.B2(n_387),
.Y(n_3269)
);

OAI21xp5_ASAP7_75t_SL g3270 ( 
.A1(n_3041),
.A2(n_388),
.B(n_389),
.Y(n_3270)
);

NOR2xp33_ASAP7_75t_SL g3271 ( 
.A(n_3035),
.B(n_390),
.Y(n_3271)
);

AOI221xp5_ASAP7_75t_SL g3272 ( 
.A1(n_3084),
.A2(n_394),
.B1(n_390),
.B2(n_393),
.C(n_395),
.Y(n_3272)
);

NAND2xp5_ASAP7_75t_SL g3273 ( 
.A(n_3102),
.B(n_395),
.Y(n_3273)
);

NAND2xp5_ASAP7_75t_L g3274 ( 
.A(n_3060),
.B(n_396),
.Y(n_3274)
);

NAND2xp5_ASAP7_75t_L g3275 ( 
.A(n_3061),
.B(n_396),
.Y(n_3275)
);

INVx1_ASAP7_75t_L g3276 ( 
.A(n_3154),
.Y(n_3276)
);

NOR2xp33_ASAP7_75t_L g3277 ( 
.A(n_3071),
.B(n_397),
.Y(n_3277)
);

NAND2xp5_ASAP7_75t_L g3278 ( 
.A(n_3063),
.B(n_397),
.Y(n_3278)
);

INVx1_ASAP7_75t_L g3279 ( 
.A(n_3156),
.Y(n_3279)
);

NAND2xp5_ASAP7_75t_L g3280 ( 
.A(n_3067),
.B(n_3069),
.Y(n_3280)
);

AOI22xp5_ASAP7_75t_L g3281 ( 
.A1(n_3186),
.A2(n_400),
.B1(n_398),
.B2(n_399),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3160),
.Y(n_3282)
);

NOR2xp67_ASAP7_75t_L g3283 ( 
.A(n_3086),
.B(n_399),
.Y(n_3283)
);

OAI221xp5_ASAP7_75t_L g3284 ( 
.A1(n_3079),
.A2(n_402),
.B1(n_400),
.B2(n_401),
.C(n_403),
.Y(n_3284)
);

NAND2xp5_ASAP7_75t_L g3285 ( 
.A(n_3070),
.B(n_401),
.Y(n_3285)
);

INVx1_ASAP7_75t_SL g3286 ( 
.A(n_2999),
.Y(n_3286)
);

INVx2_ASAP7_75t_L g3287 ( 
.A(n_3192),
.Y(n_3287)
);

OAI32xp33_ASAP7_75t_L g3288 ( 
.A1(n_3095),
.A2(n_405),
.A3(n_402),
.B1(n_404),
.B2(n_406),
.Y(n_3288)
);

NAND2xp5_ASAP7_75t_L g3289 ( 
.A(n_3076),
.B(n_407),
.Y(n_3289)
);

INVx2_ASAP7_75t_L g3290 ( 
.A(n_3009),
.Y(n_3290)
);

NAND2xp5_ASAP7_75t_L g3291 ( 
.A(n_3054),
.B(n_407),
.Y(n_3291)
);

INVx1_ASAP7_75t_L g3292 ( 
.A(n_3166),
.Y(n_3292)
);

NAND3xp33_ASAP7_75t_L g3293 ( 
.A(n_3132),
.B(n_408),
.C(n_409),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_SL g3294 ( 
.A(n_3171),
.B(n_3013),
.Y(n_3294)
);

NOR2xp33_ASAP7_75t_R g3295 ( 
.A(n_3062),
.B(n_408),
.Y(n_3295)
);

OAI321xp33_ASAP7_75t_L g3296 ( 
.A1(n_3137),
.A2(n_3109),
.A3(n_3100),
.B1(n_3121),
.B2(n_3122),
.C(n_3123),
.Y(n_3296)
);

OAI21xp33_ASAP7_75t_SL g3297 ( 
.A1(n_3195),
.A2(n_409),
.B(n_410),
.Y(n_3297)
);

NAND3xp33_ASAP7_75t_SL g3298 ( 
.A(n_3133),
.B(n_411),
.C(n_412),
.Y(n_3298)
);

AOI22xp5_ASAP7_75t_L g3299 ( 
.A1(n_3111),
.A2(n_3106),
.B1(n_3124),
.B2(n_3117),
.Y(n_3299)
);

NAND2xp5_ASAP7_75t_L g3300 ( 
.A(n_3056),
.B(n_412),
.Y(n_3300)
);

AOI222xp33_ASAP7_75t_L g3301 ( 
.A1(n_3131),
.A2(n_415),
.B1(n_417),
.B2(n_413),
.C1(n_414),
.C2(n_416),
.Y(n_3301)
);

NAND2xp33_ASAP7_75t_L g3302 ( 
.A(n_3170),
.B(n_413),
.Y(n_3302)
);

AOI21xp33_ASAP7_75t_L g3303 ( 
.A1(n_3036),
.A2(n_415),
.B(n_416),
.Y(n_3303)
);

INVx1_ASAP7_75t_L g3304 ( 
.A(n_3167),
.Y(n_3304)
);

AND2x2_ASAP7_75t_L g3305 ( 
.A(n_3044),
.B(n_417),
.Y(n_3305)
);

INVx2_ASAP7_75t_L g3306 ( 
.A(n_3051),
.Y(n_3306)
);

NAND2xp5_ASAP7_75t_L g3307 ( 
.A(n_3046),
.B(n_3042),
.Y(n_3307)
);

NAND2xp5_ASAP7_75t_L g3308 ( 
.A(n_3043),
.B(n_418),
.Y(n_3308)
);

NAND2xp5_ASAP7_75t_L g3309 ( 
.A(n_3050),
.B(n_418),
.Y(n_3309)
);

INVxp67_ASAP7_75t_L g3310 ( 
.A(n_3149),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3168),
.Y(n_3311)
);

OAI21xp33_ASAP7_75t_L g3312 ( 
.A1(n_3018),
.A2(n_419),
.B(n_420),
.Y(n_3312)
);

OAI21xp5_ASAP7_75t_L g3313 ( 
.A1(n_3077),
.A2(n_419),
.B(n_420),
.Y(n_3313)
);

AOI22xp33_ASAP7_75t_L g3314 ( 
.A1(n_3125),
.A2(n_423),
.B1(n_421),
.B2(n_422),
.Y(n_3314)
);

NAND2xp5_ASAP7_75t_L g3315 ( 
.A(n_2997),
.B(n_421),
.Y(n_3315)
);

A2O1A1Ixp33_ASAP7_75t_L g3316 ( 
.A1(n_3087),
.A2(n_424),
.B(n_422),
.C(n_423),
.Y(n_3316)
);

OAI31xp33_ASAP7_75t_L g3317 ( 
.A1(n_3087),
.A2(n_426),
.A3(n_424),
.B(n_425),
.Y(n_3317)
);

INVxp67_ASAP7_75t_L g3318 ( 
.A(n_3149),
.Y(n_3318)
);

INVxp67_ASAP7_75t_L g3319 ( 
.A(n_3055),
.Y(n_3319)
);

INVx1_ASAP7_75t_L g3320 ( 
.A(n_3173),
.Y(n_3320)
);

O2A1O1Ixp33_ASAP7_75t_SL g3321 ( 
.A1(n_3004),
.A2(n_3169),
.B(n_3177),
.C(n_3162),
.Y(n_3321)
);

AOI21xp33_ASAP7_75t_L g3322 ( 
.A1(n_3085),
.A2(n_426),
.B(n_427),
.Y(n_3322)
);

AND2x2_ASAP7_75t_L g3323 ( 
.A(n_3011),
.B(n_428),
.Y(n_3323)
);

INVx2_ASAP7_75t_L g3324 ( 
.A(n_3048),
.Y(n_3324)
);

OAI21xp33_ASAP7_75t_SL g3325 ( 
.A1(n_3026),
.A2(n_428),
.B(n_429),
.Y(n_3325)
);

OAI21xp5_ASAP7_75t_SL g3326 ( 
.A1(n_3037),
.A2(n_429),
.B(n_430),
.Y(n_3326)
);

INVxp67_ASAP7_75t_L g3327 ( 
.A(n_3057),
.Y(n_3327)
);

INVx3_ASAP7_75t_L g3328 ( 
.A(n_3024),
.Y(n_3328)
);

NAND2xp33_ASAP7_75t_SL g3329 ( 
.A(n_3142),
.B(n_430),
.Y(n_3329)
);

INVxp33_ASAP7_75t_L g3330 ( 
.A(n_3064),
.Y(n_3330)
);

AOI22xp5_ASAP7_75t_L g3331 ( 
.A1(n_3027),
.A2(n_433),
.B1(n_431),
.B2(n_432),
.Y(n_3331)
);

OAI22xp5_ASAP7_75t_L g3332 ( 
.A1(n_3030),
.A2(n_436),
.B1(n_434),
.B2(n_435),
.Y(n_3332)
);

INVx1_ASAP7_75t_L g3333 ( 
.A(n_3175),
.Y(n_3333)
);

OAI22xp33_ASAP7_75t_SL g3334 ( 
.A1(n_3187),
.A2(n_437),
.B1(n_434),
.B2(n_436),
.Y(n_3334)
);

AOI322xp5_ASAP7_75t_L g3335 ( 
.A1(n_3039),
.A2(n_443),
.A3(n_442),
.B1(n_440),
.B2(n_438),
.C1(n_439),
.C2(n_441),
.Y(n_3335)
);

INVx1_ASAP7_75t_L g3336 ( 
.A(n_3176),
.Y(n_3336)
);

INVx1_ASAP7_75t_SL g3337 ( 
.A(n_3144),
.Y(n_3337)
);

OR2x2_ASAP7_75t_L g3338 ( 
.A(n_3019),
.B(n_3139),
.Y(n_3338)
);

AOI22xp5_ASAP7_75t_L g3339 ( 
.A1(n_3103),
.A2(n_443),
.B1(n_438),
.B2(n_442),
.Y(n_3339)
);

NAND2xp5_ASAP7_75t_L g3340 ( 
.A(n_3148),
.B(n_444),
.Y(n_3340)
);

AOI21xp5_ASAP7_75t_L g3341 ( 
.A1(n_3194),
.A2(n_444),
.B(n_445),
.Y(n_3341)
);

INVx1_ASAP7_75t_SL g3342 ( 
.A(n_3295),
.Y(n_3342)
);

INVx1_ASAP7_75t_L g3343 ( 
.A(n_3268),
.Y(n_3343)
);

INVxp67_ASAP7_75t_L g3344 ( 
.A(n_3207),
.Y(n_3344)
);

OR2x2_ASAP7_75t_L g3345 ( 
.A(n_3223),
.B(n_3147),
.Y(n_3345)
);

AND2x2_ASAP7_75t_L g3346 ( 
.A(n_3215),
.B(n_3158),
.Y(n_3346)
);

INVx1_ASAP7_75t_L g3347 ( 
.A(n_3202),
.Y(n_3347)
);

INVx1_ASAP7_75t_L g3348 ( 
.A(n_3196),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_L g3349 ( 
.A(n_3203),
.B(n_3153),
.Y(n_3349)
);

INVx3_ASAP7_75t_L g3350 ( 
.A(n_3215),
.Y(n_3350)
);

AND2x2_ASAP7_75t_L g3351 ( 
.A(n_3328),
.B(n_3091),
.Y(n_3351)
);

INVxp67_ASAP7_75t_L g3352 ( 
.A(n_3271),
.Y(n_3352)
);

NOR2xp33_ASAP7_75t_L g3353 ( 
.A(n_3235),
.B(n_3155),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3310),
.B(n_3318),
.Y(n_3354)
);

INVx1_ASAP7_75t_L g3355 ( 
.A(n_3197),
.Y(n_3355)
);

AND2x2_ASAP7_75t_L g3356 ( 
.A(n_3328),
.B(n_3001),
.Y(n_3356)
);

NOR3xp33_ASAP7_75t_L g3357 ( 
.A(n_3296),
.B(n_3010),
.C(n_3023),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3198),
.Y(n_3358)
);

AOI22xp33_ASAP7_75t_L g3359 ( 
.A1(n_3229),
.A2(n_3165),
.B1(n_3190),
.B2(n_3184),
.Y(n_3359)
);

NAND2xp5_ASAP7_75t_L g3360 ( 
.A(n_3255),
.B(n_3159),
.Y(n_3360)
);

INVx1_ASAP7_75t_L g3361 ( 
.A(n_3205),
.Y(n_3361)
);

INVx1_ASAP7_75t_L g3362 ( 
.A(n_3208),
.Y(n_3362)
);

INVx1_ASAP7_75t_L g3363 ( 
.A(n_3222),
.Y(n_3363)
);

INVx1_ASAP7_75t_L g3364 ( 
.A(n_3225),
.Y(n_3364)
);

NAND2xp5_ASAP7_75t_L g3365 ( 
.A(n_3244),
.B(n_3164),
.Y(n_3365)
);

AND2x2_ASAP7_75t_L g3366 ( 
.A(n_3216),
.B(n_3178),
.Y(n_3366)
);

INVx1_ASAP7_75t_SL g3367 ( 
.A(n_3329),
.Y(n_3367)
);

AOI22xp33_ASAP7_75t_L g3368 ( 
.A1(n_3227),
.A2(n_3032),
.B1(n_3185),
.B2(n_3181),
.Y(n_3368)
);

NAND2xp5_ASAP7_75t_L g3369 ( 
.A(n_3281),
.B(n_3180),
.Y(n_3369)
);

AND2x2_ASAP7_75t_L g3370 ( 
.A(n_3330),
.B(n_3193),
.Y(n_3370)
);

INVx1_ASAP7_75t_L g3371 ( 
.A(n_3232),
.Y(n_3371)
);

INVx1_ASAP7_75t_L g3372 ( 
.A(n_3239),
.Y(n_3372)
);

INVx1_ASAP7_75t_SL g3373 ( 
.A(n_3286),
.Y(n_3373)
);

NOR2xp33_ASAP7_75t_L g3374 ( 
.A(n_3248),
.B(n_3052),
.Y(n_3374)
);

INVxp67_ASAP7_75t_L g3375 ( 
.A(n_3212),
.Y(n_3375)
);

AND2x2_ASAP7_75t_L g3376 ( 
.A(n_3306),
.B(n_3089),
.Y(n_3376)
);

NAND2x1_ASAP7_75t_L g3377 ( 
.A(n_3240),
.B(n_3188),
.Y(n_3377)
);

AOI22xp33_ASAP7_75t_L g3378 ( 
.A1(n_3253),
.A2(n_3191),
.B1(n_3090),
.B2(n_3047),
.Y(n_3378)
);

INVx2_ASAP7_75t_SL g3379 ( 
.A(n_3237),
.Y(n_3379)
);

AND2x2_ASAP7_75t_L g3380 ( 
.A(n_3337),
.B(n_3008),
.Y(n_3380)
);

NOR2xp33_ASAP7_75t_L g3381 ( 
.A(n_3294),
.B(n_3083),
.Y(n_3381)
);

INVx1_ASAP7_75t_L g3382 ( 
.A(n_3246),
.Y(n_3382)
);

NOR2xp33_ASAP7_75t_SL g3383 ( 
.A(n_3283),
.B(n_3075),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3262),
.Y(n_3384)
);

INVx1_ASAP7_75t_L g3385 ( 
.A(n_3276),
.Y(n_3385)
);

AND2x2_ASAP7_75t_L g3386 ( 
.A(n_3324),
.B(n_3092),
.Y(n_3386)
);

INVx1_ASAP7_75t_SL g3387 ( 
.A(n_3302),
.Y(n_3387)
);

OA21x2_ASAP7_75t_L g3388 ( 
.A1(n_3226),
.A2(n_3068),
.B(n_3017),
.Y(n_3388)
);

NAND2xp5_ASAP7_75t_L g3389 ( 
.A(n_3206),
.B(n_3021),
.Y(n_3389)
);

OR2x2_ASAP7_75t_L g3390 ( 
.A(n_3338),
.B(n_3040),
.Y(n_3390)
);

AND2x2_ASAP7_75t_L g3391 ( 
.A(n_3319),
.B(n_445),
.Y(n_3391)
);

NAND2xp5_ASAP7_75t_L g3392 ( 
.A(n_3299),
.B(n_446),
.Y(n_3392)
);

INVx1_ASAP7_75t_L g3393 ( 
.A(n_3279),
.Y(n_3393)
);

INVx1_ASAP7_75t_L g3394 ( 
.A(n_3282),
.Y(n_3394)
);

INVx1_ASAP7_75t_L g3395 ( 
.A(n_3292),
.Y(n_3395)
);

AOI222xp33_ASAP7_75t_SL g3396 ( 
.A1(n_3327),
.A2(n_448),
.B1(n_450),
.B2(n_446),
.C1(n_447),
.C2(n_449),
.Y(n_3396)
);

OR2x2_ASAP7_75t_L g3397 ( 
.A(n_3233),
.B(n_447),
.Y(n_3397)
);

INVxp67_ASAP7_75t_L g3398 ( 
.A(n_3240),
.Y(n_3398)
);

NAND2xp5_ASAP7_75t_L g3399 ( 
.A(n_3297),
.B(n_448),
.Y(n_3399)
);

NAND2x1_ASAP7_75t_L g3400 ( 
.A(n_3290),
.B(n_449),
.Y(n_3400)
);

INVx1_ASAP7_75t_SL g3401 ( 
.A(n_3200),
.Y(n_3401)
);

NAND2xp5_ASAP7_75t_L g3402 ( 
.A(n_3211),
.B(n_3341),
.Y(n_3402)
);

INVx1_ASAP7_75t_L g3403 ( 
.A(n_3304),
.Y(n_3403)
);

INVx1_ASAP7_75t_L g3404 ( 
.A(n_3311),
.Y(n_3404)
);

AND2x2_ASAP7_75t_L g3405 ( 
.A(n_3252),
.B(n_450),
.Y(n_3405)
);

NAND2xp5_ASAP7_75t_L g3406 ( 
.A(n_3238),
.B(n_451),
.Y(n_3406)
);

NAND2xp5_ASAP7_75t_L g3407 ( 
.A(n_3220),
.B(n_452),
.Y(n_3407)
);

NAND2xp5_ASAP7_75t_L g3408 ( 
.A(n_3287),
.B(n_452),
.Y(n_3408)
);

NAND2xp5_ASAP7_75t_L g3409 ( 
.A(n_3221),
.B(n_453),
.Y(n_3409)
);

AND2x2_ASAP7_75t_L g3410 ( 
.A(n_3234),
.B(n_453),
.Y(n_3410)
);

INVx1_ASAP7_75t_L g3411 ( 
.A(n_3320),
.Y(n_3411)
);

NOR2xp33_ASAP7_75t_L g3412 ( 
.A(n_3218),
.B(n_454),
.Y(n_3412)
);

NAND2xp5_ASAP7_75t_L g3413 ( 
.A(n_3254),
.B(n_454),
.Y(n_3413)
);

INVxp67_ASAP7_75t_L g3414 ( 
.A(n_3273),
.Y(n_3414)
);

NOR2xp33_ASAP7_75t_L g3415 ( 
.A(n_3267),
.B(n_455),
.Y(n_3415)
);

OR2x2_ASAP7_75t_L g3416 ( 
.A(n_3280),
.B(n_456),
.Y(n_3416)
);

NOR2xp33_ASAP7_75t_L g3417 ( 
.A(n_3247),
.B(n_456),
.Y(n_3417)
);

INVx1_ASAP7_75t_SL g3418 ( 
.A(n_3256),
.Y(n_3418)
);

OR2x2_ASAP7_75t_L g3419 ( 
.A(n_3307),
.B(n_457),
.Y(n_3419)
);

INVx1_ASAP7_75t_L g3420 ( 
.A(n_3333),
.Y(n_3420)
);

INVx1_ASAP7_75t_L g3421 ( 
.A(n_3336),
.Y(n_3421)
);

INVx3_ASAP7_75t_L g3422 ( 
.A(n_3230),
.Y(n_3422)
);

INVx1_ASAP7_75t_SL g3423 ( 
.A(n_3236),
.Y(n_3423)
);

INVx1_ASAP7_75t_SL g3424 ( 
.A(n_3315),
.Y(n_3424)
);

CKINVDCx20_ASAP7_75t_R g3425 ( 
.A(n_3242),
.Y(n_3425)
);

AND2x2_ASAP7_75t_SL g3426 ( 
.A(n_3217),
.B(n_3314),
.Y(n_3426)
);

INVx1_ASAP7_75t_L g3427 ( 
.A(n_3323),
.Y(n_3427)
);

NAND2xp5_ASAP7_75t_L g3428 ( 
.A(n_3326),
.B(n_457),
.Y(n_3428)
);

OAI31xp33_ASAP7_75t_L g3429 ( 
.A1(n_3243),
.A2(n_460),
.A3(n_458),
.B(n_459),
.Y(n_3429)
);

OR2x2_ASAP7_75t_L g3430 ( 
.A(n_3250),
.B(n_460),
.Y(n_3430)
);

AOI22xp33_ASAP7_75t_L g3431 ( 
.A1(n_3231),
.A2(n_463),
.B1(n_461),
.B2(n_462),
.Y(n_3431)
);

NOR2xp33_ASAP7_75t_SL g3432 ( 
.A(n_3317),
.B(n_462),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3258),
.Y(n_3433)
);

INVx2_ASAP7_75t_L g3434 ( 
.A(n_3305),
.Y(n_3434)
);

INVx1_ASAP7_75t_L g3435 ( 
.A(n_3261),
.Y(n_3435)
);

NAND2xp5_ASAP7_75t_L g3436 ( 
.A(n_3272),
.B(n_3325),
.Y(n_3436)
);

NOR2xp33_ASAP7_75t_L g3437 ( 
.A(n_3199),
.B(n_464),
.Y(n_3437)
);

INVx2_ASAP7_75t_SL g3438 ( 
.A(n_3340),
.Y(n_3438)
);

INVx2_ASAP7_75t_L g3439 ( 
.A(n_3350),
.Y(n_3439)
);

INVx1_ASAP7_75t_SL g3440 ( 
.A(n_3342),
.Y(n_3440)
);

INVx1_ASAP7_75t_L g3441 ( 
.A(n_3347),
.Y(n_3441)
);

INVx5_ASAP7_75t_L g3442 ( 
.A(n_3350),
.Y(n_3442)
);

INVx1_ASAP7_75t_L g3443 ( 
.A(n_3343),
.Y(n_3443)
);

INVx1_ASAP7_75t_L g3444 ( 
.A(n_3344),
.Y(n_3444)
);

INVx2_ASAP7_75t_L g3445 ( 
.A(n_3346),
.Y(n_3445)
);

INVx2_ASAP7_75t_L g3446 ( 
.A(n_3356),
.Y(n_3446)
);

INVx2_ASAP7_75t_L g3447 ( 
.A(n_3351),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3383),
.B(n_3321),
.Y(n_3448)
);

INVx1_ASAP7_75t_L g3449 ( 
.A(n_3354),
.Y(n_3449)
);

BUFx2_ASAP7_75t_L g3450 ( 
.A(n_3379),
.Y(n_3450)
);

INVx1_ASAP7_75t_L g3451 ( 
.A(n_3397),
.Y(n_3451)
);

INVx1_ASAP7_75t_L g3452 ( 
.A(n_3348),
.Y(n_3452)
);

BUFx6f_ASAP7_75t_L g3453 ( 
.A(n_3410),
.Y(n_3453)
);

NAND2xp5_ASAP7_75t_L g3454 ( 
.A(n_3367),
.B(n_3265),
.Y(n_3454)
);

INVx1_ASAP7_75t_L g3455 ( 
.A(n_3355),
.Y(n_3455)
);

INVx1_ASAP7_75t_L g3456 ( 
.A(n_3358),
.Y(n_3456)
);

HB1xp67_ASAP7_75t_L g3457 ( 
.A(n_3373),
.Y(n_3457)
);

INVx1_ASAP7_75t_L g3458 ( 
.A(n_3361),
.Y(n_3458)
);

INVx1_ASAP7_75t_L g3459 ( 
.A(n_3362),
.Y(n_3459)
);

INVx1_ASAP7_75t_SL g3460 ( 
.A(n_3387),
.Y(n_3460)
);

INVx1_ASAP7_75t_L g3461 ( 
.A(n_3363),
.Y(n_3461)
);

BUFx12f_ASAP7_75t_L g3462 ( 
.A(n_3430),
.Y(n_3462)
);

NOR2xp33_ASAP7_75t_L g3463 ( 
.A(n_3352),
.B(n_3375),
.Y(n_3463)
);

INVx1_ASAP7_75t_L g3464 ( 
.A(n_3364),
.Y(n_3464)
);

INVx1_ASAP7_75t_L g3465 ( 
.A(n_3371),
.Y(n_3465)
);

INVxp33_ASAP7_75t_SL g3466 ( 
.A(n_3353),
.Y(n_3466)
);

INVx2_ASAP7_75t_L g3467 ( 
.A(n_3380),
.Y(n_3467)
);

INVxp33_ASAP7_75t_SL g3468 ( 
.A(n_3374),
.Y(n_3468)
);

INVx1_ASAP7_75t_L g3469 ( 
.A(n_3372),
.Y(n_3469)
);

INVxp67_ASAP7_75t_L g3470 ( 
.A(n_3432),
.Y(n_3470)
);

INVx1_ASAP7_75t_L g3471 ( 
.A(n_3382),
.Y(n_3471)
);

NOR2xp33_ASAP7_75t_L g3472 ( 
.A(n_3414),
.B(n_3204),
.Y(n_3472)
);

INVx1_ASAP7_75t_L g3473 ( 
.A(n_3384),
.Y(n_3473)
);

INVx1_ASAP7_75t_L g3474 ( 
.A(n_3385),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3393),
.Y(n_3475)
);

INVx1_ASAP7_75t_SL g3476 ( 
.A(n_3418),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3394),
.Y(n_3477)
);

HB1xp67_ASAP7_75t_L g3478 ( 
.A(n_3377),
.Y(n_3478)
);

INVx1_ASAP7_75t_L g3479 ( 
.A(n_3395),
.Y(n_3479)
);

INVxp67_ASAP7_75t_L g3480 ( 
.A(n_3381),
.Y(n_3480)
);

INVx1_ASAP7_75t_L g3481 ( 
.A(n_3403),
.Y(n_3481)
);

INVx2_ASAP7_75t_L g3482 ( 
.A(n_3366),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3404),
.Y(n_3483)
);

INVxp33_ASAP7_75t_L g3484 ( 
.A(n_3365),
.Y(n_3484)
);

INVx1_ASAP7_75t_L g3485 ( 
.A(n_3411),
.Y(n_3485)
);

CKINVDCx20_ASAP7_75t_R g3486 ( 
.A(n_3425),
.Y(n_3486)
);

INVx2_ASAP7_75t_L g3487 ( 
.A(n_3376),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3420),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3421),
.Y(n_3489)
);

INVx2_ASAP7_75t_L g3490 ( 
.A(n_3434),
.Y(n_3490)
);

INVx1_ASAP7_75t_L g3491 ( 
.A(n_3427),
.Y(n_3491)
);

NOR2xp33_ASAP7_75t_L g3492 ( 
.A(n_3401),
.B(n_3209),
.Y(n_3492)
);

HB1xp67_ASAP7_75t_L g3493 ( 
.A(n_3422),
.Y(n_3493)
);

INVx1_ASAP7_75t_SL g3494 ( 
.A(n_3370),
.Y(n_3494)
);

BUFx2_ASAP7_75t_L g3495 ( 
.A(n_3422),
.Y(n_3495)
);

INVx1_ASAP7_75t_L g3496 ( 
.A(n_3391),
.Y(n_3496)
);

NAND2xp5_ASAP7_75t_L g3497 ( 
.A(n_3426),
.B(n_3277),
.Y(n_3497)
);

INVx1_ASAP7_75t_L g3498 ( 
.A(n_3405),
.Y(n_3498)
);

INVx2_ASAP7_75t_L g3499 ( 
.A(n_3400),
.Y(n_3499)
);

INVx2_ASAP7_75t_L g3500 ( 
.A(n_3345),
.Y(n_3500)
);

INVx2_ASAP7_75t_L g3501 ( 
.A(n_3390),
.Y(n_3501)
);

NOR2xp33_ASAP7_75t_L g3502 ( 
.A(n_3423),
.B(n_3274),
.Y(n_3502)
);

INVx1_ASAP7_75t_L g3503 ( 
.A(n_3408),
.Y(n_3503)
);

INVx1_ASAP7_75t_L g3504 ( 
.A(n_3398),
.Y(n_3504)
);

INVx2_ASAP7_75t_SL g3505 ( 
.A(n_3386),
.Y(n_3505)
);

INVx2_ASAP7_75t_L g3506 ( 
.A(n_3438),
.Y(n_3506)
);

INVx1_ASAP7_75t_L g3507 ( 
.A(n_3416),
.Y(n_3507)
);

INVx1_ASAP7_75t_L g3508 ( 
.A(n_3419),
.Y(n_3508)
);

INVx1_ASAP7_75t_L g3509 ( 
.A(n_3433),
.Y(n_3509)
);

INVx1_ASAP7_75t_L g3510 ( 
.A(n_3435),
.Y(n_3510)
);

INVx1_ASAP7_75t_L g3511 ( 
.A(n_3407),
.Y(n_3511)
);

INVx1_ASAP7_75t_L g3512 ( 
.A(n_3406),
.Y(n_3512)
);

INVx5_ASAP7_75t_L g3513 ( 
.A(n_3396),
.Y(n_3513)
);

INVx1_ASAP7_75t_L g3514 ( 
.A(n_3424),
.Y(n_3514)
);

INVx1_ASAP7_75t_L g3515 ( 
.A(n_3399),
.Y(n_3515)
);

INVx2_ASAP7_75t_SL g3516 ( 
.A(n_3388),
.Y(n_3516)
);

INVx1_ASAP7_75t_L g3517 ( 
.A(n_3392),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3412),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3388),
.Y(n_3519)
);

INVx1_ASAP7_75t_L g3520 ( 
.A(n_3413),
.Y(n_3520)
);

INVx1_ASAP7_75t_SL g3521 ( 
.A(n_3360),
.Y(n_3521)
);

INVx2_ASAP7_75t_L g3522 ( 
.A(n_3369),
.Y(n_3522)
);

INVx1_ASAP7_75t_L g3523 ( 
.A(n_3436),
.Y(n_3523)
);

INVx2_ASAP7_75t_L g3524 ( 
.A(n_3389),
.Y(n_3524)
);

INVx1_ASAP7_75t_L g3525 ( 
.A(n_3409),
.Y(n_3525)
);

INVx2_ASAP7_75t_L g3526 ( 
.A(n_3402),
.Y(n_3526)
);

INVx1_ASAP7_75t_L g3527 ( 
.A(n_3415),
.Y(n_3527)
);

NAND2xp5_ASAP7_75t_L g3528 ( 
.A(n_3368),
.B(n_3334),
.Y(n_3528)
);

AND2x4_ASAP7_75t_L g3529 ( 
.A(n_3357),
.B(n_3228),
.Y(n_3529)
);

INVx1_ASAP7_75t_SL g3530 ( 
.A(n_3428),
.Y(n_3530)
);

INVx1_ASAP7_75t_L g3531 ( 
.A(n_3417),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3437),
.Y(n_3532)
);

INVx8_ASAP7_75t_L g3533 ( 
.A(n_3429),
.Y(n_3533)
);

INVx1_ASAP7_75t_L g3534 ( 
.A(n_3349),
.Y(n_3534)
);

INVx2_ASAP7_75t_L g3535 ( 
.A(n_3378),
.Y(n_3535)
);

OR2x2_ASAP7_75t_L g3536 ( 
.A(n_3359),
.B(n_3298),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3431),
.Y(n_3537)
);

CKINVDCx20_ASAP7_75t_R g3538 ( 
.A(n_3425),
.Y(n_3538)
);

BUFx2_ASAP7_75t_L g3539 ( 
.A(n_3350),
.Y(n_3539)
);

INVx3_ASAP7_75t_SL g3540 ( 
.A(n_3373),
.Y(n_3540)
);

OAI21xp33_ASAP7_75t_SL g3541 ( 
.A1(n_3448),
.A2(n_3335),
.B(n_3201),
.Y(n_3541)
);

NOR3xp33_ASAP7_75t_SL g3542 ( 
.A(n_3463),
.B(n_3284),
.C(n_3269),
.Y(n_3542)
);

OAI221xp5_ASAP7_75t_SL g3543 ( 
.A1(n_3536),
.A2(n_3241),
.B1(n_3224),
.B2(n_3260),
.C(n_3245),
.Y(n_3543)
);

NOR2xp33_ASAP7_75t_L g3544 ( 
.A(n_3466),
.B(n_3259),
.Y(n_3544)
);

NOR2xp33_ASAP7_75t_L g3545 ( 
.A(n_3540),
.B(n_3275),
.Y(n_3545)
);

NAND2xp5_ASAP7_75t_L g3546 ( 
.A(n_3513),
.B(n_3308),
.Y(n_3546)
);

AOI211x1_ASAP7_75t_L g3547 ( 
.A1(n_3528),
.A2(n_3313),
.B(n_3210),
.C(n_3213),
.Y(n_3547)
);

NOR3xp33_ASAP7_75t_L g3548 ( 
.A(n_3497),
.B(n_3263),
.C(n_3322),
.Y(n_3548)
);

NOR2x1_ASAP7_75t_L g3549 ( 
.A(n_3486),
.B(n_3214),
.Y(n_3549)
);

OAI322xp33_ASAP7_75t_L g3550 ( 
.A1(n_3534),
.A2(n_3219),
.A3(n_3339),
.B1(n_3331),
.B2(n_3332),
.C1(n_3293),
.C2(n_3257),
.Y(n_3550)
);

AND4x1_ASAP7_75t_L g3551 ( 
.A(n_3523),
.B(n_3266),
.C(n_3301),
.D(n_3316),
.Y(n_3551)
);

AOI22xp5_ASAP7_75t_L g3552 ( 
.A1(n_3529),
.A2(n_3264),
.B1(n_3270),
.B2(n_3249),
.Y(n_3552)
);

AOI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_3533),
.A2(n_3251),
.B(n_3303),
.Y(n_3553)
);

NAND4xp25_ASAP7_75t_L g3554 ( 
.A(n_3476),
.B(n_3312),
.C(n_3289),
.D(n_3285),
.Y(n_3554)
);

NAND3xp33_ASAP7_75t_SL g3555 ( 
.A(n_3454),
.B(n_3309),
.C(n_3291),
.Y(n_3555)
);

NOR3xp33_ASAP7_75t_L g3556 ( 
.A(n_3480),
.B(n_3300),
.C(n_3278),
.Y(n_3556)
);

INVx1_ASAP7_75t_L g3557 ( 
.A(n_3493),
.Y(n_3557)
);

NOR4xp25_ASAP7_75t_L g3558 ( 
.A(n_3504),
.B(n_3288),
.C(n_467),
.D(n_465),
.Y(n_3558)
);

NOR2x1_ASAP7_75t_L g3559 ( 
.A(n_3538),
.B(n_465),
.Y(n_3559)
);

AOI21xp33_ASAP7_75t_L g3560 ( 
.A1(n_3484),
.A2(n_466),
.B(n_467),
.Y(n_3560)
);

NAND2xp5_ASAP7_75t_L g3561 ( 
.A(n_3513),
.B(n_466),
.Y(n_3561)
);

NAND4xp25_ASAP7_75t_L g3562 ( 
.A(n_3460),
.B(n_470),
.C(n_468),
.D(n_469),
.Y(n_3562)
);

HB1xp67_ASAP7_75t_L g3563 ( 
.A(n_3478),
.Y(n_3563)
);

INVx1_ASAP7_75t_L g3564 ( 
.A(n_3495),
.Y(n_3564)
);

NAND3xp33_ASAP7_75t_L g3565 ( 
.A(n_3457),
.B(n_468),
.C(n_469),
.Y(n_3565)
);

NAND3xp33_ASAP7_75t_L g3566 ( 
.A(n_3519),
.B(n_470),
.C(n_471),
.Y(n_3566)
);

NOR4xp25_ASAP7_75t_L g3567 ( 
.A(n_3521),
.B(n_473),
.C(n_471),
.D(n_472),
.Y(n_3567)
);

NAND3xp33_ASAP7_75t_SL g3568 ( 
.A(n_3440),
.B(n_472),
.C(n_474),
.Y(n_3568)
);

AO21x1_ASAP7_75t_L g3569 ( 
.A1(n_3537),
.A2(n_474),
.B(n_476),
.Y(n_3569)
);

OAI211xp5_ASAP7_75t_SL g3570 ( 
.A1(n_3526),
.A2(n_479),
.B(n_476),
.C(n_478),
.Y(n_3570)
);

INVx1_ASAP7_75t_L g3571 ( 
.A(n_3539),
.Y(n_3571)
);

NAND2xp5_ASAP7_75t_L g3572 ( 
.A(n_3450),
.B(n_478),
.Y(n_3572)
);

NAND5xp2_ASAP7_75t_L g3573 ( 
.A(n_3468),
.B(n_483),
.C(n_481),
.D(n_482),
.E(n_484),
.Y(n_3573)
);

AO21x1_ASAP7_75t_L g3574 ( 
.A1(n_3525),
.A2(n_481),
.B(n_482),
.Y(n_3574)
);

NAND3xp33_ASAP7_75t_L g3575 ( 
.A(n_3442),
.B(n_3516),
.C(n_3470),
.Y(n_3575)
);

NAND2xp5_ASAP7_75t_L g3576 ( 
.A(n_3445),
.B(n_483),
.Y(n_3576)
);

NAND2xp5_ASAP7_75t_SL g3577 ( 
.A(n_3442),
.B(n_484),
.Y(n_3577)
);

NAND4xp75_ASAP7_75t_L g3578 ( 
.A(n_3514),
.B(n_489),
.C(n_487),
.D(n_488),
.Y(n_3578)
);

AND2x2_ASAP7_75t_L g3579 ( 
.A(n_3447),
.B(n_489),
.Y(n_3579)
);

NOR2x1_ASAP7_75t_L g3580 ( 
.A(n_3439),
.B(n_490),
.Y(n_3580)
);

NAND4xp75_ASAP7_75t_L g3581 ( 
.A(n_3444),
.B(n_492),
.C(n_490),
.D(n_491),
.Y(n_3581)
);

NOR3xp33_ASAP7_75t_L g3582 ( 
.A(n_3449),
.B(n_3517),
.C(n_3530),
.Y(n_3582)
);

OAI211xp5_ASAP7_75t_L g3583 ( 
.A1(n_3533),
.A2(n_493),
.B(n_491),
.C(n_492),
.Y(n_3583)
);

NAND2xp5_ASAP7_75t_L g3584 ( 
.A(n_3494),
.B(n_494),
.Y(n_3584)
);

NAND3xp33_ASAP7_75t_L g3585 ( 
.A(n_3522),
.B(n_496),
.C(n_497),
.Y(n_3585)
);

AOI21xp5_ASAP7_75t_L g3586 ( 
.A1(n_3524),
.A2(n_496),
.B(n_497),
.Y(n_3586)
);

NOR2x1_ASAP7_75t_L g3587 ( 
.A(n_3499),
.B(n_498),
.Y(n_3587)
);

OAI211xp5_ASAP7_75t_L g3588 ( 
.A1(n_3535),
.A2(n_500),
.B(n_498),
.C(n_499),
.Y(n_3588)
);

NOR2x1_ASAP7_75t_L g3589 ( 
.A(n_3506),
.B(n_499),
.Y(n_3589)
);

NAND4xp25_ASAP7_75t_SL g3590 ( 
.A(n_3515),
.B(n_3446),
.C(n_3467),
.D(n_3496),
.Y(n_3590)
);

INVx1_ASAP7_75t_L g3591 ( 
.A(n_3500),
.Y(n_3591)
);

O2A1O1Ixp33_ASAP7_75t_L g3592 ( 
.A1(n_3520),
.A2(n_3443),
.B(n_3502),
.C(n_3441),
.Y(n_3592)
);

AOI21xp33_ASAP7_75t_SL g3593 ( 
.A1(n_3505),
.A2(n_501),
.B(n_503),
.Y(n_3593)
);

AOI211xp5_ASAP7_75t_SL g3594 ( 
.A1(n_3492),
.A2(n_505),
.B(n_503),
.C(n_504),
.Y(n_3594)
);

NAND4xp75_ASAP7_75t_L g3595 ( 
.A(n_3491),
.B(n_506),
.C(n_504),
.D(n_505),
.Y(n_3595)
);

OAI211xp5_ASAP7_75t_L g3596 ( 
.A1(n_3472),
.A2(n_508),
.B(n_506),
.C(n_507),
.Y(n_3596)
);

NAND4xp25_ASAP7_75t_L g3597 ( 
.A(n_3482),
.B(n_3487),
.C(n_3501),
.D(n_3507),
.Y(n_3597)
);

NOR2xp33_ASAP7_75t_L g3598 ( 
.A(n_3453),
.B(n_507),
.Y(n_3598)
);

OAI22xp33_ASAP7_75t_SL g3599 ( 
.A1(n_3451),
.A2(n_512),
.B1(n_509),
.B2(n_510),
.Y(n_3599)
);

NOR3x1_ASAP7_75t_L g3600 ( 
.A(n_3498),
.B(n_509),
.C(n_510),
.Y(n_3600)
);

NAND4xp25_ASAP7_75t_L g3601 ( 
.A(n_3508),
.B(n_514),
.C(n_512),
.D(n_513),
.Y(n_3601)
);

NOR4xp25_ASAP7_75t_L g3602 ( 
.A(n_3509),
.B(n_516),
.C(n_513),
.D(n_515),
.Y(n_3602)
);

A2O1A1Ixp33_ASAP7_75t_L g3603 ( 
.A1(n_3527),
.A2(n_517),
.B(n_515),
.C(n_516),
.Y(n_3603)
);

O2A1O1Ixp33_ASAP7_75t_L g3604 ( 
.A1(n_3531),
.A2(n_519),
.B(n_517),
.C(n_518),
.Y(n_3604)
);

NAND3xp33_ASAP7_75t_SL g3605 ( 
.A(n_3532),
.B(n_518),
.C(n_519),
.Y(n_3605)
);

NOR2xp67_ASAP7_75t_SL g3606 ( 
.A(n_3462),
.B(n_520),
.Y(n_3606)
);

NOR2xp33_ASAP7_75t_L g3607 ( 
.A(n_3453),
.B(n_521),
.Y(n_3607)
);

INVx1_ASAP7_75t_L g3608 ( 
.A(n_3490),
.Y(n_3608)
);

NAND4xp25_ASAP7_75t_L g3609 ( 
.A(n_3549),
.B(n_3518),
.C(n_3511),
.D(n_3512),
.Y(n_3609)
);

OAI322xp33_ASAP7_75t_L g3610 ( 
.A1(n_3546),
.A2(n_3458),
.A3(n_3455),
.B1(n_3459),
.B2(n_3461),
.C1(n_3456),
.C2(n_3452),
.Y(n_3610)
);

NAND2xp5_ASAP7_75t_L g3611 ( 
.A(n_3567),
.B(n_3503),
.Y(n_3611)
);

INVx1_ASAP7_75t_L g3612 ( 
.A(n_3557),
.Y(n_3612)
);

NAND2xp5_ASAP7_75t_L g3613 ( 
.A(n_3564),
.B(n_3510),
.Y(n_3613)
);

AOI21xp5_ASAP7_75t_L g3614 ( 
.A1(n_3561),
.A2(n_3465),
.B(n_3464),
.Y(n_3614)
);

AOI222xp33_ASAP7_75t_L g3615 ( 
.A1(n_3541),
.A2(n_3474),
.B1(n_3471),
.B2(n_3475),
.C1(n_3473),
.C2(n_3469),
.Y(n_3615)
);

NAND3xp33_ASAP7_75t_L g3616 ( 
.A(n_3548),
.B(n_3479),
.C(n_3477),
.Y(n_3616)
);

NAND4xp25_ASAP7_75t_L g3617 ( 
.A(n_3575),
.B(n_3483),
.C(n_3485),
.D(n_3481),
.Y(n_3617)
);

AOI22xp5_ASAP7_75t_L g3618 ( 
.A1(n_3552),
.A2(n_3489),
.B1(n_3488),
.B2(n_523),
.Y(n_3618)
);

AOI221xp5_ASAP7_75t_L g3619 ( 
.A1(n_3547),
.A2(n_524),
.B1(n_521),
.B2(n_522),
.C(n_525),
.Y(n_3619)
);

AOI21xp33_ASAP7_75t_L g3620 ( 
.A1(n_3544),
.A2(n_522),
.B(n_524),
.Y(n_3620)
);

OAI22xp5_ASAP7_75t_L g3621 ( 
.A1(n_3543),
.A2(n_527),
.B1(n_525),
.B2(n_526),
.Y(n_3621)
);

HB1xp67_ASAP7_75t_L g3622 ( 
.A(n_3587),
.Y(n_3622)
);

OAI22xp33_ASAP7_75t_SL g3623 ( 
.A1(n_3571),
.A2(n_529),
.B1(n_526),
.B2(n_527),
.Y(n_3623)
);

A2O1A1Ixp33_ASAP7_75t_L g3624 ( 
.A1(n_3583),
.A2(n_532),
.B(n_529),
.C(n_530),
.Y(n_3624)
);

O2A1O1Ixp33_ASAP7_75t_L g3625 ( 
.A1(n_3568),
.A2(n_533),
.B(n_530),
.C(n_532),
.Y(n_3625)
);

INVx2_ASAP7_75t_L g3626 ( 
.A(n_3580),
.Y(n_3626)
);

OAI221xp5_ASAP7_75t_L g3627 ( 
.A1(n_3551),
.A2(n_537),
.B1(n_535),
.B2(n_536),
.C(n_538),
.Y(n_3627)
);

OA22x2_ASAP7_75t_L g3628 ( 
.A1(n_3563),
.A2(n_3591),
.B1(n_3608),
.B2(n_3577),
.Y(n_3628)
);

OAI211xp5_ASAP7_75t_SL g3629 ( 
.A1(n_3553),
.A2(n_537),
.B(n_535),
.C(n_536),
.Y(n_3629)
);

AOI221xp5_ASAP7_75t_L g3630 ( 
.A1(n_3558),
.A2(n_540),
.B1(n_538),
.B2(n_539),
.C(n_541),
.Y(n_3630)
);

AOI21xp5_ASAP7_75t_L g3631 ( 
.A1(n_3550),
.A2(n_540),
.B(n_542),
.Y(n_3631)
);

O2A1O1Ixp33_ASAP7_75t_L g3632 ( 
.A1(n_3599),
.A2(n_545),
.B(n_543),
.C(n_544),
.Y(n_3632)
);

OAI211xp5_ASAP7_75t_L g3633 ( 
.A1(n_3602),
.A2(n_546),
.B(n_543),
.C(n_544),
.Y(n_3633)
);

OAI221xp5_ASAP7_75t_L g3634 ( 
.A1(n_3542),
.A2(n_550),
.B1(n_546),
.B2(n_547),
.C(n_551),
.Y(n_3634)
);

INVx1_ASAP7_75t_L g3635 ( 
.A(n_3572),
.Y(n_3635)
);

OAI311xp33_ASAP7_75t_L g3636 ( 
.A1(n_3597),
.A2(n_553),
.A3(n_551),
.B1(n_552),
.C1(n_554),
.Y(n_3636)
);

AOI321xp33_ASAP7_75t_L g3637 ( 
.A1(n_3582),
.A2(n_555),
.A3(n_558),
.B1(n_552),
.B2(n_554),
.C(n_557),
.Y(n_3637)
);

OAI21xp5_ASAP7_75t_SL g3638 ( 
.A1(n_3545),
.A2(n_555),
.B(n_558),
.Y(n_3638)
);

NAND3xp33_ASAP7_75t_SL g3639 ( 
.A(n_3569),
.B(n_3574),
.C(n_3594),
.Y(n_3639)
);

AOI221xp5_ASAP7_75t_L g3640 ( 
.A1(n_3592),
.A2(n_561),
.B1(n_559),
.B2(n_560),
.C(n_562),
.Y(n_3640)
);

NOR2xp33_ASAP7_75t_L g3641 ( 
.A(n_3606),
.B(n_561),
.Y(n_3641)
);

NAND2xp5_ASAP7_75t_L g3642 ( 
.A(n_3559),
.B(n_3593),
.Y(n_3642)
);

AOI22xp33_ASAP7_75t_L g3643 ( 
.A1(n_3555),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_3643)
);

AOI22xp5_ASAP7_75t_L g3644 ( 
.A1(n_3590),
.A2(n_568),
.B1(n_566),
.B2(n_567),
.Y(n_3644)
);

XOR2x2_ASAP7_75t_L g3645 ( 
.A(n_3578),
.B(n_569),
.Y(n_3645)
);

AOI22xp5_ASAP7_75t_L g3646 ( 
.A1(n_3556),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3646)
);

AOI22xp5_ASAP7_75t_L g3647 ( 
.A1(n_3554),
.A2(n_572),
.B1(n_570),
.B2(n_571),
.Y(n_3647)
);

INVx1_ASAP7_75t_SL g3648 ( 
.A(n_3589),
.Y(n_3648)
);

XNOR2xp5_ASAP7_75t_L g3649 ( 
.A(n_3562),
.B(n_573),
.Y(n_3649)
);

AOI21xp5_ASAP7_75t_L g3650 ( 
.A1(n_3586),
.A2(n_574),
.B(n_576),
.Y(n_3650)
);

AOI221xp5_ASAP7_75t_L g3651 ( 
.A1(n_3560),
.A2(n_584),
.B1(n_582),
.B2(n_583),
.C(n_586),
.Y(n_3651)
);

OAI21xp5_ASAP7_75t_L g3652 ( 
.A1(n_3566),
.A2(n_582),
.B(n_583),
.Y(n_3652)
);

OAI31xp33_ASAP7_75t_L g3653 ( 
.A1(n_3588),
.A2(n_3596),
.A3(n_3570),
.B(n_3573),
.Y(n_3653)
);

AOI21xp5_ASAP7_75t_L g3654 ( 
.A1(n_3605),
.A2(n_584),
.B(n_586),
.Y(n_3654)
);

OAI311xp33_ASAP7_75t_L g3655 ( 
.A1(n_3601),
.A2(n_589),
.A3(n_587),
.B1(n_588),
.C1(n_590),
.Y(n_3655)
);

AOI21xp5_ASAP7_75t_L g3656 ( 
.A1(n_3565),
.A2(n_587),
.B(n_588),
.Y(n_3656)
);

BUFx6f_ASAP7_75t_L g3657 ( 
.A(n_3579),
.Y(n_3657)
);

OAI311xp33_ASAP7_75t_L g3658 ( 
.A1(n_3585),
.A2(n_595),
.A3(n_591),
.B1(n_594),
.C1(n_596),
.Y(n_3658)
);

AOI22xp5_ASAP7_75t_L g3659 ( 
.A1(n_3598),
.A2(n_597),
.B1(n_595),
.B2(n_596),
.Y(n_3659)
);

AOI21xp33_ASAP7_75t_SL g3660 ( 
.A1(n_3584),
.A2(n_598),
.B(n_600),
.Y(n_3660)
);

A2O1A1Ixp33_ASAP7_75t_L g3661 ( 
.A1(n_3604),
.A2(n_601),
.B(n_598),
.C(n_600),
.Y(n_3661)
);

AOI22xp5_ASAP7_75t_L g3662 ( 
.A1(n_3607),
.A2(n_604),
.B1(n_602),
.B2(n_603),
.Y(n_3662)
);

AOI211xp5_ASAP7_75t_L g3663 ( 
.A1(n_3603),
.A2(n_604),
.B(n_602),
.C(n_603),
.Y(n_3663)
);

INVx1_ASAP7_75t_L g3664 ( 
.A(n_3622),
.Y(n_3664)
);

AND2x4_ASAP7_75t_L g3665 ( 
.A(n_3626),
.B(n_3600),
.Y(n_3665)
);

NAND2x1p5_ASAP7_75t_L g3666 ( 
.A(n_3648),
.B(n_3576),
.Y(n_3666)
);

NAND2x1p5_ASAP7_75t_L g3667 ( 
.A(n_3657),
.B(n_3581),
.Y(n_3667)
);

AO22x2_ASAP7_75t_L g3668 ( 
.A1(n_3621),
.A2(n_3595),
.B1(n_609),
.B2(n_605),
.Y(n_3668)
);

INVx1_ASAP7_75t_SL g3669 ( 
.A(n_3642),
.Y(n_3669)
);

HB1xp67_ASAP7_75t_L g3670 ( 
.A(n_3657),
.Y(n_3670)
);

INVx1_ASAP7_75t_L g3671 ( 
.A(n_3657),
.Y(n_3671)
);

XNOR2xp5_ASAP7_75t_L g3672 ( 
.A(n_3649),
.B(n_605),
.Y(n_3672)
);

NOR2x1_ASAP7_75t_L g3673 ( 
.A(n_3639),
.B(n_606),
.Y(n_3673)
);

INVx1_ASAP7_75t_L g3674 ( 
.A(n_3613),
.Y(n_3674)
);

NOR2x1_ASAP7_75t_L g3675 ( 
.A(n_3638),
.B(n_606),
.Y(n_3675)
);

XNOR2x1_ASAP7_75t_L g3676 ( 
.A(n_3645),
.B(n_609),
.Y(n_3676)
);

AND2x2_ASAP7_75t_SL g3677 ( 
.A(n_3611),
.B(n_610),
.Y(n_3677)
);

AND2x4_ASAP7_75t_L g3678 ( 
.A(n_3612),
.B(n_611),
.Y(n_3678)
);

INVx1_ASAP7_75t_L g3679 ( 
.A(n_3628),
.Y(n_3679)
);

INVx2_ASAP7_75t_L g3680 ( 
.A(n_3635),
.Y(n_3680)
);

AND2x2_ASAP7_75t_L g3681 ( 
.A(n_3615),
.B(n_611),
.Y(n_3681)
);

AOI22xp5_ASAP7_75t_L g3682 ( 
.A1(n_3630),
.A2(n_614),
.B1(n_612),
.B2(n_613),
.Y(n_3682)
);

NAND4xp75_ASAP7_75t_L g3683 ( 
.A(n_3631),
.B(n_615),
.C(n_612),
.D(n_614),
.Y(n_3683)
);

XOR2x2_ASAP7_75t_L g3684 ( 
.A(n_3619),
.B(n_616),
.Y(n_3684)
);

XNOR2x1_ASAP7_75t_L g3685 ( 
.A(n_3618),
.B(n_618),
.Y(n_3685)
);

OR2x2_ASAP7_75t_L g3686 ( 
.A(n_3609),
.B(n_618),
.Y(n_3686)
);

NAND4xp75_ASAP7_75t_L g3687 ( 
.A(n_3614),
.B(n_621),
.C(n_619),
.D(n_620),
.Y(n_3687)
);

XNOR2xp5_ASAP7_75t_L g3688 ( 
.A(n_3644),
.B(n_619),
.Y(n_3688)
);

INVxp67_ASAP7_75t_SL g3689 ( 
.A(n_3641),
.Y(n_3689)
);

INVx1_ASAP7_75t_L g3690 ( 
.A(n_3610),
.Y(n_3690)
);

OAI21xp33_ASAP7_75t_L g3691 ( 
.A1(n_3617),
.A2(n_622),
.B(n_623),
.Y(n_3691)
);

XOR2xp5_ASAP7_75t_L g3692 ( 
.A(n_3616),
.B(n_622),
.Y(n_3692)
);

AND2x2_ASAP7_75t_L g3693 ( 
.A(n_3652),
.B(n_623),
.Y(n_3693)
);

NAND4xp75_ASAP7_75t_L g3694 ( 
.A(n_3640),
.B(n_627),
.C(n_624),
.D(n_626),
.Y(n_3694)
);

INVx1_ASAP7_75t_SL g3695 ( 
.A(n_3654),
.Y(n_3695)
);

NOR2xp33_ASAP7_75t_R g3696 ( 
.A(n_3671),
.B(n_3643),
.Y(n_3696)
);

NAND2xp33_ASAP7_75t_SL g3697 ( 
.A(n_3670),
.B(n_3636),
.Y(n_3697)
);

NAND2xp5_ASAP7_75t_L g3698 ( 
.A(n_3665),
.B(n_3653),
.Y(n_3698)
);

NOR2xp33_ASAP7_75t_R g3699 ( 
.A(n_3664),
.B(n_3623),
.Y(n_3699)
);

NOR2xp33_ASAP7_75t_R g3700 ( 
.A(n_3672),
.B(n_3660),
.Y(n_3700)
);

NAND2xp5_ASAP7_75t_SL g3701 ( 
.A(n_3673),
.B(n_3637),
.Y(n_3701)
);

XNOR2xp5_ASAP7_75t_L g3702 ( 
.A(n_3676),
.B(n_3627),
.Y(n_3702)
);

NAND2xp5_ASAP7_75t_SL g3703 ( 
.A(n_3677),
.B(n_3625),
.Y(n_3703)
);

NAND2xp5_ASAP7_75t_L g3704 ( 
.A(n_3681),
.B(n_3624),
.Y(n_3704)
);

NAND2xp5_ASAP7_75t_SL g3705 ( 
.A(n_3667),
.B(n_3632),
.Y(n_3705)
);

NAND2xp5_ASAP7_75t_L g3706 ( 
.A(n_3669),
.B(n_3633),
.Y(n_3706)
);

NAND3xp33_ASAP7_75t_L g3707 ( 
.A(n_3690),
.B(n_3629),
.C(n_3663),
.Y(n_3707)
);

NOR2xp33_ASAP7_75t_R g3708 ( 
.A(n_3679),
.B(n_3620),
.Y(n_3708)
);

NOR2xp33_ASAP7_75t_R g3709 ( 
.A(n_3688),
.B(n_3634),
.Y(n_3709)
);

NOR3xp33_ASAP7_75t_SL g3710 ( 
.A(n_3691),
.B(n_3661),
.C(n_3658),
.Y(n_3710)
);

NAND2xp5_ASAP7_75t_L g3711 ( 
.A(n_3668),
.B(n_3656),
.Y(n_3711)
);

NAND2xp33_ASAP7_75t_L g3712 ( 
.A(n_3699),
.B(n_3687),
.Y(n_3712)
);

INVx1_ASAP7_75t_L g3713 ( 
.A(n_3698),
.Y(n_3713)
);

OAI221xp5_ASAP7_75t_L g3714 ( 
.A1(n_3697),
.A2(n_3686),
.B1(n_3695),
.B2(n_3692),
.C(n_3666),
.Y(n_3714)
);

NAND2xp5_ASAP7_75t_L g3715 ( 
.A(n_3702),
.B(n_3668),
.Y(n_3715)
);

INVxp67_ASAP7_75t_SL g3716 ( 
.A(n_3703),
.Y(n_3716)
);

OAI22xp5_ASAP7_75t_L g3717 ( 
.A1(n_3707),
.A2(n_3647),
.B1(n_3682),
.B2(n_3706),
.Y(n_3717)
);

INVx1_ASAP7_75t_L g3718 ( 
.A(n_3716),
.Y(n_3718)
);

AOI21xp5_ASAP7_75t_L g3719 ( 
.A1(n_3712),
.A2(n_3701),
.B(n_3705),
.Y(n_3719)
);

AOI22xp33_ASAP7_75t_L g3720 ( 
.A1(n_3713),
.A2(n_3708),
.B1(n_3696),
.B2(n_3704),
.Y(n_3720)
);

INVx1_ASAP7_75t_L g3721 ( 
.A(n_3718),
.Y(n_3721)
);

INVx2_ASAP7_75t_L g3722 ( 
.A(n_3719),
.Y(n_3722)
);

XNOR2xp5_ASAP7_75t_L g3723 ( 
.A(n_3720),
.B(n_3684),
.Y(n_3723)
);

AOI31xp33_ASAP7_75t_L g3724 ( 
.A1(n_3723),
.A2(n_3715),
.A3(n_3689),
.B(n_3711),
.Y(n_3724)
);

AOI31xp33_ASAP7_75t_L g3725 ( 
.A1(n_3721),
.A2(n_3722),
.A3(n_3674),
.B(n_3680),
.Y(n_3725)
);

AOI22xp33_ASAP7_75t_L g3726 ( 
.A1(n_3722),
.A2(n_3714),
.B1(n_3717),
.B2(n_3709),
.Y(n_3726)
);

NAND2xp5_ASAP7_75t_L g3727 ( 
.A(n_3724),
.B(n_3675),
.Y(n_3727)
);

OAI22xp5_ASAP7_75t_L g3728 ( 
.A1(n_3726),
.A2(n_3683),
.B1(n_3710),
.B2(n_3685),
.Y(n_3728)
);

O2A1O1Ixp33_ASAP7_75t_L g3729 ( 
.A1(n_3725),
.A2(n_3655),
.B(n_3678),
.C(n_3693),
.Y(n_3729)
);

AOI21xp5_ASAP7_75t_L g3730 ( 
.A1(n_3727),
.A2(n_3650),
.B(n_3651),
.Y(n_3730)
);

OAI21xp5_ASAP7_75t_L g3731 ( 
.A1(n_3729),
.A2(n_3728),
.B(n_3646),
.Y(n_3731)
);

OAI21xp5_ASAP7_75t_L g3732 ( 
.A1(n_3729),
.A2(n_3694),
.B(n_3662),
.Y(n_3732)
);

HB1xp67_ASAP7_75t_L g3733 ( 
.A(n_3732),
.Y(n_3733)
);

INVx1_ASAP7_75t_L g3734 ( 
.A(n_3731),
.Y(n_3734)
);

AOI221xp5_ASAP7_75t_L g3735 ( 
.A1(n_3734),
.A2(n_3730),
.B1(n_3733),
.B2(n_3700),
.C(n_3659),
.Y(n_3735)
);

AOI211xp5_ASAP7_75t_L g3736 ( 
.A1(n_3735),
.A2(n_630),
.B(n_628),
.C(n_629),
.Y(n_3736)
);


endmodule