module fake_netlist_6_4041_n_191 (n_16, n_1, n_9, n_8, n_18, n_10, n_21, n_24, n_6, n_15, n_27, n_3, n_14, n_0, n_4, n_22, n_26, n_13, n_11, n_28, n_17, n_23, n_12, n_20, n_7, n_30, n_2, n_5, n_19, n_29, n_31, n_25, n_191);

input n_16;
input n_1;
input n_9;
input n_8;
input n_18;
input n_10;
input n_21;
input n_24;
input n_6;
input n_15;
input n_27;
input n_3;
input n_14;
input n_0;
input n_4;
input n_22;
input n_26;
input n_13;
input n_11;
input n_28;
input n_17;
input n_23;
input n_12;
input n_20;
input n_7;
input n_30;
input n_2;
input n_5;
input n_19;
input n_29;
input n_31;
input n_25;

output n_191;

wire n_52;
wire n_91;
wire n_119;
wire n_46;
wire n_146;
wire n_163;
wire n_147;
wire n_154;
wire n_88;
wire n_98;
wire n_113;
wire n_39;
wire n_63;
wire n_73;
wire n_148;
wire n_138;
wire n_161;
wire n_68;
wire n_166;
wire n_184;
wire n_50;
wire n_158;
wire n_49;
wire n_83;
wire n_101;
wire n_167;
wire n_144;
wire n_174;
wire n_127;
wire n_125;
wire n_168;
wire n_153;
wire n_178;
wire n_77;
wire n_156;
wire n_149;
wire n_152;
wire n_106;
wire n_92;
wire n_145;
wire n_42;
wire n_133;
wire n_96;
wire n_90;
wire n_160;
wire n_105;
wire n_131;
wire n_54;
wire n_132;
wire n_188;
wire n_102;
wire n_186;
wire n_87;
wire n_189;
wire n_32;
wire n_66;
wire n_85;
wire n_99;
wire n_78;
wire n_84;
wire n_130;
wire n_164;
wire n_100;
wire n_129;
wire n_121;
wire n_137;
wire n_142;
wire n_143;
wire n_180;
wire n_47;
wire n_62;
wire n_155;
wire n_75;
wire n_109;
wire n_150;
wire n_122;
wire n_45;
wire n_34;
wire n_140;
wire n_70;
wire n_120;
wire n_37;
wire n_67;
wire n_33;
wire n_82;
wire n_38;
wire n_110;
wire n_151;
wire n_61;
wire n_112;
wire n_172;
wire n_81;
wire n_59;
wire n_181;
wire n_76;
wire n_36;
wire n_182;
wire n_124;
wire n_55;
wire n_126;
wire n_94;
wire n_97;
wire n_108;
wire n_58;
wire n_116;
wire n_64;
wire n_117;
wire n_118;
wire n_175;
wire n_48;
wire n_65;
wire n_40;
wire n_93;
wire n_80;
wire n_141;
wire n_135;
wire n_165;
wire n_139;
wire n_41;
wire n_134;
wire n_177;
wire n_176;
wire n_114;
wire n_86;
wire n_104;
wire n_95;
wire n_179;
wire n_107;
wire n_71;
wire n_74;
wire n_190;
wire n_123;
wire n_136;
wire n_72;
wire n_187;
wire n_89;
wire n_173;
wire n_103;
wire n_111;
wire n_60;
wire n_159;
wire n_157;
wire n_162;
wire n_170;
wire n_185;
wire n_35;
wire n_183;
wire n_115;
wire n_69;
wire n_128;
wire n_79;
wire n_43;
wire n_171;
wire n_57;
wire n_169;
wire n_53;
wire n_51;
wire n_44;
wire n_56;

INVx2_ASAP7_75t_L g32 ( 
.A(n_26),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_6),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVxp67_ASAP7_75t_SL g35 ( 
.A(n_10),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_3),
.Y(n_37)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

INVxp67_ASAP7_75t_SL g41 ( 
.A(n_22),
.Y(n_41)
);

CKINVDCx5p33_ASAP7_75t_R g42 ( 
.A(n_14),
.Y(n_42)
);

INVxp67_ASAP7_75t_SL g43 ( 
.A(n_24),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_12),
.Y(n_44)
);

INVxp33_ASAP7_75t_L g45 ( 
.A(n_21),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_6),
.Y(n_46)
);

CKINVDCx5p33_ASAP7_75t_R g47 ( 
.A(n_8),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_1),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_15),
.Y(n_49)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_7),
.Y(n_50)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_11),
.Y(n_51)
);

INVx1_ASAP7_75t_SL g52 ( 
.A(n_9),
.Y(n_52)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_27),
.Y(n_53)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_32),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_37),
.Y(n_55)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_37),
.Y(n_56)
);

INVx2_ASAP7_75t_L g57 ( 
.A(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_32),
.B(n_0),
.Y(n_58)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_40),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_34),
.B(n_0),
.Y(n_61)
);

CKINVDCx5p33_ASAP7_75t_R g62 ( 
.A(n_42),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

OAI22xp33_ASAP7_75t_L g64 ( 
.A1(n_52),
.A2(n_1),
.B1(n_2),
.B2(n_3),
.Y(n_64)
);

OR2x6_ASAP7_75t_L g65 ( 
.A(n_34),
.B(n_2),
.Y(n_65)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_38),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_39),
.B(n_4),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g68 ( 
.A(n_45),
.B(n_4),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_39),
.B(n_5),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_33),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_70)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_53),
.Y(n_71)
);

INVx2_ASAP7_75t_L g72 ( 
.A(n_53),
.Y(n_72)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_44),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_44),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_62),
.B(n_47),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_55),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_SL g77 ( 
.A(n_68),
.B(n_52),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_61),
.B(n_51),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g79 ( 
.A(n_58),
.B(n_51),
.Y(n_79)
);

INVx2_ASAP7_75t_L g80 ( 
.A(n_57),
.Y(n_80)
);

INVx2_ASAP7_75t_SL g81 ( 
.A(n_66),
.Y(n_81)
);

INVx2_ASAP7_75t_L g82 ( 
.A(n_57),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_R g83 ( 
.A(n_59),
.B(n_36),
.Y(n_83)
);

AND2x4_ASAP7_75t_L g84 ( 
.A(n_66),
.B(n_43),
.Y(n_84)
);

INVx3_ASAP7_75t_L g85 ( 
.A(n_57),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g86 ( 
.A(n_65),
.Y(n_86)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_54),
.Y(n_87)
);

CKINVDCx5p33_ASAP7_75t_R g88 ( 
.A(n_65),
.Y(n_88)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_54),
.Y(n_89)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_66),
.Y(n_90)
);

BUFx2_ASAP7_75t_L g91 ( 
.A(n_65),
.Y(n_91)
);

OAI21x1_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_59),
.B(n_54),
.Y(n_92)
);

INVx3_ASAP7_75t_L g93 ( 
.A(n_80),
.Y(n_93)
);

OAI22x1_ASAP7_75t_L g94 ( 
.A1(n_88),
.A2(n_70),
.B1(n_35),
.B2(n_50),
.Y(n_94)
);

AOI31xp67_ASAP7_75t_L g95 ( 
.A1(n_78),
.A2(n_72),
.A3(n_71),
.B(n_67),
.Y(n_95)
);

INVx5_ASAP7_75t_L g96 ( 
.A(n_85),
.Y(n_96)
);

AND2x2_ASAP7_75t_SL g97 ( 
.A(n_91),
.B(n_69),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_84),
.B(n_59),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_84),
.B(n_59),
.Y(n_99)
);

INVxp67_ASAP7_75t_SL g100 ( 
.A(n_85),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_84),
.B(n_72),
.Y(n_101)
);

AOI221xp5_ASAP7_75t_L g102 ( 
.A1(n_77),
.A2(n_64),
.B1(n_70),
.B2(n_46),
.C(n_48),
.Y(n_102)
);

BUFx2_ASAP7_75t_L g103 ( 
.A(n_83),
.Y(n_103)
);

AOI21xp5_ASAP7_75t_SL g104 ( 
.A1(n_98),
.A2(n_84),
.B(n_81),
.Y(n_104)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_98),
.Y(n_105)
);

A2O1A1Ixp33_ASAP7_75t_SL g106 ( 
.A1(n_100),
.A2(n_41),
.B(n_71),
.C(n_72),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_94),
.A2(n_65),
.B1(n_86),
.B2(n_91),
.Y(n_107)
);

NOR2x1_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_65),
.Y(n_108)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_93),
.Y(n_109)
);

A2O1A1Ixp33_ASAP7_75t_L g110 ( 
.A1(n_99),
.A2(n_92),
.B(n_102),
.C(n_97),
.Y(n_110)
);

CKINVDCx5p33_ASAP7_75t_R g111 ( 
.A(n_103),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_105),
.B(n_103),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_111),
.B(n_94),
.Y(n_113)
);

INVx3_ASAP7_75t_L g114 ( 
.A(n_109),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_L g115 ( 
.A(n_105),
.B(n_97),
.Y(n_115)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_109),
.Y(n_116)
);

NAND2x1p5_ASAP7_75t_L g117 ( 
.A(n_108),
.B(n_92),
.Y(n_117)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_110),
.Y(n_118)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_116),
.Y(n_119)
);

INVx2_ASAP7_75t_L g120 ( 
.A(n_116),
.Y(n_120)
);

AO21x2_ASAP7_75t_L g121 ( 
.A1(n_118),
.A2(n_104),
.B(n_106),
.Y(n_121)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_114),
.Y(n_122)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_114),
.Y(n_123)
);

INVx1_ASAP7_75t_SL g124 ( 
.A(n_119),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g125 ( 
.A(n_120),
.B(n_115),
.Y(n_125)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_119),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_120),
.B(n_97),
.Y(n_127)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_122),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g129 ( 
.A1(n_122),
.A2(n_118),
.B1(n_112),
.B2(n_113),
.Y(n_129)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_123),
.Y(n_130)
);

NOR2x1_ASAP7_75t_L g131 ( 
.A(n_123),
.B(n_104),
.Y(n_131)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_121),
.B(n_113),
.Y(n_132)
);

AND2x2_ASAP7_75t_L g133 ( 
.A(n_121),
.B(n_108),
.Y(n_133)
);

HB1xp67_ASAP7_75t_L g134 ( 
.A(n_121),
.Y(n_134)
);

OAI221xp5_ASAP7_75t_SL g135 ( 
.A1(n_132),
.A2(n_107),
.B1(n_49),
.B2(n_48),
.C(n_46),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_L g136 ( 
.A1(n_131),
.A2(n_117),
.B(n_114),
.Y(n_136)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_126),
.Y(n_137)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_132),
.Y(n_138)
);

AND2x2_ASAP7_75t_L g139 ( 
.A(n_130),
.B(n_127),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g140 ( 
.A1(n_129),
.A2(n_86),
.B1(n_49),
.B2(n_50),
.Y(n_140)
);

AOI221xp5_ASAP7_75t_L g141 ( 
.A1(n_124),
.A2(n_75),
.B1(n_73),
.B2(n_63),
.C(n_55),
.Y(n_141)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_128),
.Y(n_142)
);

NOR4xp25_ASAP7_75t_L g143 ( 
.A(n_135),
.B(n_133),
.C(n_128),
.D(n_125),
.Y(n_143)
);

NOR3x1_ASAP7_75t_L g144 ( 
.A(n_137),
.B(n_73),
.C(n_63),
.Y(n_144)
);

INVx3_ASAP7_75t_SL g145 ( 
.A(n_138),
.Y(n_145)
);

OAI22xp33_ASAP7_75t_L g146 ( 
.A1(n_140),
.A2(n_131),
.B1(n_117),
.B2(n_134),
.Y(n_146)
);

NAND4xp25_ASAP7_75t_L g147 ( 
.A(n_141),
.B(n_60),
.C(n_56),
.D(n_76),
.Y(n_147)
);

AOI221x1_ASAP7_75t_L g148 ( 
.A1(n_136),
.A2(n_133),
.B1(n_130),
.B2(n_71),
.C(n_60),
.Y(n_148)
);

AOI221xp5_ASAP7_75t_L g149 ( 
.A1(n_139),
.A2(n_56),
.B1(n_76),
.B2(n_74),
.C(n_54),
.Y(n_149)
);

AOI211xp5_ASAP7_75t_L g150 ( 
.A1(n_139),
.A2(n_74),
.B(n_81),
.C(n_13),
.Y(n_150)
);

NAND2xp5_ASAP7_75t_SL g151 ( 
.A(n_142),
.B(n_117),
.Y(n_151)
);

AO22x1_ASAP7_75t_L g152 ( 
.A1(n_142),
.A2(n_74),
.B1(n_114),
.B2(n_13),
.Y(n_152)
);

NOR2x1p5_ASAP7_75t_L g153 ( 
.A(n_147),
.B(n_90),
.Y(n_153)
);

INVx1_ASAP7_75t_SL g154 ( 
.A(n_145),
.Y(n_154)
);

NAND3xp33_ASAP7_75t_L g155 ( 
.A(n_150),
.B(n_90),
.C(n_87),
.Y(n_155)
);

AND2x2_ASAP7_75t_L g156 ( 
.A(n_151),
.B(n_10),
.Y(n_156)
);

INVx2_ASAP7_75t_SL g157 ( 
.A(n_152),
.Y(n_157)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_149),
.Y(n_158)
);

NAND2xp33_ASAP7_75t_SL g159 ( 
.A(n_144),
.B(n_11),
.Y(n_159)
);

HB1xp67_ASAP7_75t_L g160 ( 
.A(n_143),
.Y(n_160)
);

NOR2xp67_ASAP7_75t_L g161 ( 
.A(n_148),
.B(n_14),
.Y(n_161)
);

NOR2x1p5_ASAP7_75t_L g162 ( 
.A(n_155),
.B(n_143),
.Y(n_162)
);

NAND3x1_ASAP7_75t_SL g163 ( 
.A(n_156),
.B(n_15),
.C(n_146),
.Y(n_163)
);

AND2x4_ASAP7_75t_L g164 ( 
.A(n_154),
.B(n_17),
.Y(n_164)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_156),
.Y(n_165)
);

OR2x2_ASAP7_75t_L g166 ( 
.A(n_160),
.B(n_87),
.Y(n_166)
);

AND2x2_ASAP7_75t_SL g167 ( 
.A(n_157),
.B(n_87),
.Y(n_167)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_157),
.Y(n_168)
);

OR2x2_ASAP7_75t_L g169 ( 
.A(n_161),
.B(n_89),
.Y(n_169)
);

AOI22xp33_ASAP7_75t_L g170 ( 
.A1(n_158),
.A2(n_89),
.B1(n_82),
.B2(n_80),
.Y(n_170)
);

AOI32xp33_ASAP7_75t_L g171 ( 
.A1(n_168),
.A2(n_159),
.A3(n_161),
.B1(n_153),
.B2(n_28),
.Y(n_171)
);

OAI322xp33_ASAP7_75t_L g172 ( 
.A1(n_165),
.A2(n_89),
.A3(n_82),
.B1(n_80),
.B2(n_153),
.C1(n_85),
.C2(n_31),
.Y(n_172)
);

OAI22xp5_ASAP7_75t_L g173 ( 
.A1(n_162),
.A2(n_167),
.B1(n_165),
.B2(n_163),
.Y(n_173)
);

A2O1A1Ixp33_ASAP7_75t_L g174 ( 
.A1(n_167),
.A2(n_19),
.B(n_20),
.C(n_25),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_166),
.Y(n_175)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_164),
.A2(n_29),
.B(n_30),
.C(n_95),
.Y(n_176)
);

AOI322xp5_ASAP7_75t_L g177 ( 
.A1(n_164),
.A2(n_85),
.A3(n_93),
.B1(n_95),
.B2(n_96),
.C1(n_163),
.C2(n_170),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g178 ( 
.A(n_175),
.B(n_169),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_173),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g180 ( 
.A(n_177),
.B(n_170),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_L g181 ( 
.A1(n_174),
.A2(n_93),
.B(n_96),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_172),
.Y(n_182)
);

INVx2_ASAP7_75t_L g183 ( 
.A(n_171),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_176),
.B(n_93),
.Y(n_184)
);

OAI22xp33_ASAP7_75t_L g185 ( 
.A1(n_183),
.A2(n_96),
.B1(n_180),
.B2(n_179),
.Y(n_185)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_178),
.Y(n_186)
);

INVx2_ASAP7_75t_L g187 ( 
.A(n_178),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_183),
.A2(n_96),
.B1(n_182),
.B2(n_181),
.Y(n_188)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_186),
.Y(n_189)
);

AOI21xp5_ASAP7_75t_L g190 ( 
.A1(n_185),
.A2(n_184),
.B(n_96),
.Y(n_190)
);

AOI221xp5_ASAP7_75t_L g191 ( 
.A1(n_189),
.A2(n_96),
.B1(n_187),
.B2(n_188),
.C(n_190),
.Y(n_191)
);


endmodule