module fake_jpeg_120_n_116 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_116);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_116;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

BUFx3_ASAP7_75t_L g12 ( 
.A(n_2),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_5),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_2),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_6),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_1),
.B(n_4),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_11),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

INVxp67_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

INVx11_ASAP7_75t_L g21 ( 
.A(n_7),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_3),
.B(n_8),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_10),
.B(n_4),
.Y(n_24)
);

BUFx12f_ASAP7_75t_L g25 ( 
.A(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_3),
.Y(n_26)
);

OR2x2_ASAP7_75t_L g57 ( 
.A(n_26),
.B(n_32),
.Y(n_57)
);

INVx13_ASAP7_75t_L g27 ( 
.A(n_21),
.Y(n_27)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_27),
.Y(n_59)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_19),
.Y(n_28)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_28),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_25),
.Y(n_29)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_29),
.Y(n_45)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_25),
.Y(n_30)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_30),
.Y(n_58)
);

INVx5_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g32 ( 
.A(n_24),
.B(n_5),
.Y(n_32)
);

INVx13_ASAP7_75t_L g33 ( 
.A(n_21),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_33),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g34 ( 
.A1(n_19),
.A2(n_12),
.B1(n_23),
.B2(n_15),
.Y(n_34)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_34),
.A2(n_37),
.B1(n_28),
.B2(n_33),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_35),
.Y(n_62)
);

INVx8_ASAP7_75t_L g36 ( 
.A(n_16),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_36),
.B(n_0),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_25),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_37),
.B(n_12),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_18),
.B(n_9),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_38),
.B(n_39),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_17),
.B(n_10),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_20),
.B(n_0),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_40),
.B(n_17),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g41 ( 
.A(n_15),
.B(n_0),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_SL g50 ( 
.A(n_41),
.B(n_32),
.Y(n_50)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_42),
.Y(n_64)
);

AOI22xp33_ASAP7_75t_SL g43 ( 
.A1(n_30),
.A2(n_13),
.B1(n_14),
.B2(n_20),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_43),
.B(n_46),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_13),
.B1(n_14),
.B2(n_23),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_44),
.B(n_49),
.Y(n_66)
);

MAJIxp5_ASAP7_75t_L g47 ( 
.A(n_29),
.B(n_1),
.C(n_35),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_47),
.B(n_48),
.C(n_61),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_26),
.B(n_1),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_50),
.B(n_51),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_31),
.B(n_29),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_35),
.B(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g68 ( 
.A(n_52),
.B(n_53),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_28),
.B(n_36),
.Y(n_53)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_28),
.B(n_27),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_55),
.B(n_60),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_50),
.Y(n_74)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_42),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_69),
.B(n_72),
.Y(n_85)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_62),
.Y(n_70)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_70),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_52),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_60),
.Y(n_73)
);

INVx4_ASAP7_75t_L g84 ( 
.A(n_73),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_74),
.B(n_78),
.Y(n_80)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_62),
.Y(n_75)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_75),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_61),
.B(n_49),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_76),
.B(n_79),
.C(n_59),
.Y(n_83)
);

INVxp67_ASAP7_75t_L g90 ( 
.A(n_77),
.Y(n_90)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_48),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_68),
.B(n_56),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_81),
.B(n_88),
.Y(n_94)
);

AOI22xp5_ASAP7_75t_L g82 ( 
.A1(n_67),
.A2(n_51),
.B1(n_47),
.B2(n_59),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_82),
.A2(n_86),
.B1(n_69),
.B2(n_71),
.Y(n_96)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_83),
.B(n_89),
.C(n_79),
.Y(n_93)
);

AOI22xp5_ASAP7_75t_L g86 ( 
.A1(n_67),
.A2(n_58),
.B1(n_45),
.B2(n_57),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_76),
.Y(n_88)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_64),
.B(n_58),
.C(n_57),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_85),
.B(n_64),
.Y(n_92)
);

AND2x2_ASAP7_75t_L g101 ( 
.A(n_92),
.B(n_97),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g103 ( 
.A(n_93),
.B(n_83),
.C(n_89),
.Y(n_103)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_87),
.Y(n_95)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g100 ( 
.A1(n_96),
.A2(n_98),
.B1(n_90),
.B2(n_66),
.Y(n_100)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_91),
.Y(n_97)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_80),
.Y(n_98)
);

NAND3xp33_ASAP7_75t_L g99 ( 
.A(n_90),
.B(n_66),
.C(n_78),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_SL g104 ( 
.A(n_99),
.B(n_82),
.Y(n_104)
);

XNOR2xp5_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_104),
.Y(n_107)
);

MAJIxp5_ASAP7_75t_L g108 ( 
.A(n_103),
.B(n_93),
.C(n_96),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_92),
.A2(n_86),
.B1(n_70),
.B2(n_75),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_105),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_108),
.B(n_109),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_103),
.B(n_94),
.C(n_97),
.Y(n_109)
);

BUFx24_ASAP7_75t_SL g110 ( 
.A(n_107),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_110),
.B(n_112),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_106),
.B(n_101),
.Y(n_112)
);

A2O1A1Ixp33_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_101),
.B(n_102),
.C(n_84),
.Y(n_113)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_113),
.B(n_84),
.C(n_73),
.Y(n_115)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_115),
.B(n_114),
.Y(n_116)
);


endmodule