module fake_jpeg_2138_n_230 (n_13, n_21, n_53, n_33, n_1, n_45, n_10, n_23, n_27, n_6, n_22, n_47, n_51, n_14, n_40, n_19, n_18, n_20, n_35, n_48, n_52, n_46, n_41, n_4, n_34, n_30, n_39, n_42, n_16, n_49, n_3, n_0, n_24, n_28, n_38, n_26, n_44, n_9, n_5, n_36, n_11, n_17, n_25, n_31, n_2, n_29, n_37, n_43, n_50, n_12, n_32, n_8, n_15, n_7, n_230);

input n_13;
input n_21;
input n_53;
input n_33;
input n_1;
input n_45;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_47;
input n_51;
input n_14;
input n_40;
input n_19;
input n_18;
input n_20;
input n_35;
input n_48;
input n_52;
input n_46;
input n_41;
input n_4;
input n_34;
input n_30;
input n_39;
input n_42;
input n_16;
input n_49;
input n_3;
input n_0;
input n_24;
input n_28;
input n_38;
input n_26;
input n_44;
input n_9;
input n_5;
input n_36;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_37;
input n_43;
input n_50;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_230;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_228;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_155;
wire n_207;
wire n_103;
wire n_150;
wire n_160;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_223;
wire n_171;
wire n_119;
wire n_69;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_143;
wire n_202;
wire n_122;
wire n_75;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_145;
wire n_108;
wire n_68;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_211;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_91;
wire n_54;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_149;
wire n_157;
wire n_87;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_18),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_24),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_42),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx3_ASAP7_75t_L g58 ( 
.A(n_53),
.Y(n_58)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_32),
.Y(n_59)
);

INVx6_ASAP7_75t_SL g60 ( 
.A(n_37),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_5),
.Y(n_61)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_25),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_39),
.Y(n_64)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_29),
.Y(n_65)
);

BUFx3_ASAP7_75t_L g66 ( 
.A(n_28),
.Y(n_66)
);

BUFx12_ASAP7_75t_L g67 ( 
.A(n_36),
.Y(n_67)
);

INVx6_ASAP7_75t_L g68 ( 
.A(n_2),
.Y(n_68)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_30),
.Y(n_69)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_34),
.Y(n_70)
);

CKINVDCx20_ASAP7_75t_R g71 ( 
.A(n_31),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_23),
.Y(n_72)
);

BUFx5_ASAP7_75t_L g73 ( 
.A(n_40),
.Y(n_73)
);

INVx1_ASAP7_75t_L g74 ( 
.A(n_52),
.Y(n_74)
);

CKINVDCx20_ASAP7_75t_R g75 ( 
.A(n_26),
.Y(n_75)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_10),
.Y(n_76)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_46),
.Y(n_77)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_15),
.Y(n_78)
);

BUFx12_ASAP7_75t_L g79 ( 
.A(n_50),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_51),
.Y(n_80)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_81),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_56),
.Y(n_82)
);

INVx6_ASAP7_75t_L g101 ( 
.A(n_82),
.Y(n_101)
);

BUFx6f_ASAP7_75t_L g83 ( 
.A(n_56),
.Y(n_83)
);

INVx3_ASAP7_75t_SL g93 ( 
.A(n_83),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g84 ( 
.A(n_59),
.Y(n_84)
);

INVx2_ASAP7_75t_SL g99 ( 
.A(n_84),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g85 ( 
.A(n_59),
.Y(n_85)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_85),
.Y(n_94)
);

INVx2_ASAP7_75t_L g86 ( 
.A(n_63),
.Y(n_86)
);

INVxp67_ASAP7_75t_L g100 ( 
.A(n_86),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g87 ( 
.A(n_65),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_87),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_SL g88 ( 
.A(n_54),
.B(n_0),
.Y(n_88)
);

AOI21xp33_ASAP7_75t_L g98 ( 
.A1(n_88),
.A2(n_60),
.B(n_62),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g89 ( 
.A(n_65),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g90 ( 
.A(n_89),
.B(n_57),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_98),
.Y(n_109)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_82),
.A2(n_57),
.B1(n_76),
.B2(n_78),
.Y(n_91)
);

OAI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_91),
.A2(n_89),
.B1(n_87),
.B2(n_80),
.Y(n_113)
);

AND2x2_ASAP7_75t_SL g92 ( 
.A(n_81),
.B(n_66),
.Y(n_92)
);

XNOR2xp5_ASAP7_75t_L g110 ( 
.A(n_92),
.B(n_102),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g96 ( 
.A1(n_83),
.A2(n_58),
.B1(n_55),
.B2(n_69),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_96),
.A2(n_97),
.B1(n_60),
.B2(n_69),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_L g97 ( 
.A1(n_84),
.A2(n_68),
.B1(n_58),
.B2(n_66),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g102 ( 
.A1(n_85),
.A2(n_78),
.B1(n_62),
.B2(n_76),
.Y(n_102)
);

INVx4_ASAP7_75t_L g104 ( 
.A(n_99),
.Y(n_104)
);

INVx3_ASAP7_75t_L g131 ( 
.A(n_104),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g105 ( 
.A(n_101),
.Y(n_105)
);

INVx2_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

INVx6_ASAP7_75t_L g106 ( 
.A(n_99),
.Y(n_106)
);

INVx2_ASAP7_75t_L g136 ( 
.A(n_106),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_100),
.B(n_55),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g127 ( 
.A(n_107),
.B(n_113),
.Y(n_127)
);

INVx4_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

HB1xp67_ASAP7_75t_L g126 ( 
.A(n_108),
.Y(n_126)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_94),
.Y(n_111)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_111),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g112 ( 
.A(n_96),
.B(n_80),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_112),
.B(n_115),
.Y(n_124)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_94),
.Y(n_114)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_100),
.Y(n_115)
);

INVx5_ASAP7_75t_L g116 ( 
.A(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_116),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_123),
.Y(n_129)
);

AOI22xp5_ASAP7_75t_L g118 ( 
.A1(n_90),
.A2(n_95),
.B1(n_103),
.B2(n_93),
.Y(n_118)
);

OAI22xp33_ASAP7_75t_SL g145 ( 
.A1(n_118),
.A2(n_71),
.B1(n_68),
.B2(n_73),
.Y(n_145)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_93),
.Y(n_119)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_92),
.Y(n_120)
);

INVxp67_ASAP7_75t_L g138 ( 
.A(n_120),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_SL g121 ( 
.A(n_95),
.B(n_61),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_121),
.B(n_122),
.Y(n_142)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_92),
.B(n_64),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_103),
.B(n_74),
.Y(n_123)
);

AOI21xp33_ASAP7_75t_L g128 ( 
.A1(n_109),
.A2(n_74),
.B(n_102),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_SL g147 ( 
.A(n_128),
.B(n_0),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_120),
.B(n_77),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g161 ( 
.A(n_130),
.B(n_137),
.Y(n_161)
);

XNOR2xp5_ASAP7_75t_L g133 ( 
.A(n_110),
.B(n_93),
.Y(n_133)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_133),
.B(n_79),
.C(n_67),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_106),
.Y(n_137)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_139),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g141 ( 
.A(n_110),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g148 ( 
.A(n_141),
.B(n_108),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_75),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_SL g166 ( 
.A(n_143),
.B(n_2),
.Y(n_166)
);

OAI21xp33_ASAP7_75t_L g144 ( 
.A1(n_105),
.A2(n_70),
.B(n_72),
.Y(n_144)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_144),
.A2(n_79),
.B(n_67),
.Y(n_152)
);

AOI22xp5_ASAP7_75t_L g170 ( 
.A1(n_145),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_170)
);

MAJx2_ASAP7_75t_L g146 ( 
.A(n_141),
.B(n_73),
.C(n_67),
.Y(n_146)
);

MAJIxp5_ASAP7_75t_L g174 ( 
.A(n_146),
.B(n_153),
.C(n_168),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_147),
.B(n_149),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_SL g176 ( 
.A(n_148),
.B(n_4),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_142),
.B(n_116),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_SL g150 ( 
.A1(n_138),
.A2(n_104),
.B(n_79),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g180 ( 
.A1(n_150),
.A2(n_6),
.B(n_7),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g151 ( 
.A1(n_127),
.A2(n_129),
.B1(n_124),
.B2(n_138),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g190 ( 
.A1(n_151),
.A2(n_9),
.B1(n_11),
.B2(n_12),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_158),
.Y(n_172)
);

CKINVDCx16_ASAP7_75t_R g154 ( 
.A(n_126),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_154),
.B(n_155),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g155 ( 
.A(n_144),
.B(n_1),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g156 ( 
.A(n_133),
.B(n_49),
.Y(n_156)
);

NAND2xp5_ASAP7_75t_L g171 ( 
.A(n_156),
.B(n_168),
.Y(n_171)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_125),
.Y(n_157)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_157),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_134),
.B(n_132),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g160 ( 
.A(n_140),
.B(n_1),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g189 ( 
.A(n_160),
.B(n_164),
.Y(n_189)
);

O2A1O1Ixp33_ASAP7_75t_SL g162 ( 
.A1(n_140),
.A2(n_48),
.B(n_47),
.C(n_45),
.Y(n_162)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_162),
.A2(n_27),
.B(n_7),
.Y(n_179)
);

AOI22xp5_ASAP7_75t_L g163 ( 
.A1(n_135),
.A2(n_44),
.B1(n_43),
.B2(n_41),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_L g177 ( 
.A1(n_163),
.A2(n_166),
.B1(n_170),
.B2(n_6),
.Y(n_177)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_131),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_131),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_3),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g187 ( 
.A(n_167),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_136),
.B(n_38),
.Y(n_168)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_136),
.Y(n_169)
);

INVxp33_ASAP7_75t_L g173 ( 
.A(n_169),
.Y(n_173)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_171),
.B(n_176),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g194 ( 
.A1(n_177),
.A2(n_179),
.B1(n_152),
.B2(n_162),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_150),
.A2(n_35),
.B(n_33),
.Y(n_178)
);

A2O1A1Ixp33_ASAP7_75t_SL g198 ( 
.A1(n_178),
.A2(n_188),
.B(n_12),
.C(n_13),
.Y(n_198)
);

CKINVDCx14_ASAP7_75t_R g193 ( 
.A(n_180),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_156),
.B(n_8),
.Y(n_181)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_181),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g182 ( 
.A(n_161),
.Y(n_182)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_182),
.Y(n_202)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_151),
.B(n_8),
.Y(n_185)
);

HB1xp67_ASAP7_75t_L g195 ( 
.A(n_185),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g186 ( 
.A(n_153),
.B(n_9),
.C(n_11),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g199 ( 
.A(n_186),
.B(n_13),
.C(n_14),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_157),
.A2(n_146),
.B(n_159),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_190),
.A2(n_17),
.B1(n_18),
.B2(n_19),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_185),
.A2(n_170),
.B1(n_169),
.B2(n_163),
.Y(n_192)
);

AOI22xp5_ASAP7_75t_L g211 ( 
.A1(n_192),
.A2(n_200),
.B1(n_203),
.B2(n_179),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g204 ( 
.A(n_194),
.B(n_198),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_199),
.B(n_180),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_L g200 ( 
.A1(n_190),
.A2(n_14),
.B1(n_15),
.B2(n_16),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_174),
.B(n_16),
.C(n_17),
.Y(n_201)
);

MAJIxp5_ASAP7_75t_L g206 ( 
.A(n_201),
.B(n_178),
.C(n_186),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_196),
.B(n_188),
.Y(n_205)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_205),
.B(n_206),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_207),
.B(n_208),
.Y(n_217)
);

AOI21xp5_ASAP7_75t_L g208 ( 
.A1(n_193),
.A2(n_172),
.B(n_202),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_195),
.B(n_175),
.Y(n_209)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_209),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_189),
.Y(n_210)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_210),
.A2(n_211),
.B1(n_193),
.B2(n_183),
.Y(n_215)
);

XOR2xp5_ASAP7_75t_L g212 ( 
.A(n_197),
.B(n_174),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_212),
.B(n_171),
.C(n_176),
.Y(n_218)
);

OAI22xp5_ASAP7_75t_L g222 ( 
.A1(n_215),
.A2(n_216),
.B1(n_198),
.B2(n_173),
.Y(n_222)
);

AOI22xp5_ASAP7_75t_L g216 ( 
.A1(n_204),
.A2(n_187),
.B1(n_184),
.B2(n_173),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_218),
.B(n_206),
.Y(n_220)
);

AOI22xp33_ASAP7_75t_SL g219 ( 
.A1(n_213),
.A2(n_198),
.B1(n_191),
.B2(n_205),
.Y(n_219)
);

OAI22xp5_ASAP7_75t_SL g224 ( 
.A1(n_219),
.A2(n_221),
.B1(n_222),
.B2(n_19),
.Y(n_224)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_220),
.B(n_214),
.C(n_218),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_217),
.A2(n_198),
.B1(n_212),
.B2(n_181),
.Y(n_221)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_223),
.A2(n_224),
.B(n_219),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_225),
.B(n_223),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_226),
.B(n_22),
.Y(n_227)
);

NAND2xp5_ASAP7_75t_SL g228 ( 
.A(n_227),
.B(n_20),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g229 ( 
.A(n_228),
.B(n_20),
.C(n_21),
.Y(n_229)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_229),
.B(n_22),
.Y(n_230)
);


endmodule