module fake_jpeg_1914_n_192 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_192);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_192;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_24;
wire n_44;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_91;
wire n_54;
wire n_93;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_189;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_1),
.Y(n_15)
);

BUFx12f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

BUFx2_ASAP7_75t_L g18 ( 
.A(n_6),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_5),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

INVx6_ASAP7_75t_L g21 ( 
.A(n_3),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_10),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_1),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_14),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_0),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_14),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_6),
.Y(n_32)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_6),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_18),
.Y(n_34)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_24),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_35),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_24),
.Y(n_36)
);

INVx6_ASAP7_75t_L g58 ( 
.A(n_36),
.Y(n_58)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_26),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_37),
.B(n_45),
.Y(n_54)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_18),
.Y(n_38)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_38),
.Y(n_77)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_24),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g74 ( 
.A(n_39),
.Y(n_74)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx11_ASAP7_75t_L g70 ( 
.A(n_40),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_41),
.Y(n_69)
);

INVx6_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_42),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_L g43 ( 
.A(n_20),
.B(n_0),
.C(n_2),
.Y(n_43)
);

AND2x2_ASAP7_75t_L g56 ( 
.A(n_43),
.B(n_47),
.Y(n_56)
);

BUFx3_ASAP7_75t_L g44 ( 
.A(n_18),
.Y(n_44)
);

NAND2xp33_ASAP7_75t_SL g61 ( 
.A(n_44),
.B(n_48),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_3),
.Y(n_45)
);

INVx5_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_46),
.Y(n_75)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_20),
.Y(n_47)
);

INVx2_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_26),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_49),
.B(n_51),
.Y(n_60)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_16),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_SL g57 ( 
.A(n_50),
.B(n_52),
.Y(n_57)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_18),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_16),
.Y(n_52)
);

CKINVDCx14_ASAP7_75t_SL g53 ( 
.A(n_34),
.Y(n_53)
);

BUFx2_ASAP7_75t_L g93 ( 
.A(n_53),
.Y(n_93)
);

NAND2x2_ASAP7_75t_SL g55 ( 
.A(n_43),
.B(n_29),
.Y(n_55)
);

A2O1A1Ixp33_ASAP7_75t_L g81 ( 
.A1(n_55),
.A2(n_29),
.B(n_25),
.C(n_23),
.Y(n_81)
);

OAI22xp33_ASAP7_75t_L g59 ( 
.A1(n_35),
.A2(n_21),
.B1(n_27),
.B2(n_33),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_L g90 ( 
.A1(n_59),
.A2(n_68),
.B1(n_25),
.B2(n_19),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_50),
.B(n_30),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_62),
.B(n_63),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_52),
.B(n_30),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_46),
.B(n_28),
.Y(n_64)
);

NOR2xp33_ASAP7_75t_L g101 ( 
.A(n_64),
.B(n_4),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_41),
.B(n_31),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_65),
.B(n_67),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_36),
.B(n_22),
.Y(n_67)
);

AOI22xp33_ASAP7_75t_L g68 ( 
.A1(n_39),
.A2(n_15),
.B1(n_19),
.B2(n_23),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g71 ( 
.A(n_38),
.B(n_22),
.Y(n_71)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_71),
.B(n_56),
.Y(n_86)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_44),
.A2(n_33),
.B1(n_27),
.B2(n_16),
.Y(n_72)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_72),
.A2(n_33),
.B1(n_27),
.B2(n_29),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_42),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g87 ( 
.A(n_76),
.B(n_78),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_SL g78 ( 
.A(n_40),
.B(n_15),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_40),
.A2(n_21),
.B1(n_17),
.B2(n_29),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_SL g91 ( 
.A1(n_79),
.A2(n_17),
.B1(n_32),
.B2(n_29),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_81),
.B(n_95),
.Y(n_126)
);

INVxp67_ASAP7_75t_L g115 ( 
.A(n_82),
.Y(n_115)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx1_ASAP7_75t_L g109 ( 
.A(n_83),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_56),
.B(n_32),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_SL g111 ( 
.A(n_85),
.B(n_76),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_86),
.B(n_102),
.Y(n_114)
);

BUFx12_ASAP7_75t_L g89 ( 
.A(n_70),
.Y(n_89)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_90),
.A2(n_91),
.B1(n_92),
.B2(n_100),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g92 ( 
.A1(n_79),
.A2(n_59),
.B1(n_55),
.B2(n_67),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g94 ( 
.A(n_56),
.B(n_3),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_94),
.B(n_105),
.Y(n_106)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_55),
.B(n_65),
.C(n_71),
.Y(n_95)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_60),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_96),
.B(n_101),
.Y(n_116)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_73),
.Y(n_97)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_97),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_66),
.Y(n_98)
);

INVx3_ASAP7_75t_L g108 ( 
.A(n_98),
.Y(n_108)
);

INVx1_ASAP7_75t_SL g99 ( 
.A(n_61),
.Y(n_99)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_99),
.Y(n_107)
);

AOI22xp33_ASAP7_75t_SL g100 ( 
.A1(n_55),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_57),
.Y(n_102)
);

INVxp67_ASAP7_75t_L g103 ( 
.A(n_75),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_80),
.Y(n_118)
);

OAI22x1_ASAP7_75t_SL g104 ( 
.A1(n_61),
.A2(n_4),
.B1(n_5),
.B2(n_7),
.Y(n_104)
);

AO21x1_ASAP7_75t_L g117 ( 
.A1(n_104),
.A2(n_75),
.B(n_9),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_54),
.B(n_7),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_111),
.B(n_117),
.Y(n_130)
);

OAI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_84),
.A2(n_69),
.B1(n_58),
.B2(n_66),
.Y(n_112)
);

AOI22xp5_ASAP7_75t_L g128 ( 
.A1(n_112),
.A2(n_113),
.B1(n_123),
.B2(n_81),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_84),
.A2(n_69),
.B1(n_58),
.B2(n_66),
.Y(n_113)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_118),
.Y(n_132)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_83),
.Y(n_119)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_119),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_95),
.B(n_80),
.Y(n_121)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_121),
.B(n_87),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g123 ( 
.A1(n_86),
.A2(n_74),
.B1(n_77),
.B2(n_70),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_96),
.B(n_77),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_124),
.B(n_93),
.Y(n_141)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_74),
.Y(n_125)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_125),
.B(n_104),
.C(n_97),
.Y(n_133)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_114),
.A2(n_99),
.B1(n_102),
.B2(n_91),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g145 ( 
.A1(n_127),
.A2(n_135),
.B1(n_123),
.B2(n_113),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_128),
.Y(n_146)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_107),
.A2(n_87),
.B(n_85),
.Y(n_129)
);

AOI21xp5_ASAP7_75t_L g155 ( 
.A1(n_129),
.A2(n_112),
.B(n_108),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g151 ( 
.A(n_131),
.B(n_133),
.Y(n_151)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_121),
.B(n_88),
.Y(n_134)
);

A2O1A1O1Ixp25_ASAP7_75t_L g149 ( 
.A1(n_134),
.A2(n_143),
.B(n_106),
.C(n_125),
.D(n_111),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g135 ( 
.A1(n_120),
.A2(n_98),
.B1(n_103),
.B2(n_93),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_109),
.Y(n_137)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_137),
.Y(n_152)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_109),
.Y(n_138)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_138),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_110),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_139),
.B(n_141),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g140 ( 
.A1(n_126),
.A2(n_105),
.B(n_93),
.Y(n_140)
);

OAI21xp5_ASAP7_75t_L g147 ( 
.A1(n_140),
.A2(n_142),
.B(n_117),
.Y(n_147)
);

OAI21xp33_ASAP7_75t_SL g142 ( 
.A1(n_115),
.A2(n_89),
.B(n_74),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g143 ( 
.A(n_126),
.B(n_98),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_141),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_144),
.B(n_148),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_139),
.B1(n_132),
.B2(n_130),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g160 ( 
.A(n_147),
.Y(n_160)
);

INVxp67_ASAP7_75t_L g148 ( 
.A(n_136),
.Y(n_148)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

OAI32xp33_ASAP7_75t_L g150 ( 
.A1(n_131),
.A2(n_117),
.A3(n_106),
.B1(n_115),
.B2(n_110),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g163 ( 
.A(n_150),
.Y(n_163)
);

AO221x1_ASAP7_75t_L g153 ( 
.A1(n_135),
.A2(n_122),
.B1(n_89),
.B2(n_116),
.C(n_119),
.Y(n_153)
);

INVxp67_ASAP7_75t_L g167 ( 
.A(n_153),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g158 ( 
.A1(n_155),
.A2(n_157),
.B1(n_128),
.B2(n_129),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_134),
.B(n_108),
.Y(n_157)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_158),
.B(n_162),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_151),
.B(n_143),
.C(n_140),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_166),
.C(n_147),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_146),
.A2(n_130),
.B1(n_132),
.B2(n_133),
.Y(n_164)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_164),
.Y(n_173)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_151),
.B(n_127),
.C(n_138),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g168 ( 
.A(n_159),
.B(n_146),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g175 ( 
.A(n_168),
.B(n_170),
.C(n_172),
.Y(n_175)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_169),
.B(n_167),
.Y(n_179)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_161),
.B(n_154),
.C(n_152),
.Y(n_170)
);

AOI21xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_156),
.B(n_155),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_171),
.A2(n_160),
.B1(n_167),
.B2(n_163),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g172 ( 
.A(n_166),
.B(n_150),
.Y(n_172)
);

NOR2xp67_ASAP7_75t_SL g176 ( 
.A(n_168),
.B(n_165),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g182 ( 
.A1(n_176),
.A2(n_177),
.B(n_174),
.Y(n_182)
);

AND2x2_ASAP7_75t_SL g178 ( 
.A(n_174),
.B(n_163),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_178),
.B(n_180),
.Y(n_181)
);

OAI21xp5_ASAP7_75t_L g183 ( 
.A1(n_179),
.A2(n_175),
.B(n_172),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_173),
.B(n_148),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_182),
.B(n_183),
.Y(n_187)
);

AOI22xp33_ASAP7_75t_L g184 ( 
.A1(n_178),
.A2(n_137),
.B1(n_149),
.B2(n_145),
.Y(n_184)
);

O2A1O1Ixp33_ASAP7_75t_SL g185 ( 
.A1(n_184),
.A2(n_178),
.B(n_175),
.C(n_136),
.Y(n_185)
);

OAI21xp5_ASAP7_75t_L g188 ( 
.A1(n_185),
.A2(n_186),
.B(n_8),
.Y(n_188)
);

AOI31xp67_ASAP7_75t_SL g186 ( 
.A1(n_181),
.A2(n_8),
.A3(n_9),
.B(n_10),
.Y(n_186)
);

OAI321xp33_ASAP7_75t_L g190 ( 
.A1(n_188),
.A2(n_189),
.A3(n_8),
.B1(n_10),
.B2(n_11),
.C(n_12),
.Y(n_190)
);

AOI21xp5_ASAP7_75t_SL g189 ( 
.A1(n_187),
.A2(n_89),
.B(n_9),
.Y(n_189)
);

OAI21xp5_ASAP7_75t_L g191 ( 
.A1(n_190),
.A2(n_12),
.B(n_74),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g192 ( 
.A(n_191),
.B(n_12),
.Y(n_192)
);


endmodule