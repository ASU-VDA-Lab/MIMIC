module fake_jpeg_23634_n_48 (n_3, n_2, n_1, n_0, n_4, n_6, n_5, n_48);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_6;
input n_5;

output n_48;

wire n_13;
wire n_21;
wire n_33;
wire n_45;
wire n_23;
wire n_10;
wire n_27;
wire n_22;
wire n_47;
wire n_14;
wire n_40;
wire n_19;
wire n_20;
wire n_18;
wire n_35;
wire n_46;
wire n_41;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_16;
wire n_24;
wire n_28;
wire n_38;
wire n_26;
wire n_44;
wire n_9;
wire n_36;
wire n_11;
wire n_17;
wire n_31;
wire n_25;
wire n_29;
wire n_37;
wire n_43;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

INVx1_ASAP7_75t_L g7 ( 
.A(n_4),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

CKINVDCx20_ASAP7_75t_R g10 ( 
.A(n_1),
.Y(n_10)
);

NOR2xp33_ASAP7_75t_L g11 ( 
.A(n_5),
.B(n_2),
.Y(n_11)
);

BUFx2_ASAP7_75t_L g12 ( 
.A(n_4),
.Y(n_12)
);

INVx11_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_2),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g30 ( 
.A(n_15),
.B(n_19),
.Y(n_30)
);

INVx8_ASAP7_75t_L g16 ( 
.A(n_12),
.Y(n_16)
);

INVx5_ASAP7_75t_L g25 ( 
.A(n_16),
.Y(n_25)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_SL g24 ( 
.A1(n_17),
.A2(n_20),
.B1(n_22),
.B2(n_9),
.Y(n_24)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_12),
.Y(n_18)
);

INVxp67_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_7),
.B(n_0),
.Y(n_19)
);

AOI22xp33_ASAP7_75t_SL g20 ( 
.A1(n_13),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_7),
.B(n_3),
.Y(n_21)
);

OAI21xp5_ASAP7_75t_SL g23 ( 
.A1(n_21),
.A2(n_7),
.B(n_9),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_L g22 ( 
.A1(n_8),
.A2(n_3),
.B1(n_5),
.B2(n_13),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_21),
.Y(n_32)
);

NAND2xp33_ASAP7_75t_SL g35 ( 
.A(n_24),
.B(n_20),
.Y(n_35)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_19),
.Y(n_26)
);

INVx1_ASAP7_75t_L g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g27 ( 
.A1(n_17),
.A2(n_8),
.B1(n_10),
.B2(n_14),
.Y(n_27)
);

XOR2xp5_ASAP7_75t_L g31 ( 
.A(n_27),
.B(n_22),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g29 ( 
.A1(n_19),
.A2(n_11),
.B(n_10),
.Y(n_29)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_29),
.A2(n_21),
.B(n_11),
.Y(n_36)
);

XNOR2xp5_ASAP7_75t_L g37 ( 
.A(n_31),
.B(n_32),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_30),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_SL g40 ( 
.A(n_34),
.B(n_14),
.Y(n_40)
);

MAJIxp5_ASAP7_75t_L g41 ( 
.A(n_35),
.B(n_24),
.C(n_27),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_9),
.Y(n_39)
);

MAJIxp5_ASAP7_75t_L g38 ( 
.A(n_31),
.B(n_15),
.C(n_29),
.Y(n_38)
);

OAI21xp5_ASAP7_75t_SL g45 ( 
.A1(n_38),
.A2(n_39),
.B(n_41),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_L g44 ( 
.A1(n_40),
.A2(n_8),
.B1(n_28),
.B2(n_16),
.Y(n_44)
);

OAI321xp33_ASAP7_75t_L g42 ( 
.A1(n_37),
.A2(n_32),
.A3(n_36),
.B1(n_33),
.B2(n_25),
.C(n_18),
.Y(n_42)
);

AOI21xp5_ASAP7_75t_L g47 ( 
.A1(n_42),
.A2(n_44),
.B(n_45),
.Y(n_47)
);

AOI322xp5_ASAP7_75t_L g43 ( 
.A1(n_38),
.A2(n_33),
.A3(n_16),
.B1(n_12),
.B2(n_15),
.C1(n_18),
.C2(n_25),
.Y(n_43)
);

MAJIxp5_ASAP7_75t_L g46 ( 
.A(n_43),
.B(n_16),
.C(n_28),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g48 ( 
.A(n_46),
.B(n_47),
.Y(n_48)
);


endmodule