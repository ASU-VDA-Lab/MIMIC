module fake_jpeg_4633_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_145;
wire n_20;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g16 ( 
.A(n_10),
.Y(n_16)
);

HB1xp67_ASAP7_75t_L g17 ( 
.A(n_1),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_8),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_14),
.Y(n_20)
);

INVx6_ASAP7_75t_SL g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_13),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_11),
.Y(n_24)
);

HB1xp67_ASAP7_75t_L g25 ( 
.A(n_14),
.Y(n_25)
);

INVx4_ASAP7_75t_L g26 ( 
.A(n_11),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_15),
.Y(n_27)
);

CKINVDCx16_ASAP7_75t_R g28 ( 
.A(n_6),
.Y(n_28)
);

INVx4_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_11),
.Y(n_31)
);

INVx8_ASAP7_75t_SL g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_15),
.Y(n_33)
);

INVxp67_ASAP7_75t_L g34 ( 
.A(n_0),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_25),
.B(n_14),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_35),
.B(n_38),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_32),
.Y(n_36)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_36),
.Y(n_56)
);

BUFx5_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

BUFx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

INVx1_ASAP7_75t_L g38 ( 
.A(n_21),
.Y(n_38)
);

BUFx2_ASAP7_75t_L g39 ( 
.A(n_21),
.Y(n_39)
);

INVx2_ASAP7_75t_L g53 ( 
.A(n_39),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_16),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_40),
.B(n_41),
.Y(n_55)
);

INVx8_ASAP7_75t_L g41 ( 
.A(n_21),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_22),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_42),
.B(n_43),
.Y(n_58)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_22),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_16),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_44),
.B(n_45),
.Y(n_64)
);

INVx2_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_17),
.Y(n_46)
);

INVx2_ASAP7_75t_SL g60 ( 
.A(n_46),
.Y(n_60)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g63 ( 
.A(n_47),
.B(n_24),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g48 ( 
.A(n_37),
.B(n_23),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_SL g72 ( 
.A(n_48),
.B(n_43),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_43),
.A2(n_19),
.B1(n_31),
.B2(n_34),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_50),
.A2(n_59),
.B1(n_67),
.B2(n_38),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g51 ( 
.A1(n_41),
.A2(n_19),
.B1(n_31),
.B2(n_29),
.Y(n_51)
);

AOI22xp33_ASAP7_75t_SL g91 ( 
.A1(n_51),
.A2(n_62),
.B1(n_65),
.B2(n_71),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_41),
.A2(n_29),
.B1(n_26),
.B2(n_31),
.Y(n_52)
);

A2O1A1Ixp33_ASAP7_75t_L g79 ( 
.A1(n_52),
.A2(n_70),
.B(n_35),
.C(n_39),
.Y(n_79)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_37),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_54),
.B(n_68),
.Y(n_83)
);

AND2x2_ASAP7_75t_SL g57 ( 
.A(n_37),
.B(n_19),
.Y(n_57)
);

AND2x2_ASAP7_75t_SL g76 ( 
.A(n_57),
.B(n_36),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_L g59 ( 
.A1(n_43),
.A2(n_31),
.B1(n_26),
.B2(n_29),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_41),
.A2(n_26),
.B1(n_28),
.B2(n_16),
.Y(n_62)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_63),
.B(n_66),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g65 ( 
.A1(n_41),
.A2(n_28),
.B1(n_24),
.B2(n_30),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g66 ( 
.A(n_45),
.B(n_23),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g67 ( 
.A1(n_45),
.A2(n_18),
.B1(n_30),
.B2(n_27),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_35),
.Y(n_68)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_39),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_69),
.B(n_36),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g70 ( 
.A1(n_46),
.A2(n_33),
.B1(n_27),
.B2(n_18),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_43),
.A2(n_24),
.B1(n_33),
.B2(n_23),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_72),
.B(n_74),
.Y(n_106)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

BUFx2_ASAP7_75t_L g132 ( 
.A(n_73),
.Y(n_132)
);

CKINVDCx14_ASAP7_75t_R g74 ( 
.A(n_55),
.Y(n_74)
);

BUFx3_ASAP7_75t_L g75 ( 
.A(n_57),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_75),
.B(n_77),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g110 ( 
.A(n_76),
.B(n_48),
.Y(n_110)
);

INVx2_ASAP7_75t_L g77 ( 
.A(n_61),
.Y(n_77)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_58),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_78),
.B(n_81),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_79),
.A2(n_88),
.B1(n_93),
.B2(n_104),
.Y(n_105)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_63),
.Y(n_81)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_63),
.Y(n_82)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_82),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g84 ( 
.A(n_55),
.Y(n_84)
);

HB1xp67_ASAP7_75t_L g107 ( 
.A(n_84),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g85 ( 
.A(n_68),
.B(n_44),
.Y(n_85)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_85),
.Y(n_115)
);

INVx4_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g114 ( 
.A(n_86),
.Y(n_114)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_67),
.Y(n_87)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_87),
.Y(n_119)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_89),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_64),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_L g112 ( 
.A1(n_90),
.A2(n_56),
.B1(n_46),
.B2(n_69),
.Y(n_112)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_64),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_92),
.Y(n_108)
);

OAI22xp33_ASAP7_75t_SL g93 ( 
.A1(n_57),
.A2(n_47),
.B1(n_38),
.B2(n_44),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g94 ( 
.A(n_56),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_94),
.Y(n_125)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_70),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_L g122 ( 
.A(n_95),
.B(n_96),
.Y(n_122)
);

AND2x2_ASAP7_75t_L g96 ( 
.A(n_66),
.B(n_48),
.Y(n_96)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_70),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_98),
.B(n_99),
.Y(n_126)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_58),
.Y(n_99)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_61),
.Y(n_100)
);

BUFx6f_ASAP7_75t_L g131 ( 
.A(n_100),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_66),
.B(n_47),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_101),
.B(n_103),
.Y(n_128)
);

AO22x1_ASAP7_75t_SL g102 ( 
.A1(n_50),
.A2(n_42),
.B1(n_36),
.B2(n_46),
.Y(n_102)
);

OAI22xp5_ASAP7_75t_SL g109 ( 
.A1(n_102),
.A2(n_59),
.B1(n_56),
.B2(n_50),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_49),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g104 ( 
.A(n_48),
.B(n_40),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_109),
.A2(n_118),
.B1(n_133),
.B2(n_72),
.Y(n_150)
);

XOR2xp5_ASAP7_75t_L g140 ( 
.A(n_110),
.B(n_120),
.Y(n_140)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_102),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_111),
.B(n_112),
.Y(n_157)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_87),
.A2(n_52),
.B1(n_51),
.B2(n_71),
.Y(n_118)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_73),
.B(n_52),
.C(n_54),
.Y(n_120)
);

AOI22xp33_ASAP7_75t_L g121 ( 
.A1(n_89),
.A2(n_95),
.B1(n_98),
.B2(n_102),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g160 ( 
.A1(n_121),
.A2(n_88),
.B1(n_91),
.B2(n_83),
.Y(n_160)
);

INVx2_ASAP7_75t_L g123 ( 
.A(n_102),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_123),
.B(n_127),
.Y(n_145)
);

INVx3_ASAP7_75t_L g127 ( 
.A(n_76),
.Y(n_127)
);

BUFx3_ASAP7_75t_L g129 ( 
.A(n_76),
.Y(n_129)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_129),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_79),
.A2(n_65),
.B1(n_68),
.B2(n_62),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g134 ( 
.A(n_110),
.B(n_76),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g178 ( 
.A(n_134),
.B(n_162),
.Y(n_178)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_128),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g167 ( 
.A(n_135),
.B(n_138),
.Y(n_167)
);

A2O1A1O1Ixp25_ASAP7_75t_L g136 ( 
.A1(n_106),
.A2(n_96),
.B(n_86),
.C(n_75),
.D(n_80),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_SL g172 ( 
.A(n_136),
.B(n_163),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_108),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_137),
.Y(n_173)
);

NAND3xp33_ASAP7_75t_SL g138 ( 
.A(n_119),
.B(n_103),
.C(n_82),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g139 ( 
.A1(n_122),
.A2(n_92),
.B(n_90),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g191 ( 
.A1(n_139),
.A2(n_144),
.B(n_39),
.Y(n_191)
);

CKINVDCx14_ASAP7_75t_R g141 ( 
.A(n_124),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_141),
.B(n_143),
.Y(n_175)
);

XOR2xp5_ASAP7_75t_L g142 ( 
.A(n_122),
.B(n_101),
.Y(n_142)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_142),
.B(n_115),
.C(n_114),
.Y(n_176)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_128),
.Y(n_143)
);

OAI21xp5_ASAP7_75t_SL g144 ( 
.A1(n_126),
.A2(n_75),
.B(n_81),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_108),
.Y(n_146)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_146),
.Y(n_193)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_107),
.B(n_74),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g180 ( 
.A(n_147),
.Y(n_180)
);

AOI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_126),
.A2(n_80),
.B(n_96),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_148),
.A2(n_164),
.B(n_77),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g149 ( 
.A(n_116),
.B(n_84),
.Y(n_149)
);

CKINVDCx16_ASAP7_75t_R g197 ( 
.A(n_149),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_150),
.A2(n_161),
.B1(n_127),
.B2(n_111),
.Y(n_169)
);

OR2x2_ASAP7_75t_L g151 ( 
.A(n_119),
.B(n_104),
.Y(n_151)
);

OAI21xp5_ASAP7_75t_L g195 ( 
.A1(n_151),
.A2(n_60),
.B(n_61),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g152 ( 
.A(n_125),
.Y(n_152)
);

NOR3xp33_ASAP7_75t_L g192 ( 
.A(n_152),
.B(n_165),
.C(n_131),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_116),
.B(n_99),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_SL g179 ( 
.A(n_153),
.B(n_158),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_113),
.B(n_80),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g189 ( 
.A(n_154),
.B(n_159),
.Y(n_189)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_132),
.Y(n_156)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_156),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_130),
.B(n_85),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_113),
.B(n_83),
.Y(n_159)
);

AOI22xp5_ASAP7_75t_L g171 ( 
.A1(n_160),
.A2(n_118),
.B1(n_105),
.B2(n_109),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_48),
.B1(n_104),
.B2(n_56),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_129),
.B(n_49),
.Y(n_162)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_117),
.Y(n_163)
);

AOI21xp5_ASAP7_75t_L g164 ( 
.A1(n_120),
.A2(n_53),
.B(n_69),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_125),
.Y(n_165)
);

INVxp67_ASAP7_75t_L g166 ( 
.A(n_164),
.Y(n_166)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_166),
.B(n_170),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g201 ( 
.A1(n_169),
.A2(n_181),
.B1(n_183),
.B2(n_190),
.Y(n_201)
);

INVxp67_ASAP7_75t_L g170 ( 
.A(n_145),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_171),
.A2(n_174),
.B1(n_184),
.B2(n_185),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g174 ( 
.A1(n_145),
.A2(n_130),
.B1(n_114),
.B2(n_132),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_176),
.B(n_177),
.C(n_182),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_140),
.B(n_114),
.C(n_132),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g181 ( 
.A1(n_150),
.A2(n_115),
.B1(n_53),
.B2(n_97),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_140),
.B(n_54),
.C(n_53),
.Y(n_182)
);

OA22x2_ASAP7_75t_L g183 ( 
.A1(n_161),
.A2(n_94),
.B1(n_36),
.B2(n_60),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g184 ( 
.A1(n_160),
.A2(n_60),
.B1(n_94),
.B2(n_100),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_L g185 ( 
.A1(n_156),
.A2(n_155),
.B1(n_139),
.B2(n_163),
.Y(n_185)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_151),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_186),
.B(n_165),
.Y(n_209)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_188),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_134),
.B(n_39),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g190 ( 
.A1(n_157),
.A2(n_42),
.B1(n_40),
.B2(n_60),
.Y(n_190)
);

OAI22xp5_ASAP7_75t_L g219 ( 
.A1(n_191),
.A2(n_198),
.B1(n_199),
.B2(n_153),
.Y(n_219)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_192),
.Y(n_210)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_148),
.A2(n_61),
.B(n_60),
.Y(n_194)
);

XOR2xp5_ASAP7_75t_L g207 ( 
.A(n_194),
.B(n_144),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_195),
.B(n_149),
.Y(n_203)
);

NAND2x1_ASAP7_75t_SL g196 ( 
.A(n_151),
.B(n_155),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g202 ( 
.A(n_196),
.B(n_200),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_135),
.A2(n_42),
.B1(n_22),
.B2(n_23),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_143),
.A2(n_154),
.B1(n_162),
.B2(n_136),
.Y(n_199)
);

OR2x2_ASAP7_75t_L g200 ( 
.A(n_137),
.B(n_22),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g253 ( 
.A1(n_203),
.A2(n_0),
.B(n_2),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g205 ( 
.A(n_199),
.B(n_142),
.Y(n_205)
);

MAJIxp5_ASAP7_75t_L g233 ( 
.A(n_205),
.B(n_224),
.C(n_228),
.Y(n_233)
);

BUFx24_ASAP7_75t_SL g206 ( 
.A(n_175),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g238 ( 
.A(n_206),
.B(n_213),
.Y(n_238)
);

XOR2xp5_ASAP7_75t_L g245 ( 
.A(n_207),
.B(n_188),
.Y(n_245)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_209),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_189),
.B(n_159),
.Y(n_212)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_212),
.Y(n_252)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_174),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_167),
.B(n_146),
.Y(n_214)
);

CKINVDCx16_ASAP7_75t_R g230 ( 
.A(n_214),
.Y(n_230)
);

XOR2x1_ASAP7_75t_L g215 ( 
.A(n_196),
.B(n_158),
.Y(n_215)
);

XNOR2xp5_ASAP7_75t_SL g240 ( 
.A(n_215),
.B(n_187),
.Y(n_240)
);

INVx1_ASAP7_75t_L g217 ( 
.A(n_198),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_217),
.B(n_222),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_179),
.B(n_147),
.Y(n_218)
);

CKINVDCx20_ASAP7_75t_R g254 ( 
.A(n_218),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_219),
.A2(n_166),
.B1(n_183),
.B2(n_195),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g220 ( 
.A1(n_169),
.A2(n_152),
.B1(n_42),
.B2(n_131),
.Y(n_220)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_220),
.A2(n_221),
.B1(n_0),
.B2(n_3),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_181),
.A2(n_131),
.B1(n_23),
.B2(n_20),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_189),
.B(n_23),
.Y(n_222)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_179),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g239 ( 
.A(n_223),
.B(n_225),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g224 ( 
.A(n_178),
.B(n_20),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_173),
.B(n_13),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_173),
.B(n_13),
.Y(n_226)
);

NAND3xp33_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_12),
.C(n_10),
.Y(n_244)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g237 ( 
.A1(n_227),
.A2(n_229),
.B(n_194),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_182),
.B(n_20),
.C(n_1),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g229 ( 
.A(n_184),
.Y(n_229)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_215),
.A2(n_196),
.B(n_183),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_232),
.B(n_249),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_170),
.B1(n_191),
.B2(n_186),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_L g263 ( 
.A1(n_234),
.A2(n_242),
.B1(n_243),
.B2(n_246),
.Y(n_263)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_235),
.Y(n_266)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_208),
.A2(n_172),
.B1(n_183),
.B2(n_193),
.Y(n_236)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_236),
.Y(n_273)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_237),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g258 ( 
.A(n_240),
.B(n_247),
.Y(n_258)
);

OAI22xp5_ASAP7_75t_L g242 ( 
.A1(n_229),
.A2(n_193),
.B1(n_171),
.B2(n_197),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_L g243 ( 
.A1(n_201),
.A2(n_180),
.B1(n_177),
.B2(n_200),
.Y(n_243)
);

MAJIxp5_ASAP7_75t_SL g256 ( 
.A(n_244),
.B(n_247),
.C(n_222),
.Y(n_256)
);

XOR2xp5_ASAP7_75t_L g262 ( 
.A(n_245),
.B(n_204),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_176),
.B1(n_178),
.B2(n_168),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_SL g247 ( 
.A(n_205),
.B(n_20),
.Y(n_247)
);

AOI22xp5_ASAP7_75t_L g248 ( 
.A1(n_202),
.A2(n_227),
.B1(n_211),
.B2(n_203),
.Y(n_248)
);

CKINVDCx20_ASAP7_75t_R g259 ( 
.A(n_248),
.Y(n_259)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_202),
.A2(n_168),
.B1(n_20),
.B2(n_2),
.Y(n_249)
);

AO21x1_ASAP7_75t_L g250 ( 
.A1(n_202),
.A2(n_20),
.B(n_1),
.Y(n_250)
);

OA21x2_ASAP7_75t_L g269 ( 
.A1(n_250),
.A2(n_3),
.B(n_4),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g251 ( 
.A1(n_201),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g276 ( 
.A(n_251),
.B(n_253),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_255),
.B(n_223),
.Y(n_257)
);

OAI21xp33_ASAP7_75t_L g291 ( 
.A1(n_256),
.A2(n_9),
.B(n_12),
.Y(n_291)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_257),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_258),
.B(n_268),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_233),
.B(n_216),
.C(n_224),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_260),
.B(n_262),
.C(n_264),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g264 ( 
.A(n_245),
.B(n_204),
.Y(n_264)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_233),
.B(n_216),
.C(n_207),
.Y(n_265)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_267),
.C(n_270),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_240),
.B(n_228),
.C(n_212),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_248),
.B(n_221),
.Y(n_268)
);

OAI22xp33_ASAP7_75t_SL g277 ( 
.A1(n_269),
.A2(n_254),
.B1(n_250),
.B2(n_232),
.Y(n_277)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_243),
.B(n_12),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g271 ( 
.A(n_230),
.B(n_3),
.Y(n_271)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_271),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g272 ( 
.A(n_235),
.B(n_3),
.C(n_4),
.Y(n_272)
);

NOR2xp33_ASAP7_75t_L g292 ( 
.A(n_272),
.B(n_5),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_241),
.B(n_4),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_274),
.B(n_5),
.Y(n_290)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_277),
.Y(n_301)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_266),
.A2(n_236),
.B1(n_252),
.B2(n_251),
.Y(n_278)
);

INVx1_ASAP7_75t_L g303 ( 
.A(n_278),
.Y(n_303)
);

AOI22xp5_ASAP7_75t_L g279 ( 
.A1(n_275),
.A2(n_241),
.B1(n_252),
.B2(n_231),
.Y(n_279)
);

OAI22xp5_ASAP7_75t_L g302 ( 
.A1(n_279),
.A2(n_285),
.B1(n_287),
.B2(n_269),
.Y(n_302)
);

INVxp33_ASAP7_75t_L g281 ( 
.A(n_261),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_281),
.B(n_289),
.Y(n_296)
);

AOI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_273),
.A2(n_254),
.B1(n_237),
.B2(n_249),
.Y(n_284)
);

CKINVDCx14_ASAP7_75t_R g294 ( 
.A(n_284),
.Y(n_294)
);

AOI22xp5_ASAP7_75t_L g285 ( 
.A1(n_259),
.A2(n_231),
.B1(n_255),
.B2(n_253),
.Y(n_285)
);

AOI22xp5_ASAP7_75t_L g287 ( 
.A1(n_268),
.A2(n_239),
.B1(n_238),
.B2(n_7),
.Y(n_287)
);

OAI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_263),
.A2(n_239),
.B1(n_9),
.B2(n_10),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_290),
.B(n_292),
.Y(n_299)
);

NOR2xp33_ASAP7_75t_L g306 ( 
.A(n_291),
.B(n_293),
.Y(n_306)
);

INVxp67_ASAP7_75t_SL g293 ( 
.A(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_280),
.B(n_276),
.Y(n_295)
);

AOI21xp5_ASAP7_75t_L g310 ( 
.A1(n_295),
.A2(n_278),
.B(n_288),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g297 ( 
.A(n_282),
.B(n_260),
.C(n_265),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g319 ( 
.A(n_297),
.B(n_298),
.C(n_300),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_282),
.B(n_286),
.C(n_262),
.Y(n_298)
);

MAJIxp5_ASAP7_75t_L g300 ( 
.A(n_286),
.B(n_264),
.C(n_267),
.Y(n_300)
);

INVx1_ASAP7_75t_L g314 ( 
.A(n_302),
.Y(n_314)
);

MAJIxp5_ASAP7_75t_L g304 ( 
.A(n_279),
.B(n_270),
.C(n_258),
.Y(n_304)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_304),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g305 ( 
.A(n_283),
.B(n_269),
.Y(n_305)
);

XNOR2xp5_ASAP7_75t_L g312 ( 
.A(n_305),
.B(n_283),
.Y(n_312)
);

HB1xp67_ASAP7_75t_L g307 ( 
.A(n_281),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_307),
.B(n_287),
.Y(n_308)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_308),
.Y(n_327)
);

NOR2xp67_ASAP7_75t_L g309 ( 
.A(n_305),
.B(n_304),
.Y(n_309)
);

OAI22xp33_ASAP7_75t_SL g323 ( 
.A1(n_309),
.A2(n_318),
.B1(n_297),
.B2(n_298),
.Y(n_323)
);

AOI21xp5_ASAP7_75t_L g326 ( 
.A1(n_310),
.A2(n_315),
.B(n_6),
.Y(n_326)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_301),
.B(n_285),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g320 ( 
.A(n_311),
.B(n_313),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g322 ( 
.A(n_312),
.B(n_300),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_L g313 ( 
.A(n_303),
.B(n_284),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_295),
.B(n_5),
.Y(n_315)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_296),
.B(n_9),
.Y(n_317)
);

OAI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_317),
.A2(n_299),
.B(n_306),
.Y(n_321)
);

INVx11_ASAP7_75t_L g318 ( 
.A(n_294),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_321),
.B(n_324),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_SL g333 ( 
.A(n_322),
.B(n_325),
.Y(n_333)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_323),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_315),
.B(n_6),
.Y(n_324)
);

INVxp67_ASAP7_75t_L g325 ( 
.A(n_310),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_326),
.B(n_328),
.Y(n_329)
);

NOR2xp33_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_6),
.Y(n_328)
);

OR2x2_ASAP7_75t_L g331 ( 
.A(n_320),
.B(n_314),
.Y(n_331)
);

NOR3xp33_ASAP7_75t_L g337 ( 
.A(n_331),
.B(n_326),
.C(n_7),
.Y(n_337)
);

A2O1A1Ixp33_ASAP7_75t_SL g332 ( 
.A1(n_325),
.A2(n_316),
.B(n_312),
.C(n_319),
.Y(n_332)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_332),
.Y(n_336)
);

OAI21xp5_ASAP7_75t_SL g335 ( 
.A1(n_333),
.A2(n_319),
.B(n_327),
.Y(n_335)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_335),
.B(n_337),
.Y(n_338)
);

AOI21x1_ASAP7_75t_L g339 ( 
.A1(n_338),
.A2(n_330),
.B(n_336),
.Y(n_339)
);

AOI221xp5_ASAP7_75t_L g340 ( 
.A1(n_339),
.A2(n_329),
.B1(n_334),
.B2(n_7),
.C(n_8),
.Y(n_340)
);

INVx1_ASAP7_75t_L g341 ( 
.A(n_340),
.Y(n_341)
);

XNOR2xp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_7),
.Y(n_342)
);


endmodule