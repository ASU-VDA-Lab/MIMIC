module fake_jpeg_3996_n_189 (n_13, n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_189);

input n_13;
input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_189;

wire n_159;
wire n_117;
wire n_144;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_14;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_178;
wire n_166;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_31;
wire n_155;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_177;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_131;
wire n_56;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_161;
wire n_22;
wire n_138;
wire n_101;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_86;
wire n_156;
wire n_115;
wire n_123;
wire n_176;
wire n_112;
wire n_95;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_135;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_140;
wire n_128;
wire n_82;
wire n_96;

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_13),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_13),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_11),
.Y(n_16)
);

INVx2_ASAP7_75t_SL g17 ( 
.A(n_6),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_8),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_6),
.Y(n_20)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_11),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_1),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_4),
.Y(n_24)
);

BUFx6f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx5_ASAP7_75t_L g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_4),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_17),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g51 ( 
.A(n_32),
.B(n_33),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_17),
.B(n_0),
.Y(n_33)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_23),
.Y(n_34)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_34),
.Y(n_74)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_30),
.Y(n_35)
);

INVx8_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

BUFx3_ASAP7_75t_L g36 ( 
.A(n_14),
.Y(n_36)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_36),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_17),
.B(n_0),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g58 ( 
.A(n_37),
.B(n_39),
.Y(n_58)
);

BUFx3_ASAP7_75t_L g38 ( 
.A(n_14),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_38),
.B(n_44),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_19),
.B(n_1),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_15),
.B(n_1),
.Y(n_40)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_40),
.B(n_29),
.Y(n_62)
);

BUFx12f_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g56 ( 
.A(n_41),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_28),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_42),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g43 ( 
.A(n_28),
.Y(n_43)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_43),
.Y(n_66)
);

INVx2_ASAP7_75t_SL g44 ( 
.A(n_28),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_14),
.Y(n_45)
);

INVx5_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

INVx8_ASAP7_75t_L g46 ( 
.A(n_16),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_25),
.Y(n_61)
);

BUFx2_ASAP7_75t_L g47 ( 
.A(n_36),
.Y(n_47)
);

INVx3_ASAP7_75t_L g103 ( 
.A(n_47),
.Y(n_103)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_38),
.Y(n_49)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_49),
.B(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_19),
.Y(n_54)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_54),
.B(n_57),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g55 ( 
.A(n_45),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g82 ( 
.A(n_55),
.Y(n_82)
);

NAND2x1_ASAP7_75t_SL g57 ( 
.A(n_32),
.B(n_21),
.Y(n_57)
);

INVx2_ASAP7_75t_L g59 ( 
.A(n_46),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_59),
.B(n_60),
.Y(n_93)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_33),
.Y(n_60)
);

CKINVDCx14_ASAP7_75t_R g95 ( 
.A(n_61),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g102 ( 
.A(n_62),
.B(n_12),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_34),
.A2(n_20),
.B1(n_27),
.B2(n_18),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_SL g88 ( 
.A1(n_63),
.A2(n_77),
.B1(n_3),
.B2(n_5),
.Y(n_88)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_37),
.B(n_29),
.Y(n_67)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_67),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_42),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_68),
.B(n_41),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_46),
.A2(n_18),
.B1(n_27),
.B2(n_20),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_69),
.A2(n_71),
.B1(n_2),
.B2(n_3),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_44),
.B(n_21),
.Y(n_70)
);

INVx1_ASAP7_75t_L g91 ( 
.A(n_70),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_35),
.A2(n_31),
.B1(n_26),
.B2(n_24),
.Y(n_71)
);

MAJIxp5_ASAP7_75t_L g72 ( 
.A(n_42),
.B(n_15),
.C(n_31),
.Y(n_72)
);

MAJIxp5_ASAP7_75t_L g83 ( 
.A(n_72),
.B(n_25),
.C(n_16),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_42),
.B(n_26),
.Y(n_73)
);

AND2x2_ASAP7_75t_L g99 ( 
.A(n_73),
.B(n_76),
.Y(n_99)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_44),
.B(n_22),
.Y(n_75)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_75),
.Y(n_92)
);

OR2x2_ASAP7_75t_L g76 ( 
.A(n_43),
.B(n_24),
.Y(n_76)
);

OAI22xp5_ASAP7_75t_SL g77 ( 
.A1(n_43),
.A2(n_22),
.B1(n_23),
.B2(n_25),
.Y(n_77)
);

NAND2x1_ASAP7_75t_SL g78 ( 
.A(n_43),
.B(n_28),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_SL g85 ( 
.A1(n_78),
.A2(n_16),
.B1(n_23),
.B2(n_41),
.Y(n_85)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_41),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_79),
.B(n_5),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_81),
.B(n_90),
.Y(n_111)
);

AND2x2_ASAP7_75t_L g126 ( 
.A(n_83),
.B(n_88),
.Y(n_126)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_85),
.A2(n_78),
.B(n_57),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_SL g118 ( 
.A(n_86),
.B(n_77),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_73),
.B(n_2),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g113 ( 
.A(n_87),
.B(n_89),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_60),
.B(n_3),
.Y(n_89)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_50),
.Y(n_90)
);

INVx4_ASAP7_75t_L g94 ( 
.A(n_50),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_94),
.B(n_104),
.Y(n_124)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_96),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_56),
.B(n_6),
.Y(n_97)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_97),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_58),
.B(n_7),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g114 ( 
.A(n_100),
.B(n_102),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_63),
.A2(n_7),
.B1(n_9),
.B2(n_10),
.Y(n_101)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_101),
.B(n_54),
.Y(n_108)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_53),
.Y(n_104)
);

BUFx24_ASAP7_75t_SL g105 ( 
.A(n_84),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_105),
.B(n_106),
.Y(n_136)
);

CKINVDCx12_ASAP7_75t_R g106 ( 
.A(n_104),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_L g128 ( 
.A1(n_107),
.A2(n_108),
.B1(n_118),
.B2(n_100),
.Y(n_128)
);

INVxp67_ASAP7_75t_L g109 ( 
.A(n_80),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g129 ( 
.A(n_109),
.B(n_119),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g112 ( 
.A(n_87),
.B(n_72),
.Y(n_112)
);

XOR2xp5_ASAP7_75t_L g137 ( 
.A(n_112),
.B(n_125),
.Y(n_137)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_93),
.Y(n_115)
);

CKINVDCx20_ASAP7_75t_R g139 ( 
.A(n_115),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_88),
.B(n_76),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_117),
.B(n_122),
.Y(n_131)
);

INVxp67_ASAP7_75t_L g119 ( 
.A(n_81),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_89),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_120),
.B(n_108),
.Y(n_140)
);

AND2x6_ASAP7_75t_L g121 ( 
.A(n_99),
.B(n_68),
.Y(n_121)
);

NOR3xp33_ASAP7_75t_SL g135 ( 
.A(n_121),
.B(n_92),
.C(n_91),
.Y(n_135)
);

OAI21xp5_ASAP7_75t_L g122 ( 
.A1(n_99),
.A2(n_51),
.B(n_66),
.Y(n_122)
);

OR2x4_ASAP7_75t_L g123 ( 
.A(n_99),
.B(n_48),
.Y(n_123)
);

OAI21xp5_ASAP7_75t_L g142 ( 
.A1(n_123),
.A2(n_56),
.B(n_64),
.Y(n_142)
);

XOR2xp5_ASAP7_75t_L g125 ( 
.A(n_98),
.B(n_66),
.Y(n_125)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_121),
.A2(n_85),
.B1(n_95),
.B2(n_59),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g145 ( 
.A(n_127),
.B(n_132),
.Y(n_145)
);

NOR3xp33_ASAP7_75t_L g154 ( 
.A(n_128),
.B(n_116),
.C(n_110),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_113),
.B(n_98),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_143),
.Y(n_152)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_124),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_118),
.A2(n_92),
.B1(n_101),
.B2(n_91),
.Y(n_133)
);

NAND2xp5_ASAP7_75t_SL g146 ( 
.A(n_133),
.B(n_144),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_126),
.A2(n_98),
.B1(n_83),
.B2(n_74),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_134),
.B(n_135),
.Y(n_153)
);

CKINVDCx16_ASAP7_75t_R g138 ( 
.A(n_111),
.Y(n_138)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_138),
.B(n_141),
.Y(n_157)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_140),
.Y(n_147)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_123),
.Y(n_141)
);

AO21x1_ASAP7_75t_L g148 ( 
.A1(n_142),
.A2(n_119),
.B(n_125),
.Y(n_148)
);

OAI32xp33_ASAP7_75t_L g143 ( 
.A1(n_126),
.A2(n_82),
.A3(n_84),
.B1(n_48),
.B2(n_52),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_122),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_148),
.B(n_154),
.Y(n_164)
);

INVx1_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx1_ASAP7_75t_L g161 ( 
.A(n_149),
.Y(n_161)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_137),
.B(n_112),
.C(n_64),
.Y(n_150)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_150),
.B(n_151),
.C(n_131),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g151 ( 
.A(n_137),
.B(n_126),
.C(n_117),
.Y(n_151)
);

A2O1A1O1Ixp25_ASAP7_75t_L g155 ( 
.A1(n_142),
.A2(n_109),
.B(n_114),
.C(n_79),
.D(n_49),
.Y(n_155)
);

A2O1A1O1Ixp25_ASAP7_75t_L g160 ( 
.A1(n_155),
.A2(n_156),
.B(n_143),
.C(n_127),
.D(n_141),
.Y(n_160)
);

NOR3xp33_ASAP7_75t_SL g156 ( 
.A(n_135),
.B(n_103),
.C(n_65),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g158 ( 
.A(n_157),
.Y(n_158)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_158),
.B(n_166),
.Y(n_171)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_150),
.B(n_131),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_159),
.B(n_163),
.C(n_162),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g170 ( 
.A1(n_160),
.A2(n_136),
.B(n_47),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_152),
.A2(n_144),
.B1(n_134),
.B2(n_130),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_162),
.Y(n_173)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_145),
.A2(n_152),
.B1(n_146),
.B2(n_153),
.Y(n_165)
);

CKINVDCx20_ASAP7_75t_R g175 ( 
.A(n_165),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g166 ( 
.A1(n_156),
.A2(n_148),
.B1(n_151),
.B2(n_155),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_147),
.A2(n_139),
.B1(n_132),
.B2(n_65),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g174 ( 
.A(n_167),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g168 ( 
.A1(n_145),
.A2(n_74),
.B1(n_103),
.B2(n_94),
.Y(n_168)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_168),
.B(n_7),
.C(n_9),
.Y(n_172)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_169),
.B(n_170),
.C(n_163),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g176 ( 
.A(n_172),
.B(n_164),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g183 ( 
.A(n_176),
.B(n_178),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_177),
.B(n_159),
.Y(n_182)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_173),
.B(n_161),
.Y(n_178)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_175),
.B(n_168),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g184 ( 
.A(n_179),
.B(n_180),
.Y(n_184)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_171),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_174),
.B(n_164),
.Y(n_181)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_182),
.B(n_166),
.C(n_181),
.Y(n_185)
);

NOR2xp33_ASAP7_75t_SL g188 ( 
.A(n_185),
.B(n_182),
.Y(n_188)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_184),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_SL g187 ( 
.A1(n_186),
.A2(n_183),
.B(n_160),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_187),
.B(n_188),
.Y(n_189)
);


endmodule