module fake_jpeg_20575_n_20 (n_3, n_2, n_1, n_0, n_4, n_20);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;

output n_20;

wire n_13;
wire n_10;
wire n_6;
wire n_14;
wire n_19;
wire n_18;
wire n_16;
wire n_9;
wire n_5;
wire n_11;
wire n_17;
wire n_12;
wire n_8;
wire n_15;
wire n_7;

INVx2_ASAP7_75t_L g5 ( 
.A(n_0),
.Y(n_5)
);

NAND2xp5_ASAP7_75t_L g6 ( 
.A(n_3),
.B(n_4),
.Y(n_6)
);

NAND2xp5_ASAP7_75t_L g7 ( 
.A(n_4),
.B(n_1),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_0),
.Y(n_8)
);

INVx1_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

NAND2xp5_ASAP7_75t_SL g13 ( 
.A(n_9),
.B(n_10),
.Y(n_13)
);

INVx3_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

AOI221xp5_ASAP7_75t_L g11 ( 
.A1(n_6),
.A2(n_2),
.B1(n_3),
.B2(n_0),
.C(n_1),
.Y(n_11)
);

NAND2xp5_ASAP7_75t_SL g16 ( 
.A(n_11),
.B(n_12),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g12 ( 
.A(n_7),
.B(n_1),
.Y(n_12)
);

OAI22xp5_ASAP7_75t_L g14 ( 
.A1(n_9),
.A2(n_5),
.B1(n_6),
.B2(n_8),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g18 ( 
.A(n_14),
.B(n_15),
.Y(n_18)
);

OAI22xp5_ASAP7_75t_L g15 ( 
.A1(n_12),
.A2(n_2),
.B1(n_8),
.B2(n_10),
.Y(n_15)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_13),
.Y(n_17)
);

AOI22xp33_ASAP7_75t_L g19 ( 
.A1(n_17),
.A2(n_14),
.B1(n_16),
.B2(n_18),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_SL g20 ( 
.A(n_19),
.B(n_17),
.Y(n_20)
);


endmodule