module real_jpeg_25192_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_38;
wire n_35;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_247;
wire n_146;
wire n_78;
wire n_83;
wire n_249;
wire n_166;
wire n_176;
wire n_221;
wire n_215;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_255;
wire n_243;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_200;
wire n_48;
wire n_164;
wire n_184;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_178;
wire n_67;
wire n_79;
wire n_238;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_222;
wire n_19;
wire n_148;
wire n_262;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_159;
wire n_72;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_192;
wire n_203;
wire n_100;
wire n_198;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_110;
wire n_61;
wire n_195;
wire n_258;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_228;
wire n_150;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_259;
wire n_225;
wire n_232;
wire n_43;
wire n_57;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_185;
wire n_125;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_97;
wire n_75;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_167;
wire n_202;
wire n_179;
wire n_213;
wire n_216;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_256;
wire n_182;
wire n_269;
wire n_96;
wire n_253;
wire n_89;

INVx3_ASAP7_75t_L g68 ( 
.A(n_0),
.Y(n_68)
);

INVx6_ASAP7_75t_L g73 ( 
.A(n_0),
.Y(n_73)
);

INVx6_ASAP7_75t_L g121 ( 
.A(n_0),
.Y(n_121)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_0),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g233 ( 
.A1(n_0),
.A2(n_117),
.B1(n_234),
.B2(n_236),
.Y(n_233)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_1),
.Y(n_40)
);

OAI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_2),
.A2(n_38),
.B1(n_41),
.B2(n_56),
.Y(n_55)
);

CKINVDCx16_ASAP7_75t_R g56 ( 
.A(n_2),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_L g100 ( 
.A1(n_2),
.A2(n_30),
.B1(n_56),
.B2(n_101),
.Y(n_100)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_2),
.A2(n_49),
.B1(n_50),
.B2(n_56),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g192 ( 
.A1(n_2),
.A2(n_56),
.B1(n_65),
.B2(n_66),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_3),
.A2(n_65),
.B1(n_66),
.B2(n_88),
.Y(n_87)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_3),
.Y(n_88)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_4),
.A2(n_65),
.B1(n_66),
.B2(n_70),
.Y(n_69)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_4),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_4),
.A2(n_49),
.B1(n_50),
.B2(n_70),
.Y(n_127)
);

BUFx12f_ASAP7_75t_L g79 ( 
.A(n_5),
.Y(n_79)
);

BUFx10_ASAP7_75t_L g65 ( 
.A(n_6),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g26 ( 
.A1(n_7),
.A2(n_27),
.B1(n_28),
.B2(n_30),
.Y(n_26)
);

CKINVDCx16_ASAP7_75t_R g27 ( 
.A(n_7),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_L g153 ( 
.A1(n_7),
.A2(n_27),
.B1(n_38),
.B2(n_41),
.Y(n_153)
);

AOI22xp33_ASAP7_75t_L g195 ( 
.A1(n_7),
.A2(n_27),
.B1(n_49),
.B2(n_50),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_7),
.A2(n_27),
.B1(n_65),
.B2(n_66),
.Y(n_235)
);

BUFx10_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_9),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_9),
.B(n_37),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_9),
.B(n_50),
.C(n_52),
.Y(n_185)
);

AOI22xp33_ASAP7_75t_L g199 ( 
.A1(n_9),
.A2(n_38),
.B1(n_41),
.B2(n_111),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_9),
.B(n_106),
.Y(n_217)
);

AOI22xp33_ASAP7_75t_L g228 ( 
.A1(n_9),
.A2(n_49),
.B1(n_50),
.B2(n_111),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g230 ( 
.A(n_9),
.B(n_65),
.C(n_78),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_L g248 ( 
.A1(n_9),
.A2(n_67),
.B(n_222),
.Y(n_248)
);

AOI22xp33_ASAP7_75t_SL g83 ( 
.A1(n_10),
.A2(n_49),
.B1(n_50),
.B2(n_84),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_10),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_10),
.A2(n_65),
.B1(n_66),
.B2(n_84),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g135 ( 
.A1(n_10),
.A2(n_38),
.B1(n_41),
.B2(n_84),
.Y(n_135)
);

BUFx12f_ASAP7_75t_L g52 ( 
.A(n_11),
.Y(n_52)
);

OAI22xp5_ASAP7_75t_L g63 ( 
.A1(n_12),
.A2(n_64),
.B1(n_65),
.B2(n_66),
.Y(n_63)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_12),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_L g91 ( 
.A1(n_12),
.A2(n_49),
.B1(n_50),
.B2(n_64),
.Y(n_91)
);

INVx13_ASAP7_75t_L g29 ( 
.A(n_13),
.Y(n_29)
);

AOI22xp33_ASAP7_75t_SL g46 ( 
.A1(n_14),
.A2(n_38),
.B1(n_41),
.B2(n_47),
.Y(n_46)
);

CKINVDCx20_ASAP7_75t_R g47 ( 
.A(n_14),
.Y(n_47)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_14),
.A2(n_47),
.B1(n_49),
.B2(n_50),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_L g169 ( 
.A1(n_14),
.A2(n_47),
.B1(n_65),
.B2(n_66),
.Y(n_169)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_15),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g42 ( 
.A1(n_16),
.A2(n_30),
.B1(n_31),
.B2(n_43),
.Y(n_42)
);

CKINVDCx16_ASAP7_75t_R g43 ( 
.A(n_16),
.Y(n_43)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_16),
.A2(n_38),
.B1(n_41),
.B2(n_43),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_16),
.A2(n_43),
.B1(n_49),
.B2(n_50),
.Y(n_196)
);

AOI22xp5_ASAP7_75t_SL g221 ( 
.A1(n_16),
.A2(n_43),
.B1(n_65),
.B2(n_66),
.Y(n_221)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_145),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_143),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_122),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_20),
.B(n_122),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_85),
.C(n_95),
.Y(n_20)
);

AOI22xp5_ASAP7_75t_L g269 ( 
.A1(n_21),
.A2(n_22),
.B1(n_85),
.B2(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g21 ( 
.A(n_22),
.Y(n_21)
);

XOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_60),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_44),
.B2(n_45),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_25),
.B(n_44),
.C(n_60),
.Y(n_142)
);

AOI22xp5_ASAP7_75t_L g25 ( 
.A1(n_26),
.A2(n_32),
.B1(n_37),
.B2(n_42),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g97 ( 
.A(n_26),
.Y(n_97)
);

INVx11_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx8_ASAP7_75t_L g31 ( 
.A(n_29),
.Y(n_31)
);

OAI22xp33_ASAP7_75t_L g33 ( 
.A1(n_29),
.A2(n_31),
.B1(n_34),
.B2(n_35),
.Y(n_33)
);

INVx8_ASAP7_75t_L g101 ( 
.A(n_29),
.Y(n_101)
);

INVx6_ASAP7_75t_L g115 ( 
.A(n_29),
.Y(n_115)
);

INVx11_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_31),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_32),
.B(n_99),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g138 ( 
.A(n_32),
.Y(n_138)
);

AOI21xp5_ASAP7_75t_L g158 ( 
.A1(n_32),
.A2(n_140),
.B(n_159),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_33),
.B(n_36),
.Y(n_32)
);

INVx4_ASAP7_75t_L g35 ( 
.A(n_34),
.Y(n_35)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_34),
.A2(n_35),
.B1(n_38),
.B2(n_41),
.Y(n_37)
);

A2O1A1Ixp33_ASAP7_75t_L g109 ( 
.A1(n_34),
.A2(n_38),
.B(n_110),
.C(n_112),
.Y(n_109)
);

NAND3xp33_ASAP7_75t_SL g112 ( 
.A(n_35),
.B(n_41),
.C(n_113),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_L g96 ( 
.A1(n_36),
.A2(n_97),
.B(n_98),
.Y(n_96)
);

NOR2xp33_ASAP7_75t_L g140 ( 
.A(n_36),
.B(n_100),
.Y(n_140)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_37),
.Y(n_36)
);

INVx5_ASAP7_75t_L g41 ( 
.A(n_38),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_L g59 ( 
.A1(n_38),
.A2(n_41),
.B1(n_52),
.B2(n_53),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g184 ( 
.A(n_38),
.B(n_185),
.Y(n_184)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

INVx8_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g137 ( 
.A(n_42),
.Y(n_137)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp5_ASAP7_75t_L g45 ( 
.A1(n_46),
.A2(n_48),
.B(n_54),
.Y(n_45)
);

OAI22xp5_ASAP7_75t_SL g134 ( 
.A1(n_46),
.A2(n_48),
.B1(n_58),
.B2(n_135),
.Y(n_134)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_59),
.Y(n_58)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_48),
.Y(n_106)
);

OAI21xp5_ASAP7_75t_SL g164 ( 
.A1(n_48),
.A2(n_54),
.B(n_165),
.Y(n_164)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_49),
.A2(n_50),
.B1(n_52),
.B2(n_53),
.Y(n_48)
);

OAI22xp33_ASAP7_75t_L g77 ( 
.A1(n_49),
.A2(n_50),
.B1(n_78),
.B2(n_80),
.Y(n_77)
);

INVx3_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_50),
.B(n_230),
.Y(n_229)
);

BUFx6f_ASAP7_75t_L g50 ( 
.A(n_51),
.Y(n_50)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_52),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_55),
.B(n_57),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g105 ( 
.A(n_55),
.B(n_106),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g152 ( 
.A1(n_57),
.A2(n_104),
.B1(n_106),
.B2(n_153),
.Y(n_152)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

OAI21xp5_ASAP7_75t_SL g102 ( 
.A1(n_58),
.A2(n_103),
.B(n_105),
.Y(n_102)
);

OAI21xp33_ASAP7_75t_L g198 ( 
.A1(n_58),
.A2(n_105),
.B(n_199),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_61),
.B(n_74),
.Y(n_60)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_61),
.B(n_74),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_SL g61 ( 
.A1(n_62),
.A2(n_67),
.B1(n_69),
.B2(n_71),
.Y(n_61)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g116 ( 
.A1(n_63),
.A2(n_117),
.B1(n_118),
.B2(n_120),
.Y(n_116)
);

INVx5_ASAP7_75t_L g66 ( 
.A(n_65),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_65),
.B(n_68),
.Y(n_67)
);

OA22x2_ASAP7_75t_L g81 ( 
.A1(n_65),
.A2(n_66),
.B1(n_78),
.B2(n_80),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_66),
.B(n_247),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g86 ( 
.A1(n_67),
.A2(n_69),
.B1(n_71),
.B2(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_67),
.Y(n_117)
);

AOI21xp5_ASAP7_75t_L g129 ( 
.A1(n_67),
.A2(n_71),
.B(n_87),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_67),
.A2(n_119),
.B1(n_169),
.B2(n_170),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_67),
.B(n_192),
.Y(n_191)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_67),
.A2(n_221),
.B(n_222),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_68),
.B(n_111),
.Y(n_247)
);

INVx5_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx5_ASAP7_75t_L g72 ( 
.A(n_73),
.Y(n_72)
);

INVx2_ASAP7_75t_L g223 ( 
.A(n_73),
.Y(n_223)
);

OAI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_81),
.B1(n_82),
.B2(n_83),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_SL g208 ( 
.A1(n_75),
.A2(n_209),
.B(n_210),
.Y(n_208)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_75),
.A2(n_210),
.B(n_228),
.Y(n_227)
);

INVx1_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

AOI22xp5_ASAP7_75t_L g89 ( 
.A1(n_76),
.A2(n_90),
.B1(n_91),
.B2(n_92),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_76),
.A2(n_91),
.B1(n_92),
.B2(n_127),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g156 ( 
.A(n_76),
.B(n_157),
.Y(n_156)
);

AOI22xp5_ASAP7_75t_L g193 ( 
.A1(n_76),
.A2(n_92),
.B1(n_194),
.B2(n_196),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_77),
.B(n_81),
.Y(n_76)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_78),
.Y(n_80)
);

BUFx24_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g92 ( 
.A(n_81),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_L g155 ( 
.A1(n_81),
.A2(n_82),
.B(n_156),
.Y(n_155)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_81),
.A2(n_156),
.B(n_195),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_81),
.B(n_111),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g90 ( 
.A(n_83),
.Y(n_90)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_85),
.Y(n_270)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_86),
.A2(n_89),
.B1(n_93),
.B2(n_94),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_86),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g131 ( 
.A(n_86),
.B(n_94),
.Y(n_131)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_89),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_92),
.B(n_157),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_95),
.B(n_269),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.C(n_107),
.Y(n_95)
);

XNOR2xp5_ASAP7_75t_L g173 ( 
.A(n_96),
.B(n_102),
.Y(n_173)
);

INVxp67_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx16_ASAP7_75t_R g103 ( 
.A(n_104),
.Y(n_103)
);

XNOR2xp5_ASAP7_75t_SL g172 ( 
.A(n_107),
.B(n_173),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_108),
.B(n_116),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_108),
.A2(n_109),
.B1(n_116),
.B2(n_162),
.Y(n_161)
);

CKINVDCx14_ASAP7_75t_R g108 ( 
.A(n_109),
.Y(n_108)
);

OAI21xp33_ASAP7_75t_L g159 ( 
.A1(n_110),
.A2(n_111),
.B(n_113),
.Y(n_159)
);

INVx8_ASAP7_75t_L g113 ( 
.A(n_114),
.Y(n_113)
);

INVx8_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_116),
.Y(n_162)
);

CKINVDCx16_ASAP7_75t_R g118 ( 
.A(n_119),
.Y(n_118)
);

INVx3_ASAP7_75t_SL g120 ( 
.A(n_121),
.Y(n_120)
);

INVx8_ASAP7_75t_L g190 ( 
.A(n_121),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_142),
.Y(n_122)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_130),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_SL g124 ( 
.A1(n_125),
.A2(n_126),
.B1(n_128),
.B2(n_129),
.Y(n_124)
);

CKINVDCx20_ASAP7_75t_R g125 ( 
.A(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_129),
.Y(n_128)
);

OAI22xp5_ASAP7_75t_L g130 ( 
.A1(n_131),
.A2(n_132),
.B1(n_133),
.B2(n_141),
.Y(n_130)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_131),
.Y(n_141)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_133),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_SL g133 ( 
.A(n_134),
.B(n_136),
.Y(n_133)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_137),
.A2(n_138),
.B(n_139),
.Y(n_136)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVxp67_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

O2A1O1Ixp33_ASAP7_75t_SL g145 ( 
.A1(n_146),
.A2(n_177),
.B(n_266),
.C(n_271),
.Y(n_145)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_171),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_147),
.B(n_171),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_148),
.B(n_160),
.C(n_163),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_L g260 ( 
.A1(n_148),
.A2(n_149),
.B1(n_261),
.B2(n_262),
.Y(n_260)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

XOR2xp5_ASAP7_75t_L g149 ( 
.A(n_150),
.B(n_158),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g150 ( 
.A1(n_151),
.A2(n_152),
.B1(n_154),
.B2(n_155),
.Y(n_150)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

MAJIxp5_ASAP7_75t_L g176 ( 
.A(n_152),
.B(n_154),
.C(n_158),
.Y(n_176)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_153),
.Y(n_165)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_155),
.Y(n_154)
);

AOI22xp5_ASAP7_75t_L g262 ( 
.A1(n_160),
.A2(n_161),
.B1(n_163),
.B2(n_263),
.Y(n_262)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_161),
.Y(n_160)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_163),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_164),
.B(n_166),
.C(n_168),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g202 ( 
.A(n_164),
.B(n_203),
.Y(n_202)
);

AOI22xp5_ASAP7_75t_L g203 ( 
.A1(n_166),
.A2(n_167),
.B1(n_168),
.B2(n_204),
.Y(n_203)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_168),
.Y(n_204)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_169),
.Y(n_187)
);

BUFx2_ASAP7_75t_L g243 ( 
.A(n_170),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_174),
.Y(n_171)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_172),
.B(n_175),
.C(n_176),
.Y(n_267)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_176),
.Y(n_174)
);

NOR2xp33_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_179),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_259),
.B(n_265),
.Y(n_179)
);

OAI21xp5_ASAP7_75t_L g180 ( 
.A1(n_181),
.A2(n_211),
.B(n_258),
.Y(n_180)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_200),
.Y(n_181)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_182),
.B(n_200),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_183),
.B(n_193),
.C(n_197),
.Y(n_182)
);

XNOR2xp5_ASAP7_75t_L g253 ( 
.A(n_183),
.B(n_254),
.Y(n_253)
);

XNOR2xp5_ASAP7_75t_SL g183 ( 
.A(n_184),
.B(n_186),
.Y(n_183)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_184),
.B(n_186),
.Y(n_207)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_187),
.A2(n_188),
.B(n_191),
.Y(n_186)
);

INVx3_ASAP7_75t_L g188 ( 
.A(n_189),
.Y(n_188)
);

INVx5_ASAP7_75t_L g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_191),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g224 ( 
.A(n_192),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_193),
.A2(n_197),
.B1(n_198),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_193),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g194 ( 
.A(n_195),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_196),
.Y(n_209)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g200 ( 
.A1(n_201),
.A2(n_202),
.B1(n_205),
.B2(n_206),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_201),
.B(n_207),
.C(n_208),
.Y(n_264)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_202),
.Y(n_201)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_206),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_208),
.Y(n_206)
);

AOI21xp5_ASAP7_75t_L g211 ( 
.A1(n_212),
.A2(n_252),
.B(n_257),
.Y(n_211)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_213),
.A2(n_231),
.B(n_251),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_SL g213 ( 
.A(n_214),
.B(n_225),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g251 ( 
.A(n_214),
.B(n_225),
.Y(n_251)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_215),
.B(n_220),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_217),
.B1(n_218),
.B2(n_219),
.Y(n_215)
);

MAJIxp5_ASAP7_75t_L g256 ( 
.A(n_216),
.B(n_219),
.C(n_220),
.Y(n_256)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g218 ( 
.A(n_219),
.Y(n_218)
);

CKINVDCx16_ASAP7_75t_R g236 ( 
.A(n_221),
.Y(n_236)
);

NAND2xp5_ASAP7_75t_L g222 ( 
.A(n_223),
.B(n_224),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_226),
.B(n_229),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g237 ( 
.A1(n_226),
.A2(n_227),
.B1(n_229),
.B2(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_227),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g238 ( 
.A(n_229),
.Y(n_238)
);

AOI21xp5_ASAP7_75t_L g231 ( 
.A1(n_232),
.A2(n_239),
.B(n_250),
.Y(n_231)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_233),
.B(n_237),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g250 ( 
.A(n_233),
.B(n_237),
.Y(n_250)
);

CKINVDCx16_ASAP7_75t_R g234 ( 
.A(n_235),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_235),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_240),
.A2(n_245),
.B(n_249),
.Y(n_239)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_241),
.B(n_242),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g249 ( 
.A(n_241),
.B(n_242),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_248),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_253),
.B(n_256),
.Y(n_252)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_253),
.B(n_256),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_260),
.B(n_264),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_260),
.B(n_264),
.Y(n_265)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_262),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_267),
.B(n_268),
.Y(n_271)
);


endmodule