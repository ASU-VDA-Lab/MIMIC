module real_aes_1615_n_105 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_104, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_103, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_105);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_104;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_103;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_105;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_778;
wire n_800;
wire n_522;
wire n_838;
wire n_485;
wire n_822;
wire n_222;
wire n_750;
wire n_631;
wire n_357;
wire n_503;
wire n_287;
wire n_635;
wire n_386;
wire n_673;
wire n_792;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_841;
wire n_318;
wire n_718;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_319;
wire n_364;
wire n_555;
wire n_421;
wire n_329;
wire n_766;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_571;
wire n_549;
wire n_376;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_594;
wire n_186;
wire n_767;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_775;
wire n_161;
wire n_763;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_815;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_816;
wire n_292;
wire n_539;
wire n_400;
wire n_626;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_578;
wire n_372;
wire n_528;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_824;
wire n_467;
wire n_327;
wire n_774;
wire n_813;
wire n_106;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_174;
wire n_840;
wire n_570;
wire n_675;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_784;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_178;
wire n_409;
wire n_748;
wire n_781;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_119;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_812;
wire n_817;
wire n_443;
wire n_565;
wire n_782;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_819;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_722;
wire n_745;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_363;
wire n_417;
wire n_449;
wire n_754;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_505;
wire n_434;
wire n_502;
wire n_527;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_602;
wire n_402;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_807;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_832;
wire n_410;
wire n_120;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_768;
wire n_412;
wire n_542;
wire n_163;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_779;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_765;
wire n_826;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_233;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_107;
wire n_229;
wire n_827;
wire n_809;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_335;
wire n_177;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_740;
wire n_371;
wire n_698;
wire n_166;
wire n_541;
wire n_224;
wire n_839;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_836;
wire n_793;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_772;
wire n_450;
wire n_788;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_474;
wire n_829;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_729;
wire n_687;
wire n_646;
wire n_710;
wire n_650;
wire n_743;
wire n_823;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_802;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_842;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_798;
wire n_237;
wire n_797;
wire n_668;
NAND2xp5_ASAP7_75t_L g579 ( .A(n_0), .B(n_178), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_1), .B(n_839), .Y(n_838) );
INVx1_ASAP7_75t_L g136 ( .A(n_2), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g540 ( .A(n_3), .B(n_541), .Y(n_540) );
NAND2xp33_ASAP7_75t_SL g622 ( .A(n_4), .B(n_165), .Y(n_622) );
NAND2xp5_ASAP7_75t_SL g169 ( .A(n_5), .B(n_145), .Y(n_169) );
INVx1_ASAP7_75t_L g615 ( .A(n_6), .Y(n_615) );
INVx1_ASAP7_75t_L g191 ( .A(n_7), .Y(n_191) );
CKINVDCx16_ASAP7_75t_R g839 ( .A(n_8), .Y(n_839) );
CKINVDCx5p33_ASAP7_75t_R g207 ( .A(n_9), .Y(n_207) );
AND2x2_ASAP7_75t_L g538 ( .A(n_10), .B(n_222), .Y(n_538) );
INVx2_ASAP7_75t_L g144 ( .A(n_11), .Y(n_144) );
CKINVDCx16_ASAP7_75t_R g500 ( .A(n_12), .Y(n_500) );
NOR3xp33_ASAP7_75t_L g837 ( .A(n_12), .B(n_838), .C(n_840), .Y(n_837) );
INVx1_ASAP7_75t_L g179 ( .A(n_13), .Y(n_179) );
AOI221x1_ASAP7_75t_L g618 ( .A1(n_14), .A2(n_196), .B1(n_543), .B2(n_619), .C(n_621), .Y(n_618) );
NAND2xp5_ASAP7_75t_SL g602 ( .A(n_15), .B(n_541), .Y(n_602) );
INVx1_ASAP7_75t_L g504 ( .A(n_16), .Y(n_504) );
NOR2xp33_ASAP7_75t_SL g835 ( .A(n_16), .B(n_505), .Y(n_835) );
INVx1_ASAP7_75t_L g176 ( .A(n_17), .Y(n_176) );
INVx1_ASAP7_75t_SL g251 ( .A(n_18), .Y(n_251) );
INVxp33_ASAP7_75t_L g842 ( .A(n_19), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g155 ( .A(n_20), .B(n_156), .Y(n_155) );
AOI22xp5_ASAP7_75t_L g815 ( .A1(n_21), .A2(n_816), .B1(n_817), .B2(n_818), .Y(n_815) );
INVx1_ASAP7_75t_L g816 ( .A(n_21), .Y(n_816) );
AOI33xp33_ASAP7_75t_L g228 ( .A1(n_22), .A2(n_52), .A3(n_133), .B1(n_151), .B2(n_229), .B3(n_230), .Y(n_228) );
AOI21xp5_ASAP7_75t_L g542 ( .A1(n_23), .A2(n_543), .B(n_544), .Y(n_542) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_24), .B(n_178), .Y(n_545) );
AOI221xp5_ASAP7_75t_SL g589 ( .A1(n_25), .A2(n_41), .B1(n_541), .B2(n_543), .C(n_590), .Y(n_589) );
INVx1_ASAP7_75t_L g200 ( .A(n_26), .Y(n_200) );
OAI22x1_ASAP7_75t_R g494 ( .A1(n_27), .A2(n_65), .B1(n_495), .B2(n_496), .Y(n_494) );
INVx1_ASAP7_75t_L g496 ( .A(n_27), .Y(n_496) );
OA21x2_ASAP7_75t_L g143 ( .A1(n_28), .A2(n_93), .B(n_144), .Y(n_143) );
OR2x2_ASAP7_75t_L g146 ( .A(n_28), .B(n_93), .Y(n_146) );
NAND2xp5_ASAP7_75t_L g606 ( .A(n_29), .B(n_181), .Y(n_606) );
INVxp67_ASAP7_75t_L g617 ( .A(n_30), .Y(n_617) );
AND2x2_ASAP7_75t_L g564 ( .A(n_31), .B(n_221), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_32), .B(n_189), .Y(n_248) );
AOI21xp5_ASAP7_75t_L g577 ( .A1(n_33), .A2(n_543), .B(n_578), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g591 ( .A(n_34), .B(n_181), .Y(n_591) );
AND2x2_ASAP7_75t_L g139 ( .A(n_35), .B(n_140), .Y(n_139) );
INVx1_ASAP7_75t_L g150 ( .A(n_35), .Y(n_150) );
AND2x2_ASAP7_75t_L g165 ( .A(n_35), .B(n_136), .Y(n_165) );
OR2x6_ASAP7_75t_L g502 ( .A(n_36), .B(n_503), .Y(n_502) );
INVxp67_ASAP7_75t_L g840 ( .A(n_36), .Y(n_840) );
CKINVDCx20_ASAP7_75t_R g202 ( .A(n_37), .Y(n_202) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_38), .B(n_189), .Y(n_215) );
AOI22xp5_ASAP7_75t_L g129 ( .A1(n_39), .A2(n_130), .B1(n_142), .B2(n_145), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g161 ( .A(n_40), .B(n_162), .Y(n_161) );
AOI22xp5_ASAP7_75t_L g570 ( .A1(n_42), .A2(n_83), .B1(n_148), .B2(n_543), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g252 ( .A(n_43), .B(n_156), .Y(n_252) );
AOI22xp5_ASAP7_75t_SL g819 ( .A1(n_44), .A2(n_74), .B1(n_820), .B2(n_821), .Y(n_819) );
CKINVDCx20_ASAP7_75t_R g821 ( .A(n_44), .Y(n_821) );
CKINVDCx20_ASAP7_75t_R g825 ( .A(n_45), .Y(n_825) );
NAND2xp5_ASAP7_75t_L g562 ( .A(n_46), .B(n_178), .Y(n_562) );
NAND2xp5_ASAP7_75t_SL g193 ( .A(n_47), .B(n_167), .Y(n_193) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_48), .B(n_156), .Y(n_192) );
CKINVDCx5p33_ASAP7_75t_R g141 ( .A(n_49), .Y(n_141) );
AND2x2_ASAP7_75t_L g582 ( .A(n_50), .B(n_221), .Y(n_582) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_51), .B(n_221), .Y(n_593) );
NAND2xp5_ASAP7_75t_L g219 ( .A(n_53), .B(n_156), .Y(n_219) );
INVx1_ASAP7_75t_L g134 ( .A(n_54), .Y(n_134) );
INVx1_ASAP7_75t_L g158 ( .A(n_54), .Y(n_158) );
XOR2x2_ASAP7_75t_L g818 ( .A(n_55), .B(n_819), .Y(n_818) );
AND2x2_ASAP7_75t_L g220 ( .A(n_56), .B(n_221), .Y(n_220) );
AOI221xp5_ASAP7_75t_L g188 ( .A1(n_57), .A2(n_76), .B1(n_148), .B2(n_189), .C(n_190), .Y(n_188) );
NAND2xp5_ASAP7_75t_L g243 ( .A(n_58), .B(n_189), .Y(n_243) );
NAND2xp5_ASAP7_75t_SL g563 ( .A(n_59), .B(n_541), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g209 ( .A(n_60), .B(n_142), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g239 ( .A1(n_61), .A2(n_148), .B(n_240), .Y(n_239) );
AND2x2_ASAP7_75t_L g555 ( .A(n_62), .B(n_221), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_63), .B(n_181), .Y(n_580) );
INVx1_ASAP7_75t_L g172 ( .A(n_64), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g495 ( .A(n_65), .Y(n_495) );
AND2x2_ASAP7_75t_SL g607 ( .A(n_65), .B(n_222), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g553 ( .A(n_66), .B(n_178), .Y(n_553) );
AOI21xp5_ASAP7_75t_L g559 ( .A1(n_67), .A2(n_543), .B(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g218 ( .A(n_68), .Y(n_218) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_69), .B(n_181), .Y(n_546) );
AND2x2_ASAP7_75t_SL g571 ( .A(n_70), .B(n_167), .Y(n_571) );
AOI21xp5_ASAP7_75t_L g216 ( .A1(n_71), .A2(n_148), .B(n_217), .Y(n_216) );
AOI22xp5_ASAP7_75t_L g117 ( .A1(n_72), .A2(n_91), .B1(n_118), .B2(n_119), .Y(n_117) );
INVx1_ASAP7_75t_L g119 ( .A(n_72), .Y(n_119) );
INVx1_ASAP7_75t_L g140 ( .A(n_73), .Y(n_140) );
INVx1_ASAP7_75t_L g160 ( .A(n_73), .Y(n_160) );
CKINVDCx20_ASAP7_75t_R g820 ( .A(n_74), .Y(n_820) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_75), .B(n_189), .Y(n_231) );
AND2x2_ASAP7_75t_L g253 ( .A(n_77), .B(n_196), .Y(n_253) );
INVx1_ASAP7_75t_L g173 ( .A(n_78), .Y(n_173) );
AOI21xp5_ASAP7_75t_L g249 ( .A1(n_79), .A2(n_148), .B(n_250), .Y(n_249) );
A2O1A1Ixp33_ASAP7_75t_L g147 ( .A1(n_80), .A2(n_148), .B(n_154), .C(n_166), .Y(n_147) );
NAND2xp5_ASAP7_75t_SL g554 ( .A(n_81), .B(n_541), .Y(n_554) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_82), .A2(n_86), .B1(n_189), .B2(n_541), .Y(n_569) );
INVx1_ASAP7_75t_L g505 ( .A(n_84), .Y(n_505) );
AND2x2_ASAP7_75t_SL g237 ( .A(n_85), .B(n_196), .Y(n_237) );
AOI22xp5_ASAP7_75t_L g225 ( .A1(n_87), .A2(n_148), .B1(n_226), .B2(n_227), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g605 ( .A(n_88), .B(n_178), .Y(n_605) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_89), .B(n_178), .Y(n_592) );
OAI22xp5_ASAP7_75t_SL g115 ( .A1(n_90), .A2(n_116), .B1(n_117), .B2(n_120), .Y(n_115) );
INVx1_ASAP7_75t_L g120 ( .A(n_90), .Y(n_120) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_91), .Y(n_118) );
NOR3xp33_ASAP7_75t_L g519 ( .A(n_91), .B(n_123), .C(n_464), .Y(n_519) );
AOI21xp5_ASAP7_75t_L g550 ( .A1(n_92), .A2(n_543), .B(n_551), .Y(n_550) );
INVx1_ASAP7_75t_L g241 ( .A(n_94), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g552 ( .A(n_95), .B(n_181), .Y(n_552) );
AND2x2_ASAP7_75t_L g232 ( .A(n_96), .B(n_196), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_97), .A2(n_198), .B(n_199), .C(n_201), .Y(n_197) );
NAND2xp5_ASAP7_75t_L g581 ( .A(n_98), .B(n_541), .Y(n_581) );
INVxp67_ASAP7_75t_L g620 ( .A(n_99), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g561 ( .A(n_100), .B(n_181), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g603 ( .A1(n_101), .A2(n_543), .B(n_604), .Y(n_603) );
INVx1_ASAP7_75t_L g515 ( .A(n_102), .Y(n_515) );
BUFx2_ASAP7_75t_SL g111 ( .A(n_103), .Y(n_111) );
BUFx2_ASAP7_75t_L g506 ( .A(n_103), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_104), .B(n_156), .Y(n_242) );
AOI21xp33_ASAP7_75t_L g105 ( .A1(n_106), .A2(n_829), .B(n_841), .Y(n_105) );
AO21x2_ASAP7_75t_L g106 ( .A1(n_107), .A2(n_507), .B(n_824), .Y(n_106) );
AOI21xp5_ASAP7_75t_L g107 ( .A1(n_108), .A2(n_112), .B(n_498), .Y(n_107) );
CKINVDCx5p33_ASAP7_75t_R g108 ( .A(n_109), .Y(n_108) );
CKINVDCx11_ASAP7_75t_R g109 ( .A(n_110), .Y(n_109) );
CKINVDCx8_ASAP7_75t_R g110 ( .A(n_111), .Y(n_110) );
OAI22xp5_ASAP7_75t_L g112 ( .A1(n_113), .A2(n_493), .B1(n_494), .B2(n_497), .Y(n_112) );
INVx2_ASAP7_75t_L g497 ( .A(n_113), .Y(n_497) );
XNOR2x1_ASAP7_75t_L g113 ( .A(n_114), .B(n_121), .Y(n_113) );
CKINVDCx5p33_ASAP7_75t_R g114 ( .A(n_115), .Y(n_114) );
INVx1_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
AOI21xp5_ASAP7_75t_L g521 ( .A1(n_118), .A2(n_522), .B(n_523), .Y(n_521) );
AOI21xp5_ASAP7_75t_SL g524 ( .A1(n_118), .A2(n_525), .B(n_526), .Y(n_524) );
AND2x2_ASAP7_75t_L g121 ( .A(n_122), .B(n_427), .Y(n_121) );
NOR2xp33_ASAP7_75t_L g122 ( .A(n_123), .B(n_350), .Y(n_122) );
INVxp67_ASAP7_75t_L g523 ( .A(n_123), .Y(n_523) );
NAND3xp33_ASAP7_75t_L g123 ( .A(n_124), .B(n_297), .C(n_330), .Y(n_123) );
AOI211xp5_ASAP7_75t_L g124 ( .A1(n_125), .A2(n_254), .B(n_263), .C(n_287), .Y(n_124) );
OAI21xp33_ASAP7_75t_L g125 ( .A1(n_126), .A2(n_183), .B(n_233), .Y(n_125) );
OR2x2_ASAP7_75t_L g307 ( .A(n_126), .B(n_308), .Y(n_307) );
OR2x2_ASAP7_75t_L g462 ( .A(n_126), .B(n_463), .Y(n_462) );
INVx2_ASAP7_75t_L g126 ( .A(n_127), .Y(n_126) );
AOI22xp33_ASAP7_75t_SL g352 ( .A1(n_127), .A2(n_353), .B1(n_357), .B2(n_359), .Y(n_352) );
AND2x2_ASAP7_75t_L g389 ( .A(n_127), .B(n_390), .Y(n_389) );
AND2x2_ASAP7_75t_L g127 ( .A(n_128), .B(n_168), .Y(n_127) );
INVx1_ASAP7_75t_L g286 ( .A(n_128), .Y(n_286) );
AND2x4_ASAP7_75t_L g303 ( .A(n_128), .B(n_284), .Y(n_303) );
INVx2_ASAP7_75t_L g325 ( .A(n_128), .Y(n_325) );
HB1xp67_ASAP7_75t_L g408 ( .A(n_128), .Y(n_408) );
AND2x2_ASAP7_75t_L g479 ( .A(n_128), .B(n_236), .Y(n_479) );
AND2x2_ASAP7_75t_L g128 ( .A(n_129), .B(n_147), .Y(n_128) );
NOR3xp33_ASAP7_75t_L g130 ( .A(n_131), .B(n_137), .C(n_141), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x4_ASAP7_75t_L g189 ( .A(n_132), .B(n_138), .Y(n_189) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_135), .Y(n_132) );
OR2x6_ASAP7_75t_L g163 ( .A(n_133), .B(n_152), .Y(n_163) );
INVxp33_ASAP7_75t_L g229 ( .A(n_133), .Y(n_229) );
INVx2_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
AND2x2_ASAP7_75t_L g153 ( .A(n_134), .B(n_136), .Y(n_153) );
AND2x4_ASAP7_75t_L g181 ( .A(n_134), .B(n_159), .Y(n_181) );
HB1xp67_ASAP7_75t_L g135 ( .A(n_136), .Y(n_135) );
INVx1_ASAP7_75t_L g137 ( .A(n_138), .Y(n_137) );
BUFx3_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
AND2x6_ASAP7_75t_L g543 ( .A(n_139), .B(n_153), .Y(n_543) );
INVx2_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
AND2x6_ASAP7_75t_L g178 ( .A(n_140), .B(n_157), .Y(n_178) );
INVx4_ASAP7_75t_L g196 ( .A(n_142), .Y(n_196) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_142), .B(n_206), .Y(n_205) );
AOI21x1_ASAP7_75t_L g575 ( .A1(n_142), .A2(n_576), .B(n_582), .Y(n_575) );
INVx3_ASAP7_75t_L g142 ( .A(n_143), .Y(n_142) );
BUFx4f_ASAP7_75t_L g167 ( .A(n_143), .Y(n_167) );
AND2x4_ASAP7_75t_L g145 ( .A(n_144), .B(n_146), .Y(n_145) );
AND2x2_ASAP7_75t_SL g222 ( .A(n_144), .B(n_146), .Y(n_222) );
NOR2xp33_ASAP7_75t_L g182 ( .A(n_145), .B(n_164), .Y(n_182) );
AOI21xp5_ASAP7_75t_L g238 ( .A1(n_145), .A2(n_239), .B(n_243), .Y(n_238) );
AOI21xp5_ASAP7_75t_L g539 ( .A1(n_145), .A2(n_540), .B(n_542), .Y(n_539) );
NOR2xp33_ASAP7_75t_L g614 ( .A(n_145), .B(n_615), .Y(n_614) );
NOR2xp33_ASAP7_75t_L g616 ( .A(n_145), .B(n_617), .Y(n_616) );
NOR2xp33_ASAP7_75t_L g619 ( .A(n_145), .B(n_620), .Y(n_619) );
NOR3xp33_ASAP7_75t_L g621 ( .A(n_145), .B(n_174), .C(n_622), .Y(n_621) );
INVxp67_ASAP7_75t_L g208 ( .A(n_148), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g613 ( .A1(n_148), .A2(n_189), .B1(n_614), .B2(n_616), .Y(n_613) );
AND2x4_ASAP7_75t_L g148 ( .A(n_149), .B(n_153), .Y(n_148) );
NOR2x1p5_ASAP7_75t_L g149 ( .A(n_150), .B(n_151), .Y(n_149) );
INVx1_ASAP7_75t_L g230 ( .A(n_151), .Y(n_230) );
INVx3_ASAP7_75t_L g151 ( .A(n_152), .Y(n_151) );
AOI21xp5_ASAP7_75t_L g154 ( .A1(n_155), .A2(n_161), .B(n_164), .Y(n_154) );
INVx1_ASAP7_75t_L g174 ( .A(n_156), .Y(n_174) );
AND2x4_ASAP7_75t_L g541 ( .A(n_156), .B(n_165), .Y(n_541) );
AND2x4_ASAP7_75t_L g156 ( .A(n_157), .B(n_159), .Y(n_156) );
INVx2_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
INVx2_ASAP7_75t_L g159 ( .A(n_160), .Y(n_159) );
INVx2_ASAP7_75t_L g162 ( .A(n_163), .Y(n_162) );
OAI22xp5_ASAP7_75t_L g171 ( .A1(n_163), .A2(n_172), .B1(n_173), .B2(n_174), .Y(n_171) );
O2A1O1Ixp33_ASAP7_75t_SL g190 ( .A1(n_163), .A2(n_164), .B(n_191), .C(n_192), .Y(n_190) );
INVxp67_ASAP7_75t_L g198 ( .A(n_163), .Y(n_198) );
O2A1O1Ixp33_ASAP7_75t_L g217 ( .A1(n_163), .A2(n_164), .B(n_218), .C(n_219), .Y(n_217) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_163), .A2(n_164), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g250 ( .A1(n_163), .A2(n_164), .B(n_251), .C(n_252), .Y(n_250) );
INVx1_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_164), .A2(n_545), .B(n_546), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g551 ( .A1(n_164), .A2(n_552), .B(n_553), .Y(n_551) );
AOI21xp5_ASAP7_75t_L g560 ( .A1(n_164), .A2(n_561), .B(n_562), .Y(n_560) );
AOI21xp5_ASAP7_75t_L g578 ( .A1(n_164), .A2(n_579), .B(n_580), .Y(n_578) );
AOI21xp5_ASAP7_75t_L g590 ( .A1(n_164), .A2(n_591), .B(n_592), .Y(n_590) );
AOI21xp5_ASAP7_75t_L g604 ( .A1(n_164), .A2(n_605), .B(n_606), .Y(n_604) );
INVx5_ASAP7_75t_L g164 ( .A(n_165), .Y(n_164) );
HB1xp67_ASAP7_75t_L g201 ( .A(n_165), .Y(n_201) );
AO21x2_ASAP7_75t_L g223 ( .A1(n_166), .A2(n_224), .B(n_232), .Y(n_223) );
AO21x2_ASAP7_75t_L g268 ( .A1(n_166), .A2(n_224), .B(n_232), .Y(n_268) );
AOI21x1_ASAP7_75t_L g567 ( .A1(n_166), .A2(n_568), .B(n_571), .Y(n_567) );
INVx2_ASAP7_75t_SL g166 ( .A(n_167), .Y(n_166) );
OA21x2_ASAP7_75t_L g187 ( .A1(n_167), .A2(n_188), .B(n_193), .Y(n_187) );
AOI21xp5_ASAP7_75t_L g601 ( .A1(n_167), .A2(n_602), .B(n_603), .Y(n_601) );
AND2x2_ASAP7_75t_L g244 ( .A(n_168), .B(n_245), .Y(n_244) );
INVx2_ASAP7_75t_L g273 ( .A(n_168), .Y(n_273) );
INVx3_ASAP7_75t_L g284 ( .A(n_168), .Y(n_284) );
AND2x4_ASAP7_75t_L g168 ( .A(n_169), .B(n_170), .Y(n_168) );
OAI21xp5_ASAP7_75t_L g170 ( .A1(n_171), .A2(n_175), .B(n_182), .Y(n_170) );
NOR2xp33_ASAP7_75t_L g199 ( .A(n_174), .B(n_200), .Y(n_199) );
OAI22xp5_ASAP7_75t_L g175 ( .A1(n_176), .A2(n_177), .B1(n_179), .B2(n_180), .Y(n_175) );
INVxp67_ASAP7_75t_L g177 ( .A(n_178), .Y(n_177) );
INVxp67_ASAP7_75t_L g180 ( .A(n_181), .Y(n_180) );
OAI22xp5_ASAP7_75t_L g473 ( .A1(n_183), .A2(n_474), .B1(n_476), .B2(n_478), .Y(n_473) );
NAND2xp5_ASAP7_75t_SL g484 ( .A(n_183), .B(n_485), .Y(n_484) );
INVx2_ASAP7_75t_SL g183 ( .A(n_184), .Y(n_183) );
AND2x2_ASAP7_75t_L g184 ( .A(n_185), .B(n_211), .Y(n_184) );
INVx3_ASAP7_75t_L g257 ( .A(n_185), .Y(n_257) );
AND2x2_ASAP7_75t_L g265 ( .A(n_185), .B(n_266), .Y(n_265) );
HB1xp67_ASAP7_75t_L g295 ( .A(n_185), .Y(n_295) );
NAND2x1_ASAP7_75t_SL g489 ( .A(n_185), .B(n_256), .Y(n_489) );
AND2x4_ASAP7_75t_L g185 ( .A(n_186), .B(n_194), .Y(n_185) );
INVx2_ASAP7_75t_L g186 ( .A(n_187), .Y(n_186) );
INVx1_ASAP7_75t_L g262 ( .A(n_187), .Y(n_262) );
NAND2xp5_ASAP7_75t_L g280 ( .A(n_187), .B(n_268), .Y(n_280) );
AND2x2_ASAP7_75t_L g293 ( .A(n_187), .B(n_194), .Y(n_293) );
AND2x4_ASAP7_75t_L g300 ( .A(n_187), .B(n_301), .Y(n_300) );
HB1xp67_ASAP7_75t_L g349 ( .A(n_187), .Y(n_349) );
INVxp67_ASAP7_75t_L g356 ( .A(n_187), .Y(n_356) );
INVx1_ASAP7_75t_L g361 ( .A(n_187), .Y(n_361) );
INVx1_ASAP7_75t_L g210 ( .A(n_189), .Y(n_210) );
INVx1_ASAP7_75t_L g260 ( .A(n_194), .Y(n_260) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_194), .B(n_270), .Y(n_279) );
INVx2_ASAP7_75t_L g347 ( .A(n_194), .Y(n_347) );
INVx1_ASAP7_75t_L g386 ( .A(n_194), .Y(n_386) );
OR2x2_ASAP7_75t_L g194 ( .A(n_195), .B(n_204), .Y(n_194) );
OAI22xp5_ASAP7_75t_L g195 ( .A1(n_196), .A2(n_197), .B1(n_202), .B2(n_203), .Y(n_195) );
INVx3_ASAP7_75t_L g203 ( .A(n_196), .Y(n_203) );
AO21x2_ASAP7_75t_L g213 ( .A1(n_203), .A2(n_214), .B(n_220), .Y(n_213) );
AO21x2_ASAP7_75t_L g270 ( .A1(n_203), .A2(n_214), .B(n_220), .Y(n_270) );
OAI22xp5_ASAP7_75t_L g204 ( .A1(n_205), .A2(n_208), .B1(n_209), .B2(n_210), .Y(n_204) );
INVx1_ASAP7_75t_L g206 ( .A(n_207), .Y(n_206) );
AND2x2_ASAP7_75t_L g316 ( .A(n_211), .B(n_293), .Y(n_316) );
AND2x2_ASAP7_75t_L g384 ( .A(n_211), .B(n_385), .Y(n_384) );
AND2x2_ASAP7_75t_L g398 ( .A(n_211), .B(n_399), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_211), .B(n_413), .Y(n_412) );
AND2x4_ASAP7_75t_L g211 ( .A(n_212), .B(n_223), .Y(n_211) );
INVx2_ASAP7_75t_L g212 ( .A(n_213), .Y(n_212) );
NOR2x1_ASAP7_75t_L g261 ( .A(n_213), .B(n_262), .Y(n_261) );
AND2x2_ASAP7_75t_L g354 ( .A(n_213), .B(n_347), .Y(n_354) );
AND2x2_ASAP7_75t_L g445 ( .A(n_213), .B(n_267), .Y(n_445) );
NAND2xp5_ASAP7_75t_L g214 ( .A(n_215), .B(n_216), .Y(n_214) );
CKINVDCx5p33_ASAP7_75t_R g246 ( .A(n_221), .Y(n_246) );
OA21x2_ASAP7_75t_L g588 ( .A1(n_221), .A2(n_589), .B(n_593), .Y(n_588) );
BUFx6f_ASAP7_75t_L g221 ( .A(n_222), .Y(n_221) );
INVx1_ASAP7_75t_L g256 ( .A(n_223), .Y(n_256) );
INVx2_ASAP7_75t_L g301 ( .A(n_223), .Y(n_301) );
AND2x2_ASAP7_75t_L g346 ( .A(n_223), .B(n_347), .Y(n_346) );
NAND2xp5_ASAP7_75t_SL g224 ( .A(n_225), .B(n_231), .Y(n_224) );
INVx1_ASAP7_75t_L g227 ( .A(n_228), .Y(n_227) );
INVx1_ASAP7_75t_L g233 ( .A(n_234), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_235), .B(n_244), .Y(n_234) );
AND2x2_ASAP7_75t_L g388 ( .A(n_235), .B(n_389), .Y(n_388) );
OR2x6_ASAP7_75t_L g447 ( .A(n_235), .B(n_448), .Y(n_447) );
BUFx6f_ASAP7_75t_L g235 ( .A(n_236), .Y(n_235) );
INVx4_ASAP7_75t_L g277 ( .A(n_236), .Y(n_277) );
AND2x4_ASAP7_75t_L g285 ( .A(n_236), .B(n_286), .Y(n_285) );
OR2x2_ASAP7_75t_L g320 ( .A(n_236), .B(n_245), .Y(n_320) );
INVx2_ASAP7_75t_L g369 ( .A(n_236), .Y(n_369) );
NAND2xp5_ASAP7_75t_SL g418 ( .A(n_236), .B(n_343), .Y(n_418) );
AND2x2_ASAP7_75t_L g455 ( .A(n_236), .B(n_273), .Y(n_455) );
NAND2xp5_ASAP7_75t_L g463 ( .A(n_236), .B(n_338), .Y(n_463) );
OR2x6_ASAP7_75t_L g236 ( .A(n_237), .B(n_238), .Y(n_236) );
AND2x2_ASAP7_75t_L g296 ( .A(n_244), .B(n_285), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_244), .B(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_SL g435 ( .A(n_244), .B(n_323), .Y(n_435) );
NAND2xp5_ASAP7_75t_L g457 ( .A(n_244), .B(n_336), .Y(n_457) );
HB1xp67_ASAP7_75t_L g275 ( .A(n_245), .Y(n_275) );
AND2x2_ASAP7_75t_L g283 ( .A(n_245), .B(n_284), .Y(n_283) );
HB1xp67_ASAP7_75t_L g306 ( .A(n_245), .Y(n_306) );
INVx2_ASAP7_75t_L g309 ( .A(n_245), .Y(n_309) );
INVx1_ASAP7_75t_L g342 ( .A(n_245), .Y(n_342) );
INVx1_ASAP7_75t_L g390 ( .A(n_245), .Y(n_390) );
AO21x2_ASAP7_75t_L g245 ( .A1(n_246), .A2(n_247), .B(n_253), .Y(n_245) );
AO21x2_ASAP7_75t_L g548 ( .A1(n_246), .A2(n_549), .B(n_555), .Y(n_548) );
AO21x2_ASAP7_75t_L g557 ( .A1(n_246), .A2(n_558), .B(n_564), .Y(n_557) );
AO21x2_ASAP7_75t_L g596 ( .A1(n_246), .A2(n_558), .B(n_564), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g247 ( .A(n_248), .B(n_249), .Y(n_247) );
NAND2xp33_ASAP7_75t_L g254 ( .A(n_255), .B(n_258), .Y(n_254) );
OR2x2_ASAP7_75t_L g255 ( .A(n_256), .B(n_257), .Y(n_255) );
NAND2xp5_ASAP7_75t_L g332 ( .A(n_256), .B(n_259), .Y(n_332) );
OR2x2_ASAP7_75t_L g404 ( .A(n_256), .B(n_405), .Y(n_404) );
AND4x1_ASAP7_75t_SL g450 ( .A(n_256), .B(n_432), .C(n_451), .D(n_452), .Y(n_450) );
OR2x2_ASAP7_75t_L g474 ( .A(n_257), .B(n_475), .Y(n_474) );
INVx1_ASAP7_75t_L g258 ( .A(n_259), .Y(n_258) );
AND2x2_ASAP7_75t_L g259 ( .A(n_260), .B(n_261), .Y(n_259) );
AND2x2_ASAP7_75t_L g311 ( .A(n_260), .B(n_312), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g461 ( .A(n_260), .B(n_269), .Y(n_461) );
AND2x2_ASAP7_75t_L g486 ( .A(n_261), .B(n_346), .Y(n_486) );
OAI32xp33_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_271), .A3(n_276), .B1(n_278), .B2(n_281), .Y(n_263) );
INVx2_ASAP7_75t_L g264 ( .A(n_265), .Y(n_264) );
AND2x2_ASAP7_75t_L g359 ( .A(n_266), .B(n_360), .Y(n_359) );
AND2x2_ASAP7_75t_L g459 ( .A(n_266), .B(n_413), .Y(n_459) );
AND2x4_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
AND2x2_ASAP7_75t_L g355 ( .A(n_267), .B(n_356), .Y(n_355) );
INVx1_ASAP7_75t_L g441 ( .A(n_267), .Y(n_441) );
INVx2_ASAP7_75t_L g267 ( .A(n_268), .Y(n_267) );
NAND2xp5_ASAP7_75t_L g475 ( .A(n_268), .B(n_270), .Y(n_475) );
INVx3_ASAP7_75t_L g292 ( .A(n_269), .Y(n_292) );
NAND2x1p5_ASAP7_75t_L g470 ( .A(n_269), .B(n_397), .Y(n_470) );
INVx3_ASAP7_75t_L g269 ( .A(n_270), .Y(n_269) );
HB1xp67_ASAP7_75t_L g329 ( .A(n_270), .Y(n_329) );
AND2x2_ASAP7_75t_L g348 ( .A(n_270), .B(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g271 ( .A(n_272), .Y(n_271) );
INVx1_ASAP7_75t_L g482 ( .A(n_272), .Y(n_482) );
NAND2x1_ASAP7_75t_L g272 ( .A(n_273), .B(n_274), .Y(n_272) );
INVx1_ASAP7_75t_L g322 ( .A(n_273), .Y(n_322) );
NOR2x1_ASAP7_75t_L g423 ( .A(n_273), .B(n_424), .Y(n_423) );
INVx1_ASAP7_75t_L g274 ( .A(n_275), .Y(n_274) );
NAND2xp5_ASAP7_75t_L g381 ( .A(n_276), .B(n_382), .Y(n_381) );
HB1xp67_ASAP7_75t_L g276 ( .A(n_277), .Y(n_276) );
OR2x2_ASAP7_75t_L g314 ( .A(n_277), .B(n_282), .Y(n_314) );
AND2x4_ASAP7_75t_L g336 ( .A(n_277), .B(n_286), .Y(n_336) );
AND2x4_ASAP7_75t_SL g407 ( .A(n_277), .B(n_408), .Y(n_407) );
NOR2x1_ASAP7_75t_L g433 ( .A(n_277), .B(n_358), .Y(n_433) );
OAI22xp5_ASAP7_75t_L g400 ( .A1(n_278), .A2(n_401), .B1(n_404), .B2(n_406), .Y(n_400) );
OR2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_280), .Y(n_278) );
INVx2_ASAP7_75t_SL g420 ( .A(n_279), .Y(n_420) );
INVx2_ASAP7_75t_L g312 ( .A(n_280), .Y(n_312) );
NAND2xp5_ASAP7_75t_L g281 ( .A(n_282), .B(n_285), .Y(n_281) );
INVx1_ASAP7_75t_SL g282 ( .A(n_283), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g288 ( .A(n_283), .B(n_289), .Y(n_288) );
AOI22xp5_ASAP7_75t_L g421 ( .A1(n_283), .A2(n_419), .B1(n_422), .B2(n_425), .Y(n_421) );
INVx1_ASAP7_75t_L g343 ( .A(n_284), .Y(n_343) );
AND2x2_ASAP7_75t_L g366 ( .A(n_284), .B(n_325), .Y(n_366) );
INVx2_ASAP7_75t_L g289 ( .A(n_285), .Y(n_289) );
OAI21xp5_ASAP7_75t_SL g287 ( .A1(n_288), .A2(n_290), .B(n_294), .Y(n_287) );
INVx1_ASAP7_75t_SL g290 ( .A(n_291), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g362 ( .A1(n_291), .A2(n_363), .B1(n_367), .B2(n_368), .Y(n_362) );
AND2x2_ASAP7_75t_L g291 ( .A(n_292), .B(n_293), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_292), .B(n_306), .Y(n_305) );
NAND2xp5_ASAP7_75t_L g376 ( .A(n_292), .B(n_360), .Y(n_376) );
INVx1_ASAP7_75t_L g380 ( .A(n_292), .Y(n_380) );
NAND2xp5_ASAP7_75t_L g294 ( .A(n_295), .B(n_296), .Y(n_294) );
NOR3xp33_ASAP7_75t_L g297 ( .A(n_298), .B(n_313), .C(n_317), .Y(n_297) );
OAI22xp5_ASAP7_75t_L g298 ( .A1(n_299), .A2(n_302), .B1(n_307), .B2(n_310), .Y(n_298) );
INVx1_ASAP7_75t_L g299 ( .A(n_300), .Y(n_299) );
AND2x2_ASAP7_75t_L g327 ( .A(n_300), .B(n_328), .Y(n_327) );
AND2x2_ASAP7_75t_L g367 ( .A(n_300), .B(n_354), .Y(n_367) );
AND2x2_ASAP7_75t_L g419 ( .A(n_300), .B(n_420), .Y(n_419) );
AND2x2_ASAP7_75t_L g436 ( .A(n_300), .B(n_386), .Y(n_436) );
AND2x2_ASAP7_75t_L g491 ( .A(n_300), .B(n_385), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_303), .B(n_304), .Y(n_302) );
INVx4_ASAP7_75t_L g358 ( .A(n_303), .Y(n_358) );
AND2x2_ASAP7_75t_L g368 ( .A(n_303), .B(n_369), .Y(n_368) );
INVx1_ASAP7_75t_L g304 ( .A(n_305), .Y(n_304) );
BUFx2_ASAP7_75t_L g373 ( .A(n_306), .Y(n_373) );
AND2x2_ASAP7_75t_L g382 ( .A(n_306), .B(n_366), .Y(n_382) );
INVx1_ASAP7_75t_L g417 ( .A(n_308), .Y(n_417) );
HB1xp67_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx2_ASAP7_75t_L g338 ( .A(n_309), .Y(n_338) );
INVxp67_ASAP7_75t_L g310 ( .A(n_311), .Y(n_310) );
NAND2xp5_ASAP7_75t_L g431 ( .A(n_311), .B(n_432), .Y(n_431) );
NAND2xp5_ASAP7_75t_L g379 ( .A(n_312), .B(n_380), .Y(n_379) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_314), .B(n_315), .Y(n_313) );
INVx2_ASAP7_75t_L g315 ( .A(n_316), .Y(n_315) );
AOI21xp5_ASAP7_75t_L g317 ( .A1(n_318), .A2(n_321), .B(n_326), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_319), .B(n_358), .Y(n_467) );
INVx2_ASAP7_75t_SL g319 ( .A(n_320), .Y(n_319) );
NAND2xp5_ASAP7_75t_L g321 ( .A(n_322), .B(n_323), .Y(n_321) );
AOI21xp33_ASAP7_75t_SL g330 ( .A1(n_322), .A2(n_331), .B(n_333), .Y(n_330) );
AND2x2_ASAP7_75t_L g477 ( .A(n_322), .B(n_336), .Y(n_477) );
AND2x4_ASAP7_75t_L g340 ( .A(n_323), .B(n_341), .Y(n_340) );
INVx2_ASAP7_75t_SL g374 ( .A(n_323), .Y(n_374) );
NAND2xp5_ASAP7_75t_SL g456 ( .A(n_323), .B(n_390), .Y(n_456) );
INVx2_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g324 ( .A(n_325), .Y(n_324) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
INVx1_ASAP7_75t_L g331 ( .A(n_332), .Y(n_331) );
AOI21xp33_ASAP7_75t_L g333 ( .A1(n_334), .A2(n_339), .B(n_344), .Y(n_333) );
INVx1_ASAP7_75t_L g334 ( .A(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g335 ( .A(n_336), .B(n_337), .Y(n_335) );
HB1xp67_ASAP7_75t_L g393 ( .A(n_336), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g415 ( .A(n_336), .B(n_341), .Y(n_415) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_337), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_L g399 ( .A(n_337), .Y(n_399) );
INVx1_ASAP7_75t_L g403 ( .A(n_337), .Y(n_403) );
AND2x2_ASAP7_75t_L g487 ( .A(n_337), .B(n_455), .Y(n_487) );
AND2x2_ASAP7_75t_L g490 ( .A(n_337), .B(n_407), .Y(n_490) );
INVx3_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
INVx1_ASAP7_75t_L g339 ( .A(n_340), .Y(n_339) );
AND2x4_ASAP7_75t_SL g341 ( .A(n_342), .B(n_343), .Y(n_341) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_342), .B(n_366), .Y(n_365) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
AND2x4_ASAP7_75t_L g345 ( .A(n_346), .B(n_348), .Y(n_345) );
INVx1_ASAP7_75t_L g469 ( .A(n_346), .Y(n_469) );
AND2x2_ASAP7_75t_L g360 ( .A(n_347), .B(n_361), .Y(n_360) );
NOR2xp33_ASAP7_75t_L g520 ( .A(n_350), .B(n_428), .Y(n_520) );
INVxp67_ASAP7_75t_L g522 ( .A(n_350), .Y(n_522) );
NAND4xp75_ASAP7_75t_L g350 ( .A(n_351), .B(n_370), .C(n_391), .D(n_409), .Y(n_350) );
AND2x2_ASAP7_75t_L g351 ( .A(n_352), .B(n_362), .Y(n_351) );
AND2x2_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
NAND2x1p5_ASAP7_75t_L g440 ( .A(n_354), .B(n_441), .Y(n_440) );
NAND2x1p5_ASAP7_75t_L g426 ( .A(n_355), .B(n_420), .Y(n_426) );
NAND2xp5_ASAP7_75t_R g442 ( .A(n_358), .B(n_443), .Y(n_442) );
INVx2_ASAP7_75t_L g492 ( .A(n_358), .Y(n_492) );
INVx2_ASAP7_75t_L g405 ( .A(n_360), .Y(n_405) );
BUFx3_ASAP7_75t_L g397 ( .A(n_361), .Y(n_397) );
INVx2_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
BUFx2_ASAP7_75t_L g364 ( .A(n_365), .Y(n_364) );
INVx2_ASAP7_75t_L g448 ( .A(n_366), .Y(n_448) );
AND2x2_ASAP7_75t_L g402 ( .A(n_368), .B(n_403), .Y(n_402) );
INVx1_ASAP7_75t_L g424 ( .A(n_369), .Y(n_424) );
AOI21xp5_ASAP7_75t_L g370 ( .A1(n_371), .A2(n_375), .B(n_377), .Y(n_370) );
AND2x2_ASAP7_75t_L g371 ( .A(n_372), .B(n_374), .Y(n_371) );
INVx1_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_373), .B(n_407), .Y(n_406) );
NOR2xp33_ASAP7_75t_L g394 ( .A(n_374), .B(n_395), .Y(n_394) );
INVx1_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
HB1xp67_ASAP7_75t_L g471 ( .A(n_376), .Y(n_471) );
OAI22xp5_ASAP7_75t_L g377 ( .A1(n_378), .A2(n_381), .B1(n_383), .B2(n_387), .Y(n_377) );
HB1xp67_ASAP7_75t_L g378 ( .A(n_379), .Y(n_378) );
INVx1_ASAP7_75t_SL g383 ( .A(n_384), .Y(n_383) );
OA21x2_ASAP7_75t_L g392 ( .A1(n_385), .A2(n_393), .B(n_394), .Y(n_392) );
INVx1_ASAP7_75t_L g413 ( .A(n_385), .Y(n_413) );
INVx2_ASAP7_75t_L g385 ( .A(n_386), .Y(n_385) );
AND2x2_ASAP7_75t_L g444 ( .A(n_386), .B(n_445), .Y(n_444) );
INVx1_ASAP7_75t_L g452 ( .A(n_386), .Y(n_452) );
NAND2xp5_ASAP7_75t_L g446 ( .A(n_387), .B(n_447), .Y(n_446) );
INVx2_ASAP7_75t_L g387 ( .A(n_388), .Y(n_387) );
AND2x2_ASAP7_75t_L g422 ( .A(n_390), .B(n_423), .Y(n_422) );
AOI21xp5_ASAP7_75t_L g391 ( .A1(n_392), .A2(n_398), .B(n_400), .Y(n_391) );
INVx2_ASAP7_75t_L g395 ( .A(n_396), .Y(n_395) );
OR2x2_ASAP7_75t_L g439 ( .A(n_396), .B(n_440), .Y(n_439) );
INVx3_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx2_ASAP7_75t_L g401 ( .A(n_402), .Y(n_401) );
HB1xp67_ASAP7_75t_L g451 ( .A(n_403), .Y(n_451) );
INVx2_ASAP7_75t_SL g443 ( .A(n_407), .Y(n_443) );
AND2x2_ASAP7_75t_L g409 ( .A(n_410), .B(n_421), .Y(n_409) );
AOI22xp5_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_414), .B1(n_416), .B2(n_419), .Y(n_410) );
INVx1_ASAP7_75t_L g411 ( .A(n_412), .Y(n_411) );
INVx1_ASAP7_75t_L g414 ( .A(n_415), .Y(n_414) );
INVx1_ASAP7_75t_L g472 ( .A(n_416), .Y(n_472) );
NOR2x1_ASAP7_75t_L g416 ( .A(n_417), .B(n_418), .Y(n_416) );
INVx3_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
NOR2xp33_ASAP7_75t_L g427 ( .A(n_428), .B(n_464), .Y(n_427) );
INVxp67_ASAP7_75t_L g526 ( .A(n_428), .Y(n_526) );
NAND3xp33_ASAP7_75t_L g428 ( .A(n_429), .B(n_437), .C(n_449), .Y(n_428) );
NOR2x1_ASAP7_75t_L g429 ( .A(n_430), .B(n_434), .Y(n_429) );
INVx1_ASAP7_75t_L g430 ( .A(n_431), .Y(n_430) );
BUFx2_ASAP7_75t_L g432 ( .A(n_433), .Y(n_432) );
AND2x2_ASAP7_75t_L g434 ( .A(n_435), .B(n_436), .Y(n_434) );
AOI22xp33_ASAP7_75t_SL g437 ( .A1(n_438), .A2(n_442), .B1(n_444), .B2(n_446), .Y(n_437) );
INVx1_ASAP7_75t_L g438 ( .A(n_439), .Y(n_438) );
NOR3xp33_ASAP7_75t_L g449 ( .A(n_450), .B(n_453), .C(n_460), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g453 ( .A1(n_454), .A2(n_457), .B(n_458), .Y(n_453) );
NAND2xp5_ASAP7_75t_L g454 ( .A(n_455), .B(n_456), .Y(n_454) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
NOR2xp33_ASAP7_75t_L g460 ( .A(n_461), .B(n_462), .Y(n_460) );
INVxp67_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g464 ( .A(n_465), .B(n_483), .Y(n_464) );
NOR3xp33_ASAP7_75t_L g465 ( .A(n_466), .B(n_473), .C(n_480), .Y(n_465) );
OAI22xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_468), .B1(n_471), .B2(n_472), .Y(n_466) );
OR2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_470), .Y(n_468) );
NOR3xp33_ASAP7_75t_L g480 ( .A(n_474), .B(n_479), .C(n_481), .Y(n_480) );
INVx1_ASAP7_75t_L g476 ( .A(n_477), .Y(n_476) );
INVx1_ASAP7_75t_L g478 ( .A(n_479), .Y(n_478) );
INVxp67_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
AOI222xp33_ASAP7_75t_L g483 ( .A1(n_484), .A2(n_487), .B1(n_488), .B2(n_490), .C1(n_491), .C2(n_492), .Y(n_483) );
INVx1_ASAP7_75t_SL g485 ( .A(n_486), .Y(n_485) );
INVx2_ASAP7_75t_SL g488 ( .A(n_489), .Y(n_488) );
INVx1_ASAP7_75t_L g493 ( .A(n_494), .Y(n_493) );
NOR2x1_ASAP7_75t_R g498 ( .A(n_499), .B(n_506), .Y(n_498) );
BUFx3_ASAP7_75t_L g828 ( .A(n_499), .Y(n_828) );
NAND2xp5_ASAP7_75t_L g499 ( .A(n_500), .B(n_501), .Y(n_499) );
OR2x2_ASAP7_75t_L g514 ( .A(n_500), .B(n_502), .Y(n_514) );
AND2x6_ASAP7_75t_SL g530 ( .A(n_500), .B(n_502), .Y(n_530) );
OR2x6_ASAP7_75t_SL g814 ( .A(n_500), .B(n_501), .Y(n_814) );
CKINVDCx5p33_ASAP7_75t_R g501 ( .A(n_502), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g503 ( .A(n_504), .B(n_505), .Y(n_503) );
HB1xp67_ASAP7_75t_L g510 ( .A(n_506), .Y(n_510) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_508), .B(n_516), .Y(n_507) );
NOR2xp33_ASAP7_75t_L g508 ( .A(n_509), .B(n_511), .Y(n_508) );
CKINVDCx20_ASAP7_75t_R g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_SL g511 ( .A(n_512), .B(n_515), .Y(n_511) );
INVx1_ASAP7_75t_SL g512 ( .A(n_513), .Y(n_512) );
INVx2_ASAP7_75t_L g513 ( .A(n_514), .Y(n_513) );
AOI22xp5_ASAP7_75t_L g516 ( .A1(n_517), .A2(n_815), .B1(n_822), .B2(n_823), .Y(n_516) );
OAI22xp5_ASAP7_75t_L g517 ( .A1(n_518), .A2(n_527), .B1(n_531), .B2(n_812), .Y(n_517) );
AO22x2_ASAP7_75t_L g823 ( .A1(n_518), .A2(n_528), .B1(n_531), .B2(n_813), .Y(n_823) );
AOI211x1_ASAP7_75t_L g518 ( .A1(n_519), .A2(n_520), .B(n_521), .C(n_524), .Y(n_518) );
INVx4_ASAP7_75t_SL g527 ( .A(n_528), .Y(n_527) );
INVx3_ASAP7_75t_SL g528 ( .A(n_529), .Y(n_528) );
CKINVDCx5p33_ASAP7_75t_R g529 ( .A(n_530), .Y(n_529) );
INVx3_ASAP7_75t_SL g531 ( .A(n_532), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_533), .B(n_742), .Y(n_532) );
NOR4xp25_ASAP7_75t_SL g533 ( .A(n_534), .B(n_635), .C(n_679), .D(n_706), .Y(n_533) );
OAI221xp5_ASAP7_75t_L g534 ( .A1(n_535), .A2(n_598), .B1(n_608), .B2(n_623), .C(n_625), .Y(n_534) );
AOI32xp33_ASAP7_75t_L g535 ( .A1(n_536), .A2(n_565), .A3(n_572), .B1(n_583), .B2(n_594), .Y(n_535) );
NOR2xp33_ASAP7_75t_L g777 ( .A(n_536), .B(n_778), .Y(n_777) );
AOI22xp5_ASAP7_75t_L g805 ( .A1(n_536), .A2(n_748), .B1(n_806), .B2(n_809), .Y(n_805) );
AND2x4_ASAP7_75t_SL g536 ( .A(n_537), .B(n_547), .Y(n_536) );
INVx5_ASAP7_75t_L g597 ( .A(n_537), .Y(n_597) );
OR2x2_ASAP7_75t_L g624 ( .A(n_537), .B(n_596), .Y(n_624) );
AND2x4_ASAP7_75t_L g626 ( .A(n_537), .B(n_557), .Y(n_626) );
INVx2_ASAP7_75t_L g641 ( .A(n_537), .Y(n_641) );
OR2x2_ASAP7_75t_L g653 ( .A(n_537), .B(n_566), .Y(n_653) );
AND2x2_ASAP7_75t_L g660 ( .A(n_537), .B(n_556), .Y(n_660) );
AND2x2_ASAP7_75t_SL g702 ( .A(n_537), .B(n_585), .Y(n_702) );
HB1xp67_ASAP7_75t_L g759 ( .A(n_537), .Y(n_759) );
OR2x6_ASAP7_75t_L g537 ( .A(n_538), .B(n_539), .Y(n_537) );
INVx3_ASAP7_75t_SL g654 ( .A(n_547), .Y(n_654) );
AND2x2_ASAP7_75t_L g673 ( .A(n_547), .B(n_597), .Y(n_673) );
AOI32xp33_ASAP7_75t_L g788 ( .A1(n_547), .A2(n_659), .A3(n_689), .B1(n_719), .B2(n_754), .Y(n_788) );
AND2x4_ASAP7_75t_L g547 ( .A(n_548), .B(n_556), .Y(n_547) );
AND2x2_ASAP7_75t_L g628 ( .A(n_548), .B(n_566), .Y(n_628) );
OR2x2_ASAP7_75t_L g644 ( .A(n_548), .B(n_557), .Y(n_644) );
INVx1_ASAP7_75t_L g667 ( .A(n_548), .Y(n_667) );
INVx2_ASAP7_75t_L g683 ( .A(n_548), .Y(n_683) );
AND2x2_ASAP7_75t_L g720 ( .A(n_548), .B(n_585), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g739 ( .A(n_548), .B(n_557), .Y(n_739) );
HB1xp67_ASAP7_75t_L g808 ( .A(n_548), .Y(n_808) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_554), .Y(n_549) );
INVx2_ASAP7_75t_L g556 ( .A(n_557), .Y(n_556) );
AND2x2_ASAP7_75t_L g775 ( .A(n_557), .B(n_566), .Y(n_775) );
HB1xp67_ASAP7_75t_L g797 ( .A(n_557), .Y(n_797) );
NAND2xp5_ASAP7_75t_L g558 ( .A(n_559), .B(n_563), .Y(n_558) );
OR2x2_ASAP7_75t_L g623 ( .A(n_565), .B(n_624), .Y(n_623) );
AND2x2_ASAP7_75t_L g629 ( .A(n_565), .B(n_630), .Y(n_629) );
AND2x2_ASAP7_75t_L g642 ( .A(n_565), .B(n_643), .Y(n_642) );
AND2x2_ASAP7_75t_L g804 ( .A(n_565), .B(n_673), .Y(n_804) );
BUFx2_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AND2x2_ASAP7_75t_L g733 ( .A(n_566), .B(n_683), .Y(n_733) );
INVx2_ASAP7_75t_L g566 ( .A(n_567), .Y(n_566) );
BUFx6f_ASAP7_75t_L g585 ( .A(n_567), .Y(n_585) );
NAND2xp5_ASAP7_75t_L g568 ( .A(n_569), .B(n_570), .Y(n_568) );
NOR2xp33_ASAP7_75t_L g802 ( .A(n_572), .B(n_700), .Y(n_802) );
INVx1_ASAP7_75t_L g572 ( .A(n_573), .Y(n_572) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_573), .B(n_750), .Y(n_749) );
HB1xp67_ASAP7_75t_L g573 ( .A(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g587 ( .A(n_574), .B(n_588), .Y(n_587) );
INVx1_ASAP7_75t_L g609 ( .A(n_574), .Y(n_609) );
AND2x2_ASAP7_75t_L g633 ( .A(n_574), .B(n_634), .Y(n_633) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_574), .B(n_611), .Y(n_649) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_574), .B(n_671), .Y(n_670) );
INVx2_ASAP7_75t_L g691 ( .A(n_574), .Y(n_691) );
OR2x2_ASAP7_75t_L g710 ( .A(n_574), .B(n_637), .Y(n_710) );
INVx1_ASAP7_75t_L g717 ( .A(n_574), .Y(n_717) );
NOR2xp33_ASAP7_75t_R g769 ( .A(n_574), .B(n_600), .Y(n_769) );
NAND2xp5_ASAP7_75t_L g773 ( .A(n_574), .B(n_612), .Y(n_773) );
INVx3_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
NAND2xp5_ASAP7_75t_L g576 ( .A(n_577), .B(n_581), .Y(n_576) );
AOI32xp33_ASAP7_75t_L g796 ( .A1(n_583), .A2(n_632), .A3(n_797), .B1(n_798), .B2(n_799), .Y(n_796) );
INVx3_ASAP7_75t_L g583 ( .A(n_584), .Y(n_583) );
OR2x2_ASAP7_75t_L g584 ( .A(n_585), .B(n_586), .Y(n_584) );
INVx2_ASAP7_75t_L g663 ( .A(n_585), .Y(n_663) );
AND2x4_ASAP7_75t_L g682 ( .A(n_585), .B(n_683), .Y(n_682) );
NOR2xp33_ASAP7_75t_L g711 ( .A(n_585), .B(n_654), .Y(n_711) );
OR2x2_ASAP7_75t_L g765 ( .A(n_585), .B(n_766), .Y(n_765) );
OR2x2_ASAP7_75t_L g723 ( .A(n_586), .B(n_724), .Y(n_723) );
OR2x2_ASAP7_75t_L g781 ( .A(n_586), .B(n_782), .Y(n_781) );
INVx2_ASAP7_75t_L g586 ( .A(n_587), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g747 ( .A(n_587), .B(n_600), .Y(n_747) );
AND2x2_ASAP7_75t_L g784 ( .A(n_587), .B(n_750), .Y(n_784) );
INVx2_ASAP7_75t_L g634 ( .A(n_588), .Y(n_634) );
INVx2_ASAP7_75t_L g637 ( .A(n_588), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g657 ( .A(n_588), .B(n_600), .Y(n_657) );
INVx1_ASAP7_75t_L g688 ( .A(n_588), .Y(n_688) );
OR2x2_ASAP7_75t_L g714 ( .A(n_588), .B(n_600), .Y(n_714) );
HB1xp67_ASAP7_75t_L g766 ( .A(n_588), .Y(n_766) );
BUFx3_ASAP7_75t_L g795 ( .A(n_588), .Y(n_795) );
HB1xp67_ASAP7_75t_L g594 ( .A(n_595), .Y(n_594) );
INVx2_ASAP7_75t_L g664 ( .A(n_595), .Y(n_664) );
NAND2xp5_ASAP7_75t_L g725 ( .A(n_595), .B(n_682), .Y(n_725) );
NAND2xp5_ASAP7_75t_L g752 ( .A(n_595), .B(n_753), .Y(n_752) );
AND2x4_ASAP7_75t_L g595 ( .A(n_596), .B(n_597), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g666 ( .A(n_596), .B(n_667), .Y(n_666) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_596), .A2(n_663), .B(n_681), .Y(n_696) );
OAI32xp33_ASAP7_75t_L g718 ( .A1(n_597), .A2(n_719), .A3(n_721), .B1(n_723), .B2(n_725), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g791 ( .A(n_597), .B(n_682), .Y(n_791) );
HB1xp67_ASAP7_75t_L g598 ( .A(n_599), .Y(n_598) );
INVx1_ASAP7_75t_L g724 ( .A(n_599), .Y(n_724) );
NOR2x1p5_ASAP7_75t_L g794 ( .A(n_599), .B(n_795), .Y(n_794) );
INVx2_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x4_ASAP7_75t_L g610 ( .A(n_600), .B(n_611), .Y(n_610) );
AND2x4_ASAP7_75t_SL g632 ( .A(n_600), .B(n_612), .Y(n_632) );
OR2x2_ASAP7_75t_L g636 ( .A(n_600), .B(n_637), .Y(n_636) );
INVx2_ASAP7_75t_L g671 ( .A(n_600), .Y(n_671) );
AND2x2_ASAP7_75t_L g689 ( .A(n_600), .B(n_690), .Y(n_689) );
OR2x2_ASAP7_75t_L g700 ( .A(n_600), .B(n_612), .Y(n_700) );
OR2x2_ASAP7_75t_L g762 ( .A(n_600), .B(n_763), .Y(n_762) );
OR2x2_ASAP7_75t_L g779 ( .A(n_600), .B(n_710), .Y(n_779) );
INVx1_ASAP7_75t_L g811 ( .A(n_600), .Y(n_811) );
OR2x6_ASAP7_75t_L g600 ( .A(n_601), .B(n_607), .Y(n_600) );
NAND2xp5_ASAP7_75t_L g608 ( .A(n_609), .B(n_610), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g763 ( .A(n_609), .B(n_688), .Y(n_763) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_610), .B(n_722), .Y(n_721) );
AOI222xp33_ASAP7_75t_L g726 ( .A1(n_610), .A2(n_727), .B1(n_732), .B2(n_734), .C1(n_737), .C2(n_740), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_610), .B(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g754 ( .A(n_610), .B(n_633), .Y(n_754) );
AND2x2_ASAP7_75t_L g716 ( .A(n_611), .B(n_717), .Y(n_716) );
OR2x2_ASAP7_75t_L g731 ( .A(n_611), .B(n_636), .Y(n_731) );
INVx3_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g669 ( .A(n_612), .B(n_637), .Y(n_669) );
AND2x4_ASAP7_75t_L g690 ( .A(n_612), .B(n_691), .Y(n_690) );
AND2x2_ASAP7_75t_L g750 ( .A(n_612), .B(n_671), .Y(n_750) );
AND2x4_ASAP7_75t_L g612 ( .A(n_613), .B(n_618), .Y(n_612) );
INVx1_ASAP7_75t_SL g630 ( .A(n_624), .Y(n_630) );
NAND2xp33_ASAP7_75t_SL g799 ( .A(n_624), .B(n_654), .Y(n_799) );
A2O1A1Ixp33_ASAP7_75t_L g625 ( .A1(n_626), .A2(n_627), .B(n_629), .C(n_631), .Y(n_625) );
INVx2_ASAP7_75t_SL g676 ( .A(n_626), .Y(n_676) );
AND2x2_ASAP7_75t_L g680 ( .A(n_627), .B(n_681), .Y(n_680) );
INVx1_ASAP7_75t_L g627 ( .A(n_628), .Y(n_627) );
NAND2xp5_ASAP7_75t_L g675 ( .A(n_628), .B(n_676), .Y(n_675) );
O2A1O1Ixp33_ASAP7_75t_L g701 ( .A1(n_628), .A2(n_666), .B(n_702), .C(n_703), .Y(n_701) );
AND2x2_ASAP7_75t_L g778 ( .A(n_628), .B(n_759), .Y(n_778) );
AND2x2_ASAP7_75t_L g631 ( .A(n_632), .B(n_633), .Y(n_631) );
AND2x4_ASAP7_75t_L g677 ( .A(n_632), .B(n_678), .Y(n_677) );
INVx1_ASAP7_75t_SL g782 ( .A(n_632), .Y(n_782) );
OAI211xp5_ASAP7_75t_L g635 ( .A1(n_636), .A2(n_638), .B(n_645), .C(n_672), .Y(n_635) );
INVx2_ASAP7_75t_L g647 ( .A(n_636), .Y(n_647) );
OR2x2_ASAP7_75t_L g694 ( .A(n_636), .B(n_695), .Y(n_694) );
HB1xp67_ASAP7_75t_L g678 ( .A(n_637), .Y(n_678) );
INVx1_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
AND2x2_ASAP7_75t_L g639 ( .A(n_640), .B(n_642), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g681 ( .A(n_640), .B(n_682), .Y(n_681) );
AND2x2_ASAP7_75t_L g732 ( .A(n_640), .B(n_733), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g786 ( .A(n_640), .B(n_720), .Y(n_786) );
INVx2_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AOI222xp33_ASAP7_75t_L g744 ( .A1(n_642), .A2(n_745), .B1(n_746), .B2(n_748), .C1(n_751), .C2(n_754), .Y(n_744) );
AOI221xp5_ASAP7_75t_L g707 ( .A1(n_643), .A2(n_708), .B1(n_711), .B2(n_712), .C(n_718), .Y(n_707) );
AND2x2_ASAP7_75t_L g745 ( .A(n_643), .B(n_702), .Y(n_745) );
INVx2_ASAP7_75t_L g643 ( .A(n_644), .Y(n_643) );
NAND2xp33_ASAP7_75t_SL g658 ( .A(n_644), .B(n_659), .Y(n_658) );
AOI221x1_ASAP7_75t_L g645 ( .A1(n_646), .A2(n_650), .B1(n_655), .B2(n_658), .C(n_661), .Y(n_645) );
AND2x4_ASAP7_75t_L g646 ( .A(n_647), .B(n_648), .Y(n_646) );
AND2x2_ASAP7_75t_L g798 ( .A(n_648), .B(n_736), .Y(n_798) );
INVx1_ASAP7_75t_L g648 ( .A(n_649), .Y(n_648) );
OR2x2_ASAP7_75t_L g656 ( .A(n_649), .B(n_657), .Y(n_656) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_652), .B(n_654), .Y(n_651) );
INVx1_ASAP7_75t_SL g652 ( .A(n_653), .Y(n_652) );
OAI32xp33_ASAP7_75t_L g764 ( .A1(n_654), .A2(n_695), .A3(n_765), .B1(n_767), .B2(n_771), .Y(n_764) );
OAI21xp33_ASAP7_75t_SL g783 ( .A1(n_655), .A2(n_784), .B(n_785), .Y(n_783) );
INVx2_ASAP7_75t_L g655 ( .A(n_656), .Y(n_655) );
INVx2_ASAP7_75t_L g659 ( .A(n_660), .Y(n_659) );
AOI21xp33_ASAP7_75t_L g661 ( .A1(n_662), .A2(n_665), .B(n_668), .Y(n_661) );
OR2x2_ASAP7_75t_L g662 ( .A(n_663), .B(n_664), .Y(n_662) );
OR2x2_ASAP7_75t_L g665 ( .A(n_663), .B(n_666), .Y(n_665) );
OR2x2_ASAP7_75t_L g738 ( .A(n_663), .B(n_739), .Y(n_738) );
AOI221xp5_ASAP7_75t_L g692 ( .A1(n_667), .A2(n_693), .B1(n_696), .B2(n_697), .C(n_701), .Y(n_692) );
INVx1_ASAP7_75t_L g768 ( .A(n_667), .Y(n_768) );
HB1xp67_ASAP7_75t_L g774 ( .A(n_667), .Y(n_774) );
OR2x2_ASAP7_75t_L g668 ( .A(n_669), .B(n_670), .Y(n_668) );
OAI21xp33_ASAP7_75t_L g672 ( .A1(n_673), .A2(n_674), .B(n_677), .Y(n_672) );
INVx1_ASAP7_75t_L g674 ( .A(n_675), .Y(n_674) );
NOR2xp33_ASAP7_75t_L g740 ( .A(n_676), .B(n_741), .Y(n_740) );
OAI21xp5_ASAP7_75t_SL g679 ( .A1(n_680), .A2(n_684), .B(n_692), .Y(n_679) );
HB1xp67_ASAP7_75t_L g753 ( .A(n_683), .Y(n_753) );
INVx1_ASAP7_75t_L g684 ( .A(n_685), .Y(n_684) );
AND2x2_ASAP7_75t_L g685 ( .A(n_686), .B(n_689), .Y(n_685) );
NAND2xp5_ASAP7_75t_L g698 ( .A(n_686), .B(n_699), .Y(n_698) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVxp67_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
INVx1_ASAP7_75t_L g705 ( .A(n_688), .Y(n_705) );
INVx1_ASAP7_75t_L g695 ( .A(n_690), .Y(n_695) );
AND2x2_ASAP7_75t_SL g704 ( .A(n_690), .B(n_705), .Y(n_704) );
NAND2xp5_ASAP7_75t_L g735 ( .A(n_690), .B(n_736), .Y(n_735) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_690), .B(n_811), .Y(n_810) );
INVx1_ASAP7_75t_L g693 ( .A(n_694), .Y(n_693) );
INVx1_ASAP7_75t_SL g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g699 ( .A(n_700), .Y(n_699) );
OR2x2_ASAP7_75t_L g709 ( .A(n_700), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g703 ( .A(n_704), .Y(n_703) );
HB1xp67_ASAP7_75t_L g770 ( .A(n_705), .Y(n_770) );
NAND2xp5_ASAP7_75t_SL g706 ( .A(n_707), .B(n_726), .Y(n_706) );
INVx1_ASAP7_75t_L g708 ( .A(n_709), .Y(n_708) );
INVx1_ASAP7_75t_L g722 ( .A(n_710), .Y(n_722) );
INVx1_ASAP7_75t_SL g712 ( .A(n_713), .Y(n_712) );
OR2x2_ASAP7_75t_L g713 ( .A(n_714), .B(n_715), .Y(n_713) );
INVx1_ASAP7_75t_SL g736 ( .A(n_714), .Y(n_736) );
INVx1_ASAP7_75t_SL g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g793 ( .A(n_716), .B(n_794), .Y(n_793) );
HB1xp67_ASAP7_75t_L g730 ( .A(n_717), .Y(n_730) );
BUFx2_ASAP7_75t_L g719 ( .A(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_SL g727 ( .A(n_728), .B(n_731), .Y(n_727) );
INVxp67_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
INVx1_ASAP7_75t_L g741 ( .A(n_733), .Y(n_741) );
INVx1_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
INVx1_ASAP7_75t_SL g737 ( .A(n_738), .Y(n_737) );
INVx1_ASAP7_75t_L g760 ( .A(n_739), .Y(n_760) );
NOR4xp25_ASAP7_75t_L g742 ( .A(n_743), .B(n_776), .C(n_787), .D(n_800), .Y(n_742) );
NAND2xp5_ASAP7_75t_L g743 ( .A(n_744), .B(n_755), .Y(n_743) );
O2A1O1Ixp33_ASAP7_75t_L g755 ( .A1(n_745), .A2(n_756), .B(n_761), .C(n_764), .Y(n_755) );
INVx1_ASAP7_75t_SL g746 ( .A(n_747), .Y(n_746) );
INVx1_ASAP7_75t_L g748 ( .A(n_749), .Y(n_748) );
INVx1_ASAP7_75t_L g751 ( .A(n_752), .Y(n_751) );
INVx2_ASAP7_75t_L g756 ( .A(n_757), .Y(n_756) );
NAND2xp5_ASAP7_75t_SL g757 ( .A(n_758), .B(n_760), .Y(n_757) );
OAI211xp5_ASAP7_75t_L g767 ( .A1(n_758), .A2(n_768), .B(n_769), .C(n_770), .Y(n_767) );
INVx1_ASAP7_75t_L g758 ( .A(n_759), .Y(n_758) );
INVx1_ASAP7_75t_SL g761 ( .A(n_762), .Y(n_761) );
OAI21xp33_ASAP7_75t_SL g771 ( .A1(n_772), .A2(n_774), .B(n_775), .Y(n_771) );
INVx1_ASAP7_75t_L g772 ( .A(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_SL g806 ( .A(n_775), .B(n_807), .Y(n_806) );
OAI221xp5_ASAP7_75t_SL g776 ( .A1(n_777), .A2(n_779), .B1(n_780), .B2(n_781), .C(n_783), .Y(n_776) );
INVx1_ASAP7_75t_SL g780 ( .A(n_778), .Y(n_780) );
INVx1_ASAP7_75t_L g785 ( .A(n_786), .Y(n_785) );
NAND3xp33_ASAP7_75t_SL g787 ( .A(n_788), .B(n_789), .C(n_796), .Y(n_787) );
NAND2xp5_ASAP7_75t_L g789 ( .A(n_790), .B(n_792), .Y(n_789) );
INVx1_ASAP7_75t_L g790 ( .A(n_791), .Y(n_790) );
INVx1_ASAP7_75t_L g792 ( .A(n_793), .Y(n_792) );
OAI21xp33_ASAP7_75t_L g800 ( .A1(n_801), .A2(n_803), .B(n_805), .Y(n_800) );
INVx1_ASAP7_75t_L g801 ( .A(n_802), .Y(n_801) );
INVxp33_ASAP7_75t_L g803 ( .A(n_804), .Y(n_803) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
INVx1_ASAP7_75t_SL g809 ( .A(n_810), .Y(n_809) );
CKINVDCx20_ASAP7_75t_R g812 ( .A(n_813), .Y(n_812) );
CKINVDCx11_ASAP7_75t_R g813 ( .A(n_814), .Y(n_813) );
INVx1_ASAP7_75t_L g822 ( .A(n_815), .Y(n_822) );
CKINVDCx20_ASAP7_75t_R g817 ( .A(n_818), .Y(n_817) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_825), .B(n_826), .Y(n_824) );
CKINVDCx11_ASAP7_75t_R g826 ( .A(n_827), .Y(n_826) );
CKINVDCx20_ASAP7_75t_R g827 ( .A(n_828), .Y(n_827) );
INVx1_ASAP7_75t_SL g829 ( .A(n_830), .Y(n_829) );
CKINVDCx20_ASAP7_75t_R g830 ( .A(n_831), .Y(n_830) );
BUFx2_ASAP7_75t_L g831 ( .A(n_832), .Y(n_831) );
INVx1_ASAP7_75t_L g832 ( .A(n_833), .Y(n_832) );
INVx2_ASAP7_75t_L g843 ( .A(n_833), .Y(n_843) );
OR2x2_ASAP7_75t_SL g833 ( .A(n_834), .B(n_836), .Y(n_833) );
CKINVDCx16_ASAP7_75t_R g834 ( .A(n_835), .Y(n_834) );
INVx1_ASAP7_75t_L g836 ( .A(n_837), .Y(n_836) );
NOR2xp33_ASAP7_75t_L g841 ( .A(n_842), .B(n_843), .Y(n_841) );
endmodule