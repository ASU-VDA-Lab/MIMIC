module fake_jpeg_634_n_127 (n_13, n_21, n_33, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_34, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_127);

input n_13;
input n_21;
input n_33;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_34;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_127;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_103;
wire n_50;
wire n_124;
wire n_57;
wire n_119;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_109;
wire n_113;
wire n_106;
wire n_111;
wire n_44;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_54;
wire n_91;
wire n_93;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_100;
wire n_118;
wire n_82;
wire n_96;

INVx1_ASAP7_75t_SL g35 ( 
.A(n_34),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_0),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_10),
.Y(n_37)
);

INVx2_ASAP7_75t_L g38 ( 
.A(n_27),
.Y(n_38)
);

INVx13_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

BUFx3_ASAP7_75t_L g40 ( 
.A(n_21),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_4),
.Y(n_41)
);

CKINVDCx20_ASAP7_75t_R g42 ( 
.A(n_5),
.Y(n_42)
);

INVx8_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_25),
.Y(n_45)
);

BUFx3_ASAP7_75t_L g46 ( 
.A(n_22),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx2_ASAP7_75t_L g48 ( 
.A(n_40),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g57 ( 
.A(n_48),
.B(n_54),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_47),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_49),
.A2(n_42),
.B1(n_41),
.B2(n_44),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_47),
.B(n_33),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_50),
.B(n_38),
.Y(n_60)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_35),
.B(n_1),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g55 ( 
.A(n_52),
.B(n_53),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_35),
.B(n_2),
.Y(n_53)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_46),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_50),
.B(n_38),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_58),
.Y(n_67)
);

NOR2xp33_ASAP7_75t_L g58 ( 
.A(n_52),
.B(n_36),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g68 ( 
.A(n_60),
.B(n_61),
.Y(n_68)
);

NOR2xp33_ASAP7_75t_L g61 ( 
.A(n_53),
.B(n_36),
.Y(n_61)
);

AOI21xp33_ASAP7_75t_SL g62 ( 
.A1(n_48),
.A2(n_46),
.B(n_45),
.Y(n_62)
);

XNOR2xp5_ASAP7_75t_L g73 ( 
.A(n_62),
.B(n_49),
.Y(n_73)
);

INVx6_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_63),
.Y(n_71)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_64),
.B(n_57),
.Y(n_74)
);

AND2x6_ASAP7_75t_L g65 ( 
.A(n_62),
.B(n_55),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_65),
.B(n_75),
.Y(n_79)
);

OR2x2_ASAP7_75t_L g66 ( 
.A(n_60),
.B(n_54),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_66),
.B(n_70),
.Y(n_85)
);

INVx4_ASAP7_75t_L g69 ( 
.A(n_63),
.Y(n_69)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_69),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_56),
.B(n_55),
.Y(n_70)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_59),
.Y(n_72)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_72),
.Y(n_77)
);

OR2x2_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_76),
.Y(n_78)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_74),
.A2(n_63),
.B(n_39),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_57),
.B(n_44),
.Y(n_75)
);

AND2x2_ASAP7_75t_L g76 ( 
.A(n_57),
.B(n_54),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_68),
.B(n_45),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_80),
.B(n_81),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g81 ( 
.A1(n_73),
.A2(n_59),
.B1(n_51),
.B2(n_42),
.Y(n_81)
);

INVxp67_ASAP7_75t_L g82 ( 
.A(n_76),
.Y(n_82)
);

NAND2xp5_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_84),
.Y(n_98)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_67),
.B(n_51),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g96 ( 
.A(n_83),
.B(n_88),
.C(n_16),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_66),
.Y(n_84)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_71),
.Y(n_87)
);

INVx1_ASAP7_75t_L g93 ( 
.A(n_87),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g88 ( 
.A(n_65),
.B(n_37),
.C(n_41),
.Y(n_88)
);

AOI21x1_ASAP7_75t_L g95 ( 
.A1(n_89),
.A2(n_39),
.B(n_43),
.Y(n_95)
);

CKINVDCx16_ASAP7_75t_R g90 ( 
.A(n_86),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_90),
.B(n_91),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_85),
.B(n_71),
.Y(n_91)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_78),
.B(n_69),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g105 ( 
.A(n_92),
.B(n_100),
.C(n_14),
.Y(n_105)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_77),
.Y(n_94)
);

INVx1_ASAP7_75t_L g112 ( 
.A(n_94),
.Y(n_112)
);

OAI21xp5_ASAP7_75t_SL g107 ( 
.A1(n_95),
.A2(n_6),
.B(n_8),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_96),
.B(n_99),
.Y(n_106)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_83),
.B(n_3),
.Y(n_99)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_78),
.B(n_43),
.C(n_17),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_88),
.B(n_79),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_9),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_81),
.B(n_3),
.Y(n_102)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_102),
.B(n_8),
.Y(n_108)
);

AOI322xp5_ASAP7_75t_L g103 ( 
.A1(n_98),
.A2(n_82),
.A3(n_86),
.B1(n_18),
.B2(n_20),
.C1(n_32),
.C2(n_31),
.Y(n_103)
);

MAJIxp5_ASAP7_75t_L g116 ( 
.A(n_103),
.B(n_105),
.C(n_111),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_97),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_104),
.A2(n_110),
.B1(n_100),
.B2(n_93),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_107),
.B(n_108),
.Y(n_114)
);

AOI21xp5_ASAP7_75t_L g110 ( 
.A1(n_92),
.A2(n_95),
.B(n_96),
.Y(n_110)
);

INVx1_ASAP7_75t_L g113 ( 
.A(n_112),
.Y(n_113)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_113),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g120 ( 
.A(n_115),
.B(n_110),
.C(n_23),
.Y(n_120)
);

AOI22xp5_ASAP7_75t_L g117 ( 
.A1(n_109),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_117)
);

A2O1A1Ixp33_ASAP7_75t_SL g118 ( 
.A1(n_117),
.A2(n_105),
.B(n_106),
.C(n_107),
.Y(n_118)
);

HB1xp67_ASAP7_75t_L g121 ( 
.A(n_118),
.Y(n_121)
);

MAJx2_ASAP7_75t_L g122 ( 
.A(n_120),
.B(n_116),
.C(n_24),
.Y(n_122)
);

AOI21x1_ASAP7_75t_L g123 ( 
.A1(n_122),
.A2(n_121),
.B(n_114),
.Y(n_123)
);

AOI322xp5_ASAP7_75t_L g124 ( 
.A1(n_123),
.A2(n_114),
.A3(n_119),
.B1(n_28),
.B2(n_15),
.C1(n_19),
.C2(n_29),
.Y(n_124)
);

AOI21xp5_ASAP7_75t_L g125 ( 
.A1(n_124),
.A2(n_30),
.B(n_12),
.Y(n_125)
);

NOR3xp33_ASAP7_75t_L g126 ( 
.A(n_125),
.B(n_11),
.C(n_13),
.Y(n_126)
);

FAx1_ASAP7_75t_SL g127 ( 
.A(n_126),
.B(n_13),
.CI(n_116),
.CON(n_127),
.SN(n_127)
);


endmodule