module fake_jpeg_21446_n_136 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_136);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_136;

wire n_117;
wire n_105;
wire n_64;
wire n_55;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_134;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_124;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_81;
wire n_129;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_131;
wire n_56;
wire n_79;
wire n_132;
wire n_133;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_115;
wire n_123;
wire n_112;
wire n_95;
wire n_97;
wire n_135;
wire n_36;
wire n_62;
wire n_120;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_128;
wire n_96;

INVx1_ASAP7_75t_L g13 ( 
.A(n_0),
.Y(n_13)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_10),
.Y(n_14)
);

INVx1_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx16_ASAP7_75t_R g16 ( 
.A(n_3),
.Y(n_16)
);

NOR2xp33_ASAP7_75t_L g17 ( 
.A(n_7),
.B(n_1),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_6),
.Y(n_19)
);

INVx1_ASAP7_75t_L g20 ( 
.A(n_8),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_5),
.Y(n_21)
);

BUFx12_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx24_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

CKINVDCx20_ASAP7_75t_R g24 ( 
.A(n_10),
.Y(n_24)
);

BUFx16f_ASAP7_75t_L g25 ( 
.A(n_12),
.Y(n_25)
);

BUFx4f_ASAP7_75t_L g26 ( 
.A(n_8),
.Y(n_26)
);

INVx3_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx3_ASAP7_75t_L g28 ( 
.A(n_23),
.Y(n_28)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_28),
.Y(n_44)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_23),
.Y(n_29)
);

INVx2_ASAP7_75t_L g49 ( 
.A(n_29),
.Y(n_49)
);

INVx2_ASAP7_75t_L g30 ( 
.A(n_26),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_30),
.B(n_33),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_23),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

AND2x2_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NOR2xp33_ASAP7_75t_SL g41 ( 
.A(n_32),
.B(n_36),
.Y(n_41)
);

NOR2xp33_ASAP7_75t_L g33 ( 
.A(n_14),
.B(n_5),
.Y(n_33)
);

INVx3_ASAP7_75t_L g34 ( 
.A(n_26),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_34),
.B(n_35),
.Y(n_38)
);

CKINVDCx16_ASAP7_75t_R g35 ( 
.A(n_13),
.Y(n_35)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_26),
.B(n_1),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_36),
.B(n_22),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_39),
.B(n_41),
.Y(n_55)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_31),
.Y(n_40)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_40),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_32),
.B(n_14),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_42),
.B(n_43),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_17),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_28),
.B(n_24),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_45),
.B(n_48),
.Y(n_62)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_30),
.A2(n_27),
.B1(n_13),
.B2(n_16),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_46),
.B(n_50),
.Y(n_53)
);

AOI21xp5_ASAP7_75t_L g48 ( 
.A1(n_34),
.A2(n_1),
.B(n_2),
.Y(n_48)
);

AOI22xp5_ASAP7_75t_L g50 ( 
.A1(n_29),
.A2(n_27),
.B1(n_3),
.B2(n_4),
.Y(n_50)
);

AOI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_48),
.A2(n_18),
.B1(n_15),
.B2(n_20),
.Y(n_51)
);

XOR2xp5_ASAP7_75t_L g68 ( 
.A(n_51),
.B(n_50),
.Y(n_68)
);

INVx13_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_54),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g56 ( 
.A(n_39),
.B(n_31),
.Y(n_56)
);

NAND2xp5_ASAP7_75t_L g76 ( 
.A(n_56),
.B(n_65),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_SL g74 ( 
.A(n_57),
.B(n_59),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g58 ( 
.A(n_41),
.B(n_22),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g80 ( 
.A(n_58),
.B(n_25),
.C(n_18),
.Y(n_80)
);

INVxp67_ASAP7_75t_L g59 ( 
.A(n_38),
.Y(n_59)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_47),
.Y(n_61)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_61),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g63 ( 
.A(n_46),
.B(n_24),
.Y(n_63)
);

AND2x2_ASAP7_75t_L g66 ( 
.A(n_63),
.B(n_64),
.Y(n_66)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_38),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g65 ( 
.A(n_37),
.B(n_15),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g84 ( 
.A(n_68),
.B(n_75),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_SL g69 ( 
.A(n_60),
.B(n_43),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_SL g88 ( 
.A(n_69),
.B(n_78),
.Y(n_88)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_57),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_71),
.Y(n_86)
);

BUFx24_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx2_ASAP7_75t_SL g83 ( 
.A(n_72),
.Y(n_83)
);

OA22x2_ASAP7_75t_L g73 ( 
.A1(n_63),
.A2(n_50),
.B1(n_49),
.B2(n_44),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g90 ( 
.A1(n_73),
.A2(n_53),
.B(n_52),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_L g75 ( 
.A1(n_53),
.A2(n_37),
.B1(n_42),
.B2(n_45),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_62),
.B(n_49),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_77),
.B(n_56),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_64),
.B(n_19),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g79 ( 
.A(n_60),
.B(n_19),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_SL g91 ( 
.A(n_79),
.B(n_65),
.Y(n_91)
);

XNOR2xp5_ASAP7_75t_L g82 ( 
.A(n_80),
.B(n_62),
.Y(n_82)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_70),
.Y(n_81)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_81),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_82),
.B(n_85),
.Y(n_97)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_70),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g100 ( 
.A(n_87),
.B(n_90),
.Y(n_100)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_67),
.Y(n_89)
);

INVx1_ASAP7_75t_L g99 ( 
.A(n_89),
.Y(n_99)
);

INVx1_ASAP7_75t_L g103 ( 
.A(n_91),
.Y(n_103)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_76),
.B(n_55),
.Y(n_92)
);

INVx1_ASAP7_75t_L g104 ( 
.A(n_92),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_77),
.A2(n_63),
.B(n_52),
.Y(n_93)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_93),
.A2(n_66),
.B(n_74),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g94 ( 
.A(n_84),
.B(n_80),
.C(n_58),
.Y(n_94)
);

MAJIxp5_ASAP7_75t_L g109 ( 
.A(n_94),
.B(n_102),
.C(n_51),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_93),
.A2(n_73),
.B1(n_68),
.B2(n_76),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_95),
.A2(n_44),
.B1(n_61),
.B2(n_83),
.Y(n_113)
);

AOI21x1_ASAP7_75t_L g98 ( 
.A1(n_87),
.A2(n_73),
.B(n_66),
.Y(n_98)
);

AOI21xp5_ASAP7_75t_L g107 ( 
.A1(n_98),
.A2(n_90),
.B(n_92),
.Y(n_107)
);

XOR2xp5_ASAP7_75t_L g111 ( 
.A(n_101),
.B(n_73),
.Y(n_111)
);

MAJIxp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_66),
.C(n_55),
.Y(n_102)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_96),
.Y(n_105)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_105),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_103),
.B(n_88),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_106),
.B(n_107),
.Y(n_114)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_99),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_108),
.B(n_112),
.Y(n_119)
);

MAJIxp5_ASAP7_75t_L g115 ( 
.A(n_109),
.B(n_110),
.C(n_111),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g110 ( 
.A(n_94),
.B(n_81),
.C(n_86),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_97),
.B(n_71),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_113),
.A2(n_100),
.B1(n_83),
.B2(n_72),
.Y(n_118)
);

AOI322xp5_ASAP7_75t_L g116 ( 
.A1(n_111),
.A2(n_104),
.A3(n_98),
.B1(n_101),
.B2(n_100),
.C1(n_97),
.C2(n_102),
.Y(n_116)
);

AND2x2_ASAP7_75t_L g123 ( 
.A(n_116),
.B(n_72),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g124 ( 
.A(n_118),
.B(n_54),
.Y(n_124)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_113),
.A2(n_110),
.B1(n_109),
.B2(n_83),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_120),
.B(n_86),
.Y(n_121)
);

OAI21xp5_ASAP7_75t_L g126 ( 
.A1(n_121),
.A2(n_124),
.B(n_117),
.Y(n_126)
);

INVxp33_ASAP7_75t_L g122 ( 
.A(n_119),
.Y(n_122)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_122),
.B(n_125),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_123),
.B(n_118),
.C(n_115),
.Y(n_129)
);

AO21x2_ASAP7_75t_L g125 ( 
.A1(n_114),
.A2(n_47),
.B(n_22),
.Y(n_125)
);

AOI322xp5_ASAP7_75t_L g130 ( 
.A1(n_126),
.A2(n_127),
.A3(n_20),
.B1(n_11),
.B2(n_12),
.C1(n_9),
.C2(n_2),
.Y(n_130)
);

NAND4xp25_ASAP7_75t_L g127 ( 
.A(n_125),
.B(n_120),
.C(n_117),
.D(n_115),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_L g132 ( 
.A1(n_129),
.A2(n_25),
.B1(n_21),
.B2(n_4),
.Y(n_132)
);

MAJIxp5_ASAP7_75t_L g133 ( 
.A(n_130),
.B(n_131),
.C(n_132),
.Y(n_133)
);

XOR2xp5_ASAP7_75t_L g131 ( 
.A(n_128),
.B(n_25),
.Y(n_131)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_131),
.B(n_21),
.C(n_3),
.Y(n_134)
);

AOI21xp5_ASAP7_75t_L g135 ( 
.A1(n_134),
.A2(n_2),
.B(n_4),
.Y(n_135)
);

XOR2xp5_ASAP7_75t_L g136 ( 
.A(n_135),
.B(n_133),
.Y(n_136)
);


endmodule