module fake_jpeg_23118_n_17 (n_3, n_2, n_1, n_0, n_4, n_5, n_17);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_17;

wire n_13;
wire n_11;
wire n_14;
wire n_16;
wire n_12;
wire n_10;
wire n_8;
wire n_9;
wire n_15;
wire n_6;
wire n_7;

INVx4_ASAP7_75t_L g6 ( 
.A(n_0),
.Y(n_6)
);

INVx13_ASAP7_75t_L g7 ( 
.A(n_5),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_4),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_1),
.Y(n_9)
);

INVx2_ASAP7_75t_L g10 ( 
.A(n_0),
.Y(n_10)
);

AND2x2_ASAP7_75t_L g11 ( 
.A(n_2),
.B(n_3),
.Y(n_11)
);

AND2x6_ASAP7_75t_L g12 ( 
.A(n_11),
.B(n_1),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g15 ( 
.A(n_12),
.Y(n_15)
);

BUFx12f_ASAP7_75t_SL g13 ( 
.A(n_8),
.Y(n_13)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_9),
.A2(n_2),
.B1(n_10),
.B2(n_6),
.Y(n_14)
);

AOI21xp5_ASAP7_75t_L g16 ( 
.A1(n_15),
.A2(n_13),
.B(n_14),
.Y(n_16)
);

AOI22xp5_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_7),
.B1(n_11),
.B2(n_13),
.Y(n_17)
);


endmodule