module fake_jpeg_21941_n_242 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_242);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_242;

wire n_159;
wire n_117;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_75;
wire n_122;
wire n_37;
wire n_233;
wire n_121;
wire n_99;
wire n_102;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_172;
wire n_173;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_118;
wire n_140;
wire n_82;
wire n_128;
wire n_100;
wire n_96;

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_9),
.Y(n_16)
);

BUFx4f_ASAP7_75t_L g17 ( 
.A(n_7),
.Y(n_17)
);

INVx2_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

BUFx8_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_3),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_14),
.Y(n_23)
);

BUFx8_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_10),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g27 ( 
.A(n_3),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_9),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_8),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_4),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_12),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_6),
.Y(n_34)
);

INVx4_ASAP7_75t_SL g35 ( 
.A(n_17),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_40),
.Y(n_60)
);

INVx2_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_36),
.Y(n_59)
);

INVx11_ASAP7_75t_L g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g49 ( 
.A(n_37),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_17),
.Y(n_38)
);

INVx8_ASAP7_75t_L g65 ( 
.A(n_38),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_17),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

INVx4_ASAP7_75t_SL g40 ( 
.A(n_30),
.Y(n_40)
);

BUFx12_ASAP7_75t_L g41 ( 
.A(n_20),
.Y(n_41)
);

INVx5_ASAP7_75t_L g48 ( 
.A(n_41),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g42 ( 
.A(n_16),
.B(n_34),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g50 ( 
.A(n_42),
.B(n_34),
.Y(n_50)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_20),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g63 ( 
.A(n_44),
.B(n_47),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_20),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_45),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g46 ( 
.A(n_19),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g76 ( 
.A(n_46),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_23),
.B(n_0),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_50),
.B(n_51),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_16),
.Y(n_51)
);

INVx3_ASAP7_75t_L g52 ( 
.A(n_37),
.Y(n_52)
);

NOR2xp33_ASAP7_75t_L g82 ( 
.A(n_52),
.B(n_53),
.Y(n_82)
);

CKINVDCx5p33_ASAP7_75t_R g53 ( 
.A(n_44),
.Y(n_53)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_41),
.Y(n_54)
);

INVx6_ASAP7_75t_L g93 ( 
.A(n_54),
.Y(n_93)
);

AOI22xp33_ASAP7_75t_SL g55 ( 
.A1(n_35),
.A2(n_18),
.B1(n_29),
.B2(n_28),
.Y(n_55)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_55),
.A2(n_56),
.B1(n_57),
.B2(n_58),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g56 ( 
.A1(n_40),
.A2(n_32),
.B1(n_30),
.B2(n_15),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g57 ( 
.A1(n_35),
.A2(n_29),
.B1(n_28),
.B2(n_26),
.Y(n_57)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_38),
.A2(n_33),
.B1(n_22),
.B2(n_15),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_46),
.B(n_26),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g94 ( 
.A(n_61),
.B(n_67),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_40),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_62),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g64 ( 
.A(n_41),
.B(n_23),
.Y(n_64)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_64),
.Y(n_85)
);

BUFx12f_ASAP7_75t_L g66 ( 
.A(n_41),
.Y(n_66)
);

INVxp67_ASAP7_75t_L g96 ( 
.A(n_66),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_46),
.B(n_33),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_36),
.A2(n_25),
.B1(n_22),
.B2(n_27),
.Y(n_71)
);

O2A1O1Ixp33_ASAP7_75t_L g89 ( 
.A1(n_71),
.A2(n_74),
.B(n_32),
.C(n_30),
.Y(n_89)
);

AOI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_38),
.A2(n_27),
.B1(n_25),
.B2(n_19),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_SL g103 ( 
.A1(n_72),
.A2(n_79),
.B1(n_21),
.B2(n_31),
.Y(n_103)
);

BUFx16f_ASAP7_75t_L g73 ( 
.A(n_43),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_73),
.B(n_75),
.Y(n_109)
);

O2A1O1Ixp33_ASAP7_75t_SL g74 ( 
.A1(n_39),
.A2(n_45),
.B(n_43),
.C(n_32),
.Y(n_74)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_39),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_45),
.B(n_24),
.Y(n_77)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_77),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g78 ( 
.A(n_46),
.Y(n_78)
);

BUFx2_ASAP7_75t_L g99 ( 
.A(n_78),
.Y(n_99)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_35),
.A2(n_19),
.B1(n_24),
.B2(n_21),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g80 ( 
.A(n_47),
.B(n_24),
.Y(n_80)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_80),
.Y(n_102)
);

INVx3_ASAP7_75t_L g81 ( 
.A(n_73),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g133 ( 
.A(n_81),
.B(n_83),
.Y(n_133)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_65),
.Y(n_83)
);

INVx2_ASAP7_75t_L g84 ( 
.A(n_65),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g111 ( 
.A(n_84),
.B(n_92),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g86 ( 
.A(n_57),
.B(n_58),
.Y(n_86)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_86),
.B(n_105),
.Y(n_132)
);

AOI22xp33_ASAP7_75t_L g115 ( 
.A1(n_89),
.A2(n_59),
.B1(n_48),
.B2(n_78),
.Y(n_115)
);

AOI21xp33_ASAP7_75t_L g90 ( 
.A1(n_63),
.A2(n_24),
.B(n_21),
.Y(n_90)
);

OAI22xp5_ASAP7_75t_SL g119 ( 
.A1(n_90),
.A2(n_104),
.B1(n_52),
.B2(n_75),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_L g91 ( 
.A1(n_58),
.A2(n_24),
.B1(n_21),
.B2(n_31),
.Y(n_91)
);

OAI22xp5_ASAP7_75t_L g120 ( 
.A1(n_91),
.A2(n_59),
.B1(n_76),
.B2(n_68),
.Y(n_120)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_60),
.Y(n_92)
);

INVx1_ASAP7_75t_L g95 ( 
.A(n_56),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g112 ( 
.A(n_95),
.B(n_97),
.Y(n_112)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_55),
.Y(n_97)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_98),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g118 ( 
.A(n_103),
.B(n_76),
.Y(n_118)
);

OAI22xp5_ASAP7_75t_SL g104 ( 
.A1(n_72),
.A2(n_21),
.B1(n_31),
.B2(n_2),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_49),
.B(n_31),
.Y(n_105)
);

AOI21xp5_ASAP7_75t_SL g106 ( 
.A1(n_74),
.A2(n_0),
.B(n_1),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_SL g124 ( 
.A(n_106),
.B(n_0),
.Y(n_124)
);

INVxp67_ASAP7_75t_L g107 ( 
.A(n_79),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_107),
.B(n_108),
.Y(n_117)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_66),
.Y(n_108)
);

OR2x2_ASAP7_75t_L g110 ( 
.A(n_101),
.B(n_66),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_110),
.B(n_134),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g113 ( 
.A(n_109),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g143 ( 
.A(n_113),
.B(n_127),
.Y(n_143)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_82),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g141 ( 
.A(n_114),
.B(n_116),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_115),
.A2(n_122),
.B1(n_83),
.B2(n_84),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g116 ( 
.A(n_99),
.Y(n_116)
);

AOI22xp33_ASAP7_75t_L g145 ( 
.A1(n_118),
.A2(n_123),
.B1(n_104),
.B2(n_98),
.Y(n_145)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_119),
.A2(n_120),
.B1(n_121),
.B2(n_128),
.Y(n_160)
);

OAI22xp5_ASAP7_75t_SL g121 ( 
.A1(n_86),
.A2(n_68),
.B1(n_49),
.B2(n_70),
.Y(n_121)
);

AO22x2_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_49),
.B1(n_70),
.B2(n_69),
.Y(n_122)
);

OAI22x1_ASAP7_75t_L g123 ( 
.A1(n_107),
.A2(n_69),
.B1(n_1),
.B2(n_2),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_SL g146 ( 
.A(n_124),
.B(n_125),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g125 ( 
.A(n_94),
.B(n_1),
.Y(n_125)
);

INVx2_ASAP7_75t_L g127 ( 
.A(n_93),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_95),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_128)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_99),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g153 ( 
.A(n_129),
.B(n_135),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_102),
.B(n_5),
.Y(n_130)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_130),
.B(n_131),
.Y(n_148)
);

NOR2xp33_ASAP7_75t_L g131 ( 
.A(n_92),
.B(n_5),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g134 ( 
.A(n_87),
.B(n_6),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_105),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_85),
.B(n_8),
.Y(n_136)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_136),
.Y(n_138)
);

AOI22xp33_ASAP7_75t_SL g137 ( 
.A1(n_88),
.A2(n_8),
.B1(n_9),
.B2(n_10),
.Y(n_137)
);

AOI21xp5_ASAP7_75t_L g151 ( 
.A1(n_137),
.A2(n_106),
.B(n_124),
.Y(n_151)
);

INVx1_ASAP7_75t_L g140 ( 
.A(n_111),
.Y(n_140)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_140),
.B(n_142),
.Y(n_171)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_111),
.Y(n_142)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_133),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g164 ( 
.A(n_144),
.Y(n_164)
);

INVxp67_ASAP7_75t_L g169 ( 
.A(n_145),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_L g147 ( 
.A(n_132),
.B(n_87),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_L g166 ( 
.A(n_147),
.B(n_150),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_149),
.B(n_122),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g150 ( 
.A(n_132),
.B(n_100),
.Y(n_150)
);

OAI21xp5_ASAP7_75t_SL g176 ( 
.A1(n_151),
.A2(n_161),
.B(n_125),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g152 ( 
.A(n_135),
.B(n_103),
.C(n_96),
.Y(n_152)
);

MAJIxp5_ASAP7_75t_L g163 ( 
.A(n_152),
.B(n_159),
.C(n_123),
.Y(n_163)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_112),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_SL g165 ( 
.A(n_154),
.B(n_131),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g155 ( 
.A1(n_134),
.A2(n_89),
.B1(n_93),
.B2(n_96),
.Y(n_155)
);

OAI22xp5_ASAP7_75t_SL g173 ( 
.A1(n_155),
.A2(n_122),
.B1(n_118),
.B2(n_120),
.Y(n_173)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_116),
.Y(n_156)
);

CKINVDCx20_ASAP7_75t_R g177 ( 
.A(n_156),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g157 ( 
.A(n_114),
.B(n_81),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g170 ( 
.A(n_157),
.B(n_110),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_11),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_158),
.B(n_128),
.Y(n_175)
);

MAJIxp5_ASAP7_75t_L g159 ( 
.A(n_117),
.B(n_108),
.C(n_12),
.Y(n_159)
);

NOR4xp25_ASAP7_75t_L g161 ( 
.A(n_117),
.B(n_11),
.C(n_12),
.D(n_13),
.Y(n_161)
);

AND2x6_ASAP7_75t_L g162 ( 
.A(n_122),
.B(n_13),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g167 ( 
.A(n_162),
.B(n_123),
.Y(n_167)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_163),
.B(n_158),
.C(n_159),
.Y(n_185)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_165),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g187 ( 
.A(n_167),
.B(n_175),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g168 ( 
.A(n_147),
.B(n_121),
.Y(n_168)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_168),
.B(n_160),
.Y(n_182)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_170),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g172 ( 
.A1(n_154),
.A2(n_112),
.B(n_122),
.Y(n_172)
);

OAI21xp5_ASAP7_75t_SL g183 ( 
.A1(n_172),
.A2(n_173),
.B(n_176),
.Y(n_183)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_174),
.A2(n_180),
.B1(n_160),
.B2(n_140),
.Y(n_186)
);

OR2x2_ASAP7_75t_L g178 ( 
.A(n_153),
.B(n_110),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g190 ( 
.A(n_178),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_139),
.B(n_118),
.Y(n_179)
);

XNOR2xp5_ASAP7_75t_L g188 ( 
.A(n_179),
.B(n_181),
.Y(n_188)
);

OR2x2_ASAP7_75t_L g180 ( 
.A(n_153),
.B(n_130),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_139),
.B(n_126),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g198 ( 
.A(n_182),
.B(n_184),
.Y(n_198)
);

MAJx2_ASAP7_75t_L g184 ( 
.A(n_166),
.B(n_152),
.C(n_150),
.Y(n_184)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_185),
.B(n_192),
.C(n_163),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_SL g206 ( 
.A(n_186),
.B(n_197),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g191 ( 
.A(n_166),
.B(n_155),
.Y(n_191)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_191),
.B(n_173),
.Y(n_204)
);

XNOR2xp5_ASAP7_75t_SL g192 ( 
.A(n_168),
.B(n_141),
.Y(n_192)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_179),
.B(n_142),
.C(n_144),
.Y(n_193)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_193),
.B(n_170),
.C(n_178),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g195 ( 
.A1(n_169),
.A2(n_172),
.B1(n_162),
.B2(n_164),
.Y(n_195)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_195),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_L g196 ( 
.A1(n_164),
.A2(n_151),
.B1(n_149),
.B2(n_143),
.Y(n_196)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_196),
.Y(n_207)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_171),
.Y(n_197)
);

NOR4xp25_ASAP7_75t_L g199 ( 
.A(n_197),
.B(n_177),
.C(n_171),
.D(n_181),
.Y(n_199)
);

OAI21xp5_ASAP7_75t_L g219 ( 
.A1(n_199),
.A2(n_205),
.B(n_143),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_194),
.B(n_177),
.Y(n_200)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_200),
.Y(n_212)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_187),
.Y(n_201)
);

NAND2xp5_ASAP7_75t_SL g211 ( 
.A(n_201),
.B(n_210),
.Y(n_211)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_183),
.C(n_157),
.Y(n_218)
);

XOR2xp5_ASAP7_75t_L g215 ( 
.A(n_204),
.B(n_208),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_189),
.B(n_165),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g208 ( 
.A(n_192),
.B(n_176),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g216 ( 
.A(n_209),
.B(n_193),
.C(n_187),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_191),
.B(n_156),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_L g213 ( 
.A(n_198),
.B(n_182),
.Y(n_213)
);

MAJx2_ASAP7_75t_L g221 ( 
.A(n_213),
.B(n_218),
.C(n_204),
.Y(n_221)
);

AOI21xp5_ASAP7_75t_SL g214 ( 
.A1(n_207),
.A2(n_183),
.B(n_190),
.Y(n_214)
);

AOI21xp5_ASAP7_75t_L g223 ( 
.A1(n_214),
.A2(n_212),
.B(n_211),
.Y(n_223)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_216),
.A2(n_217),
.B(n_188),
.Y(n_227)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_198),
.B(n_185),
.C(n_184),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_219),
.B(n_148),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g220 ( 
.A1(n_206),
.A2(n_175),
.B1(n_167),
.B2(n_178),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_220),
.A2(n_202),
.B1(n_201),
.B2(n_209),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_227),
.C(n_215),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_222),
.B(n_224),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_223),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_SL g225 ( 
.A1(n_214),
.A2(n_161),
.B(n_208),
.Y(n_225)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_225),
.A2(n_224),
.B1(n_217),
.B2(n_138),
.Y(n_228)
);

OR2x2_ASAP7_75t_L g226 ( 
.A(n_216),
.B(n_136),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_226),
.B(n_148),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g234 ( 
.A(n_228),
.B(n_232),
.Y(n_234)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_231),
.B(n_146),
.C(n_126),
.Y(n_236)
);

OAI321xp33_ASAP7_75t_L g233 ( 
.A1(n_229),
.A2(n_180),
.A3(n_188),
.B1(n_146),
.B2(n_138),
.C(n_215),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_233),
.B(n_180),
.Y(n_237)
);

HB1xp67_ASAP7_75t_L g235 ( 
.A(n_230),
.Y(n_235)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_235),
.Y(n_238)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_236),
.B(n_231),
.C(n_234),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_237),
.A2(n_127),
.B(n_129),
.Y(n_241)
);

AOI21xp5_ASAP7_75t_L g240 ( 
.A1(n_239),
.A2(n_238),
.B(n_228),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_240),
.B(n_241),
.Y(n_242)
);


endmodule