module real_jpeg_13643_n_18 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_325, n_11, n_14, n_7, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_18);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_325;
input n_11;
input n_14;
input n_7;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_18;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_203;
wire n_198;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_78;
wire n_83;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_195;
wire n_110;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_176;
wire n_286;
wire n_215;
wire n_312;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_204;
wire n_158;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_273;
wire n_253;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_299;
wire n_243;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx12f_ASAP7_75t_L g100 ( 
.A(n_0),
.Y(n_100)
);

BUFx16f_ASAP7_75t_L g47 ( 
.A(n_1),
.Y(n_47)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_2),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_3),
.A2(n_59),
.B1(n_60),
.B2(n_145),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g145 ( 
.A(n_3),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g196 ( 
.A1(n_3),
.A2(n_34),
.B1(n_36),
.B2(n_145),
.Y(n_196)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_3),
.A2(n_29),
.B1(n_30),
.B2(n_145),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_3),
.A2(n_44),
.B1(n_48),
.B2(n_145),
.Y(n_247)
);

AOI22xp33_ASAP7_75t_L g37 ( 
.A1(n_4),
.A2(n_29),
.B1(n_30),
.B2(n_38),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_4),
.Y(n_38)
);

OAI22xp5_ASAP7_75t_L g81 ( 
.A1(n_4),
.A2(n_38),
.B1(n_59),
.B2(n_60),
.Y(n_81)
);

OAI22xp5_ASAP7_75t_L g105 ( 
.A1(n_4),
.A2(n_34),
.B1(n_36),
.B2(n_38),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_L g136 ( 
.A1(n_4),
.A2(n_38),
.B1(n_44),
.B2(n_48),
.Y(n_136)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_5),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g67 ( 
.A1(n_6),
.A2(n_59),
.B1(n_60),
.B2(n_68),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g68 ( 
.A(n_6),
.Y(n_68)
);

AOI22xp33_ASAP7_75t_SL g142 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_68),
.Y(n_142)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_6),
.A2(n_34),
.B1(n_36),
.B2(n_68),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_L g192 ( 
.A1(n_6),
.A2(n_44),
.B1(n_48),
.B2(n_68),
.Y(n_192)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_7),
.Y(n_30)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_8),
.A2(n_59),
.B1(n_60),
.B2(n_63),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_8),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g113 ( 
.A1(n_8),
.A2(n_29),
.B1(n_30),
.B2(n_63),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g140 ( 
.A1(n_8),
.A2(n_34),
.B1(n_36),
.B2(n_63),
.Y(n_140)
);

OAI22xp5_ASAP7_75t_L g193 ( 
.A1(n_8),
.A2(n_44),
.B1(n_48),
.B2(n_63),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g185 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_186),
.Y(n_185)
);

CKINVDCx20_ASAP7_75t_R g186 ( 
.A(n_9),
.Y(n_186)
);

AOI22xp33_ASAP7_75t_L g214 ( 
.A1(n_9),
.A2(n_59),
.B1(n_60),
.B2(n_186),
.Y(n_214)
);

OAI22xp5_ASAP7_75t_L g238 ( 
.A1(n_9),
.A2(n_34),
.B1(n_36),
.B2(n_186),
.Y(n_238)
);

OAI22xp33_ASAP7_75t_SL g259 ( 
.A1(n_9),
.A2(n_44),
.B1(n_48),
.B2(n_186),
.Y(n_259)
);

BUFx12_ASAP7_75t_L g31 ( 
.A(n_10),
.Y(n_31)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_11),
.B(n_82),
.Y(n_190)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_11),
.Y(n_203)
);

AOI21xp33_ASAP7_75t_L g211 ( 
.A1(n_11),
.A2(n_59),
.B(n_212),
.Y(n_211)
);

OAI22xp33_ASAP7_75t_L g237 ( 
.A1(n_11),
.A2(n_34),
.B1(n_36),
.B2(n_203),
.Y(n_237)
);

O2A1O1Ixp33_ASAP7_75t_L g239 ( 
.A1(n_11),
.A2(n_36),
.B(n_47),
.C(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_11),
.B(n_73),
.Y(n_243)
);

NAND2xp5_ASAP7_75t_L g261 ( 
.A(n_11),
.B(n_100),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_11),
.B(n_42),
.Y(n_264)
);

A2O1A1Ixp33_ASAP7_75t_L g273 ( 
.A1(n_11),
.A2(n_27),
.B(n_29),
.C(n_274),
.Y(n_273)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_12),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_SL g39 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_40),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g40 ( 
.A(n_13),
.Y(n_40)
);

OAI22xp5_ASAP7_75t_SL g51 ( 
.A1(n_13),
.A2(n_34),
.B1(n_36),
.B2(n_40),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g101 ( 
.A1(n_13),
.A2(n_40),
.B1(n_44),
.B2(n_48),
.Y(n_101)
);

AOI22xp33_ASAP7_75t_SL g64 ( 
.A1(n_14),
.A2(n_59),
.B1(n_60),
.B2(n_65),
.Y(n_64)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_14),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_65),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g104 ( 
.A1(n_14),
.A2(n_34),
.B1(n_36),
.B2(n_65),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g164 ( 
.A1(n_14),
.A2(n_44),
.B1(n_48),
.B2(n_65),
.Y(n_164)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_15),
.A2(n_59),
.B1(n_60),
.B2(n_108),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g108 ( 
.A(n_15),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_108),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_L g197 ( 
.A1(n_15),
.A2(n_34),
.B1(n_36),
.B2(n_108),
.Y(n_197)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_15),
.A2(n_44),
.B1(n_48),
.B2(n_108),
.Y(n_206)
);

AOI22xp33_ASAP7_75t_SL g172 ( 
.A1(n_16),
.A2(n_59),
.B1(n_60),
.B2(n_173),
.Y(n_172)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_16),
.Y(n_173)
);

AOI22xp33_ASAP7_75t_SL g188 ( 
.A1(n_16),
.A2(n_29),
.B1(n_30),
.B2(n_173),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_L g245 ( 
.A1(n_16),
.A2(n_34),
.B1(n_36),
.B2(n_173),
.Y(n_245)
);

OAI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_16),
.A2(n_44),
.B1(n_48),
.B2(n_173),
.Y(n_252)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_88),
.Y(n_18)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_86),
.Y(n_19)
);

NAND2xp5_ASAP7_75t_SL g20 ( 
.A(n_21),
.B(n_74),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_74),
.Y(n_87)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_66),
.C(n_69),
.Y(n_21)
);

AOI22xp5_ASAP7_75t_SL g149 ( 
.A1(n_22),
.A2(n_66),
.B1(n_116),
.B2(n_150),
.Y(n_149)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_22),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_53),
.Y(n_22)
);

AOI22xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_25),
.B1(n_41),
.B2(n_52),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g85 ( 
.A(n_25),
.B(n_41),
.C(n_53),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g25 ( 
.A1(n_26),
.A2(n_33),
.B1(n_37),
.B2(n_39),
.Y(n_25)
);

OAI22xp5_ASAP7_75t_SL g141 ( 
.A1(n_26),
.A2(n_33),
.B1(n_113),
.B2(n_142),
.Y(n_141)
);

OAI22xp5_ASAP7_75t_SL g169 ( 
.A1(n_26),
.A2(n_33),
.B1(n_142),
.B2(n_170),
.Y(n_169)
);

OAI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_26),
.A2(n_33),
.B1(n_188),
.B2(n_217),
.Y(n_216)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

AOI22xp5_ASAP7_75t_L g70 ( 
.A1(n_27),
.A2(n_71),
.B1(n_72),
.B2(n_73),
.Y(n_70)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_27),
.A2(n_73),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g111 ( 
.A1(n_27),
.A2(n_71),
.B1(n_73),
.B2(n_112),
.Y(n_111)
);

AOI22xp5_ASAP7_75t_L g183 ( 
.A1(n_27),
.A2(n_73),
.B1(n_184),
.B2(n_187),
.Y(n_183)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_27),
.A2(n_73),
.B1(n_296),
.B2(n_297),
.Y(n_295)
);

AND2x2_ASAP7_75t_L g27 ( 
.A(n_28),
.B(n_33),
.Y(n_27)
);

OAI22xp5_ASAP7_75t_SL g28 ( 
.A1(n_29),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g55 ( 
.A1(n_29),
.A2(n_30),
.B1(n_56),
.B2(n_57),
.Y(n_55)
);

OAI32xp33_ASAP7_75t_L g201 ( 
.A1(n_29),
.A2(n_31),
.A3(n_34),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_29),
.B(n_56),
.Y(n_227)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g202 ( 
.A(n_30),
.B(n_203),
.Y(n_202)
);

OAI32xp33_ASAP7_75t_L g226 ( 
.A1(n_30),
.A2(n_57),
.A3(n_59),
.B1(n_213),
.B2(n_227),
.Y(n_226)
);

INVx8_ASAP7_75t_L g32 ( 
.A(n_31),
.Y(n_32)
);

OA22x2_ASAP7_75t_L g33 ( 
.A1(n_31),
.A2(n_32),
.B1(n_34),
.B2(n_36),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_32),
.B(n_36),
.Y(n_204)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_33),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_L g272 ( 
.A1(n_33),
.A2(n_185),
.B(n_273),
.Y(n_272)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_34),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_34),
.A2(n_36),
.B1(n_46),
.B2(n_47),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

CKINVDCx14_ASAP7_75t_R g72 ( 
.A(n_37),
.Y(n_72)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_39),
.Y(n_77)
);

CKINVDCx16_ASAP7_75t_R g52 ( 
.A(n_41),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_41),
.B(n_66),
.C(n_70),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_41),
.A2(n_52),
.B1(n_70),
.B2(n_119),
.Y(n_118)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_49),
.B(n_51),
.Y(n_41)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_42),
.A2(n_49),
.B1(n_104),
.B2(n_105),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g114 ( 
.A1(n_42),
.A2(n_49),
.B1(n_51),
.B2(n_105),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_42),
.A2(n_49),
.B1(n_104),
.B2(n_139),
.Y(n_138)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_42),
.A2(n_49),
.B1(n_195),
.B2(n_197),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g218 ( 
.A1(n_42),
.A2(n_49),
.B1(n_167),
.B2(n_197),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_42),
.A2(n_49),
.B1(n_237),
.B2(n_238),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_42),
.A2(n_49),
.B1(n_238),
.B2(n_245),
.Y(n_244)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_43),
.B(n_50),
.Y(n_49)
);

OAI22xp5_ASAP7_75t_L g165 ( 
.A1(n_43),
.A2(n_140),
.B1(n_166),
.B2(n_168),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_SL g275 ( 
.A1(n_43),
.A2(n_168),
.B1(n_196),
.B2(n_276),
.Y(n_275)
);

OA22x2_ASAP7_75t_L g43 ( 
.A1(n_44),
.A2(n_46),
.B1(n_47),
.B2(n_48),
.Y(n_43)
);

INVx3_ASAP7_75t_SL g48 ( 
.A(n_44),
.Y(n_48)
);

AND2x2_ASAP7_75t_L g98 ( 
.A(n_44),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_44),
.B(n_261),
.Y(n_260)
);

INVx8_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

OAI21xp33_ASAP7_75t_L g240 ( 
.A1(n_46),
.A2(n_48),
.B(n_203),
.Y(n_240)
);

INVx6_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_49),
.Y(n_168)
);

OAI22xp5_ASAP7_75t_SL g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_64),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g66 ( 
.A1(n_54),
.A2(n_55),
.B1(n_62),
.B2(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g80 ( 
.A(n_54),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g106 ( 
.A1(n_54),
.A2(n_55),
.B1(n_67),
.B2(n_107),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g143 ( 
.A1(n_54),
.A2(n_55),
.B1(n_107),
.B2(n_144),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_54),
.A2(n_55),
.B1(n_144),
.B2(n_172),
.Y(n_171)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_54),
.A2(n_55),
.B1(n_211),
.B2(n_214),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g54 ( 
.A(n_55),
.B(n_58),
.Y(n_54)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_55),
.Y(n_82)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_56),
.A2(n_57),
.B1(n_59),
.B2(n_60),
.Y(n_58)
);

INVx11_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_SL g213 ( 
.A(n_60),
.B(n_203),
.Y(n_213)
);

BUFx16f_ASAP7_75t_L g60 ( 
.A(n_61),
.Y(n_60)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_64),
.Y(n_79)
);

AOI22xp5_ASAP7_75t_L g115 ( 
.A1(n_66),
.A2(n_116),
.B1(n_117),
.B2(n_118),
.Y(n_115)
);

CKINVDCx14_ASAP7_75t_R g116 ( 
.A(n_66),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g148 ( 
.A(n_69),
.B(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_70),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_75),
.B(n_85),
.Y(n_74)
);

AOI22xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_78),
.B1(n_83),
.B2(n_84),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g83 ( 
.A(n_76),
.Y(n_83)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_79),
.A2(n_80),
.B1(n_81),
.B2(n_82),
.Y(n_78)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_80),
.A2(n_82),
.B1(n_299),
.B2(n_300),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

AO21x1_ASAP7_75t_L g89 ( 
.A1(n_90),
.A2(n_151),
.B(n_321),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_146),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_122),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_92),
.B(n_122),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g92 ( 
.A(n_93),
.B(n_109),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_L g147 ( 
.A(n_93),
.B(n_115),
.C(n_120),
.Y(n_147)
);

OAI21xp5_ASAP7_75t_L g93 ( 
.A1(n_94),
.A2(n_97),
.B(n_106),
.Y(n_93)
);

OAI22xp5_ASAP7_75t_L g124 ( 
.A1(n_94),
.A2(n_95),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_95),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_102),
.Y(n_95)
);

AOI22xp5_ASAP7_75t_L g126 ( 
.A1(n_96),
.A2(n_97),
.B1(n_106),
.B2(n_127),
.Y(n_126)
);

AOI22xp5_ASAP7_75t_L g157 ( 
.A1(n_96),
.A2(n_97),
.B1(n_102),
.B2(n_103),
.Y(n_157)
);

CKINVDCx16_ASAP7_75t_R g96 ( 
.A(n_97),
.Y(n_96)
);

OAI21xp5_ASAP7_75t_SL g97 ( 
.A1(n_98),
.A2(n_100),
.B(n_101),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g134 ( 
.A1(n_98),
.A2(n_100),
.B1(n_101),
.B2(n_135),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_98),
.Y(n_162)
);

AOI22xp5_ASAP7_75t_L g191 ( 
.A1(n_98),
.A2(n_100),
.B1(n_192),
.B2(n_193),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g205 ( 
.A1(n_98),
.A2(n_100),
.B1(n_192),
.B2(n_206),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_98),
.A2(n_100),
.B1(n_164),
.B2(n_193),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g246 ( 
.A1(n_98),
.A2(n_100),
.B1(n_206),
.B2(n_247),
.Y(n_246)
);

AOI22xp5_ASAP7_75t_SL g258 ( 
.A1(n_98),
.A2(n_100),
.B1(n_203),
.B2(n_259),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_98),
.A2(n_100),
.B1(n_252),
.B2(n_259),
.Y(n_263)
);

OAI22xp5_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_136),
.B1(n_162),
.B2(n_163),
.Y(n_161)
);

OAI22xp5_ASAP7_75t_SL g250 ( 
.A1(n_99),
.A2(n_162),
.B1(n_251),
.B2(n_253),
.Y(n_250)
);

INVx4_ASAP7_75t_L g99 ( 
.A(n_100),
.Y(n_99)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_103),
.Y(n_102)
);

CKINVDCx14_ASAP7_75t_R g127 ( 
.A(n_106),
.Y(n_127)
);

AOI22xp5_ASAP7_75t_L g109 ( 
.A1(n_110),
.A2(n_115),
.B1(n_120),
.B2(n_121),
.Y(n_109)
);

CKINVDCx20_ASAP7_75t_R g120 ( 
.A(n_110),
.Y(n_120)
);

OAI21xp33_ASAP7_75t_L g129 ( 
.A1(n_110),
.A2(n_111),
.B(n_114),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_111),
.B(n_114),
.Y(n_110)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_115),
.Y(n_121)
);

INVx1_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_123),
.B(n_128),
.C(n_130),
.Y(n_122)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_123),
.A2(n_124),
.B1(n_128),
.B2(n_129),
.Y(n_175)
);

INVx1_ASAP7_75t_L g123 ( 
.A(n_124),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

INVx1_ASAP7_75t_L g128 ( 
.A(n_129),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g174 ( 
.A(n_130),
.B(n_175),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_141),
.C(n_143),
.Y(n_130)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_131),
.A2(n_132),
.B1(n_155),
.B2(n_156),
.Y(n_154)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_132),
.Y(n_131)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_137),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_133),
.A2(n_134),
.B1(n_137),
.B2(n_138),
.Y(n_306)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

INVxp67_ASAP7_75t_L g135 ( 
.A(n_136),
.Y(n_135)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

INVxp67_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

XOR2xp5_ASAP7_75t_L g156 ( 
.A(n_141),
.B(n_143),
.Y(n_156)
);

OAI21xp5_ASAP7_75t_L g321 ( 
.A1(n_146),
.A2(n_322),
.B(n_323),
.Y(n_321)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_148),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_147),
.B(n_148),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_L g151 ( 
.A1(n_152),
.A2(n_176),
.B(n_320),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_153),
.B(n_174),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g320 ( 
.A(n_153),
.B(n_174),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g153 ( 
.A(n_154),
.B(n_157),
.C(n_158),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g318 ( 
.A(n_154),
.B(n_157),
.Y(n_318)
);

INVx1_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_158),
.B(n_318),
.Y(n_317)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_159),
.B(n_169),
.C(n_171),
.Y(n_158)
);

AOI22xp5_ASAP7_75t_L g307 ( 
.A1(n_159),
.A2(n_160),
.B1(n_308),
.B2(n_309),
.Y(n_307)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_161),
.B(n_165),
.Y(n_160)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_161),
.B(n_165),
.Y(n_292)
);

CKINVDCx16_ASAP7_75t_R g163 ( 
.A(n_164),
.Y(n_163)
);

CKINVDCx16_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

XOR2xp5_ASAP7_75t_L g309 ( 
.A(n_169),
.B(n_171),
.Y(n_309)
);

INVxp67_ASAP7_75t_L g297 ( 
.A(n_170),
.Y(n_297)
);

INVxp67_ASAP7_75t_L g300 ( 
.A(n_172),
.Y(n_300)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_315),
.B(n_319),
.Y(n_176)
);

OAI221xp5_ASAP7_75t_L g177 ( 
.A1(n_178),
.A2(n_302),
.B1(n_313),
.B2(n_314),
.C(n_325),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_287),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_L g179 ( 
.A1(n_180),
.A2(n_230),
.B(n_286),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_207),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_181),
.B(n_207),
.Y(n_286)
);

MAJIxp5_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_194),
.C(n_198),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_182),
.B(n_283),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_SL g182 ( 
.A(n_183),
.B(n_189),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_183),
.B(n_190),
.C(n_191),
.Y(n_228)
);

INVxp67_ASAP7_75t_L g184 ( 
.A(n_185),
.Y(n_184)
);

INVxp67_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

XNOR2xp5_ASAP7_75t_L g189 ( 
.A(n_190),
.B(n_191),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_194),
.A2(n_198),
.B1(n_199),
.B2(n_284),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_194),
.Y(n_284)
);

INVxp67_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_199),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g199 ( 
.A(n_200),
.B(n_205),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_200),
.A2(n_201),
.B1(n_205),
.B2(n_278),
.Y(n_277)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_201),
.Y(n_200)
);

CKINVDCx16_ASAP7_75t_R g274 ( 
.A(n_202),
.Y(n_274)
);

INVx1_ASAP7_75t_L g278 ( 
.A(n_205),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g207 ( 
.A1(n_208),
.A2(n_209),
.B1(n_221),
.B2(n_229),
.Y(n_207)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_208),
.B(n_222),
.C(n_228),
.Y(n_288)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_210),
.B(n_215),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_210),
.B(n_216),
.C(n_220),
.Y(n_291)
);

CKINVDCx16_ASAP7_75t_R g212 ( 
.A(n_213),
.Y(n_212)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_214),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g215 ( 
.A1(n_216),
.A2(n_218),
.B1(n_219),
.B2(n_220),
.Y(n_215)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_216),
.Y(n_219)
);

INVxp67_ASAP7_75t_L g296 ( 
.A(n_217),
.Y(n_296)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_218),
.Y(n_220)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_221),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_SL g221 ( 
.A(n_222),
.B(n_228),
.Y(n_221)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_223),
.A2(n_224),
.B1(n_225),
.B2(n_226),
.Y(n_222)
);

NAND2xp5_ASAP7_75t_SL g301 ( 
.A(n_223),
.B(n_226),
.Y(n_301)
);

INVx1_ASAP7_75t_L g223 ( 
.A(n_224),
.Y(n_223)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g230 ( 
.A1(n_231),
.A2(n_280),
.B(n_285),
.Y(n_230)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_232),
.A2(n_268),
.B(n_279),
.Y(n_231)
);

AOI21xp5_ASAP7_75t_L g232 ( 
.A1(n_233),
.A2(n_248),
.B(n_267),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_241),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_234),
.B(n_241),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_235),
.B(n_239),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g254 ( 
.A1(n_235),
.A2(n_236),
.B1(n_239),
.B2(n_255),
.Y(n_254)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_239),
.Y(n_255)
);

XNOR2xp5_ASAP7_75t_L g241 ( 
.A(n_242),
.B(n_246),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_244),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_244),
.C(n_246),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g276 ( 
.A(n_245),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_247),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_256),
.B(n_266),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g249 ( 
.A(n_250),
.B(n_254),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_SL g266 ( 
.A(n_250),
.B(n_254),
.Y(n_266)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_257),
.A2(n_262),
.B(n_265),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_260),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_263),
.B(n_264),
.Y(n_262)
);

NOR2xp33_ASAP7_75t_SL g265 ( 
.A(n_263),
.B(n_264),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g268 ( 
.A(n_269),
.B(n_270),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g279 ( 
.A(n_269),
.B(n_270),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g270 ( 
.A(n_271),
.B(n_277),
.Y(n_270)
);

XNOR2xp5_ASAP7_75t_L g271 ( 
.A(n_272),
.B(n_275),
.Y(n_271)
);

MAJIxp5_ASAP7_75t_L g281 ( 
.A(n_272),
.B(n_275),
.C(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_281),
.B(n_282),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_SL g285 ( 
.A(n_281),
.B(n_282),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

OR2x2_ASAP7_75t_L g313 ( 
.A(n_288),
.B(n_289),
.Y(n_313)
);

XNOR2xp5_ASAP7_75t_L g289 ( 
.A(n_290),
.B(n_293),
.Y(n_289)
);

XNOR2xp5_ASAP7_75t_L g290 ( 
.A(n_291),
.B(n_292),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g303 ( 
.A(n_291),
.B(n_292),
.C(n_293),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g293 ( 
.A(n_294),
.B(n_301),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g294 ( 
.A(n_295),
.B(n_298),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_298),
.C(n_301),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_304),
.Y(n_302)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_303),
.B(n_304),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_305),
.B(n_312),
.Y(n_304)
);

AOI22xp5_ASAP7_75t_L g305 ( 
.A1(n_306),
.A2(n_307),
.B1(n_310),
.B2(n_311),
.Y(n_305)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_306),
.Y(n_310)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_306),
.B(n_311),
.C(n_312),
.Y(n_316)
);

INVx1_ASAP7_75t_L g311 ( 
.A(n_307),
.Y(n_311)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_316),
.B(n_317),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_316),
.B(n_317),
.Y(n_319)
);


endmodule