module fake_aes_3956_n_32 (n_11, n_1, n_2, n_6, n_4, n_3, n_9, n_5, n_7, n_10, n_8, n_0, n_32);
input n_11;
input n_1;
input n_2;
input n_6;
input n_4;
input n_3;
input n_9;
input n_5;
input n_7;
input n_10;
input n_8;
input n_0;
output n_32;
wire n_20;
wire n_23;
wire n_28;
wire n_31;
wire n_22;
wire n_25;
wire n_16;
wire n_26;
wire n_13;
wire n_30;
wire n_18;
wire n_12;
wire n_17;
wire n_14;
wire n_15;
wire n_24;
wire n_19;
wire n_21;
wire n_29;
wire n_27;
BUFx6f_ASAP7_75t_L g12 ( .A(n_10), .Y(n_12) );
BUFx6f_ASAP7_75t_L g13 ( .A(n_11), .Y(n_13) );
BUFx3_ASAP7_75t_L g14 ( .A(n_1), .Y(n_14) );
INVx2_ASAP7_75t_L g15 ( .A(n_5), .Y(n_15) );
CKINVDCx5p33_ASAP7_75t_R g16 ( .A(n_1), .Y(n_16) );
INVx1_ASAP7_75t_L g17 ( .A(n_4), .Y(n_17) );
INVx1_ASAP7_75t_L g18 ( .A(n_14), .Y(n_18) );
INVx1_ASAP7_75t_L g19 ( .A(n_17), .Y(n_19) );
BUFx6f_ASAP7_75t_L g20 ( .A(n_12), .Y(n_20) );
OAI22xp5_ASAP7_75t_L g21 ( .A1(n_19), .A2(n_16), .B1(n_17), .B2(n_15), .Y(n_21) );
NAND2xp5_ASAP7_75t_L g22 ( .A(n_18), .B(n_13), .Y(n_22) );
OAI22xp5_ASAP7_75t_L g23 ( .A1(n_21), .A2(n_13), .B1(n_12), .B2(n_20), .Y(n_23) );
INVx4_ASAP7_75t_L g24 ( .A(n_23), .Y(n_24) );
AND2x2_ASAP7_75t_L g25 ( .A(n_24), .B(n_22), .Y(n_25) );
INVx1_ASAP7_75t_L g26 ( .A(n_24), .Y(n_26) );
AOI322xp5_ASAP7_75t_L g27 ( .A1(n_26), .A2(n_0), .A3(n_2), .B1(n_13), .B2(n_12), .C1(n_20), .C2(n_6), .Y(n_27) );
INVx1_ASAP7_75t_SL g28 ( .A(n_25), .Y(n_28) );
OR3x2_ASAP7_75t_L g29 ( .A(n_27), .B(n_0), .C(n_2), .Y(n_29) );
NAND3xp33_ASAP7_75t_SL g30 ( .A(n_28), .B(n_25), .C(n_3), .Y(n_30) );
INVx1_ASAP7_75t_L g31 ( .A(n_29), .Y(n_31) );
AOI222xp33_ASAP7_75t_L g32 ( .A1(n_31), .A2(n_30), .B1(n_20), .B2(n_8), .C1(n_9), .C2(n_7), .Y(n_32) );
endmodule