module real_jpeg_3125_n_12 (n_5, n_4, n_8, n_0, n_1, n_11, n_2, n_6, n_7, n_3, n_10, n_9, n_12);

input n_5;
input n_4;
input n_8;
input n_0;
input n_1;
input n_11;
input n_2;
input n_6;
input n_7;
input n_3;
input n_10;
input n_9;

output n_12;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_252;
wire n_68;
wire n_260;
wire n_146;
wire n_247;
wire n_78;
wire n_83;
wire n_286;
wire n_288;
wire n_176;
wire n_166;
wire n_215;
wire n_221;
wire n_249;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_280;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_271;
wire n_281;
wire n_163;
wire n_276;
wire n_22;
wire n_287;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_173;
wire n_243;
wire n_255;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_275;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_13;
wire n_120;
wire n_113;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_141;
wire n_242;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_282;
wire n_147;
wire n_265;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_28;
wire n_44;
wire n_267;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_254;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_160;
wire n_172;
wire n_211;
wire n_45;
wire n_285;
wire n_112;
wire n_42;
wire n_268;
wire n_18;
wire n_145;
wire n_266;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_262;
wire n_118;
wire n_220;
wire n_17;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_31;
wire n_137;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_270;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_272;
wire n_192;
wire n_198;
wire n_100;
wire n_203;
wire n_23;
wire n_51;
wire n_14;
wire n_71;
wire n_90;
wire n_61;
wire n_258;
wire n_110;
wire n_195;
wire n_205;
wire n_117;
wire n_99;
wire n_193;
wire n_261;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_20;
wire n_150;
wire n_228;
wire n_30;
wire n_158;
wire n_204;
wire n_149;
wire n_15;
wire n_144;
wire n_130;
wire n_278;
wire n_241;
wire n_103;
wire n_225;
wire n_259;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_284;
wire n_277;
wire n_226;
wire n_125;
wire n_240;
wire n_185;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_264;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_190;
wire n_230;
wire n_60;
wire n_263;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_279;
wire n_128;
wire n_167;
wire n_213;
wire n_179;
wire n_216;
wire n_202;
wire n_133;
wire n_244;
wire n_138;
wire n_25;
wire n_257;
wire n_217;
wire n_53;
wire n_127;
wire n_206;
wire n_210;
wire n_224;
wire n_119;
wire n_36;
wire n_102;
wire n_81;
wire n_85;
wire n_181;
wire n_283;
wire n_101;
wire n_256;
wire n_274;
wire n_182;
wire n_253;
wire n_96;
wire n_273;
wire n_269;
wire n_89;
wire n_16;

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

AOI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_1),
.A2(n_32),
.B1(n_33),
.B2(n_36),
.Y(n_31)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_1),
.Y(n_36)
);

OAI22xp33_ASAP7_75t_SL g72 ( 
.A1(n_1),
.A2(n_36),
.B1(n_59),
.B2(n_61),
.Y(n_72)
);

AOI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_1),
.A2(n_22),
.B1(n_28),
.B2(n_36),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g27 ( 
.A1(n_2),
.A2(n_22),
.B1(n_28),
.B2(n_29),
.Y(n_27)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_2),
.A2(n_29),
.B1(n_54),
.B2(n_57),
.Y(n_63)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_2),
.A2(n_29),
.B1(n_32),
.B2(n_33),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g95 ( 
.A1(n_2),
.A2(n_29),
.B1(n_59),
.B2(n_61),
.Y(n_95)
);

MAJIxp5_ASAP7_75t_L g168 ( 
.A(n_2),
.B(n_56),
.C(n_59),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_2),
.B(n_58),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g209 ( 
.A(n_2),
.B(n_33),
.C(n_75),
.Y(n_209)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_2),
.B(n_22),
.C(n_41),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_L g244 ( 
.A(n_2),
.B(n_73),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g258 ( 
.A(n_2),
.B(n_26),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_2),
.B(n_69),
.Y(n_262)
);

BUFx3_ASAP7_75t_L g26 ( 
.A(n_3),
.Y(n_26)
);

BUFx12f_ASAP7_75t_L g75 ( 
.A(n_4),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_SL g101 ( 
.A1(n_5),
.A2(n_54),
.B1(n_57),
.B2(n_102),
.Y(n_101)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_5),
.Y(n_102)
);

OAI22xp33_ASAP7_75t_SL g164 ( 
.A1(n_5),
.A2(n_59),
.B1(n_61),
.B2(n_102),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g213 ( 
.A1(n_5),
.A2(n_32),
.B1(n_33),
.B2(n_102),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_5),
.A2(n_22),
.B1(n_28),
.B2(n_102),
.Y(n_240)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_6),
.Y(n_54)
);

BUFx16f_ASAP7_75t_L g42 ( 
.A(n_7),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g60 ( 
.A(n_8),
.Y(n_60)
);

OAI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_9),
.A2(n_32),
.B1(n_33),
.B2(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_9),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g80 ( 
.A1(n_9),
.A2(n_46),
.B1(n_59),
.B2(n_61),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_9),
.A2(n_22),
.B1(n_28),
.B2(n_46),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_9),
.A2(n_46),
.B1(n_54),
.B2(n_57),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_10),
.Y(n_56)
);

BUFx12f_ASAP7_75t_L g35 ( 
.A(n_11),
.Y(n_35)
);

XNOR2xp5_ASAP7_75t_L g12 ( 
.A(n_13),
.B(n_125),
.Y(n_12)
);

NAND2xp5_ASAP7_75t_L g13 ( 
.A(n_14),
.B(n_124),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_15),
.Y(n_14)
);

NOR2xp33_ASAP7_75t_L g15 ( 
.A(n_16),
.B(n_103),
.Y(n_15)
);

NAND2xp5_ASAP7_75t_L g124 ( 
.A(n_16),
.B(n_103),
.Y(n_124)
);

MAJIxp5_ASAP7_75t_L g16 ( 
.A(n_17),
.B(n_64),
.C(n_82),
.Y(n_16)
);

OAI22xp5_ASAP7_75t_SL g286 ( 
.A1(n_17),
.A2(n_18),
.B1(n_64),
.B2(n_287),
.Y(n_286)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_18),
.Y(n_17)
);

XOR2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_47),
.Y(n_18)
);

AOI21xp33_ASAP7_75t_L g104 ( 
.A1(n_19),
.A2(n_20),
.B(n_49),
.Y(n_104)
);

NAND2xp5_ASAP7_75t_L g19 ( 
.A(n_20),
.B(n_30),
.Y(n_19)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_20),
.A2(n_48),
.B1(n_49),
.B2(n_50),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_20),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_20),
.A2(n_30),
.B1(n_48),
.B2(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_20),
.B(n_207),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g227 ( 
.A1(n_20),
.A2(n_48),
.B1(n_207),
.B2(n_208),
.Y(n_227)
);

AOI21xp5_ASAP7_75t_L g20 ( 
.A1(n_21),
.A2(n_25),
.B(n_27),
.Y(n_20)
);

OR2x2_ASAP7_75t_L g87 ( 
.A(n_21),
.B(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g131 ( 
.A1(n_21),
.A2(n_132),
.B(n_133),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_21),
.B(n_27),
.Y(n_198)
);

NOR2xp33_ASAP7_75t_L g239 ( 
.A(n_21),
.B(n_240),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_25),
.Y(n_21)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_22),
.Y(n_28)
);

OAI22xp5_ASAP7_75t_L g43 ( 
.A1(n_22),
.A2(n_28),
.B1(n_40),
.B2(n_41),
.Y(n_43)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_22),
.B(n_258),
.Y(n_257)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_24),
.Y(n_23)
);

NOR2xp33_ASAP7_75t_SL g134 ( 
.A(n_25),
.B(n_88),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g169 ( 
.A1(n_25),
.A2(n_87),
.B(n_132),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_25),
.B(n_240),
.Y(n_254)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_26),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_SL g85 ( 
.A(n_26),
.B(n_86),
.Y(n_85)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_27),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_30),
.Y(n_149)
);

OAI21xp5_ASAP7_75t_L g30 ( 
.A1(n_31),
.A2(n_37),
.B(n_44),
.Y(n_30)
);

OAI21xp5_ASAP7_75t_L g89 ( 
.A1(n_31),
.A2(n_66),
.B(n_70),
.Y(n_89)
);

AOI22xp5_ASAP7_75t_L g39 ( 
.A1(n_32),
.A2(n_33),
.B1(n_40),
.B2(n_41),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g74 ( 
.A1(n_32),
.A2(n_33),
.B1(n_75),
.B2(n_76),
.Y(n_74)
);

INVx4_ASAP7_75t_L g32 ( 
.A(n_33),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_33),
.B(n_234),
.Y(n_233)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

BUFx12f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

AOI21x1_ASAP7_75t_SL g117 ( 
.A1(n_37),
.A2(n_70),
.B(n_118),
.Y(n_117)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_38),
.B(n_45),
.Y(n_66)
);

NAND2xp5_ASAP7_75t_L g136 ( 
.A(n_38),
.B(n_68),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_38),
.B(n_213),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_39),
.B(n_43),
.Y(n_38)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g41 ( 
.A(n_42),
.Y(n_41)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_43),
.B(n_45),
.Y(n_44)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_43),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_44),
.B(n_136),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g243 ( 
.A(n_44),
.B(n_212),
.Y(n_243)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_50),
.Y(n_49)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_62),
.B(n_63),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_SL g113 ( 
.A(n_51),
.B(n_63),
.Y(n_113)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_52),
.Y(n_51)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_52),
.B(n_101),
.Y(n_100)
);

NAND2xp5_ASAP7_75t_SL g141 ( 
.A(n_52),
.B(n_111),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_53),
.B(n_58),
.Y(n_52)
);

AOI22xp33_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_53)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g167 ( 
.A(n_54),
.B(n_168),
.Y(n_167)
);

OAI22xp5_ASAP7_75t_SL g58 ( 
.A1(n_55),
.A2(n_56),
.B1(n_59),
.B2(n_61),
.Y(n_58)
);

INVx8_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_58),
.Y(n_62)
);

NAND2xp5_ASAP7_75t_SL g98 ( 
.A(n_58),
.B(n_99),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_58),
.B(n_111),
.Y(n_110)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_58),
.B(n_101),
.Y(n_140)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_59),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g79 ( 
.A1(n_59),
.A2(n_61),
.B1(n_75),
.B2(n_76),
.Y(n_79)
);

NAND2xp5_ASAP7_75t_L g208 ( 
.A(n_59),
.B(n_209),
.Y(n_208)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

CKINVDCx16_ASAP7_75t_R g99 ( 
.A(n_63),
.Y(n_99)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_64),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_SL g64 ( 
.A1(n_65),
.A2(n_71),
.B(n_81),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_71),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g65 ( 
.A(n_66),
.B(n_67),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_66),
.B(n_225),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_67),
.B(n_212),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_SL g67 ( 
.A(n_68),
.B(n_69),
.Y(n_67)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_68),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_69),
.B(n_213),
.Y(n_225)
);

INVx1_ASAP7_75t_L g69 ( 
.A(n_70),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_72),
.A2(n_73),
.B(n_77),
.Y(n_71)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_72),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_73),
.A2(n_94),
.B(n_95),
.Y(n_137)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_73),
.B(n_95),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_73),
.B(n_164),
.Y(n_183)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_74),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_L g91 ( 
.A(n_74),
.B(n_80),
.Y(n_91)
);

INVx3_ASAP7_75t_SL g76 ( 
.A(n_75),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_SL g181 ( 
.A(n_77),
.B(n_182),
.Y(n_181)
);

NOR2xp33_ASAP7_75t_SL g77 ( 
.A(n_78),
.B(n_80),
.Y(n_77)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_78),
.Y(n_94)
);

OAI21xp5_ASAP7_75t_L g119 ( 
.A1(n_78),
.A2(n_120),
.B(n_121),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g162 ( 
.A(n_78),
.B(n_163),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_81),
.A2(n_106),
.B1(n_107),
.B2(n_123),
.Y(n_105)
);

CKINVDCx14_ASAP7_75t_R g123 ( 
.A(n_81),
.Y(n_123)
);

XNOR2xp5_ASAP7_75t_L g285 ( 
.A(n_82),
.B(n_286),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_83),
.B(n_90),
.C(n_96),
.Y(n_82)
);

XOR2xp5_ASAP7_75t_L g144 ( 
.A(n_83),
.B(n_145),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_84),
.B(n_89),
.Y(n_83)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_84),
.B(n_89),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_87),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g237 ( 
.A(n_85),
.B(n_238),
.Y(n_237)
);

NAND2xp5_ASAP7_75t_L g252 ( 
.A(n_87),
.B(n_253),
.Y(n_252)
);

OAI22xp5_ASAP7_75t_SL g145 ( 
.A1(n_90),
.A2(n_96),
.B1(n_97),
.B2(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g146 ( 
.A(n_90),
.Y(n_146)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_92),
.Y(n_90)
);

INVxp67_ASAP7_75t_L g121 ( 
.A(n_91),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_91),
.B(n_162),
.Y(n_193)
);

INVxp33_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_93),
.B(n_183),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_94),
.B(n_95),
.Y(n_93)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_100),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_110),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_L g103 ( 
.A(n_104),
.B(n_105),
.Y(n_103)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_108),
.A2(n_109),
.B1(n_114),
.B2(n_115),
.Y(n_107)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_112),
.Y(n_109)
);

INVxp67_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g179 ( 
.A(n_113),
.B(n_180),
.Y(n_179)
);

INVx1_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_116),
.A2(n_117),
.B1(n_119),
.B2(n_122),
.Y(n_115)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_116),
.B(n_179),
.C(n_181),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g188 ( 
.A1(n_116),
.A2(n_117),
.B1(n_181),
.B2(n_189),
.Y(n_188)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

CKINVDCx16_ASAP7_75t_R g122 ( 
.A(n_119),
.Y(n_122)
);

HB1xp67_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

A2O1A1O1Ixp25_ASAP7_75t_L g126 ( 
.A1(n_127),
.A2(n_171),
.B(n_282),
.C(n_283),
.D(n_288),
.Y(n_126)
);

NAND2xp5_ASAP7_75t_SL g127 ( 
.A(n_128),
.B(n_150),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g282 ( 
.A(n_128),
.B(n_150),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_129),
.B(n_142),
.Y(n_128)
);

MAJIxp5_ASAP7_75t_L g284 ( 
.A(n_129),
.B(n_143),
.C(n_148),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_137),
.C(n_138),
.Y(n_129)
);

XOR2xp5_ASAP7_75t_L g152 ( 
.A(n_130),
.B(n_153),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_135),
.Y(n_130)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_131),
.B(n_135),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g196 ( 
.A(n_133),
.B(n_197),
.Y(n_196)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g261 ( 
.A(n_134),
.B(n_239),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_136),
.B(n_225),
.Y(n_235)
);

OAI22xp5_ASAP7_75t_SL g153 ( 
.A1(n_137),
.A2(n_138),
.B1(n_139),
.B2(n_154),
.Y(n_153)
);

INVx1_ASAP7_75t_L g154 ( 
.A(n_137),
.Y(n_154)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_139),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_141),
.Y(n_139)
);

INVxp33_ASAP7_75t_L g180 ( 
.A(n_140),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g142 ( 
.A1(n_143),
.A2(n_144),
.B1(n_147),
.B2(n_148),
.Y(n_142)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g150 ( 
.A(n_151),
.B(n_155),
.C(n_170),
.Y(n_150)
);

OAI22xp5_ASAP7_75t_SL g276 ( 
.A1(n_151),
.A2(n_152),
.B1(n_170),
.B2(n_277),
.Y(n_276)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g275 ( 
.A(n_155),
.B(n_276),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_156),
.B(n_158),
.C(n_165),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g176 ( 
.A1(n_156),
.A2(n_157),
.B1(n_158),
.B2(n_159),
.Y(n_176)
);

CKINVDCx14_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g158 ( 
.A(n_159),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

INVxp67_ASAP7_75t_L g161 ( 
.A(n_162),
.Y(n_161)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g175 ( 
.A(n_165),
.B(n_176),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_L g165 ( 
.A(n_166),
.B(n_169),
.Y(n_165)
);

OAI22xp5_ASAP7_75t_L g190 ( 
.A1(n_166),
.A2(n_167),
.B1(n_169),
.B2(n_191),
.Y(n_190)
);

CKINVDCx20_ASAP7_75t_R g166 ( 
.A(n_167),
.Y(n_166)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_169),
.Y(n_191)
);

INVx1_ASAP7_75t_L g277 ( 
.A(n_170),
.Y(n_277)
);

OAI21xp5_ASAP7_75t_L g171 ( 
.A1(n_172),
.A2(n_273),
.B(n_279),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_173),
.B(n_199),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_174),
.B(n_185),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_174),
.B(n_185),
.Y(n_280)
);

XNOR2xp5_ASAP7_75t_L g174 ( 
.A(n_175),
.B(n_177),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g278 ( 
.A(n_175),
.B(n_178),
.C(n_184),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g177 ( 
.A(n_178),
.B(n_184),
.Y(n_177)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_179),
.B(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_181),
.Y(n_189)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

MAJIxp5_ASAP7_75t_L g185 ( 
.A(n_186),
.B(n_190),
.C(n_192),
.Y(n_185)
);

OAI22xp5_ASAP7_75t_SL g214 ( 
.A1(n_186),
.A2(n_187),
.B1(n_215),
.B2(n_216),
.Y(n_214)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g216 ( 
.A(n_190),
.B(n_192),
.Y(n_216)
);

MAJIxp5_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.C(n_195),
.Y(n_192)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_193),
.B(n_204),
.Y(n_203)
);

AOI22xp5_ASAP7_75t_L g204 ( 
.A1(n_194),
.A2(n_195),
.B1(n_196),
.B2(n_205),
.Y(n_204)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_194),
.Y(n_205)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_196),
.Y(n_195)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_198),
.B(n_254),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_217),
.B(n_272),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_214),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g272 ( 
.A(n_201),
.B(n_214),
.Y(n_272)
);

MAJIxp5_ASAP7_75t_L g201 ( 
.A(n_202),
.B(n_206),
.C(n_210),
.Y(n_201)
);

AOI22xp5_ASAP7_75t_L g219 ( 
.A1(n_202),
.A2(n_203),
.B1(n_220),
.B2(n_222),
.Y(n_219)
);

INVx1_ASAP7_75t_L g202 ( 
.A(n_203),
.Y(n_202)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_206),
.A2(n_210),
.B1(n_211),
.B2(n_221),
.Y(n_220)
);

INVx1_ASAP7_75t_L g221 ( 
.A(n_206),
.Y(n_221)
);

CKINVDCx20_ASAP7_75t_R g207 ( 
.A(n_208),
.Y(n_207)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_216),
.Y(n_215)
);

AOI21x1_ASAP7_75t_SL g217 ( 
.A1(n_218),
.A2(n_228),
.B(n_271),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_219),
.B(n_223),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_219),
.B(n_223),
.Y(n_271)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_220),
.Y(n_222)
);

MAJIxp5_ASAP7_75t_L g223 ( 
.A(n_224),
.B(n_226),
.C(n_227),
.Y(n_223)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_224),
.B(n_226),
.Y(n_269)
);

XOR2xp5_ASAP7_75t_L g268 ( 
.A(n_227),
.B(n_269),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_L g228 ( 
.A1(n_229),
.A2(n_266),
.B(n_270),
.Y(n_228)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_230),
.A2(n_248),
.B(n_265),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_236),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_231),
.B(n_236),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_L g231 ( 
.A(n_232),
.B(n_235),
.Y(n_231)
);

OAI22xp5_ASAP7_75t_L g250 ( 
.A1(n_232),
.A2(n_233),
.B1(n_235),
.B2(n_251),
.Y(n_250)
);

CKINVDCx20_ASAP7_75t_R g232 ( 
.A(n_233),
.Y(n_232)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_235),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_241),
.B1(n_242),
.B2(n_247),
.Y(n_236)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_237),
.Y(n_247)
);

INVxp67_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_242),
.Y(n_241)
);

OAI22xp5_ASAP7_75t_SL g242 ( 
.A1(n_243),
.A2(n_244),
.B1(n_245),
.B2(n_246),
.Y(n_242)
);

INVx1_ASAP7_75t_L g245 ( 
.A(n_243),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_244),
.Y(n_246)
);

MAJIxp5_ASAP7_75t_L g267 ( 
.A(n_244),
.B(n_245),
.C(n_247),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_SL g248 ( 
.A1(n_249),
.A2(n_255),
.B(n_264),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_250),
.B(n_252),
.Y(n_249)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_250),
.B(n_252),
.Y(n_264)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_256),
.A2(n_260),
.B(n_263),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_257),
.B(n_259),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_261),
.B(n_262),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g263 ( 
.A(n_261),
.B(n_262),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_267),
.B(n_268),
.Y(n_270)
);

INVxp67_ASAP7_75t_L g273 ( 
.A(n_274),
.Y(n_273)
);

AOI21xp5_ASAP7_75t_L g279 ( 
.A1(n_274),
.A2(n_280),
.B(n_281),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g274 ( 
.A(n_275),
.B(n_278),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_275),
.B(n_278),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_284),
.B(n_285),
.Y(n_283)
);

NOR2xp33_ASAP7_75t_L g288 ( 
.A(n_284),
.B(n_285),
.Y(n_288)
);


endmodule