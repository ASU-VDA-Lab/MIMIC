module fake_jpeg_2887_n_71 (n_13, n_21, n_1, n_10, n_6, n_14, n_19, n_18, n_20, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_71);

input n_13;
input n_21;
input n_1;
input n_10;
input n_6;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_71;

wire n_57;
wire n_53;
wire n_33;
wire n_54;
wire n_61;
wire n_45;
wire n_23;
wire n_69;
wire n_27;
wire n_55;
wire n_64;
wire n_47;
wire n_22;
wire n_51;
wire n_40;
wire n_59;
wire n_35;
wire n_48;
wire n_68;
wire n_52;
wire n_46;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_65;
wire n_34;
wire n_30;
wire n_39;
wire n_42;
wire n_49;
wire n_24;
wire n_28;
wire n_44;
wire n_26;
wire n_38;
wire n_36;
wire n_62;
wire n_25;
wire n_31;
wire n_56;
wire n_29;
wire n_37;
wire n_43;
wire n_50;
wire n_32;
wire n_70;
wire n_67;
wire n_66;

CKINVDCx20_ASAP7_75t_R g22 ( 
.A(n_7),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_11),
.B(n_2),
.Y(n_23)
);

INVx2_ASAP7_75t_L g24 ( 
.A(n_12),
.Y(n_24)
);

INVx6_ASAP7_75t_SL g25 ( 
.A(n_1),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_16),
.B(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

AND2x4_ASAP7_75t_SL g28 ( 
.A(n_23),
.B(n_21),
.Y(n_28)
);

AND2x2_ASAP7_75t_L g37 ( 
.A(n_28),
.B(n_26),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_24),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_29),
.Y(n_38)
);

BUFx4f_ASAP7_75t_SL g30 ( 
.A(n_25),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_30),
.B(n_32),
.Y(n_34)
);

INVx4_ASAP7_75t_L g31 ( 
.A(n_25),
.Y(n_31)
);

INVx4_ASAP7_75t_L g36 ( 
.A(n_31),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_26),
.Y(n_33)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_33),
.B(n_35),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g35 ( 
.A(n_28),
.B(n_22),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g39 ( 
.A(n_37),
.B(n_28),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_39),
.B(n_45),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_SL g40 ( 
.A1(n_33),
.A2(n_29),
.B1(n_24),
.B2(n_28),
.Y(n_40)
);

XOR2xp5_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_41),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g41 ( 
.A(n_37),
.B(n_27),
.Y(n_41)
);

OAI22xp5_ASAP7_75t_SL g42 ( 
.A1(n_37),
.A2(n_22),
.B1(n_27),
.B2(n_25),
.Y(n_42)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_42),
.Y(n_46)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_43),
.Y(n_51)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_36),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_41),
.B(n_34),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_48),
.B(n_3),
.Y(n_58)
);

OAI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_44),
.A2(n_38),
.B(n_30),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g59 ( 
.A(n_50),
.B(n_18),
.Y(n_59)
);

O2A1O1Ixp33_ASAP7_75t_L g52 ( 
.A1(n_40),
.A2(n_30),
.B(n_31),
.C(n_38),
.Y(n_52)
);

AOI22x1_ASAP7_75t_L g56 ( 
.A1(n_52),
.A2(n_0),
.B1(n_3),
.B2(n_4),
.Y(n_56)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_46),
.A2(n_42),
.B1(n_1),
.B2(n_2),
.Y(n_53)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_53),
.A2(n_56),
.B1(n_49),
.B2(n_52),
.Y(n_61)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_54),
.Y(n_60)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_50),
.Y(n_55)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_55),
.B(n_57),
.C(n_58),
.Y(n_63)
);

AND2x6_ASAP7_75t_L g57 ( 
.A(n_47),
.B(n_19),
.Y(n_57)
);

OAI21xp33_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_10),
.B(n_17),
.Y(n_62)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_61),
.Y(n_65)
);

MAJx2_ASAP7_75t_L g66 ( 
.A(n_62),
.B(n_64),
.C(n_63),
.Y(n_66)
);

AOI321xp33_ASAP7_75t_L g64 ( 
.A1(n_59),
.A2(n_49),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C(n_4),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_66),
.B(n_62),
.Y(n_67)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_67),
.Y(n_68)
);

OAI31xp33_ASAP7_75t_L g69 ( 
.A1(n_68),
.A2(n_65),
.A3(n_60),
.B(n_56),
.Y(n_69)
);

AOI322xp5_ASAP7_75t_SL g70 ( 
.A1(n_69),
.A2(n_5),
.A3(n_6),
.B1(n_8),
.B2(n_13),
.C1(n_14),
.C2(n_15),
.Y(n_70)
);

XNOR2xp5_ASAP7_75t_L g71 ( 
.A(n_70),
.B(n_8),
.Y(n_71)
);


endmodule