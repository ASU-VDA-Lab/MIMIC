module fake_jpeg_13825_n_98 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_32, n_8, n_15, n_7, n_98);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_32;
input n_8;
input n_15;
input n_7;

output n_98;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_84;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_88;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_89;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_35;
wire n_48;
wire n_87;
wire n_46;
wire n_86;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_82;
wire n_96;

INVx6_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_28),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_2),
.Y(n_35)
);

INVx8_ASAP7_75t_SL g36 ( 
.A(n_5),
.Y(n_36)
);

INVx1_ASAP7_75t_L g37 ( 
.A(n_9),
.Y(n_37)
);

INVx1_ASAP7_75t_SL g38 ( 
.A(n_24),
.Y(n_38)
);

BUFx5_ASAP7_75t_L g39 ( 
.A(n_31),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_23),
.Y(n_40)
);

BUFx2_ASAP7_75t_L g41 ( 
.A(n_6),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_12),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_17),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g44 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_44)
);

OR2x2_ASAP7_75t_L g58 ( 
.A(n_44),
.B(n_45),
.Y(n_58)
);

AOI22xp33_ASAP7_75t_SL g45 ( 
.A1(n_41),
.A2(n_0),
.B1(n_1),
.B2(n_3),
.Y(n_45)
);

AOI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_37),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_46),
.B(n_49),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_35),
.B(n_4),
.Y(n_47)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_47),
.B(n_48),
.Y(n_52)
);

OAI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_21),
.B1(n_32),
.B2(n_30),
.Y(n_48)
);

AOI21xp33_ASAP7_75t_L g49 ( 
.A1(n_35),
.A2(n_7),
.B(n_8),
.Y(n_49)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_38),
.B(n_7),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_50),
.B(n_51),
.Y(n_53)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_40),
.B(n_8),
.Y(n_51)
);

BUFx12f_ASAP7_75t_L g54 ( 
.A(n_51),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g65 ( 
.A(n_54),
.Y(n_65)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_46),
.Y(n_55)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_55),
.Y(n_64)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_47),
.Y(n_56)
);

INVx1_ASAP7_75t_L g66 ( 
.A(n_56),
.Y(n_66)
);

BUFx2_ASAP7_75t_L g57 ( 
.A(n_47),
.Y(n_57)
);

INVx1_ASAP7_75t_L g73 ( 
.A(n_57),
.Y(n_73)
);

INVx4_ASAP7_75t_L g59 ( 
.A(n_51),
.Y(n_59)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_59),
.B(n_61),
.Y(n_74)
);

INVx4_ASAP7_75t_L g61 ( 
.A(n_51),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_SL g62 ( 
.A1(n_58),
.A2(n_40),
.B1(n_36),
.B2(n_33),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g80 ( 
.A1(n_62),
.A2(n_25),
.B(n_26),
.Y(n_80)
);

AOI22xp5_ASAP7_75t_L g63 ( 
.A1(n_57),
.A2(n_37),
.B1(n_33),
.B2(n_42),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_SL g81 ( 
.A(n_63),
.B(n_67),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g67 ( 
.A1(n_59),
.A2(n_42),
.B1(n_43),
.B2(n_34),
.Y(n_67)
);

XNOR2xp5_ASAP7_75t_L g68 ( 
.A(n_53),
.B(n_40),
.Y(n_68)
);

MAJIxp5_ASAP7_75t_L g84 ( 
.A(n_68),
.B(n_69),
.C(n_29),
.Y(n_84)
);

OAI21xp5_ASAP7_75t_SL g69 ( 
.A1(n_58),
.A2(n_39),
.B(n_9),
.Y(n_69)
);

A2O1A1Ixp33_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_10),
.B(n_11),
.C(n_13),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_70),
.B(n_71),
.Y(n_85)
);

AOI22xp5_ASAP7_75t_L g71 ( 
.A1(n_55),
.A2(n_60),
.B1(n_52),
.B2(n_54),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_55),
.A2(n_54),
.B1(n_16),
.B2(n_18),
.Y(n_72)
);

NOR2xp33_ASAP7_75t_L g75 ( 
.A(n_72),
.B(n_15),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_75),
.A2(n_80),
.B1(n_82),
.B2(n_84),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_66),
.B(n_19),
.Y(n_76)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_76),
.Y(n_88)
);

MAJx2_ASAP7_75t_L g77 ( 
.A(n_74),
.B(n_20),
.C(n_22),
.Y(n_77)
);

MAJIxp5_ASAP7_75t_L g89 ( 
.A(n_77),
.B(n_79),
.C(n_83),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_73),
.B(n_74),
.Y(n_78)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_78),
.Y(n_87)
);

INVx1_ASAP7_75t_L g79 ( 
.A(n_62),
.Y(n_79)
);

OR2x4_ASAP7_75t_L g82 ( 
.A(n_65),
.B(n_27),
.Y(n_82)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_64),
.Y(n_83)
);

FAx1_ASAP7_75t_SL g90 ( 
.A(n_89),
.B(n_85),
.CI(n_65),
.CON(n_90),
.SN(n_90)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_90),
.B(n_91),
.C(n_92),
.Y(n_93)
);

NAND2xp5_ASAP7_75t_L g91 ( 
.A(n_87),
.B(n_76),
.Y(n_91)
);

NAND2xp5_ASAP7_75t_L g92 ( 
.A(n_87),
.B(n_70),
.Y(n_92)
);

OAI21xp5_ASAP7_75t_SL g94 ( 
.A1(n_93),
.A2(n_89),
.B(n_90),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g95 ( 
.A(n_94),
.B(n_90),
.Y(n_95)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_95),
.Y(n_96)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_96),
.A2(n_88),
.B(n_81),
.Y(n_97)
);

XOR2xp5_ASAP7_75t_L g98 ( 
.A(n_97),
.B(n_86),
.Y(n_98)
);


endmodule