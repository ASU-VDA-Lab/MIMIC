module fake_jpeg_17018_n_303 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_303);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_303;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_152;
wire n_19;
wire n_182;
wire n_84;
wire n_59;
wire n_98;
wire n_251;
wire n_252;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_278;
wire n_205;
wire n_295;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_293;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_137;
wire n_74;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_291;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_175;
wire n_187;
wire n_21;
wire n_57;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_301;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_296;
wire n_168;
wire n_298;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_44;
wire n_24;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_102;
wire n_130;
wire n_99;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_240;
wire n_212;
wire n_294;
wire n_299;
wire n_211;
wire n_300;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_302;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_297;
wire n_226;
wire n_210;
wire n_48;
wire n_35;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_256;
wire n_151;
wire n_221;
wire n_97;
wire n_169;
wire n_290;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_292;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

INVx2_ASAP7_75t_L g17 ( 
.A(n_4),
.Y(n_17)
);

BUFx24_ASAP7_75t_L g18 ( 
.A(n_4),
.Y(n_18)
);

INVx3_ASAP7_75t_L g19 ( 
.A(n_4),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_9),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_9),
.Y(n_23)
);

INVx6_ASAP7_75t_L g24 ( 
.A(n_8),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_7),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_4),
.Y(n_26)
);

BUFx12_ASAP7_75t_L g27 ( 
.A(n_14),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g28 ( 
.A(n_1),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_2),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_13),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_1),
.Y(n_31)
);

BUFx10_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_2),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_9),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_0),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_SL g36 ( 
.A(n_5),
.B(n_12),
.Y(n_36)
);

CKINVDCx14_ASAP7_75t_R g37 ( 
.A(n_0),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_12),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_40),
.Y(n_91)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_16),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_41),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_36),
.B(n_8),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g88 ( 
.A(n_42),
.B(n_46),
.Y(n_88)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_16),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g99 ( 
.A(n_43),
.Y(n_99)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_44),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_45),
.Y(n_102)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_23),
.Y(n_46)
);

BUFx12f_ASAP7_75t_L g47 ( 
.A(n_31),
.Y(n_47)
);

BUFx12f_ASAP7_75t_L g101 ( 
.A(n_47),
.Y(n_101)
);

INVx11_ASAP7_75t_L g48 ( 
.A(n_18),
.Y(n_48)
);

INVx8_ASAP7_75t_L g86 ( 
.A(n_48),
.Y(n_86)
);

INVx6_ASAP7_75t_L g49 ( 
.A(n_32),
.Y(n_49)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_49),
.Y(n_79)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_31),
.Y(n_50)
);

INVx5_ASAP7_75t_SL g95 ( 
.A(n_50),
.Y(n_95)
);

BUFx12f_ASAP7_75t_L g51 ( 
.A(n_20),
.Y(n_51)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_36),
.B(n_8),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_53),
.B(n_60),
.Y(n_74)
);

INVx11_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx2_ASAP7_75t_SL g103 ( 
.A(n_54),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g55 ( 
.A(n_20),
.Y(n_55)
);

BUFx3_ASAP7_75t_L g70 ( 
.A(n_55),
.Y(n_70)
);

BUFx12f_ASAP7_75t_L g56 ( 
.A(n_21),
.Y(n_56)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_56),
.Y(n_110)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

INVx3_ASAP7_75t_L g69 ( 
.A(n_57),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_21),
.Y(n_58)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_58),
.Y(n_81)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_30),
.Y(n_59)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_59),
.Y(n_90)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_32),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_22),
.B(n_1),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_61),
.B(n_2),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_30),
.Y(n_62)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_62),
.Y(n_94)
);

INVx2_ASAP7_75t_SL g63 ( 
.A(n_32),
.Y(n_63)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_63),
.Y(n_96)
);

INVx2_ASAP7_75t_L g64 ( 
.A(n_17),
.Y(n_64)
);

INVx6_ASAP7_75t_L g77 ( 
.A(n_64),
.Y(n_77)
);

INVx4_ASAP7_75t_L g65 ( 
.A(n_32),
.Y(n_65)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_65),
.B(n_66),
.Y(n_83)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_30),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g67 ( 
.A(n_46),
.B(n_23),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_67),
.B(n_106),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_44),
.A2(n_24),
.B1(n_26),
.B2(n_19),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_71),
.A2(n_80),
.B1(n_82),
.B2(n_87),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_61),
.B(n_26),
.Y(n_72)
);

AND2x2_ASAP7_75t_L g122 ( 
.A(n_72),
.B(n_75),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_64),
.B(n_22),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g76 ( 
.A1(n_49),
.A2(n_24),
.B1(n_19),
.B2(n_33),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_76),
.A2(n_106),
.B1(n_69),
.B2(n_73),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_L g78 ( 
.A1(n_60),
.A2(n_24),
.B1(n_37),
.B2(n_34),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g130 ( 
.A1(n_78),
.A2(n_105),
.B1(n_109),
.B2(n_56),
.Y(n_130)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_48),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_54),
.A2(n_25),
.B1(n_29),
.B2(n_35),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g84 ( 
.A(n_63),
.B(n_39),
.Y(n_84)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_84),
.Y(n_143)
);

AOI22xp33_ASAP7_75t_SL g87 ( 
.A1(n_65),
.A2(n_28),
.B1(n_34),
.B2(n_39),
.Y(n_87)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_63),
.B(n_27),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_89),
.B(n_92),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_L g92 ( 
.A(n_52),
.B(n_27),
.Y(n_92)
);

AOI21xp5_ASAP7_75t_L g93 ( 
.A1(n_51),
.A2(n_18),
.B(n_3),
.Y(n_93)
);

O2A1O1Ixp33_ASAP7_75t_L g136 ( 
.A1(n_93),
.A2(n_105),
.B(n_73),
.C(n_95),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_52),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_97),
.B(n_104),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_40),
.B(n_28),
.Y(n_100)
);

AND2x2_ASAP7_75t_L g151 ( 
.A(n_100),
.B(n_5),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_66),
.B(n_27),
.Y(n_104)
);

AOI22xp5_ASAP7_75t_SL g105 ( 
.A1(n_57),
.A2(n_38),
.B1(n_18),
.B2(n_32),
.Y(n_105)
);

AOI22xp33_ASAP7_75t_SL g107 ( 
.A1(n_66),
.A2(n_38),
.B1(n_11),
.B2(n_12),
.Y(n_107)
);

OAI22xp5_ASAP7_75t_L g117 ( 
.A1(n_107),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_117)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_58),
.B(n_15),
.Y(n_108)
);

NOR2xp33_ASAP7_75t_L g142 ( 
.A(n_108),
.B(n_2),
.Y(n_142)
);

AOI22xp33_ASAP7_75t_L g109 ( 
.A1(n_59),
.A2(n_38),
.B1(n_15),
.B2(n_10),
.Y(n_109)
);

OAI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_113),
.A2(n_117),
.B1(n_129),
.B2(n_130),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g114 ( 
.A1(n_76),
.A2(n_62),
.B1(n_45),
.B2(n_43),
.Y(n_114)
);

OAI22xp5_ASAP7_75t_SL g157 ( 
.A1(n_114),
.A2(n_139),
.B1(n_95),
.B2(n_94),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_98),
.Y(n_116)
);

INVx4_ASAP7_75t_L g161 ( 
.A(n_116),
.Y(n_161)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_72),
.B(n_50),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g168 ( 
.A(n_118),
.B(n_140),
.Y(n_168)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_103),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_119),
.B(n_120),
.Y(n_158)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_96),
.Y(n_120)
);

INVx3_ASAP7_75t_L g121 ( 
.A(n_96),
.Y(n_121)
);

INVx1_ASAP7_75t_L g163 ( 
.A(n_121),
.Y(n_163)
);

INVx5_ASAP7_75t_L g123 ( 
.A(n_86),
.Y(n_123)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_123),
.Y(n_155)
);

INVx2_ASAP7_75t_L g124 ( 
.A(n_77),
.Y(n_124)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_124),
.Y(n_184)
);

AOI22xp33_ASAP7_75t_SL g125 ( 
.A1(n_69),
.A2(n_14),
.B1(n_13),
.B2(n_11),
.Y(n_125)
);

AOI21xp5_ASAP7_75t_L g165 ( 
.A1(n_125),
.A2(n_127),
.B(n_144),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_40),
.C(n_50),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g183 ( 
.A(n_126),
.B(n_101),
.C(n_130),
.Y(n_183)
);

AOI21xp33_ASAP7_75t_L g127 ( 
.A1(n_106),
.A2(n_15),
.B(n_3),
.Y(n_127)
);

CKINVDCx14_ASAP7_75t_R g128 ( 
.A(n_67),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_128),
.B(n_131),
.Y(n_159)
);

OAI22xp33_ASAP7_75t_SL g129 ( 
.A1(n_77),
.A2(n_41),
.B1(n_56),
.B2(n_55),
.Y(n_129)
);

INVx2_ASAP7_75t_SL g131 ( 
.A(n_91),
.Y(n_131)
);

INVx1_ASAP7_75t_L g132 ( 
.A(n_75),
.Y(n_132)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_132),
.B(n_134),
.Y(n_164)
);

OAI22xp5_ASAP7_75t_L g133 ( 
.A1(n_88),
.A2(n_56),
.B1(n_55),
.B2(n_51),
.Y(n_133)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_133),
.A2(n_94),
.B1(n_90),
.B2(n_98),
.Y(n_160)
);

CKINVDCx14_ASAP7_75t_R g134 ( 
.A(n_100),
.Y(n_134)
);

INVx1_ASAP7_75t_L g135 ( 
.A(n_85),
.Y(n_135)
);

NOR2xp33_ASAP7_75t_L g166 ( 
.A(n_135),
.B(n_137),
.Y(n_166)
);

CKINVDCx14_ASAP7_75t_R g172 ( 
.A(n_136),
.Y(n_172)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_85),
.Y(n_137)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_81),
.A2(n_55),
.B1(n_51),
.B2(n_40),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_L g140 ( 
.A(n_88),
.B(n_47),
.Y(n_140)
);

INVx3_ASAP7_75t_L g141 ( 
.A(n_79),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_141),
.B(n_142),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g144 ( 
.A1(n_95),
.A2(n_3),
.B1(n_5),
.B2(n_6),
.Y(n_144)
);

NAND2xp5_ASAP7_75t_L g145 ( 
.A(n_74),
.B(n_47),
.Y(n_145)
);

NAND2xp5_ASAP7_75t_SL g153 ( 
.A(n_145),
.B(n_151),
.Y(n_153)
);

OA22x2_ASAP7_75t_L g146 ( 
.A1(n_81),
.A2(n_47),
.B1(n_50),
.B2(n_6),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g186 ( 
.A1(n_146),
.A2(n_124),
.B1(n_123),
.B2(n_148),
.Y(n_186)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_110),
.Y(n_147)
);

NOR2xp33_ASAP7_75t_L g182 ( 
.A(n_147),
.B(n_149),
.Y(n_182)
);

INVx2_ASAP7_75t_L g148 ( 
.A(n_79),
.Y(n_148)
);

INVxp67_ASAP7_75t_L g173 ( 
.A(n_148),
.Y(n_173)
);

BUFx2_ASAP7_75t_L g149 ( 
.A(n_91),
.Y(n_149)
);

NAND2xp5_ASAP7_75t_SL g150 ( 
.A(n_83),
.B(n_3),
.Y(n_150)
);

NOR2xp33_ASAP7_75t_SL g185 ( 
.A(n_150),
.B(n_112),
.Y(n_185)
);

INVx4_ASAP7_75t_L g152 ( 
.A(n_110),
.Y(n_152)
);

CKINVDCx16_ASAP7_75t_R g156 ( 
.A(n_152),
.Y(n_156)
);

OR2x2_ASAP7_75t_L g154 ( 
.A(n_132),
.B(n_86),
.Y(n_154)
);

OAI21xp5_ASAP7_75t_L g204 ( 
.A1(n_154),
.A2(n_174),
.B(n_180),
.Y(n_204)
);

OAI22xp5_ASAP7_75t_L g208 ( 
.A1(n_157),
.A2(n_160),
.B1(n_186),
.B2(n_131),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_126),
.A2(n_90),
.B1(n_102),
.B2(n_99),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_SL g192 ( 
.A1(n_162),
.A2(n_177),
.B1(n_178),
.B2(n_187),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_122),
.B(n_91),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_167),
.B(n_170),
.Y(n_197)
);

CKINVDCx16_ASAP7_75t_R g169 ( 
.A(n_135),
.Y(n_169)
);

NAND2xp5_ASAP7_75t_SL g188 ( 
.A(n_169),
.B(n_185),
.Y(n_188)
);

NAND2xp5_ASAP7_75t_SL g170 ( 
.A(n_122),
.B(n_91),
.Y(n_170)
);

AND2x2_ASAP7_75t_L g174 ( 
.A(n_118),
.B(n_5),
.Y(n_174)
);

AOI22xp5_ASAP7_75t_L g175 ( 
.A1(n_122),
.A2(n_98),
.B1(n_99),
.B2(n_102),
.Y(n_175)
);

OAI22xp5_ASAP7_75t_L g198 ( 
.A1(n_175),
.A2(n_179),
.B1(n_146),
.B2(n_120),
.Y(n_198)
);

OAI22xp5_ASAP7_75t_SL g177 ( 
.A1(n_113),
.A2(n_99),
.B1(n_102),
.B2(n_68),
.Y(n_177)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_136),
.A2(n_68),
.B1(n_70),
.B2(n_101),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g179 ( 
.A1(n_111),
.A2(n_6),
.B1(n_7),
.B2(n_70),
.Y(n_179)
);

AOI21xp5_ASAP7_75t_L g180 ( 
.A1(n_146),
.A2(n_101),
.B(n_6),
.Y(n_180)
);

OAI32xp33_ASAP7_75t_L g181 ( 
.A1(n_145),
.A2(n_7),
.A3(n_101),
.B1(n_140),
.B2(n_138),
.Y(n_181)
);

CKINVDCx14_ASAP7_75t_R g212 ( 
.A(n_181),
.Y(n_212)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_183),
.B(n_131),
.C(n_143),
.Y(n_203)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_139),
.A2(n_137),
.B1(n_146),
.B2(n_141),
.Y(n_187)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_166),
.Y(n_189)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_189),
.Y(n_224)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_166),
.Y(n_190)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_190),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_163),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g221 ( 
.A(n_191),
.B(n_211),
.Y(n_221)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_184),
.Y(n_193)
);

INVx1_ASAP7_75t_L g229 ( 
.A(n_193),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_172),
.A2(n_183),
.B1(n_171),
.B2(n_168),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g228 ( 
.A1(n_194),
.A2(n_198),
.B1(n_208),
.B2(n_210),
.Y(n_228)
);

NOR4xp25_ASAP7_75t_L g195 ( 
.A(n_168),
.B(n_115),
.C(n_151),
.D(n_152),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_SL g236 ( 
.A(n_195),
.B(n_200),
.Y(n_236)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_184),
.Y(n_196)
);

CKINVDCx16_ASAP7_75t_R g217 ( 
.A(n_196),
.Y(n_217)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_182),
.Y(n_199)
);

CKINVDCx16_ASAP7_75t_R g240 ( 
.A(n_199),
.Y(n_240)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_167),
.B(n_170),
.Y(n_200)
);

INVxp67_ASAP7_75t_L g201 ( 
.A(n_155),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g230 ( 
.A(n_201),
.B(n_205),
.Y(n_230)
);

NOR2x1_ASAP7_75t_L g202 ( 
.A(n_181),
.B(n_151),
.Y(n_202)
);

NOR2xp33_ASAP7_75t_SL g220 ( 
.A(n_202),
.B(n_154),
.Y(n_220)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_203),
.B(n_153),
.C(n_178),
.Y(n_218)
);

INVx8_ASAP7_75t_L g205 ( 
.A(n_155),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_174),
.B(n_121),
.Y(n_206)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_206),
.B(n_209),
.Y(n_233)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_182),
.Y(n_207)
);

CKINVDCx20_ASAP7_75t_R g223 ( 
.A(n_207),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g209 ( 
.A(n_174),
.B(n_154),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_SL g210 ( 
.A1(n_180),
.A2(n_116),
.B1(n_149),
.B2(n_179),
.Y(n_210)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_163),
.Y(n_211)
);

AOI22xp5_ASAP7_75t_L g213 ( 
.A1(n_187),
.A2(n_186),
.B1(n_162),
.B2(n_177),
.Y(n_213)
);

AOI22xp5_ASAP7_75t_L g232 ( 
.A1(n_213),
.A2(n_186),
.B1(n_175),
.B2(n_157),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g214 ( 
.A(n_159),
.B(n_176),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_214),
.B(n_215),
.Y(n_225)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_158),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g216 ( 
.A(n_158),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g231 ( 
.A(n_216),
.B(n_169),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g241 ( 
.A(n_218),
.B(n_219),
.C(n_226),
.Y(n_241)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_203),
.B(n_153),
.C(n_164),
.Y(n_219)
);

AOI221xp5_ASAP7_75t_L g257 ( 
.A1(n_220),
.A2(n_238),
.B1(n_233),
.B2(n_236),
.C(n_240),
.Y(n_257)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_212),
.A2(n_202),
.B1(n_165),
.B2(n_216),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_SL g251 ( 
.A1(n_222),
.A2(n_234),
.B(n_235),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g226 ( 
.A(n_200),
.B(n_164),
.C(n_165),
.Y(n_226)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_231),
.Y(n_249)
);

OAI22xp5_ASAP7_75t_L g253 ( 
.A1(n_232),
.A2(n_161),
.B1(n_239),
.B2(n_233),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_204),
.A2(n_159),
.B(n_176),
.Y(n_234)
);

AOI22xp5_ASAP7_75t_SL g235 ( 
.A1(n_198),
.A2(n_207),
.B1(n_199),
.B2(n_215),
.Y(n_235)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_194),
.A2(n_186),
.B(n_156),
.Y(n_237)
);

AOI21xp5_ASAP7_75t_L g255 ( 
.A1(n_237),
.A2(n_234),
.B(n_220),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g238 ( 
.A(n_204),
.B(n_185),
.Y(n_238)
);

INVx1_ASAP7_75t_L g252 ( 
.A(n_238),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_197),
.B(n_156),
.C(n_160),
.Y(n_239)
);

MAJIxp5_ASAP7_75t_L g248 ( 
.A(n_239),
.B(n_191),
.C(n_201),
.Y(n_248)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_235),
.B(n_189),
.Y(n_242)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_242),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_228),
.A2(n_213),
.B1(n_192),
.B2(n_210),
.Y(n_243)
);

OAI22xp5_ASAP7_75t_L g260 ( 
.A1(n_243),
.A2(n_244),
.B1(n_255),
.B2(n_232),
.Y(n_260)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_228),
.A2(n_192),
.B1(n_197),
.B2(n_209),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g245 ( 
.A(n_236),
.B(n_206),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_245),
.B(n_248),
.C(n_218),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_L g246 ( 
.A(n_223),
.B(n_190),
.Y(n_246)
);

CKINVDCx14_ASAP7_75t_R g266 ( 
.A(n_246),
.Y(n_266)
);

AOI322xp5_ASAP7_75t_L g247 ( 
.A1(n_237),
.A2(n_195),
.A3(n_188),
.B1(n_186),
.B2(n_211),
.C1(n_193),
.C2(n_196),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_247),
.B(n_256),
.Y(n_261)
);

AO221x1_ASAP7_75t_L g250 ( 
.A1(n_230),
.A2(n_161),
.B1(n_173),
.B2(n_205),
.C(n_221),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

AOI22xp5_ASAP7_75t_L g267 ( 
.A1(n_253),
.A2(n_217),
.B1(n_229),
.B2(n_248),
.Y(n_267)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_223),
.B(n_161),
.Y(n_254)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

AOI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_240),
.A2(n_224),
.B1(n_227),
.B2(n_222),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g271 ( 
.A(n_257),
.B(n_258),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g258 ( 
.A(n_225),
.Y(n_258)
);

NAND2xp5_ASAP7_75t_SL g259 ( 
.A(n_224),
.B(n_227),
.Y(n_259)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_259),
.B(n_246),
.Y(n_272)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_260),
.Y(n_273)
);

XNOR2xp5_ASAP7_75t_L g283 ( 
.A(n_263),
.B(n_251),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_241),
.B(n_226),
.C(n_219),
.Y(n_264)
);

XOR2xp5_ASAP7_75t_L g280 ( 
.A(n_264),
.B(n_265),
.Y(n_280)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_241),
.B(n_229),
.C(n_217),
.Y(n_265)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_267),
.B(n_243),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g270 ( 
.A(n_245),
.B(n_253),
.C(n_244),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g282 ( 
.A(n_270),
.B(n_251),
.Y(n_282)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_272),
.Y(n_274)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_266),
.B(n_249),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_SL g288 ( 
.A(n_275),
.B(n_276),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g276 ( 
.A1(n_262),
.A2(n_242),
.B(n_255),
.Y(n_276)
);

OAI21xp5_ASAP7_75t_L g277 ( 
.A1(n_262),
.A2(n_256),
.B(n_252),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g285 ( 
.A1(n_277),
.A2(n_278),
.B1(n_273),
.B2(n_267),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g278 ( 
.A(n_268),
.B(n_259),
.Y(n_278)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_278),
.Y(n_287)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_279),
.B(n_281),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_269),
.B(n_249),
.Y(n_281)
);

NOR2xp33_ASAP7_75t_L g286 ( 
.A(n_282),
.B(n_283),
.Y(n_286)
);

OAI322xp33_ASAP7_75t_L g284 ( 
.A1(n_274),
.A2(n_252),
.A3(n_271),
.B1(n_261),
.B2(n_264),
.C1(n_265),
.C2(n_263),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g294 ( 
.A1(n_284),
.A2(n_283),
.B(n_280),
.Y(n_294)
);

A2O1A1Ixp33_ASAP7_75t_SL g292 ( 
.A1(n_285),
.A2(n_291),
.B(n_269),
.C(n_250),
.Y(n_292)
);

HB1xp67_ASAP7_75t_L g289 ( 
.A(n_277),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g296 ( 
.A(n_289),
.B(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g291 ( 
.A(n_276),
.Y(n_291)
);

AOI31xp67_ASAP7_75t_SL g298 ( 
.A1(n_292),
.A2(n_295),
.A3(n_296),
.B(n_285),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_288),
.B(n_270),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g299 ( 
.A(n_293),
.B(n_294),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g295 ( 
.A1(n_291),
.A2(n_254),
.B1(n_282),
.B2(n_280),
.Y(n_295)
);

OAI21xp5_ASAP7_75t_SL g297 ( 
.A1(n_292),
.A2(n_286),
.B(n_290),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_297),
.B(n_298),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g301 ( 
.A(n_299),
.Y(n_301)
);

NAND2xp5_ASAP7_75t_L g302 ( 
.A(n_301),
.B(n_287),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g303 ( 
.A(n_302),
.B(n_300),
.Y(n_303)
);


endmodule