module real_jpeg_27646_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;

output n_17;

wire n_108;
wire n_54;
wire n_37;
wire n_233;
wire n_168;
wire n_73;
wire n_35;
wire n_38;
wire n_29;
wire n_91;
wire n_49;
wire n_114;
wire n_201;
wire n_68;
wire n_146;
wire n_247;
wire n_83;
wire n_78;
wire n_249;
wire n_215;
wire n_166;
wire n_176;
wire n_221;
wire n_104;
wire n_153;
wire n_194;
wire n_161;
wire n_207;
wire n_64;
wire n_177;
wire n_236;
wire n_47;
wire n_131;
wire n_163;
wire n_22;
wire n_174;
wire n_237;
wire n_87;
wire n_197;
wire n_40;
wire n_105;
wire n_243;
wire n_173;
wire n_115;
wire n_98;
wire n_27;
wire n_56;
wire n_184;
wire n_48;
wire n_164;
wire n_200;
wire n_140;
wire n_227;
wire n_126;
wire n_229;
wire n_214;
wire n_113;
wire n_120;
wire n_155;
wire n_199;
wire n_251;
wire n_93;
wire n_95;
wire n_242;
wire n_141;
wire n_65;
wire n_33;
wire n_139;
wire n_188;
wire n_142;
wire n_175;
wire n_76;
wire n_238;
wire n_67;
wire n_79;
wire n_178;
wire n_235;
wire n_107;
wire n_156;
wire n_147;
wire n_189;
wire n_170;
wire n_66;
wire n_231;
wire n_136;
wire n_44;
wire n_28;
wire n_208;
wire n_62;
wire n_162;
wire n_239;
wire n_245;
wire n_250;
wire n_121;
wire n_234;
wire n_106;
wire n_172;
wire n_211;
wire n_160;
wire n_45;
wire n_112;
wire n_42;
wire n_18;
wire n_145;
wire n_77;
wire n_109;
wire n_39;
wire n_219;
wire n_122;
wire n_94;
wire n_26;
wire n_19;
wire n_148;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_116;
wire n_246;
wire n_21;
wire n_50;
wire n_143;
wire n_196;
wire n_69;
wire n_186;
wire n_137;
wire n_31;
wire n_129;
wire n_154;
wire n_135;
wire n_152;
wire n_218;
wire n_165;
wire n_134;
wire n_223;
wire n_72;
wire n_159;
wire n_171;
wire n_151;
wire n_183;
wire n_248;
wire n_198;
wire n_203;
wire n_100;
wire n_192;
wire n_23;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_195;
wire n_110;
wire n_205;
wire n_117;
wire n_193;
wire n_99;
wire n_86;
wire n_150;
wire n_41;
wire n_80;
wire n_74;
wire n_32;
wire n_20;
wire n_70;
wire n_228;
wire n_30;
wire n_204;
wire n_158;
wire n_149;
wire n_144;
wire n_130;
wire n_241;
wire n_103;
wire n_225;
wire n_232;
wire n_57;
wire n_43;
wire n_157;
wire n_84;
wire n_212;
wire n_82;
wire n_111;
wire n_132;
wire n_226;
wire n_125;
wire n_185;
wire n_240;
wire n_55;
wire n_209;
wire n_180;
wire n_58;
wire n_52;
wire n_191;
wire n_63;
wire n_124;
wire n_24;
wire n_92;
wire n_75;
wire n_97;
wire n_187;
wire n_34;
wire n_230;
wire n_190;
wire n_60;
wire n_46;
wire n_88;
wire n_169;
wire n_59;
wire n_128;
wire n_202;
wire n_167;
wire n_244;
wire n_179;
wire n_216;
wire n_133;
wire n_213;
wire n_138;
wire n_25;
wire n_217;
wire n_53;
wire n_210;
wire n_127;
wire n_206;
wire n_224;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_181;
wire n_101;
wire n_182;
wire n_96;
wire n_89;

OAI22xp5_ASAP7_75t_SL g65 ( 
.A1(n_0),
.A2(n_56),
.B1(n_57),
.B2(n_66),
.Y(n_65)
);

CKINVDCx16_ASAP7_75t_R g66 ( 
.A(n_0),
.Y(n_66)
);

OAI22xp5_ASAP7_75t_L g113 ( 
.A1(n_0),
.A2(n_62),
.B1(n_63),
.B2(n_66),
.Y(n_113)
);

AOI22xp33_ASAP7_75t_SL g195 ( 
.A1(n_0),
.A2(n_26),
.B1(n_33),
.B2(n_66),
.Y(n_195)
);

OAI22xp5_ASAP7_75t_SL g227 ( 
.A1(n_0),
.A2(n_39),
.B1(n_40),
.B2(n_66),
.Y(n_227)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_1),
.Y(n_29)
);

INVx11_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

AOI22xp33_ASAP7_75t_L g48 ( 
.A1(n_2),
.A2(n_39),
.B1(n_40),
.B2(n_49),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_2),
.Y(n_49)
);

AOI22xp33_ASAP7_75t_SL g106 ( 
.A1(n_2),
.A2(n_26),
.B1(n_33),
.B2(n_49),
.Y(n_106)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_2),
.A2(n_49),
.B1(n_62),
.B2(n_63),
.Y(n_134)
);

CKINVDCx20_ASAP7_75t_R g100 ( 
.A(n_3),
.Y(n_100)
);

AOI21xp5_ASAP7_75t_L g101 ( 
.A1(n_3),
.A2(n_61),
.B(n_62),
.Y(n_101)
);

OAI22xp33_ASAP7_75t_SL g153 ( 
.A1(n_3),
.A2(n_56),
.B1(n_57),
.B2(n_100),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g183 ( 
.A(n_3),
.B(n_39),
.Y(n_183)
);

A2O1A1O1Ixp25_ASAP7_75t_L g185 ( 
.A1(n_3),
.A2(n_39),
.B(n_43),
.C(n_183),
.D(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_3),
.B(n_71),
.Y(n_190)
);

OAI21xp33_ASAP7_75t_L g213 ( 
.A1(n_3),
.A2(n_25),
.B(n_196),
.Y(n_213)
);

A2O1A1O1Ixp25_ASAP7_75t_L g223 ( 
.A1(n_3),
.A2(n_63),
.B(n_76),
.C(n_115),
.D(n_224),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_3),
.B(n_63),
.Y(n_224)
);

OAI22xp5_ASAP7_75t_L g54 ( 
.A1(n_4),
.A2(n_55),
.B1(n_56),
.B2(n_57),
.Y(n_54)
);

INVx1_ASAP7_75t_L g55 ( 
.A(n_4),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_L g157 ( 
.A1(n_4),
.A2(n_55),
.B1(n_62),
.B2(n_63),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g193 ( 
.A1(n_4),
.A2(n_39),
.B1(n_40),
.B2(n_55),
.Y(n_193)
);

AOI22xp33_ASAP7_75t_SL g203 ( 
.A1(n_4),
.A2(n_26),
.B1(n_33),
.B2(n_55),
.Y(n_203)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g38 ( 
.A1(n_6),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_SL g69 ( 
.A1(n_6),
.A2(n_41),
.B1(n_62),
.B2(n_63),
.Y(n_69)
);

AOI22xp33_ASAP7_75t_L g172 ( 
.A1(n_6),
.A2(n_26),
.B1(n_33),
.B2(n_41),
.Y(n_172)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_7),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g79 ( 
.A1(n_8),
.A2(n_62),
.B1(n_63),
.B2(n_80),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g80 ( 
.A(n_8),
.Y(n_80)
);

OAI22xp5_ASAP7_75t_SL g96 ( 
.A1(n_8),
.A2(n_56),
.B1(n_57),
.B2(n_80),
.Y(n_96)
);

AOI22xp33_ASAP7_75t_L g151 ( 
.A1(n_8),
.A2(n_39),
.B1(n_40),
.B2(n_80),
.Y(n_151)
);

AOI22xp5_ASAP7_75t_L g198 ( 
.A1(n_8),
.A2(n_26),
.B1(n_33),
.B2(n_80),
.Y(n_198)
);

BUFx3_ASAP7_75t_L g56 ( 
.A(n_9),
.Y(n_56)
);

AOI22xp33_ASAP7_75t_SL g85 ( 
.A1(n_10),
.A2(n_26),
.B1(n_33),
.B2(n_86),
.Y(n_85)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_10),
.Y(n_86)
);

O2A1O1Ixp33_ASAP7_75t_L g43 ( 
.A1(n_11),
.A2(n_39),
.B(n_44),
.C(n_47),
.Y(n_43)
);

INVx11_ASAP7_75t_L g46 ( 
.A(n_11),
.Y(n_46)
);

AOI22xp33_ASAP7_75t_L g35 ( 
.A1(n_12),
.A2(n_26),
.B1(n_33),
.B2(n_36),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_12),
.Y(n_36)
);

OAI22xp5_ASAP7_75t_L g122 ( 
.A1(n_12),
.A2(n_36),
.B1(n_39),
.B2(n_40),
.Y(n_122)
);

BUFx24_ASAP7_75t_L g62 ( 
.A(n_13),
.Y(n_62)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_14),
.Y(n_72)
);

INVx4_ASAP7_75t_L g74 ( 
.A(n_14),
.Y(n_74)
);

OAI22xp5_ASAP7_75t_SL g31 ( 
.A1(n_15),
.A2(n_26),
.B1(n_32),
.B2(n_33),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_15),
.Y(n_32)
);

AOI22xp33_ASAP7_75t_L g88 ( 
.A1(n_15),
.A2(n_32),
.B1(n_39),
.B2(n_40),
.Y(n_88)
);

INVx11_ASAP7_75t_SL g28 ( 
.A(n_16),
.Y(n_28)
);

XNOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_138),
.Y(n_17)
);

NAND2xp5_ASAP7_75t_L g18 ( 
.A(n_19),
.B(n_137),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_20),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_116),
.Y(n_20)
);

NAND2xp5_ASAP7_75t_SL g137 ( 
.A(n_21),
.B(n_116),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_81),
.C(n_89),
.Y(n_21)
);

XNOR2xp5_ASAP7_75t_SL g159 ( 
.A(n_22),
.B(n_81),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_SL g22 ( 
.A(n_23),
.B(n_51),
.Y(n_22)
);

MAJIxp5_ASAP7_75t_L g136 ( 
.A(n_23),
.B(n_53),
.C(n_67),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_37),
.Y(n_23)
);

XOR2xp5_ASAP7_75t_L g145 ( 
.A(n_24),
.B(n_37),
.Y(n_145)
);

OAI22xp5_ASAP7_75t_L g24 ( 
.A1(n_25),
.A2(n_30),
.B1(n_34),
.B2(n_35),
.Y(n_24)
);

OAI22xp5_ASAP7_75t_L g82 ( 
.A1(n_25),
.A2(n_35),
.B1(n_83),
.B2(n_85),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_25),
.Y(n_104)
);

AOI21xp5_ASAP7_75t_L g124 ( 
.A1(n_25),
.A2(n_85),
.B(n_108),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_25),
.A2(n_106),
.B1(n_108),
.B2(n_172),
.Y(n_171)
);

OAI21xp5_ASAP7_75t_L g194 ( 
.A1(n_25),
.A2(n_195),
.B(n_196),
.Y(n_194)
);

NOR2xp33_ASAP7_75t_L g211 ( 
.A(n_25),
.B(n_198),
.Y(n_211)
);

NAND2x1_ASAP7_75t_SL g25 ( 
.A(n_26),
.B(n_29),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_26),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_26),
.A2(n_33),
.B1(n_45),
.B2(n_46),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g184 ( 
.A(n_26),
.B(n_45),
.Y(n_184)
);

BUFx2_ASAP7_75t_L g26 ( 
.A(n_27),
.Y(n_26)
);

INVx11_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_31),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_L g103 ( 
.A1(n_31),
.A2(n_104),
.B1(n_105),
.B2(n_107),
.Y(n_103)
);

AOI32xp33_ASAP7_75t_L g182 ( 
.A1(n_33),
.A2(n_40),
.A3(n_46),
.B1(n_183),
.B2(n_184),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_33),
.B(n_215),
.Y(n_214)
);

INVx11_ASAP7_75t_L g84 ( 
.A(n_34),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_34),
.B(n_100),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_48),
.B2(n_50),
.Y(n_37)
);

OAI21xp5_ASAP7_75t_SL g148 ( 
.A1(n_38),
.A2(n_50),
.B(n_149),
.Y(n_148)
);

NAND2xp5_ASAP7_75t_SL g44 ( 
.A(n_39),
.B(n_45),
.Y(n_44)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_39),
.A2(n_40),
.B1(n_72),
.B2(n_73),
.Y(n_71)
);

AOI32xp33_ASAP7_75t_L g231 ( 
.A1(n_39),
.A2(n_62),
.A3(n_224),
.B1(n_232),
.B2(n_233),
.Y(n_231)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_40),
.Y(n_39)
);

NAND2xp33_ASAP7_75t_SL g233 ( 
.A(n_40),
.B(n_73),
.Y(n_233)
);

OAI22xp5_ASAP7_75t_L g87 ( 
.A1(n_42),
.A2(n_48),
.B1(n_50),
.B2(n_88),
.Y(n_87)
);

OAI21xp5_ASAP7_75t_SL g241 ( 
.A1(n_42),
.A2(n_242),
.B(n_243),
.Y(n_241)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_43),
.Y(n_42)
);

AOI22xp5_ASAP7_75t_L g120 ( 
.A1(n_43),
.A2(n_47),
.B1(n_121),
.B2(n_122),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_43),
.B(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_L g225 ( 
.A1(n_43),
.A2(n_47),
.B1(n_226),
.B2(n_227),
.Y(n_225)
);

INVx11_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_47),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g186 ( 
.A(n_50),
.B(n_151),
.Y(n_186)
);

OAI21xp5_ASAP7_75t_L g192 ( 
.A1(n_50),
.A2(n_149),
.B(n_193),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g208 ( 
.A(n_50),
.B(n_100),
.Y(n_208)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_53),
.B1(n_67),
.B2(n_68),
.Y(n_51)
);

CKINVDCx14_ASAP7_75t_R g52 ( 
.A(n_53),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g53 ( 
.A1(n_54),
.A2(n_58),
.B1(n_59),
.B2(n_65),
.Y(n_53)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g57 ( 
.A(n_56),
.Y(n_57)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_56),
.A2(n_57),
.B1(n_60),
.B2(n_61),
.Y(n_64)
);

A2O1A1Ixp33_ASAP7_75t_L g99 ( 
.A1(n_56),
.A2(n_60),
.B(n_100),
.C(n_101),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_58),
.B(n_96),
.Y(n_95)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_58),
.Y(n_130)
);

AOI21xp5_ASAP7_75t_L g152 ( 
.A1(n_58),
.A2(n_153),
.B(n_154),
.Y(n_152)
);

NOR2xp33_ASAP7_75t_SL g58 ( 
.A(n_59),
.B(n_64),
.Y(n_58)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_59),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g132 ( 
.A(n_59),
.B(n_96),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g59 ( 
.A1(n_60),
.A2(n_61),
.B1(n_62),
.B2(n_63),
.Y(n_59)
);

CKINVDCx14_ASAP7_75t_R g60 ( 
.A(n_61),
.Y(n_60)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_62),
.Y(n_63)
);

AOI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_62),
.A2(n_63),
.B1(n_73),
.B2(n_74),
.Y(n_77)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_65),
.Y(n_131)
);

CKINVDCx16_ASAP7_75t_R g67 ( 
.A(n_68),
.Y(n_67)
);

OAI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_70),
.B(n_75),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g133 ( 
.A1(n_69),
.A2(n_70),
.B1(n_111),
.B2(n_134),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_70),
.B(n_79),
.Y(n_115)
);

OAI21xp5_ASAP7_75t_L g170 ( 
.A1(n_70),
.A2(n_75),
.B(n_157),
.Y(n_170)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_SL g76 ( 
.A(n_71),
.B(n_77),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g155 ( 
.A1(n_71),
.A2(n_76),
.B1(n_113),
.B2(n_156),
.Y(n_155)
);

INVx6_ASAP7_75t_L g232 ( 
.A(n_73),
.Y(n_232)
);

INVx8_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_76),
.B(n_78),
.Y(n_75)
);

INVx1_ASAP7_75t_L g111 ( 
.A(n_76),
.Y(n_111)
);

INVxp67_ASAP7_75t_L g78 ( 
.A(n_79),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_87),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g126 ( 
.A(n_82),
.B(n_87),
.Y(n_126)
);

INVx5_ASAP7_75t_SL g83 ( 
.A(n_84),
.Y(n_83)
);

INVx11_ASAP7_75t_L g108 ( 
.A(n_84),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g196 ( 
.A(n_84),
.B(n_197),
.Y(n_196)
);

AOI21xp5_ASAP7_75t_L g229 ( 
.A1(n_84),
.A2(n_211),
.B(n_230),
.Y(n_229)
);

CKINVDCx20_ASAP7_75t_R g121 ( 
.A(n_88),
.Y(n_121)
);

AOI22xp5_ASAP7_75t_SL g158 ( 
.A1(n_89),
.A2(n_90),
.B1(n_159),
.B2(n_160),
.Y(n_158)
);

INVx1_ASAP7_75t_L g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g90 ( 
.A(n_91),
.B(n_97),
.C(n_109),
.Y(n_90)
);

AOI22xp5_ASAP7_75t_L g144 ( 
.A1(n_91),
.A2(n_92),
.B1(n_109),
.B2(n_110),
.Y(n_144)
);

CKINVDCx20_ASAP7_75t_R g91 ( 
.A(n_92),
.Y(n_91)
);

OAI21xp5_ASAP7_75t_L g92 ( 
.A1(n_93),
.A2(n_94),
.B(n_95),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_SL g173 ( 
.A(n_94),
.B(n_100),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g143 ( 
.A(n_97),
.B(n_144),
.Y(n_143)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_102),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_SL g168 ( 
.A1(n_98),
.A2(n_99),
.B1(n_102),
.B2(n_103),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_103),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_104),
.A2(n_107),
.B1(n_202),
.B2(n_204),
.Y(n_201)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_106),
.Y(n_105)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_108),
.Y(n_107)
);

OAI21xp5_ASAP7_75t_SL g209 ( 
.A1(n_108),
.A2(n_203),
.B(n_210),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g109 ( 
.A(n_110),
.Y(n_109)
);

OAI21xp5_ASAP7_75t_SL g110 ( 
.A1(n_111),
.A2(n_112),
.B(n_114),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

INVxp67_ASAP7_75t_L g114 ( 
.A(n_115),
.Y(n_114)
);

XNOR2xp5_ASAP7_75t_L g116 ( 
.A(n_117),
.B(n_136),
.Y(n_116)
);

XNOR2xp5_ASAP7_75t_L g117 ( 
.A(n_118),
.B(n_125),
.Y(n_117)
);

OAI22xp5_ASAP7_75t_SL g118 ( 
.A1(n_119),
.A2(n_120),
.B1(n_123),
.B2(n_124),
.Y(n_118)
);

CKINVDCx14_ASAP7_75t_R g119 ( 
.A(n_120),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_124),
.Y(n_123)
);

OAI22xp5_ASAP7_75t_L g125 ( 
.A1(n_126),
.A2(n_127),
.B1(n_128),
.B2(n_135),
.Y(n_125)
);

CKINVDCx16_ASAP7_75t_R g135 ( 
.A(n_126),
.Y(n_135)
);

INVx1_ASAP7_75t_L g127 ( 
.A(n_128),
.Y(n_127)
);

XNOR2xp5_ASAP7_75t_SL g128 ( 
.A(n_129),
.B(n_133),
.Y(n_128)
);

OAI21xp5_ASAP7_75t_SL g129 ( 
.A1(n_130),
.A2(n_131),
.B(n_132),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_175),
.Y(n_138)
);

INVxp33_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

AOI21xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_161),
.B(n_174),
.Y(n_140)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_141),
.Y(n_250)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_158),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_SL g174 ( 
.A(n_142),
.B(n_158),
.Y(n_174)
);

MAJIxp5_ASAP7_75t_L g142 ( 
.A(n_143),
.B(n_145),
.C(n_146),
.Y(n_142)
);

XNOR2xp5_ASAP7_75t_L g162 ( 
.A(n_143),
.B(n_163),
.Y(n_162)
);

XNOR2xp5_ASAP7_75t_L g163 ( 
.A(n_145),
.B(n_146),
.Y(n_163)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_147),
.B(n_152),
.C(n_155),
.Y(n_146)
);

AOI22xp5_ASAP7_75t_L g166 ( 
.A1(n_147),
.A2(n_148),
.B1(n_155),
.B2(n_167),
.Y(n_166)
);

CKINVDCx20_ASAP7_75t_R g147 ( 
.A(n_148),
.Y(n_147)
);

CKINVDCx16_ASAP7_75t_R g150 ( 
.A(n_151),
.Y(n_150)
);

XNOR2xp5_ASAP7_75t_SL g165 ( 
.A(n_152),
.B(n_166),
.Y(n_165)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_155),
.Y(n_167)
);

CKINVDCx20_ASAP7_75t_R g156 ( 
.A(n_157),
.Y(n_156)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_159),
.Y(n_160)
);

AND2x2_ASAP7_75t_L g161 ( 
.A(n_162),
.B(n_164),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g251 ( 
.A(n_162),
.B(n_164),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g164 ( 
.A(n_165),
.B(n_168),
.C(n_169),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_L g247 ( 
.A(n_165),
.B(n_248),
.Y(n_247)
);

XNOR2xp5_ASAP7_75t_L g248 ( 
.A(n_168),
.B(n_169),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g169 ( 
.A(n_170),
.B(n_171),
.C(n_173),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_170),
.B(n_238),
.Y(n_237)
);

XNOR2xp5_ASAP7_75t_L g238 ( 
.A(n_171),
.B(n_173),
.Y(n_238)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

NOR3xp33_ASAP7_75t_L g175 ( 
.A(n_176),
.B(n_250),
.C(n_251),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_177),
.A2(n_245),
.B(n_249),
.Y(n_176)
);

OAI21xp5_ASAP7_75t_SL g177 ( 
.A1(n_178),
.A2(n_235),
.B(n_244),
.Y(n_177)
);

AOI21xp5_ASAP7_75t_L g178 ( 
.A1(n_179),
.A2(n_219),
.B(n_234),
.Y(n_178)
);

OAI21xp5_ASAP7_75t_SL g179 ( 
.A1(n_180),
.A2(n_199),
.B(n_218),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g180 ( 
.A(n_181),
.B(n_187),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_181),
.B(n_187),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_182),
.B(n_185),
.Y(n_181)
);

XNOR2xp5_ASAP7_75t_L g205 ( 
.A(n_182),
.B(n_185),
.Y(n_205)
);

INVxp67_ASAP7_75t_L g243 ( 
.A(n_186),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g187 ( 
.A(n_188),
.B(n_194),
.Y(n_187)
);

AOI22xp5_ASAP7_75t_L g188 ( 
.A1(n_189),
.A2(n_190),
.B1(n_191),
.B2(n_192),
.Y(n_188)
);

MAJIxp5_ASAP7_75t_L g220 ( 
.A(n_189),
.B(n_192),
.C(n_194),
.Y(n_220)
);

CKINVDCx20_ASAP7_75t_R g189 ( 
.A(n_190),
.Y(n_189)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

CKINVDCx20_ASAP7_75t_R g226 ( 
.A(n_193),
.Y(n_226)
);

CKINVDCx20_ASAP7_75t_R g204 ( 
.A(n_195),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

AOI21xp5_ASAP7_75t_L g199 ( 
.A1(n_200),
.A2(n_206),
.B(n_217),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_205),
.Y(n_200)
);

NOR2xp33_ASAP7_75t_SL g217 ( 
.A(n_201),
.B(n_205),
.Y(n_217)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_203),
.Y(n_202)
);

OAI21xp5_ASAP7_75t_SL g206 ( 
.A1(n_207),
.A2(n_212),
.B(n_216),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_209),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_208),
.B(n_209),
.Y(n_216)
);

INVxp67_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

NAND2xp5_ASAP7_75t_SL g212 ( 
.A(n_213),
.B(n_214),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g219 ( 
.A(n_220),
.B(n_221),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_220),
.B(n_221),
.Y(n_234)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_222),
.Y(n_221)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_222),
.B(n_236),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_222),
.B(n_236),
.Y(n_244)
);

FAx1_ASAP7_75t_SL g222 ( 
.A(n_223),
.B(n_225),
.CI(n_228),
.CON(n_222),
.SN(n_222)
);

INVxp67_ASAP7_75t_L g242 ( 
.A(n_227),
.Y(n_242)
);

XNOR2xp5_ASAP7_75t_SL g228 ( 
.A(n_229),
.B(n_231),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g240 ( 
.A(n_229),
.B(n_231),
.Y(n_240)
);

XOR2xp5_ASAP7_75t_L g236 ( 
.A(n_237),
.B(n_239),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_237),
.B(n_240),
.C(n_241),
.Y(n_246)
);

XOR2xp5_ASAP7_75t_L g239 ( 
.A(n_240),
.B(n_241),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

NOR2xp33_ASAP7_75t_SL g249 ( 
.A(n_246),
.B(n_247),
.Y(n_249)
);


endmodule