module fake_netlist_6_335_n_846 (n_52, n_16, n_1, n_91, n_119, n_46, n_146, n_163, n_18, n_21, n_147, n_154, n_88, n_3, n_98, n_113, n_39, n_63, n_73, n_4, n_148, n_138, n_22, n_161, n_68, n_166, n_28, n_50, n_158, n_49, n_7, n_83, n_5, n_101, n_167, n_144, n_127, n_125, n_153, n_168, n_77, n_156, n_149, n_152, n_106, n_92, n_145, n_42, n_133, n_96, n_8, n_90, n_160, n_24, n_105, n_131, n_54, n_132, n_102, n_0, n_87, n_32, n_66, n_85, n_99, n_78, n_84, n_130, n_164, n_100, n_129, n_13, n_121, n_11, n_137, n_17, n_23, n_142, n_20, n_143, n_2, n_19, n_47, n_62, n_29, n_155, n_75, n_109, n_150, n_122, n_45, n_34, n_140, n_70, n_120, n_37, n_15, n_67, n_33, n_82, n_27, n_38, n_110, n_151, n_61, n_112, n_81, n_59, n_76, n_36, n_26, n_124, n_55, n_126, n_94, n_97, n_108, n_58, n_116, n_64, n_117, n_118, n_48, n_65, n_25, n_40, n_93, n_80, n_141, n_135, n_165, n_139, n_41, n_134, n_114, n_86, n_104, n_95, n_9, n_107, n_10, n_71, n_74, n_6, n_14, n_123, n_136, n_72, n_89, n_103, n_111, n_60, n_159, n_157, n_162, n_170, n_35, n_115, n_12, n_69, n_128, n_30, n_79, n_43, n_171, n_31, n_57, n_169, n_53, n_51, n_44, n_56, n_846);

input n_52;
input n_16;
input n_1;
input n_91;
input n_119;
input n_46;
input n_146;
input n_163;
input n_18;
input n_21;
input n_147;
input n_154;
input n_88;
input n_3;
input n_98;
input n_113;
input n_39;
input n_63;
input n_73;
input n_4;
input n_148;
input n_138;
input n_22;
input n_161;
input n_68;
input n_166;
input n_28;
input n_50;
input n_158;
input n_49;
input n_7;
input n_83;
input n_5;
input n_101;
input n_167;
input n_144;
input n_127;
input n_125;
input n_153;
input n_168;
input n_77;
input n_156;
input n_149;
input n_152;
input n_106;
input n_92;
input n_145;
input n_42;
input n_133;
input n_96;
input n_8;
input n_90;
input n_160;
input n_24;
input n_105;
input n_131;
input n_54;
input n_132;
input n_102;
input n_0;
input n_87;
input n_32;
input n_66;
input n_85;
input n_99;
input n_78;
input n_84;
input n_130;
input n_164;
input n_100;
input n_129;
input n_13;
input n_121;
input n_11;
input n_137;
input n_17;
input n_23;
input n_142;
input n_20;
input n_143;
input n_2;
input n_19;
input n_47;
input n_62;
input n_29;
input n_155;
input n_75;
input n_109;
input n_150;
input n_122;
input n_45;
input n_34;
input n_140;
input n_70;
input n_120;
input n_37;
input n_15;
input n_67;
input n_33;
input n_82;
input n_27;
input n_38;
input n_110;
input n_151;
input n_61;
input n_112;
input n_81;
input n_59;
input n_76;
input n_36;
input n_26;
input n_124;
input n_55;
input n_126;
input n_94;
input n_97;
input n_108;
input n_58;
input n_116;
input n_64;
input n_117;
input n_118;
input n_48;
input n_65;
input n_25;
input n_40;
input n_93;
input n_80;
input n_141;
input n_135;
input n_165;
input n_139;
input n_41;
input n_134;
input n_114;
input n_86;
input n_104;
input n_95;
input n_9;
input n_107;
input n_10;
input n_71;
input n_74;
input n_6;
input n_14;
input n_123;
input n_136;
input n_72;
input n_89;
input n_103;
input n_111;
input n_60;
input n_159;
input n_157;
input n_162;
input n_170;
input n_35;
input n_115;
input n_12;
input n_69;
input n_128;
input n_30;
input n_79;
input n_43;
input n_171;
input n_31;
input n_57;
input n_169;
input n_53;
input n_51;
input n_44;
input n_56;

output n_846;

wire n_591;
wire n_435;
wire n_793;
wire n_326;
wire n_801;
wire n_256;
wire n_440;
wire n_587;
wire n_695;
wire n_507;
wire n_580;
wire n_762;
wire n_209;
wire n_367;
wire n_465;
wire n_680;
wire n_741;
wire n_760;
wire n_590;
wire n_625;
wire n_661;
wire n_223;
wire n_278;
wire n_362;
wire n_341;
wire n_226;
wire n_828;
wire n_208;
wire n_462;
wire n_607;
wire n_726;
wire n_671;
wire n_316;
wire n_419;
wire n_304;
wire n_212;
wire n_700;
wire n_694;
wire n_740;
wire n_578;
wire n_703;
wire n_365;
wire n_384;
wire n_297;
wire n_595;
wire n_627;
wire n_524;
wire n_342;
wire n_820;
wire n_783;
wire n_725;
wire n_358;
wire n_751;
wire n_449;
wire n_749;
wire n_798;
wire n_188;
wire n_310;
wire n_509;
wire n_186;
wire n_245;
wire n_368;
wire n_575;
wire n_677;
wire n_805;
wire n_396;
wire n_495;
wire n_815;
wire n_350;
wire n_585;
wire n_732;
wire n_568;
wire n_392;
wire n_840;
wire n_442;
wire n_480;
wire n_724;
wire n_382;
wire n_673;
wire n_180;
wire n_628;
wire n_557;
wire n_823;
wire n_349;
wire n_643;
wire n_233;
wire n_617;
wire n_698;
wire n_845;
wire n_255;
wire n_807;
wire n_739;
wire n_284;
wire n_400;
wire n_337;
wire n_214;
wire n_485;
wire n_443;
wire n_246;
wire n_768;
wire n_471;
wire n_289;
wire n_421;
wire n_781;
wire n_424;
wire n_789;
wire n_615;
wire n_181;
wire n_182;
wire n_238;
wire n_573;
wire n_769;
wire n_202;
wire n_320;
wire n_639;
wire n_676;
wire n_327;
wire n_794;
wire n_727;
wire n_369;
wire n_597;
wire n_685;
wire n_280;
wire n_287;
wire n_832;
wire n_353;
wire n_610;
wire n_555;
wire n_389;
wire n_814;
wire n_415;
wire n_830;
wire n_230;
wire n_605;
wire n_461;
wire n_383;
wire n_826;
wire n_669;
wire n_200;
wire n_447;
wire n_176;
wire n_198;
wire n_300;
wire n_222;
wire n_179;
wire n_248;
wire n_517;
wire n_718;
wire n_747;
wire n_667;
wire n_229;
wire n_542;
wire n_644;
wire n_682;
wire n_621;
wire n_305;
wire n_721;
wire n_750;
wire n_532;
wire n_742;
wire n_173;
wire n_535;
wire n_691;
wire n_250;
wire n_372;
wire n_468;
wire n_544;
wire n_504;
wire n_314;
wire n_378;
wire n_413;
wire n_377;
wire n_791;
wire n_183;
wire n_510;
wire n_837;
wire n_836;
wire n_375;
wire n_601;
wire n_338;
wire n_522;
wire n_466;
wire n_704;
wire n_748;
wire n_506;
wire n_763;
wire n_360;
wire n_603;
wire n_235;
wire n_536;
wire n_622;
wire n_191;
wire n_340;
wire n_710;
wire n_387;
wire n_452;
wire n_616;
wire n_658;
wire n_744;
wire n_344;
wire n_581;
wire n_428;
wire n_785;
wire n_761;
wire n_746;
wire n_609;
wire n_765;
wire n_432;
wire n_641;
wire n_822;
wire n_693;
wire n_631;
wire n_174;
wire n_516;
wire n_720;
wire n_525;
wire n_758;
wire n_842;
wire n_611;
wire n_491;
wire n_656;
wire n_772;
wire n_843;
wire n_797;
wire n_666;
wire n_371;
wire n_795;
wire n_770;
wire n_567;
wire n_189;
wire n_738;
wire n_405;
wire n_213;
wire n_538;
wire n_294;
wire n_302;
wire n_499;
wire n_380;
wire n_838;
wire n_705;
wire n_647;
wire n_197;
wire n_343;
wire n_844;
wire n_448;
wire n_494;
wire n_539;
wire n_493;
wire n_397;
wire n_614;
wire n_529;
wire n_445;
wire n_425;
wire n_684;
wire n_454;
wire n_218;
wire n_638;
wire n_234;
wire n_486;
wire n_381;
wire n_236;
wire n_653;
wire n_752;
wire n_172;
wire n_713;
wire n_648;
wire n_657;
wire n_576;
wire n_472;
wire n_270;
wire n_239;
wire n_414;
wire n_563;
wire n_782;
wire n_490;
wire n_803;
wire n_290;
wire n_220;
wire n_809;
wire n_224;
wire n_839;
wire n_734;
wire n_708;
wire n_196;
wire n_402;
wire n_352;
wire n_668;
wire n_478;
wire n_626;
wire n_574;
wire n_779;
wire n_800;
wire n_460;
wire n_417;
wire n_446;
wire n_498;
wire n_662;
wire n_374;
wire n_659;
wire n_709;
wire n_366;
wire n_777;
wire n_407;
wire n_450;
wire n_808;
wire n_272;
wire n_526;
wire n_185;
wire n_712;
wire n_348;
wire n_711;
wire n_579;
wire n_376;
wire n_390;
wire n_473;
wire n_293;
wire n_334;
wire n_559;
wire n_370;
wire n_458;
wire n_232;
wire n_650;
wire n_717;
wire n_330;
wire n_771;
wire n_470;
wire n_475;
wire n_298;
wire n_492;
wire n_281;
wire n_258;
wire n_551;
wire n_699;
wire n_456;
wire n_564;
wire n_265;
wire n_260;
wire n_313;
wire n_451;
wire n_624;
wire n_824;
wire n_279;
wire n_686;
wire n_796;
wire n_252;
wire n_757;
wire n_228;
wire n_565;
wire n_594;
wire n_719;
wire n_356;
wire n_577;
wire n_184;
wire n_552;
wire n_619;
wire n_216;
wire n_455;
wire n_521;
wire n_363;
wire n_572;
wire n_395;
wire n_813;
wire n_592;
wire n_745;
wire n_654;
wire n_323;
wire n_829;
wire n_606;
wire n_393;
wire n_818;
wire n_411;
wire n_503;
wire n_716;
wire n_623;
wire n_599;
wire n_513;
wire n_776;
wire n_321;
wire n_645;
wire n_331;
wire n_227;
wire n_570;
wire n_731;
wire n_406;
wire n_483;
wire n_735;
wire n_204;
wire n_482;
wire n_755;
wire n_474;
wire n_527;
wire n_261;
wire n_608;
wire n_620;
wire n_420;
wire n_683;
wire n_630;
wire n_312;
wire n_394;
wire n_519;
wire n_541;
wire n_512;
wire n_292;
wire n_307;
wire n_469;
wire n_433;
wire n_500;
wire n_792;
wire n_476;
wire n_714;
wire n_291;
wire n_219;
wire n_543;
wire n_357;
wire n_264;
wire n_263;
wire n_589;
wire n_481;
wire n_788;
wire n_819;
wire n_821;
wire n_325;
wire n_767;
wire n_804;
wire n_329;
wire n_464;
wire n_600;
wire n_831;
wire n_802;
wire n_561;
wire n_477;
wire n_549;
wire n_533;
wire n_408;
wire n_806;
wire n_237;
wire n_584;
wire n_244;
wire n_399;
wire n_243;
wire n_548;
wire n_282;
wire n_436;
wire n_833;
wire n_211;
wire n_523;
wire n_175;
wire n_322;
wire n_707;
wire n_345;
wire n_409;
wire n_231;
wire n_354;
wire n_689;
wire n_799;
wire n_505;
wire n_240;
wire n_756;
wire n_319;
wire n_547;
wire n_537;
wire n_273;
wire n_558;
wire n_810;
wire n_635;
wire n_787;
wire n_311;
wire n_403;
wire n_723;
wire n_253;
wire n_634;
wire n_583;
wire n_596;
wire n_546;
wire n_562;
wire n_249;
wire n_201;
wire n_386;
wire n_764;
wire n_556;
wire n_692;
wire n_733;
wire n_754;
wire n_487;
wire n_550;
wire n_241;
wire n_275;
wire n_553;
wire n_652;
wire n_560;
wire n_753;
wire n_642;
wire n_276;
wire n_569;
wire n_441;
wire n_221;
wire n_811;
wire n_444;
wire n_586;
wire n_423;
wire n_737;
wire n_318;
wire n_303;
wire n_511;
wire n_715;
wire n_467;
wire n_306;
wire n_193;
wire n_269;
wire n_359;
wire n_346;
wire n_416;
wire n_530;
wire n_277;
wire n_520;
wire n_418;
wire n_618;
wire n_790;
wire n_582;
wire n_199;
wire n_266;
wire n_296;
wire n_674;
wire n_775;
wire n_571;
wire n_268;
wire n_271;
wire n_404;
wire n_651;
wire n_439;
wire n_217;
wire n_210;
wire n_299;
wire n_518;
wire n_206;
wire n_679;
wire n_453;
wire n_612;
wire n_633;
wire n_665;
wire n_333;
wire n_588;
wire n_215;
wire n_178;
wire n_247;
wire n_225;
wire n_308;
wire n_309;
wire n_759;
wire n_355;
wire n_426;
wire n_317;
wire n_632;
wire n_702;
wire n_431;
wire n_347;
wire n_812;
wire n_459;
wire n_502;
wire n_328;
wire n_672;
wire n_534;
wire n_488;
wire n_429;
wire n_373;
wire n_195;
wire n_285;
wire n_497;
wire n_780;
wire n_773;
wire n_675;
wire n_257;
wire n_730;
wire n_655;
wire n_706;
wire n_786;
wire n_670;
wire n_203;
wire n_286;
wire n_254;
wire n_207;
wire n_834;
wire n_242;
wire n_835;
wire n_690;
wire n_401;
wire n_324;
wire n_743;
wire n_766;
wire n_816;
wire n_335;
wire n_430;
wire n_463;
wire n_545;
wire n_489;
wire n_205;
wire n_604;
wire n_251;
wire n_301;
wire n_274;
wire n_636;
wire n_825;
wire n_728;
wire n_681;
wire n_729;
wire n_774;
wire n_412;
wire n_640;
wire n_660;
wire n_267;
wire n_438;
wire n_339;
wire n_784;
wire n_315;
wire n_434;
wire n_515;
wire n_288;
wire n_427;
wire n_479;
wire n_496;
wire n_598;
wire n_422;
wire n_696;
wire n_722;
wire n_688;
wire n_351;
wire n_437;
wire n_259;
wire n_177;
wire n_540;
wire n_593;
wire n_514;
wire n_646;
wire n_528;
wire n_391;
wire n_457;
wire n_687;
wire n_697;
wire n_364;
wire n_637;
wire n_295;
wire n_385;
wire n_817;
wire n_701;
wire n_629;
wire n_388;
wire n_190;
wire n_262;
wire n_484;
wire n_613;
wire n_736;
wire n_187;
wire n_501;
wire n_841;
wire n_531;
wire n_827;
wire n_508;
wire n_361;
wire n_663;
wire n_379;
wire n_778;
wire n_332;
wire n_336;
wire n_398;
wire n_410;
wire n_566;
wire n_554;
wire n_602;
wire n_194;
wire n_664;
wire n_678;
wire n_192;
wire n_649;
wire n_283;

CKINVDCx16_ASAP7_75t_R g172 ( 
.A(n_102),
.Y(n_172)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_156),
.Y(n_173)
);

CKINVDCx5p33_ASAP7_75t_R g174 ( 
.A(n_103),
.Y(n_174)
);

CKINVDCx5p33_ASAP7_75t_R g175 ( 
.A(n_25),
.Y(n_175)
);

CKINVDCx5p33_ASAP7_75t_R g176 ( 
.A(n_82),
.Y(n_176)
);

CKINVDCx5p33_ASAP7_75t_R g177 ( 
.A(n_136),
.Y(n_177)
);

BUFx3_ASAP7_75t_L g178 ( 
.A(n_167),
.Y(n_178)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

CKINVDCx5p33_ASAP7_75t_R g180 ( 
.A(n_85),
.Y(n_180)
);

CKINVDCx5p33_ASAP7_75t_R g181 ( 
.A(n_71),
.Y(n_181)
);

CKINVDCx5p33_ASAP7_75t_R g182 ( 
.A(n_39),
.Y(n_182)
);

CKINVDCx5p33_ASAP7_75t_R g183 ( 
.A(n_70),
.Y(n_183)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_4),
.Y(n_184)
);

INVx1_ASAP7_75t_L g185 ( 
.A(n_142),
.Y(n_185)
);

CKINVDCx5p33_ASAP7_75t_R g186 ( 
.A(n_131),
.Y(n_186)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_101),
.Y(n_187)
);

CKINVDCx5p33_ASAP7_75t_R g188 ( 
.A(n_72),
.Y(n_188)
);

CKINVDCx5p33_ASAP7_75t_R g189 ( 
.A(n_75),
.Y(n_189)
);

BUFx2_ASAP7_75t_L g190 ( 
.A(n_165),
.Y(n_190)
);

CKINVDCx5p33_ASAP7_75t_R g191 ( 
.A(n_160),
.Y(n_191)
);

CKINVDCx16_ASAP7_75t_R g192 ( 
.A(n_61),
.Y(n_192)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_20),
.Y(n_193)
);

CKINVDCx5p33_ASAP7_75t_R g194 ( 
.A(n_163),
.Y(n_194)
);

CKINVDCx5p33_ASAP7_75t_R g195 ( 
.A(n_169),
.Y(n_195)
);

CKINVDCx5p33_ASAP7_75t_R g196 ( 
.A(n_139),
.Y(n_196)
);

CKINVDCx5p33_ASAP7_75t_R g197 ( 
.A(n_4),
.Y(n_197)
);

CKINVDCx20_ASAP7_75t_R g198 ( 
.A(n_133),
.Y(n_198)
);

CKINVDCx20_ASAP7_75t_R g199 ( 
.A(n_117),
.Y(n_199)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_79),
.Y(n_200)
);

CKINVDCx5p33_ASAP7_75t_R g201 ( 
.A(n_55),
.Y(n_201)
);

CKINVDCx5p33_ASAP7_75t_R g202 ( 
.A(n_86),
.Y(n_202)
);

INVx1_ASAP7_75t_SL g203 ( 
.A(n_96),
.Y(n_203)
);

CKINVDCx5p33_ASAP7_75t_R g204 ( 
.A(n_99),
.Y(n_204)
);

CKINVDCx20_ASAP7_75t_R g205 ( 
.A(n_50),
.Y(n_205)
);

INVx1_ASAP7_75t_L g206 ( 
.A(n_64),
.Y(n_206)
);

CKINVDCx5p33_ASAP7_75t_R g207 ( 
.A(n_6),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_125),
.Y(n_208)
);

CKINVDCx5p33_ASAP7_75t_R g209 ( 
.A(n_42),
.Y(n_209)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_135),
.Y(n_210)
);

CKINVDCx5p33_ASAP7_75t_R g211 ( 
.A(n_143),
.Y(n_211)
);

CKINVDCx5p33_ASAP7_75t_R g212 ( 
.A(n_132),
.Y(n_212)
);

CKINVDCx5p33_ASAP7_75t_R g213 ( 
.A(n_35),
.Y(n_213)
);

CKINVDCx5p33_ASAP7_75t_R g214 ( 
.A(n_106),
.Y(n_214)
);

CKINVDCx5p33_ASAP7_75t_R g215 ( 
.A(n_25),
.Y(n_215)
);

CKINVDCx11_ASAP7_75t_R g216 ( 
.A(n_58),
.Y(n_216)
);

CKINVDCx5p33_ASAP7_75t_R g217 ( 
.A(n_40),
.Y(n_217)
);

CKINVDCx5p33_ASAP7_75t_R g218 ( 
.A(n_118),
.Y(n_218)
);

CKINVDCx5p33_ASAP7_75t_R g219 ( 
.A(n_67),
.Y(n_219)
);

CKINVDCx5p33_ASAP7_75t_R g220 ( 
.A(n_89),
.Y(n_220)
);

CKINVDCx5p33_ASAP7_75t_R g221 ( 
.A(n_93),
.Y(n_221)
);

INVx1_ASAP7_75t_L g222 ( 
.A(n_87),
.Y(n_222)
);

CKINVDCx5p33_ASAP7_75t_R g223 ( 
.A(n_124),
.Y(n_223)
);

CKINVDCx5p33_ASAP7_75t_R g224 ( 
.A(n_68),
.Y(n_224)
);

INVx1_ASAP7_75t_SL g225 ( 
.A(n_59),
.Y(n_225)
);

CKINVDCx5p33_ASAP7_75t_R g226 ( 
.A(n_110),
.Y(n_226)
);

CKINVDCx5p33_ASAP7_75t_R g227 ( 
.A(n_0),
.Y(n_227)
);

INVxp67_ASAP7_75t_L g228 ( 
.A(n_151),
.Y(n_228)
);

CKINVDCx5p33_ASAP7_75t_R g229 ( 
.A(n_121),
.Y(n_229)
);

CKINVDCx5p33_ASAP7_75t_R g230 ( 
.A(n_141),
.Y(n_230)
);

INVx2_ASAP7_75t_L g231 ( 
.A(n_164),
.Y(n_231)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_36),
.Y(n_232)
);

BUFx6f_ASAP7_75t_L g233 ( 
.A(n_38),
.Y(n_233)
);

CKINVDCx5p33_ASAP7_75t_R g234 ( 
.A(n_155),
.Y(n_234)
);

INVx1_ASAP7_75t_SL g235 ( 
.A(n_108),
.Y(n_235)
);

CKINVDCx5p33_ASAP7_75t_R g236 ( 
.A(n_34),
.Y(n_236)
);

BUFx6f_ASAP7_75t_L g237 ( 
.A(n_187),
.Y(n_237)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_193),
.Y(n_238)
);

CKINVDCx20_ASAP7_75t_R g239 ( 
.A(n_184),
.Y(n_239)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_178),
.Y(n_240)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_178),
.Y(n_241)
);

CKINVDCx20_ASAP7_75t_R g242 ( 
.A(n_216),
.Y(n_242)
);

INVxp67_ASAP7_75t_SL g243 ( 
.A(n_190),
.Y(n_243)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_173),
.Y(n_244)
);

INVx1_ASAP7_75t_SL g245 ( 
.A(n_175),
.Y(n_245)
);

INVx1_ASAP7_75t_L g246 ( 
.A(n_179),
.Y(n_246)
);

INVx1_ASAP7_75t_L g247 ( 
.A(n_185),
.Y(n_247)
);

CKINVDCx5p33_ASAP7_75t_R g248 ( 
.A(n_216),
.Y(n_248)
);

CKINVDCx5p33_ASAP7_75t_R g249 ( 
.A(n_197),
.Y(n_249)
);

CKINVDCx5p33_ASAP7_75t_R g250 ( 
.A(n_174),
.Y(n_250)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_200),
.Y(n_251)
);

HB1xp67_ASAP7_75t_L g252 ( 
.A(n_207),
.Y(n_252)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_206),
.Y(n_253)
);

INVx2_ASAP7_75t_L g254 ( 
.A(n_187),
.Y(n_254)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_208),
.Y(n_255)
);

INVxp67_ASAP7_75t_SL g256 ( 
.A(n_228),
.Y(n_256)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_210),
.Y(n_257)
);

CKINVDCx5p33_ASAP7_75t_R g258 ( 
.A(n_215),
.Y(n_258)
);

CKINVDCx5p33_ASAP7_75t_R g259 ( 
.A(n_227),
.Y(n_259)
);

NOR2xp67_ASAP7_75t_L g260 ( 
.A(n_231),
.B(n_0),
.Y(n_260)
);

INVx1_ASAP7_75t_L g261 ( 
.A(n_222),
.Y(n_261)
);

INVx1_ASAP7_75t_L g262 ( 
.A(n_232),
.Y(n_262)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_231),
.Y(n_263)
);

INVxp67_ASAP7_75t_SL g264 ( 
.A(n_187),
.Y(n_264)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_187),
.Y(n_265)
);

CKINVDCx5p33_ASAP7_75t_R g266 ( 
.A(n_198),
.Y(n_266)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_233),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_233),
.Y(n_268)
);

CKINVDCx5p33_ASAP7_75t_R g269 ( 
.A(n_198),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_203),
.B(n_225),
.Y(n_270)
);

INVx2_ASAP7_75t_L g271 ( 
.A(n_233),
.Y(n_271)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_233),
.Y(n_272)
);

CKINVDCx5p33_ASAP7_75t_R g273 ( 
.A(n_199),
.Y(n_273)
);

CKINVDCx5p33_ASAP7_75t_R g274 ( 
.A(n_199),
.Y(n_274)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_176),
.Y(n_275)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_177),
.Y(n_276)
);

INVxp67_ASAP7_75t_L g277 ( 
.A(n_235),
.Y(n_277)
);

NOR2xp33_ASAP7_75t_L g278 ( 
.A(n_172),
.B(n_1),
.Y(n_278)
);

INVxp33_ASAP7_75t_L g279 ( 
.A(n_205),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g280 ( 
.A(n_192),
.Y(n_280)
);

CKINVDCx5p33_ASAP7_75t_R g281 ( 
.A(n_205),
.Y(n_281)
);

INVx1_ASAP7_75t_L g282 ( 
.A(n_180),
.Y(n_282)
);

INVx1_ASAP7_75t_L g283 ( 
.A(n_181),
.Y(n_283)
);

CKINVDCx5p33_ASAP7_75t_R g284 ( 
.A(n_182),
.Y(n_284)
);

AND2x4_ASAP7_75t_L g285 ( 
.A(n_264),
.B(n_236),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_240),
.B(n_241),
.Y(n_286)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_265),
.Y(n_287)
);

INVx1_ASAP7_75t_L g288 ( 
.A(n_267),
.Y(n_288)
);

INVx1_ASAP7_75t_L g289 ( 
.A(n_268),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_SL g290 ( 
.A(n_277),
.B(n_183),
.Y(n_290)
);

OAI21x1_ASAP7_75t_L g291 ( 
.A1(n_254),
.A2(n_188),
.B(n_186),
.Y(n_291)
);

INVx2_ASAP7_75t_L g292 ( 
.A(n_254),
.Y(n_292)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_272),
.Y(n_293)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

INVx1_ASAP7_75t_L g295 ( 
.A(n_271),
.Y(n_295)
);

BUFx8_ASAP7_75t_L g296 ( 
.A(n_275),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_237),
.Y(n_297)
);

INVx2_ASAP7_75t_L g298 ( 
.A(n_237),
.Y(n_298)
);

BUFx6f_ASAP7_75t_L g299 ( 
.A(n_237),
.Y(n_299)
);

HB1xp67_ASAP7_75t_L g300 ( 
.A(n_249),
.Y(n_300)
);

INVx1_ASAP7_75t_L g301 ( 
.A(n_237),
.Y(n_301)
);

INVx2_ASAP7_75t_L g302 ( 
.A(n_237),
.Y(n_302)
);

OAI22xp5_ASAP7_75t_SL g303 ( 
.A1(n_239),
.A2(n_234),
.B1(n_230),
.B2(n_229),
.Y(n_303)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_238),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_L g305 ( 
.A(n_270),
.B(n_189),
.Y(n_305)
);

INVx1_ASAP7_75t_L g306 ( 
.A(n_263),
.Y(n_306)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_244),
.Y(n_307)
);

INVx1_ASAP7_75t_L g308 ( 
.A(n_246),
.Y(n_308)
);

INVx1_ASAP7_75t_L g309 ( 
.A(n_247),
.Y(n_309)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_251),
.Y(n_310)
);

BUFx6f_ASAP7_75t_L g311 ( 
.A(n_253),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g312 ( 
.A(n_256),
.B(n_191),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_L g313 ( 
.A(n_250),
.B(n_276),
.Y(n_313)
);

INVx2_ASAP7_75t_L g314 ( 
.A(n_255),
.Y(n_314)
);

BUFx3_ASAP7_75t_L g315 ( 
.A(n_257),
.Y(n_315)
);

AND2x4_ASAP7_75t_L g316 ( 
.A(n_261),
.B(n_194),
.Y(n_316)
);

NAND2xp5_ASAP7_75t_SL g317 ( 
.A(n_280),
.B(n_195),
.Y(n_317)
);

NAND2xp33_ASAP7_75t_L g318 ( 
.A(n_249),
.B(n_196),
.Y(n_318)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_262),
.Y(n_319)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_260),
.Y(n_320)
);

INVx2_ASAP7_75t_L g321 ( 
.A(n_282),
.Y(n_321)
);

NAND2xp5_ASAP7_75t_L g322 ( 
.A(n_283),
.B(n_226),
.Y(n_322)
);

INVx1_ASAP7_75t_L g323 ( 
.A(n_243),
.Y(n_323)
);

INVx2_ASAP7_75t_L g324 ( 
.A(n_252),
.Y(n_324)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_245),
.Y(n_325)
);

INVx3_ASAP7_75t_L g326 ( 
.A(n_284),
.Y(n_326)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_284),
.Y(n_327)
);

AND2x2_ASAP7_75t_L g328 ( 
.A(n_258),
.B(n_201),
.Y(n_328)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_278),
.Y(n_329)
);

INVx1_ASAP7_75t_L g330 ( 
.A(n_258),
.Y(n_330)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_259),
.B(n_224),
.Y(n_331)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_259),
.Y(n_332)
);

BUFx2_ASAP7_75t_L g333 ( 
.A(n_239),
.Y(n_333)
);

CKINVDCx16_ASAP7_75t_R g334 ( 
.A(n_242),
.Y(n_334)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_248),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_308),
.Y(n_336)
);

OR2x2_ASAP7_75t_L g337 ( 
.A(n_325),
.B(n_266),
.Y(n_337)
);

NAND2xp5_ASAP7_75t_SL g338 ( 
.A(n_325),
.B(n_329),
.Y(n_338)
);

AND2x6_ASAP7_75t_L g339 ( 
.A(n_321),
.B(n_27),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_308),
.Y(n_340)
);

INVx3_ASAP7_75t_L g341 ( 
.A(n_299),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_321),
.B(n_248),
.Y(n_342)
);

NOR2xp33_ASAP7_75t_L g343 ( 
.A(n_305),
.B(n_202),
.Y(n_343)
);

AND2x2_ASAP7_75t_L g344 ( 
.A(n_324),
.B(n_279),
.Y(n_344)
);

INVx1_ASAP7_75t_L g345 ( 
.A(n_309),
.Y(n_345)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_285),
.B(n_204),
.Y(n_346)
);

NAND2xp5_ASAP7_75t_SL g347 ( 
.A(n_329),
.B(n_209),
.Y(n_347)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_309),
.Y(n_348)
);

INVx3_ASAP7_75t_L g349 ( 
.A(n_299),
.Y(n_349)
);

NAND2x1p5_ASAP7_75t_L g350 ( 
.A(n_326),
.B(n_211),
.Y(n_350)
);

INVx1_ASAP7_75t_L g351 ( 
.A(n_310),
.Y(n_351)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_310),
.Y(n_352)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_285),
.B(n_212),
.Y(n_353)
);

NOR3xp33_ASAP7_75t_L g354 ( 
.A(n_330),
.B(n_281),
.C(n_274),
.Y(n_354)
);

BUFx10_ASAP7_75t_L g355 ( 
.A(n_316),
.Y(n_355)
);

INVx3_ASAP7_75t_L g356 ( 
.A(n_299),
.Y(n_356)
);

HB1xp67_ASAP7_75t_L g357 ( 
.A(n_320),
.Y(n_357)
);

BUFx6f_ASAP7_75t_L g358 ( 
.A(n_299),
.Y(n_358)
);

INVx2_ASAP7_75t_L g359 ( 
.A(n_292),
.Y(n_359)
);

BUFx4f_ASAP7_75t_L g360 ( 
.A(n_335),
.Y(n_360)
);

INVx2_ASAP7_75t_L g361 ( 
.A(n_292),
.Y(n_361)
);

INVx2_ASAP7_75t_L g362 ( 
.A(n_294),
.Y(n_362)
);

INVx2_ASAP7_75t_L g363 ( 
.A(n_294),
.Y(n_363)
);

AND2x2_ASAP7_75t_SL g364 ( 
.A(n_318),
.B(n_1),
.Y(n_364)
);

INVx2_ASAP7_75t_L g365 ( 
.A(n_295),
.Y(n_365)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_319),
.Y(n_366)
);

INVx2_ASAP7_75t_SL g367 ( 
.A(n_324),
.Y(n_367)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_319),
.Y(n_368)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_304),
.Y(n_369)
);

INVx1_ASAP7_75t_L g370 ( 
.A(n_304),
.Y(n_370)
);

INVx1_ASAP7_75t_L g371 ( 
.A(n_315),
.Y(n_371)
);

BUFx2_ASAP7_75t_L g372 ( 
.A(n_333),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g373 ( 
.A(n_315),
.Y(n_373)
);

INVx1_ASAP7_75t_L g374 ( 
.A(n_311),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_L g375 ( 
.A(n_285),
.B(n_213),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_L g376 ( 
.A(n_285),
.B(n_214),
.Y(n_376)
);

AND2x4_ASAP7_75t_L g377 ( 
.A(n_286),
.B(n_217),
.Y(n_377)
);

AO22x2_ASAP7_75t_L g378 ( 
.A1(n_330),
.A2(n_2),
.B1(n_3),
.B2(n_5),
.Y(n_378)
);

AND2x2_ASAP7_75t_L g379 ( 
.A(n_312),
.B(n_266),
.Y(n_379)
);

NAND2xp5_ASAP7_75t_L g380 ( 
.A(n_312),
.B(n_218),
.Y(n_380)
);

AND2x2_ASAP7_75t_L g381 ( 
.A(n_323),
.B(n_269),
.Y(n_381)
);

OR2x2_ASAP7_75t_L g382 ( 
.A(n_323),
.B(n_269),
.Y(n_382)
);

AND2x2_ASAP7_75t_L g383 ( 
.A(n_328),
.B(n_273),
.Y(n_383)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_311),
.Y(n_384)
);

INVx2_ASAP7_75t_SL g385 ( 
.A(n_316),
.Y(n_385)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_299),
.Y(n_386)
);

OAI22xp33_ASAP7_75t_SL g387 ( 
.A1(n_313),
.A2(n_223),
.B1(n_221),
.B2(n_220),
.Y(n_387)
);

NAND3xp33_ASAP7_75t_SL g388 ( 
.A(n_332),
.B(n_281),
.C(n_274),
.Y(n_388)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_322),
.B(n_219),
.Y(n_389)
);

INVx2_ASAP7_75t_L g390 ( 
.A(n_295),
.Y(n_390)
);

AND2x4_ASAP7_75t_L g391 ( 
.A(n_286),
.B(n_28),
.Y(n_391)
);

OAI221xp5_ASAP7_75t_L g392 ( 
.A1(n_306),
.A2(n_273),
.B1(n_3),
.B2(n_5),
.C(n_6),
.Y(n_392)
);

NAND2xp33_ASAP7_75t_R g393 ( 
.A(n_332),
.B(n_2),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_311),
.Y(n_394)
);

INVx1_ASAP7_75t_L g395 ( 
.A(n_311),
.Y(n_395)
);

AND3x2_ASAP7_75t_L g396 ( 
.A(n_300),
.B(n_242),
.C(n_8),
.Y(n_396)
);

AND2x4_ASAP7_75t_L g397 ( 
.A(n_316),
.B(n_29),
.Y(n_397)
);

INVx3_ASAP7_75t_L g398 ( 
.A(n_298),
.Y(n_398)
);

NAND3xp33_ASAP7_75t_L g399 ( 
.A(n_327),
.B(n_320),
.C(n_290),
.Y(n_399)
);

INVx2_ASAP7_75t_L g400 ( 
.A(n_298),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_316),
.B(n_30),
.Y(n_401)
);

INVx3_ASAP7_75t_L g402 ( 
.A(n_311),
.Y(n_402)
);

INVx1_ASAP7_75t_L g403 ( 
.A(n_307),
.Y(n_403)
);

NOR2xp33_ASAP7_75t_L g404 ( 
.A(n_327),
.B(n_7),
.Y(n_404)
);

NAND2xp5_ASAP7_75t_L g405 ( 
.A(n_331),
.B(n_31),
.Y(n_405)
);

INVx1_ASAP7_75t_L g406 ( 
.A(n_307),
.Y(n_406)
);

NAND2xp5_ASAP7_75t_SL g407 ( 
.A(n_367),
.B(n_326),
.Y(n_407)
);

NOR2xp67_ASAP7_75t_L g408 ( 
.A(n_388),
.B(n_326),
.Y(n_408)
);

NAND3xp33_ASAP7_75t_SL g409 ( 
.A(n_354),
.B(n_333),
.C(n_335),
.Y(n_409)
);

INVx1_ASAP7_75t_L g410 ( 
.A(n_362),
.Y(n_410)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_362),
.Y(n_411)
);

INVxp67_ASAP7_75t_L g412 ( 
.A(n_344),
.Y(n_412)
);

INVx1_ASAP7_75t_L g413 ( 
.A(n_336),
.Y(n_413)
);

AO22x2_ASAP7_75t_L g414 ( 
.A1(n_378),
.A2(n_382),
.B1(n_338),
.B2(n_379),
.Y(n_414)
);

AO22x2_ASAP7_75t_L g415 ( 
.A1(n_378),
.A2(n_328),
.B1(n_317),
.B2(n_303),
.Y(n_415)
);

INVx2_ASAP7_75t_L g416 ( 
.A(n_359),
.Y(n_416)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_343),
.B(n_296),
.Y(n_417)
);

AO22x2_ASAP7_75t_L g418 ( 
.A1(n_378),
.A2(n_7),
.B1(n_8),
.B2(n_9),
.Y(n_418)
);

INVx1_ASAP7_75t_L g419 ( 
.A(n_340),
.Y(n_419)
);

INVx1_ASAP7_75t_L g420 ( 
.A(n_345),
.Y(n_420)
);

AND2x2_ASAP7_75t_L g421 ( 
.A(n_367),
.B(n_314),
.Y(n_421)
);

NAND2xp33_ASAP7_75t_L g422 ( 
.A(n_385),
.B(n_314),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_385),
.A2(n_296),
.B1(n_291),
.B2(n_306),
.Y(n_423)
);

NAND2xp33_ASAP7_75t_L g424 ( 
.A(n_401),
.B(n_287),
.Y(n_424)
);

INVx4_ASAP7_75t_L g425 ( 
.A(n_373),
.Y(n_425)
);

HB1xp67_ASAP7_75t_L g426 ( 
.A(n_372),
.Y(n_426)
);

NAND2x1p5_ASAP7_75t_L g427 ( 
.A(n_373),
.B(n_291),
.Y(n_427)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_348),
.Y(n_428)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_343),
.B(n_296),
.Y(n_429)
);

AO22x2_ASAP7_75t_L g430 ( 
.A1(n_338),
.A2(n_9),
.B1(n_10),
.B2(n_11),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_351),
.Y(n_431)
);

OAI22xp5_ASAP7_75t_SL g432 ( 
.A1(n_364),
.A2(n_334),
.B1(n_293),
.B2(n_289),
.Y(n_432)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_352),
.Y(n_433)
);

INVx1_ASAP7_75t_L g434 ( 
.A(n_366),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_SL g435 ( 
.A(n_360),
.B(n_296),
.Y(n_435)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_368),
.Y(n_436)
);

INVx1_ASAP7_75t_L g437 ( 
.A(n_369),
.Y(n_437)
);

AND2x4_ASAP7_75t_L g438 ( 
.A(n_371),
.B(n_287),
.Y(n_438)
);

BUFx8_ASAP7_75t_L g439 ( 
.A(n_337),
.Y(n_439)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_370),
.Y(n_440)
);

INVx1_ASAP7_75t_L g441 ( 
.A(n_403),
.Y(n_441)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_347),
.B(n_334),
.Y(n_442)
);

AO22x2_ASAP7_75t_L g443 ( 
.A1(n_347),
.A2(n_10),
.B1(n_11),
.B2(n_12),
.Y(n_443)
);

INVx1_ASAP7_75t_L g444 ( 
.A(n_363),
.Y(n_444)
);

INVx1_ASAP7_75t_L g445 ( 
.A(n_406),
.Y(n_445)
);

AO22x2_ASAP7_75t_L g446 ( 
.A1(n_381),
.A2(n_383),
.B1(n_364),
.B2(n_393),
.Y(n_446)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_342),
.Y(n_447)
);

INVx2_ASAP7_75t_L g448 ( 
.A(n_359),
.Y(n_448)
);

AND2x2_ASAP7_75t_L g449 ( 
.A(n_357),
.B(n_288),
.Y(n_449)
);

INVx1_ASAP7_75t_L g450 ( 
.A(n_363),
.Y(n_450)
);

AO22x2_ASAP7_75t_L g451 ( 
.A1(n_393),
.A2(n_12),
.B1(n_13),
.B2(n_14),
.Y(n_451)
);

INVx1_ASAP7_75t_L g452 ( 
.A(n_365),
.Y(n_452)
);

INVx2_ASAP7_75t_L g453 ( 
.A(n_361),
.Y(n_453)
);

OAI221xp5_ASAP7_75t_L g454 ( 
.A1(n_404),
.A2(n_293),
.B1(n_289),
.B2(n_288),
.C(n_301),
.Y(n_454)
);

INVx2_ASAP7_75t_L g455 ( 
.A(n_361),
.Y(n_455)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_365),
.Y(n_456)
);

INVx1_ASAP7_75t_L g457 ( 
.A(n_390),
.Y(n_457)
);

INVx1_ASAP7_75t_L g458 ( 
.A(n_390),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_357),
.Y(n_459)
);

INVx1_ASAP7_75t_L g460 ( 
.A(n_400),
.Y(n_460)
);

INVx2_ASAP7_75t_L g461 ( 
.A(n_400),
.Y(n_461)
);

NAND2x1p5_ASAP7_75t_L g462 ( 
.A(n_397),
.B(n_302),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g463 ( 
.A1(n_397),
.A2(n_301),
.B1(n_297),
.B2(n_302),
.Y(n_463)
);

INVx2_ASAP7_75t_L g464 ( 
.A(n_398),
.Y(n_464)
);

INVx1_ASAP7_75t_L g465 ( 
.A(n_398),
.Y(n_465)
);

AO22x2_ASAP7_75t_L g466 ( 
.A1(n_399),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_466)
);

AO22x2_ASAP7_75t_L g467 ( 
.A1(n_397),
.A2(n_392),
.B1(n_391),
.B2(n_396),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g468 ( 
.A(n_391),
.B(n_297),
.Y(n_468)
);

AOI22xp5_ASAP7_75t_L g469 ( 
.A1(n_380),
.A2(n_92),
.B1(n_170),
.B2(n_168),
.Y(n_469)
);

AO22x2_ASAP7_75t_L g470 ( 
.A1(n_391),
.A2(n_15),
.B1(n_16),
.B2(n_17),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g471 ( 
.A1(n_346),
.A2(n_91),
.B1(n_166),
.B2(n_162),
.Y(n_471)
);

BUFx3_ASAP7_75t_L g472 ( 
.A(n_360),
.Y(n_472)
);

NOR2xp33_ASAP7_75t_L g473 ( 
.A(n_342),
.B(n_16),
.Y(n_473)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_398),
.Y(n_474)
);

INVx1_ASAP7_75t_L g475 ( 
.A(n_377),
.Y(n_475)
);

INVx2_ASAP7_75t_L g476 ( 
.A(n_341),
.Y(n_476)
);

INVx1_ASAP7_75t_L g477 ( 
.A(n_374),
.Y(n_477)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_384),
.Y(n_478)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_404),
.Y(n_479)
);

INVx1_ASAP7_75t_L g480 ( 
.A(n_377),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g481 ( 
.A(n_447),
.B(n_355),
.Y(n_481)
);

NAND2xp5_ASAP7_75t_SL g482 ( 
.A(n_472),
.B(n_417),
.Y(n_482)
);

NAND2xp33_ASAP7_75t_SL g483 ( 
.A(n_435),
.B(n_353),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g484 ( 
.A(n_429),
.B(n_355),
.Y(n_484)
);

XOR2xp5_ASAP7_75t_L g485 ( 
.A(n_446),
.B(n_387),
.Y(n_485)
);

AND2x2_ASAP7_75t_L g486 ( 
.A(n_412),
.B(n_377),
.Y(n_486)
);

NAND2xp33_ASAP7_75t_SL g487 ( 
.A(n_432),
.B(n_375),
.Y(n_487)
);

AND2x2_ASAP7_75t_L g488 ( 
.A(n_479),
.B(n_350),
.Y(n_488)
);

NAND2xp5_ASAP7_75t_L g489 ( 
.A(n_421),
.B(n_389),
.Y(n_489)
);

NAND2xp5_ASAP7_75t_L g490 ( 
.A(n_413),
.B(n_350),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g491 ( 
.A(n_408),
.B(n_473),
.Y(n_491)
);

NAND2xp5_ASAP7_75t_L g492 ( 
.A(n_419),
.B(n_376),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g493 ( 
.A(n_420),
.B(n_355),
.Y(n_493)
);

NAND2xp33_ASAP7_75t_SL g494 ( 
.A(n_475),
.B(n_405),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_SL g495 ( 
.A(n_425),
.B(n_402),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g496 ( 
.A(n_425),
.B(n_402),
.Y(n_496)
);

NAND2xp5_ASAP7_75t_SL g497 ( 
.A(n_480),
.B(n_394),
.Y(n_497)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_459),
.B(n_395),
.Y(n_498)
);

NAND2xp33_ASAP7_75t_SL g499 ( 
.A(n_449),
.B(n_358),
.Y(n_499)
);

NAND2xp5_ASAP7_75t_SL g500 ( 
.A(n_407),
.B(n_428),
.Y(n_500)
);

NAND2xp33_ASAP7_75t_SL g501 ( 
.A(n_426),
.B(n_358),
.Y(n_501)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_431),
.B(n_349),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_SL g503 ( 
.A(n_433),
.B(n_358),
.Y(n_503)
);

NAND2xp33_ASAP7_75t_SL g504 ( 
.A(n_434),
.B(n_358),
.Y(n_504)
);

NAND2xp5_ASAP7_75t_SL g505 ( 
.A(n_436),
.B(n_437),
.Y(n_505)
);

NAND2xp33_ASAP7_75t_SL g506 ( 
.A(n_440),
.B(n_396),
.Y(n_506)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_438),
.B(n_349),
.Y(n_507)
);

NAND2xp5_ASAP7_75t_SL g508 ( 
.A(n_438),
.B(n_349),
.Y(n_508)
);

AND2x4_ASAP7_75t_L g509 ( 
.A(n_441),
.B(n_339),
.Y(n_509)
);

NAND2xp5_ASAP7_75t_SL g510 ( 
.A(n_442),
.B(n_356),
.Y(n_510)
);

NAND2xp5_ASAP7_75t_SL g511 ( 
.A(n_445),
.B(n_468),
.Y(n_511)
);

NAND2xp5_ASAP7_75t_SL g512 ( 
.A(n_423),
.B(n_356),
.Y(n_512)
);

NAND2xp33_ASAP7_75t_SL g513 ( 
.A(n_446),
.B(n_356),
.Y(n_513)
);

NAND2xp33_ASAP7_75t_SL g514 ( 
.A(n_478),
.B(n_386),
.Y(n_514)
);

NAND2xp5_ASAP7_75t_L g515 ( 
.A(n_410),
.B(n_386),
.Y(n_515)
);

NAND2xp5_ASAP7_75t_SL g516 ( 
.A(n_410),
.B(n_386),
.Y(n_516)
);

NAND2xp5_ASAP7_75t_SL g517 ( 
.A(n_411),
.B(n_341),
.Y(n_517)
);

NAND2xp5_ASAP7_75t_SL g518 ( 
.A(n_411),
.B(n_339),
.Y(n_518)
);

NAND2xp33_ASAP7_75t_SL g519 ( 
.A(n_478),
.B(n_477),
.Y(n_519)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_444),
.B(n_450),
.Y(n_520)
);

NAND2xp5_ASAP7_75t_SL g521 ( 
.A(n_444),
.B(n_339),
.Y(n_521)
);

NAND2xp33_ASAP7_75t_SL g522 ( 
.A(n_477),
.B(n_339),
.Y(n_522)
);

NAND2xp5_ASAP7_75t_SL g523 ( 
.A(n_452),
.B(n_456),
.Y(n_523)
);

NAND2xp5_ASAP7_75t_SL g524 ( 
.A(n_457),
.B(n_339),
.Y(n_524)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_458),
.B(n_17),
.Y(n_525)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_416),
.B(n_18),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_SL g527 ( 
.A(n_463),
.B(n_32),
.Y(n_527)
);

NAND2xp5_ASAP7_75t_SL g528 ( 
.A(n_471),
.B(n_469),
.Y(n_528)
);

NAND2xp33_ASAP7_75t_SL g529 ( 
.A(n_476),
.B(n_18),
.Y(n_529)
);

NAND2xp5_ASAP7_75t_SL g530 ( 
.A(n_448),
.B(n_33),
.Y(n_530)
);

AND2x4_ASAP7_75t_L g531 ( 
.A(n_453),
.B(n_37),
.Y(n_531)
);

NAND2xp33_ASAP7_75t_SL g532 ( 
.A(n_467),
.B(n_19),
.Y(n_532)
);

NAND2xp33_ASAP7_75t_SL g533 ( 
.A(n_467),
.B(n_19),
.Y(n_533)
);

NAND2xp33_ASAP7_75t_SL g534 ( 
.A(n_415),
.B(n_20),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_SL g535 ( 
.A(n_427),
.B(n_41),
.Y(n_535)
);

NAND2xp33_ASAP7_75t_SL g536 ( 
.A(n_415),
.B(n_21),
.Y(n_536)
);

NOR2xp33_ASAP7_75t_SL g537 ( 
.A(n_488),
.B(n_439),
.Y(n_537)
);

AOI21xp5_ASAP7_75t_L g538 ( 
.A1(n_489),
.A2(n_422),
.B(n_462),
.Y(n_538)
);

OAI21x1_ASAP7_75t_L g539 ( 
.A1(n_515),
.A2(n_474),
.B(n_465),
.Y(n_539)
);

NAND2xp5_ASAP7_75t_SL g540 ( 
.A(n_490),
.B(n_439),
.Y(n_540)
);

NOR2xp33_ASAP7_75t_L g541 ( 
.A(n_492),
.B(n_409),
.Y(n_541)
);

OAI21xp5_ASAP7_75t_L g542 ( 
.A1(n_528),
.A2(n_454),
.B(n_460),
.Y(n_542)
);

AOI22xp5_ASAP7_75t_L g543 ( 
.A1(n_487),
.A2(n_414),
.B1(n_424),
.B2(n_470),
.Y(n_543)
);

INVx2_ASAP7_75t_L g544 ( 
.A(n_520),
.Y(n_544)
);

BUFx3_ASAP7_75t_L g545 ( 
.A(n_486),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_L g546 ( 
.A(n_511),
.B(n_414),
.Y(n_546)
);

AO31x2_ASAP7_75t_L g547 ( 
.A1(n_525),
.A2(n_526),
.A3(n_502),
.B(n_461),
.Y(n_547)
);

AOI21x1_ASAP7_75t_L g548 ( 
.A1(n_510),
.A2(n_464),
.B(n_455),
.Y(n_548)
);

OAI22xp5_ASAP7_75t_L g549 ( 
.A1(n_485),
.A2(n_470),
.B1(n_451),
.B2(n_418),
.Y(n_549)
);

INVx2_ASAP7_75t_L g550 ( 
.A(n_523),
.Y(n_550)
);

OAI21x1_ASAP7_75t_L g551 ( 
.A1(n_518),
.A2(n_105),
.B(n_157),
.Y(n_551)
);

OAI21x1_ASAP7_75t_L g552 ( 
.A1(n_521),
.A2(n_104),
.B(n_154),
.Y(n_552)
);

AOI21xp5_ASAP7_75t_L g553 ( 
.A1(n_494),
.A2(n_430),
.B(n_443),
.Y(n_553)
);

INVx1_ASAP7_75t_L g554 ( 
.A(n_505),
.Y(n_554)
);

OAI21x1_ASAP7_75t_L g555 ( 
.A1(n_524),
.A2(n_100),
.B(n_153),
.Y(n_555)
);

NAND3xp33_ASAP7_75t_L g556 ( 
.A(n_534),
.B(n_451),
.C(n_443),
.Y(n_556)
);

CKINVDCx5p33_ASAP7_75t_R g557 ( 
.A(n_506),
.Y(n_557)
);

AND2x4_ASAP7_75t_L g558 ( 
.A(n_481),
.B(n_43),
.Y(n_558)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_516),
.Y(n_559)
);

OAI21x1_ASAP7_75t_L g560 ( 
.A1(n_517),
.A2(n_512),
.B(n_497),
.Y(n_560)
);

INVx1_ASAP7_75t_L g561 ( 
.A(n_507),
.Y(n_561)
);

NAND2xp5_ASAP7_75t_L g562 ( 
.A(n_491),
.B(n_482),
.Y(n_562)
);

INVx2_ASAP7_75t_SL g563 ( 
.A(n_498),
.Y(n_563)
);

INVx1_ASAP7_75t_L g564 ( 
.A(n_508),
.Y(n_564)
);

NOR2xp33_ASAP7_75t_SL g565 ( 
.A(n_531),
.B(n_418),
.Y(n_565)
);

AND2x2_ASAP7_75t_L g566 ( 
.A(n_531),
.B(n_466),
.Y(n_566)
);

AOI21xp5_ASAP7_75t_L g567 ( 
.A1(n_522),
.A2(n_430),
.B(n_466),
.Y(n_567)
);

AND2x4_ASAP7_75t_L g568 ( 
.A(n_500),
.B(n_44),
.Y(n_568)
);

O2A1O1Ixp5_ASAP7_75t_SL g569 ( 
.A1(n_484),
.A2(n_21),
.B(n_22),
.C(n_23),
.Y(n_569)
);

AO21x1_ASAP7_75t_L g570 ( 
.A1(n_536),
.A2(n_22),
.B(n_23),
.Y(n_570)
);

BUFx6f_ASAP7_75t_L g571 ( 
.A(n_531),
.Y(n_571)
);

OAI21x1_ASAP7_75t_L g572 ( 
.A1(n_503),
.A2(n_98),
.B(n_161),
.Y(n_572)
);

AOI21xp5_ASAP7_75t_L g573 ( 
.A1(n_493),
.A2(n_97),
.B(n_158),
.Y(n_573)
);

OAI21xp33_ASAP7_75t_L g574 ( 
.A1(n_527),
.A2(n_24),
.B(n_26),
.Y(n_574)
);

O2A1O1Ixp33_ASAP7_75t_SL g575 ( 
.A1(n_530),
.A2(n_535),
.B(n_495),
.C(n_496),
.Y(n_575)
);

INVx5_ASAP7_75t_L g576 ( 
.A(n_509),
.Y(n_576)
);

NAND2xp5_ASAP7_75t_L g577 ( 
.A(n_513),
.B(n_95),
.Y(n_577)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_519),
.Y(n_578)
);

AOI21xp5_ASAP7_75t_L g579 ( 
.A1(n_499),
.A2(n_483),
.B(n_514),
.Y(n_579)
);

NAND2xp5_ASAP7_75t_L g580 ( 
.A(n_532),
.B(n_94),
.Y(n_580)
);

AND2x2_ASAP7_75t_L g581 ( 
.A(n_509),
.B(n_24),
.Y(n_581)
);

OAI22xp5_ASAP7_75t_SL g582 ( 
.A1(n_549),
.A2(n_533),
.B1(n_509),
.B2(n_529),
.Y(n_582)
);

OAI21x1_ASAP7_75t_L g583 ( 
.A1(n_539),
.A2(n_530),
.B(n_504),
.Y(n_583)
);

OAI21x1_ASAP7_75t_L g584 ( 
.A1(n_548),
.A2(n_501),
.B(n_45),
.Y(n_584)
);

AND2x2_ASAP7_75t_L g585 ( 
.A(n_545),
.B(n_26),
.Y(n_585)
);

OAI21x1_ASAP7_75t_L g586 ( 
.A1(n_560),
.A2(n_46),
.B(n_47),
.Y(n_586)
);

AOI21xp5_ASAP7_75t_L g587 ( 
.A1(n_538),
.A2(n_579),
.B(n_575),
.Y(n_587)
);

INVx2_ASAP7_75t_SL g588 ( 
.A(n_540),
.Y(n_588)
);

OAI21x1_ASAP7_75t_L g589 ( 
.A1(n_579),
.A2(n_48),
.B(n_49),
.Y(n_589)
);

INVx3_ASAP7_75t_L g590 ( 
.A(n_571),
.Y(n_590)
);

OAI21x1_ASAP7_75t_L g591 ( 
.A1(n_551),
.A2(n_51),
.B(n_52),
.Y(n_591)
);

OAI21x1_ASAP7_75t_L g592 ( 
.A1(n_552),
.A2(n_53),
.B(n_54),
.Y(n_592)
);

OAI21x1_ASAP7_75t_L g593 ( 
.A1(n_555),
.A2(n_56),
.B(n_57),
.Y(n_593)
);

OAI21x1_ASAP7_75t_L g594 ( 
.A1(n_572),
.A2(n_60),
.B(n_62),
.Y(n_594)
);

OR2x6_ASAP7_75t_L g595 ( 
.A(n_571),
.B(n_63),
.Y(n_595)
);

CKINVDCx5p33_ASAP7_75t_R g596 ( 
.A(n_557),
.Y(n_596)
);

INVx3_ASAP7_75t_L g597 ( 
.A(n_571),
.Y(n_597)
);

AOI21xp33_ASAP7_75t_R g598 ( 
.A1(n_580),
.A2(n_65),
.B(n_66),
.Y(n_598)
);

OAI21x1_ASAP7_75t_L g599 ( 
.A1(n_542),
.A2(n_69),
.B(n_73),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_L g600 ( 
.A1(n_541),
.A2(n_74),
.B(n_76),
.Y(n_600)
);

OAI21x1_ASAP7_75t_L g601 ( 
.A1(n_542),
.A2(n_77),
.B(n_78),
.Y(n_601)
);

OAI22xp33_ASAP7_75t_L g602 ( 
.A1(n_565),
.A2(n_80),
.B1(n_81),
.B2(n_83),
.Y(n_602)
);

O2A1O1Ixp33_ASAP7_75t_SL g603 ( 
.A1(n_553),
.A2(n_84),
.B(n_88),
.C(n_90),
.Y(n_603)
);

INVx1_ASAP7_75t_L g604 ( 
.A(n_554),
.Y(n_604)
);

INVx2_ASAP7_75t_L g605 ( 
.A(n_544),
.Y(n_605)
);

NAND2xp5_ASAP7_75t_L g606 ( 
.A(n_566),
.B(n_107),
.Y(n_606)
);

NOR2xp67_ASAP7_75t_L g607 ( 
.A(n_563),
.B(n_171),
.Y(n_607)
);

BUFx6f_ASAP7_75t_L g608 ( 
.A(n_576),
.Y(n_608)
);

NOR2x1_ASAP7_75t_SL g609 ( 
.A(n_578),
.B(n_109),
.Y(n_609)
);

BUFx10_ASAP7_75t_L g610 ( 
.A(n_558),
.Y(n_610)
);

INVx2_ASAP7_75t_L g611 ( 
.A(n_559),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_SL g612 ( 
.A(n_537),
.B(n_111),
.Y(n_612)
);

INVx1_ASAP7_75t_L g613 ( 
.A(n_550),
.Y(n_613)
);

NOR2xp33_ASAP7_75t_L g614 ( 
.A(n_549),
.B(n_112),
.Y(n_614)
);

AOI22xp33_ASAP7_75t_L g615 ( 
.A1(n_556),
.A2(n_113),
.B1(n_114),
.B2(n_115),
.Y(n_615)
);

OAI21x1_ASAP7_75t_SL g616 ( 
.A1(n_567),
.A2(n_116),
.B(n_119),
.Y(n_616)
);

INVx1_ASAP7_75t_L g617 ( 
.A(n_561),
.Y(n_617)
);

INVx3_ASAP7_75t_L g618 ( 
.A(n_576),
.Y(n_618)
);

O2A1O1Ixp33_ASAP7_75t_SL g619 ( 
.A1(n_580),
.A2(n_120),
.B(n_122),
.C(n_123),
.Y(n_619)
);

AOI221xp5_ASAP7_75t_L g620 ( 
.A1(n_574),
.A2(n_126),
.B1(n_127),
.B2(n_128),
.C(n_129),
.Y(n_620)
);

NOR2xp33_ASAP7_75t_L g621 ( 
.A(n_562),
.B(n_130),
.Y(n_621)
);

OR2x2_ASAP7_75t_L g622 ( 
.A(n_562),
.B(n_134),
.Y(n_622)
);

NOR2xp33_ASAP7_75t_R g623 ( 
.A(n_537),
.B(n_137),
.Y(n_623)
);

OR2x2_ASAP7_75t_L g624 ( 
.A(n_546),
.B(n_138),
.Y(n_624)
);

OAI21x1_ASAP7_75t_L g625 ( 
.A1(n_587),
.A2(n_573),
.B(n_577),
.Y(n_625)
);

OR2x2_ASAP7_75t_L g626 ( 
.A(n_624),
.B(n_546),
.Y(n_626)
);

INVx3_ASAP7_75t_L g627 ( 
.A(n_608),
.Y(n_627)
);

INVx1_ASAP7_75t_L g628 ( 
.A(n_605),
.Y(n_628)
);

AND2x6_ASAP7_75t_L g629 ( 
.A(n_614),
.B(n_543),
.Y(n_629)
);

AOI322xp5_ASAP7_75t_L g630 ( 
.A1(n_614),
.A2(n_565),
.A3(n_602),
.B1(n_615),
.B2(n_621),
.C1(n_612),
.C2(n_620),
.Y(n_630)
);

INVx2_ASAP7_75t_L g631 ( 
.A(n_605),
.Y(n_631)
);

INVx1_ASAP7_75t_L g632 ( 
.A(n_611),
.Y(n_632)
);

INVx1_ASAP7_75t_L g633 ( 
.A(n_611),
.Y(n_633)
);

INVx2_ASAP7_75t_L g634 ( 
.A(n_604),
.Y(n_634)
);

OAI211xp5_ASAP7_75t_SL g635 ( 
.A1(n_615),
.A2(n_577),
.B(n_564),
.C(n_570),
.Y(n_635)
);

AOI21xp5_ASAP7_75t_L g636 ( 
.A1(n_600),
.A2(n_568),
.B(n_558),
.Y(n_636)
);

INVx1_ASAP7_75t_L g637 ( 
.A(n_617),
.Y(n_637)
);

INVx3_ASAP7_75t_L g638 ( 
.A(n_608),
.Y(n_638)
);

INVx1_ASAP7_75t_L g639 ( 
.A(n_589),
.Y(n_639)
);

INVx1_ASAP7_75t_L g640 ( 
.A(n_589),
.Y(n_640)
);

NAND2xp5_ASAP7_75t_L g641 ( 
.A(n_621),
.B(n_568),
.Y(n_641)
);

BUFx6f_ASAP7_75t_L g642 ( 
.A(n_608),
.Y(n_642)
);

OR2x2_ASAP7_75t_L g643 ( 
.A(n_622),
.B(n_547),
.Y(n_643)
);

AOI21xp5_ASAP7_75t_L g644 ( 
.A1(n_602),
.A2(n_576),
.B(n_581),
.Y(n_644)
);

INVx3_ASAP7_75t_L g645 ( 
.A(n_608),
.Y(n_645)
);

AO21x2_ASAP7_75t_L g646 ( 
.A1(n_583),
.A2(n_547),
.B(n_569),
.Y(n_646)
);

INVx1_ASAP7_75t_L g647 ( 
.A(n_613),
.Y(n_647)
);

BUFx2_ASAP7_75t_L g648 ( 
.A(n_618),
.Y(n_648)
);

INVx1_ASAP7_75t_L g649 ( 
.A(n_586),
.Y(n_649)
);

INVx1_ASAP7_75t_L g650 ( 
.A(n_590),
.Y(n_650)
);

INVx1_ASAP7_75t_L g651 ( 
.A(n_590),
.Y(n_651)
);

INVx2_ASAP7_75t_L g652 ( 
.A(n_618),
.Y(n_652)
);

INVx2_ASAP7_75t_L g653 ( 
.A(n_584),
.Y(n_653)
);

INVx1_ASAP7_75t_L g654 ( 
.A(n_599),
.Y(n_654)
);

NAND2xp5_ASAP7_75t_L g655 ( 
.A(n_588),
.B(n_610),
.Y(n_655)
);

INVx3_ASAP7_75t_L g656 ( 
.A(n_601),
.Y(n_656)
);

INVx2_ASAP7_75t_SL g657 ( 
.A(n_610),
.Y(n_657)
);

INVx2_ASAP7_75t_L g658 ( 
.A(n_592),
.Y(n_658)
);

OAI21x1_ASAP7_75t_L g659 ( 
.A1(n_594),
.A2(n_547),
.B(n_576),
.Y(n_659)
);

INVx1_ASAP7_75t_L g660 ( 
.A(n_597),
.Y(n_660)
);

CKINVDCx6p67_ASAP7_75t_R g661 ( 
.A(n_595),
.Y(n_661)
);

INVx1_ASAP7_75t_L g662 ( 
.A(n_597),
.Y(n_662)
);

INVx1_ASAP7_75t_L g663 ( 
.A(n_606),
.Y(n_663)
);

NOR2xp33_ASAP7_75t_L g664 ( 
.A(n_596),
.B(n_140),
.Y(n_664)
);

INVx1_ASAP7_75t_L g665 ( 
.A(n_603),
.Y(n_665)
);

INVx2_ASAP7_75t_SL g666 ( 
.A(n_595),
.Y(n_666)
);

INVx1_ASAP7_75t_L g667 ( 
.A(n_595),
.Y(n_667)
);

AND2x2_ASAP7_75t_L g668 ( 
.A(n_609),
.B(n_585),
.Y(n_668)
);

BUFx3_ASAP7_75t_L g669 ( 
.A(n_596),
.Y(n_669)
);

INVx1_ASAP7_75t_L g670 ( 
.A(n_582),
.Y(n_670)
);

INVx2_ASAP7_75t_L g671 ( 
.A(n_592),
.Y(n_671)
);

AO21x2_ASAP7_75t_L g672 ( 
.A1(n_616),
.A2(n_144),
.B(n_145),
.Y(n_672)
);

INVx2_ASAP7_75t_SL g673 ( 
.A(n_623),
.Y(n_673)
);

INVx2_ASAP7_75t_L g674 ( 
.A(n_593),
.Y(n_674)
);

INVx1_ASAP7_75t_L g675 ( 
.A(n_603),
.Y(n_675)
);

OAI21xp5_ASAP7_75t_L g676 ( 
.A1(n_607),
.A2(n_146),
.B(n_147),
.Y(n_676)
);

OAI21x1_ASAP7_75t_L g677 ( 
.A1(n_594),
.A2(n_148),
.B(n_149),
.Y(n_677)
);

INVx1_ASAP7_75t_L g678 ( 
.A(n_593),
.Y(n_678)
);

AO21x2_ASAP7_75t_L g679 ( 
.A1(n_619),
.A2(n_150),
.B(n_152),
.Y(n_679)
);

HB1xp67_ASAP7_75t_L g680 ( 
.A(n_623),
.Y(n_680)
);

BUFx3_ASAP7_75t_L g681 ( 
.A(n_669),
.Y(n_681)
);

NAND2xp5_ASAP7_75t_L g682 ( 
.A(n_663),
.B(n_598),
.Y(n_682)
);

NAND2xp33_ASAP7_75t_R g683 ( 
.A(n_668),
.B(n_591),
.Y(n_683)
);

BUFx10_ASAP7_75t_L g684 ( 
.A(n_664),
.Y(n_684)
);

AND2x4_ASAP7_75t_L g685 ( 
.A(n_666),
.B(n_619),
.Y(n_685)
);

INVx1_ASAP7_75t_L g686 ( 
.A(n_637),
.Y(n_686)
);

NOR2xp33_ASAP7_75t_R g687 ( 
.A(n_673),
.B(n_661),
.Y(n_687)
);

NAND2xp33_ASAP7_75t_R g688 ( 
.A(n_668),
.B(n_641),
.Y(n_688)
);

NOR2xp33_ASAP7_75t_R g689 ( 
.A(n_673),
.B(n_661),
.Y(n_689)
);

AND2x4_ASAP7_75t_L g690 ( 
.A(n_666),
.B(n_667),
.Y(n_690)
);

AND2x2_ASAP7_75t_L g691 ( 
.A(n_670),
.B(n_680),
.Y(n_691)
);

NAND2xp33_ASAP7_75t_R g692 ( 
.A(n_655),
.B(n_627),
.Y(n_692)
);

BUFx3_ASAP7_75t_L g693 ( 
.A(n_669),
.Y(n_693)
);

NAND2xp33_ASAP7_75t_R g694 ( 
.A(n_627),
.B(n_645),
.Y(n_694)
);

INVx1_ASAP7_75t_L g695 ( 
.A(n_632),
.Y(n_695)
);

NAND2xp33_ASAP7_75t_R g696 ( 
.A(n_627),
.B(n_645),
.Y(n_696)
);

CKINVDCx8_ASAP7_75t_R g697 ( 
.A(n_642),
.Y(n_697)
);

NOR2xp33_ASAP7_75t_R g698 ( 
.A(n_638),
.B(n_645),
.Y(n_698)
);

XNOR2xp5_ASAP7_75t_L g699 ( 
.A(n_657),
.B(n_636),
.Y(n_699)
);

NOR2xp33_ASAP7_75t_R g700 ( 
.A(n_638),
.B(n_657),
.Y(n_700)
);

NOR2xp33_ASAP7_75t_R g701 ( 
.A(n_638),
.B(n_642),
.Y(n_701)
);

AND2x4_ASAP7_75t_L g702 ( 
.A(n_648),
.B(n_652),
.Y(n_702)
);

XOR2xp5_ASAP7_75t_L g703 ( 
.A(n_626),
.B(n_643),
.Y(n_703)
);

NAND2xp33_ASAP7_75t_R g704 ( 
.A(n_626),
.B(n_648),
.Y(n_704)
);

NAND2xp5_ASAP7_75t_L g705 ( 
.A(n_629),
.B(n_634),
.Y(n_705)
);

AND2x2_ASAP7_75t_L g706 ( 
.A(n_634),
.B(n_628),
.Y(n_706)
);

AND2x4_ASAP7_75t_L g707 ( 
.A(n_652),
.B(n_642),
.Y(n_707)
);

BUFx3_ASAP7_75t_L g708 ( 
.A(n_642),
.Y(n_708)
);

NOR2xp33_ASAP7_75t_SL g709 ( 
.A(n_676),
.B(n_644),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_632),
.Y(n_710)
);

NOR2xp33_ASAP7_75t_R g711 ( 
.A(n_642),
.B(n_660),
.Y(n_711)
);

NAND2xp5_ASAP7_75t_L g712 ( 
.A(n_629),
.B(n_647),
.Y(n_712)
);

BUFx2_ASAP7_75t_L g713 ( 
.A(n_650),
.Y(n_713)
);

INVxp67_ASAP7_75t_L g714 ( 
.A(n_637),
.Y(n_714)
);

NOR2xp33_ASAP7_75t_L g715 ( 
.A(n_651),
.B(n_662),
.Y(n_715)
);

OR2x6_ASAP7_75t_L g716 ( 
.A(n_631),
.B(n_633),
.Y(n_716)
);

AND2x4_ASAP7_75t_L g717 ( 
.A(n_633),
.B(n_631),
.Y(n_717)
);

NAND2xp5_ASAP7_75t_SL g718 ( 
.A(n_630),
.B(n_643),
.Y(n_718)
);

BUFx3_ASAP7_75t_L g719 ( 
.A(n_647),
.Y(n_719)
);

INVx2_ASAP7_75t_L g720 ( 
.A(n_678),
.Y(n_720)
);

AND2x2_ASAP7_75t_L g721 ( 
.A(n_629),
.B(n_672),
.Y(n_721)
);

INVxp67_ASAP7_75t_L g722 ( 
.A(n_629),
.Y(n_722)
);

NAND2xp5_ASAP7_75t_L g723 ( 
.A(n_629),
.B(n_675),
.Y(n_723)
);

BUFx10_ASAP7_75t_L g724 ( 
.A(n_654),
.Y(n_724)
);

HB1xp67_ASAP7_75t_L g725 ( 
.A(n_704),
.Y(n_725)
);

OR2x2_ASAP7_75t_L g726 ( 
.A(n_703),
.B(n_646),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_686),
.Y(n_727)
);

BUFx2_ASAP7_75t_L g728 ( 
.A(n_712),
.Y(n_728)
);

INVxp67_ASAP7_75t_SL g729 ( 
.A(n_719),
.Y(n_729)
);

AND2x2_ASAP7_75t_L g730 ( 
.A(n_721),
.B(n_639),
.Y(n_730)
);

AND2x2_ASAP7_75t_L g731 ( 
.A(n_705),
.B(n_639),
.Y(n_731)
);

INVx1_ASAP7_75t_L g732 ( 
.A(n_720),
.Y(n_732)
);

AND2x2_ASAP7_75t_L g733 ( 
.A(n_695),
.B(n_640),
.Y(n_733)
);

INVxp67_ASAP7_75t_L g734 ( 
.A(n_691),
.Y(n_734)
);

INVx1_ASAP7_75t_L g735 ( 
.A(n_695),
.Y(n_735)
);

AND2x2_ASAP7_75t_L g736 ( 
.A(n_710),
.B(n_640),
.Y(n_736)
);

INVx2_ASAP7_75t_L g737 ( 
.A(n_710),
.Y(n_737)
);

AOI22xp5_ASAP7_75t_L g738 ( 
.A1(n_718),
.A2(n_629),
.B1(n_635),
.B2(n_679),
.Y(n_738)
);

BUFx2_ASAP7_75t_L g739 ( 
.A(n_716),
.Y(n_739)
);

AND2x4_ASAP7_75t_L g740 ( 
.A(n_717),
.B(n_654),
.Y(n_740)
);

INVx1_ASAP7_75t_L g741 ( 
.A(n_714),
.Y(n_741)
);

INVx2_ASAP7_75t_L g742 ( 
.A(n_717),
.Y(n_742)
);

OR2x2_ASAP7_75t_L g743 ( 
.A(n_723),
.B(n_646),
.Y(n_743)
);

INVx1_ASAP7_75t_L g744 ( 
.A(n_724),
.Y(n_744)
);

AOI22xp33_ASAP7_75t_L g745 ( 
.A1(n_709),
.A2(n_672),
.B1(n_679),
.B2(n_665),
.Y(n_745)
);

INVx2_ASAP7_75t_L g746 ( 
.A(n_706),
.Y(n_746)
);

INVx2_ASAP7_75t_SL g747 ( 
.A(n_690),
.Y(n_747)
);

INVx1_ASAP7_75t_L g748 ( 
.A(n_724),
.Y(n_748)
);

AND2x4_ASAP7_75t_SL g749 ( 
.A(n_702),
.B(n_656),
.Y(n_749)
);

AND2x4_ASAP7_75t_L g750 ( 
.A(n_722),
.B(n_656),
.Y(n_750)
);

AND2x2_ASAP7_75t_L g751 ( 
.A(n_716),
.B(n_646),
.Y(n_751)
);

INVx2_ASAP7_75t_L g752 ( 
.A(n_702),
.Y(n_752)
);

INVx1_ASAP7_75t_L g753 ( 
.A(n_682),
.Y(n_753)
);

INVx2_ASAP7_75t_L g754 ( 
.A(n_713),
.Y(n_754)
);

INVx2_ASAP7_75t_L g755 ( 
.A(n_690),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_699),
.B(n_656),
.Y(n_756)
);

AOI221xp5_ASAP7_75t_SL g757 ( 
.A1(n_715),
.A2(n_675),
.B1(n_665),
.B2(n_649),
.C(n_658),
.Y(n_757)
);

AND2x2_ASAP7_75t_L g758 ( 
.A(n_728),
.B(n_707),
.Y(n_758)
);

AND2x2_ASAP7_75t_L g759 ( 
.A(n_728),
.B(n_707),
.Y(n_759)
);

AND2x2_ASAP7_75t_L g760 ( 
.A(n_730),
.B(n_685),
.Y(n_760)
);

AND2x2_ASAP7_75t_L g761 ( 
.A(n_730),
.B(n_685),
.Y(n_761)
);

OR2x2_ASAP7_75t_L g762 ( 
.A(n_726),
.B(n_671),
.Y(n_762)
);

AND2x2_ASAP7_75t_L g763 ( 
.A(n_751),
.B(n_671),
.Y(n_763)
);

AND2x2_ASAP7_75t_L g764 ( 
.A(n_751),
.B(n_674),
.Y(n_764)
);

OR2x2_ASAP7_75t_L g765 ( 
.A(n_726),
.B(n_674),
.Y(n_765)
);

INVx1_ASAP7_75t_L g766 ( 
.A(n_735),
.Y(n_766)
);

INVxp67_ASAP7_75t_SL g767 ( 
.A(n_725),
.Y(n_767)
);

AOI211xp5_ASAP7_75t_L g768 ( 
.A1(n_738),
.A2(n_689),
.B(n_687),
.C(n_693),
.Y(n_768)
);

INVx2_ASAP7_75t_L g769 ( 
.A(n_737),
.Y(n_769)
);

AND2x2_ASAP7_75t_L g770 ( 
.A(n_731),
.B(n_658),
.Y(n_770)
);

AND2x2_ASAP7_75t_L g771 ( 
.A(n_731),
.B(n_681),
.Y(n_771)
);

INVx2_ASAP7_75t_L g772 ( 
.A(n_737),
.Y(n_772)
);

AND2x2_ASAP7_75t_L g773 ( 
.A(n_752),
.B(n_708),
.Y(n_773)
);

BUFx2_ASAP7_75t_L g774 ( 
.A(n_739),
.Y(n_774)
);

INVxp67_ASAP7_75t_L g775 ( 
.A(n_753),
.Y(n_775)
);

AND2x2_ASAP7_75t_L g776 ( 
.A(n_752),
.B(n_679),
.Y(n_776)
);

OR2x2_ASAP7_75t_L g777 ( 
.A(n_762),
.B(n_743),
.Y(n_777)
);

AND2x2_ASAP7_75t_L g778 ( 
.A(n_758),
.B(n_754),
.Y(n_778)
);

AND2x4_ASAP7_75t_L g779 ( 
.A(n_774),
.B(n_748),
.Y(n_779)
);

AND2x2_ASAP7_75t_L g780 ( 
.A(n_758),
.B(n_754),
.Y(n_780)
);

NAND2xp5_ASAP7_75t_L g781 ( 
.A(n_775),
.B(n_753),
.Y(n_781)
);

AND2x2_ASAP7_75t_L g782 ( 
.A(n_759),
.B(n_756),
.Y(n_782)
);

AND2x2_ASAP7_75t_L g783 ( 
.A(n_759),
.B(n_756),
.Y(n_783)
);

OR2x2_ASAP7_75t_L g784 ( 
.A(n_762),
.B(n_743),
.Y(n_784)
);

NAND2xp5_ASAP7_75t_L g785 ( 
.A(n_770),
.B(n_741),
.Y(n_785)
);

OR2x2_ASAP7_75t_L g786 ( 
.A(n_765),
.B(n_742),
.Y(n_786)
);

AND2x2_ASAP7_75t_L g787 ( 
.A(n_771),
.B(n_734),
.Y(n_787)
);

NOR2x1_ASAP7_75t_L g788 ( 
.A(n_781),
.B(n_774),
.Y(n_788)
);

AOI22xp5_ASAP7_75t_L g789 ( 
.A1(n_782),
.A2(n_768),
.B1(n_738),
.B2(n_688),
.Y(n_789)
);

OAI221xp5_ASAP7_75t_L g790 ( 
.A1(n_781),
.A2(n_767),
.B1(n_729),
.B2(n_692),
.C(n_765),
.Y(n_790)
);

NAND2xp5_ASAP7_75t_L g791 ( 
.A(n_785),
.B(n_771),
.Y(n_791)
);

NOR2xp33_ASAP7_75t_R g792 ( 
.A(n_787),
.B(n_684),
.Y(n_792)
);

AO221x2_ASAP7_75t_L g793 ( 
.A1(n_785),
.A2(n_748),
.B1(n_744),
.B2(n_766),
.C(n_741),
.Y(n_793)
);

AO221x2_ASAP7_75t_L g794 ( 
.A1(n_779),
.A2(n_744),
.B1(n_766),
.B2(n_746),
.C(n_755),
.Y(n_794)
);

NOR2xp33_ASAP7_75t_L g795 ( 
.A(n_790),
.B(n_684),
.Y(n_795)
);

AND2x2_ASAP7_75t_L g796 ( 
.A(n_794),
.B(n_783),
.Y(n_796)
);

OR2x2_ASAP7_75t_L g797 ( 
.A(n_791),
.B(n_784),
.Y(n_797)
);

OR2x2_ASAP7_75t_L g798 ( 
.A(n_793),
.B(n_777),
.Y(n_798)
);

NAND2xp5_ASAP7_75t_L g799 ( 
.A(n_795),
.B(n_788),
.Y(n_799)
);

NAND2xp5_ASAP7_75t_L g800 ( 
.A(n_796),
.B(n_789),
.Y(n_800)
);

NAND2xp5_ASAP7_75t_L g801 ( 
.A(n_798),
.B(n_797),
.Y(n_801)
);

INVx1_ASAP7_75t_L g802 ( 
.A(n_797),
.Y(n_802)
);

HB1xp67_ASAP7_75t_L g803 ( 
.A(n_802),
.Y(n_803)
);

NAND2xp5_ASAP7_75t_L g804 ( 
.A(n_800),
.B(n_779),
.Y(n_804)
);

AND2x2_ASAP7_75t_L g805 ( 
.A(n_801),
.B(n_792),
.Y(n_805)
);

INVx2_ASAP7_75t_L g806 ( 
.A(n_803),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_804),
.Y(n_807)
);

INVx1_ASAP7_75t_L g808 ( 
.A(n_805),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_803),
.Y(n_809)
);

INVx1_ASAP7_75t_L g810 ( 
.A(n_806),
.Y(n_810)
);

NAND3xp33_ASAP7_75t_L g811 ( 
.A(n_809),
.B(n_799),
.C(n_745),
.Y(n_811)
);

NAND3xp33_ASAP7_75t_L g812 ( 
.A(n_806),
.B(n_683),
.C(n_739),
.Y(n_812)
);

NOR2x1_ASAP7_75t_SL g813 ( 
.A(n_808),
.B(n_780),
.Y(n_813)
);

NAND4xp25_ASAP7_75t_L g814 ( 
.A(n_807),
.B(n_757),
.C(n_773),
.D(n_694),
.Y(n_814)
);

AOI221xp5_ASAP7_75t_L g815 ( 
.A1(n_811),
.A2(n_773),
.B1(n_763),
.B2(n_764),
.C(n_740),
.Y(n_815)
);

OAI21xp5_ASAP7_75t_L g816 ( 
.A1(n_812),
.A2(n_625),
.B(n_677),
.Y(n_816)
);

OAI22xp5_ASAP7_75t_L g817 ( 
.A1(n_810),
.A2(n_786),
.B1(n_763),
.B2(n_764),
.Y(n_817)
);

NAND2xp5_ASAP7_75t_SL g818 ( 
.A(n_813),
.B(n_700),
.Y(n_818)
);

NAND2xp5_ASAP7_75t_L g819 ( 
.A(n_814),
.B(n_778),
.Y(n_819)
);

INVx1_ASAP7_75t_L g820 ( 
.A(n_819),
.Y(n_820)
);

AND2x2_ASAP7_75t_L g821 ( 
.A(n_818),
.B(n_761),
.Y(n_821)
);

AOI22xp5_ASAP7_75t_L g822 ( 
.A1(n_815),
.A2(n_750),
.B1(n_761),
.B2(n_760),
.Y(n_822)
);

AND2x2_ASAP7_75t_L g823 ( 
.A(n_817),
.B(n_760),
.Y(n_823)
);

AOI22xp5_ASAP7_75t_L g824 ( 
.A1(n_816),
.A2(n_750),
.B1(n_696),
.B2(n_747),
.Y(n_824)
);

NOR2xp33_ASAP7_75t_R g825 ( 
.A(n_820),
.B(n_697),
.Y(n_825)
);

NAND2xp5_ASAP7_75t_SL g826 ( 
.A(n_824),
.B(n_711),
.Y(n_826)
);

NAND3xp33_ASAP7_75t_L g827 ( 
.A(n_821),
.B(n_727),
.C(n_732),
.Y(n_827)
);

NOR2xp33_ASAP7_75t_R g828 ( 
.A(n_823),
.B(n_747),
.Y(n_828)
);

NAND3xp33_ASAP7_75t_L g829 ( 
.A(n_822),
.B(n_727),
.C(n_732),
.Y(n_829)
);

HB1xp67_ASAP7_75t_L g830 ( 
.A(n_825),
.Y(n_830)
);

AOI22xp5_ASAP7_75t_L g831 ( 
.A1(n_826),
.A2(n_750),
.B1(n_770),
.B2(n_740),
.Y(n_831)
);

AND2x2_ASAP7_75t_L g832 ( 
.A(n_828),
.B(n_829),
.Y(n_832)
);

AOI22xp5_ASAP7_75t_L g833 ( 
.A1(n_827),
.A2(n_750),
.B1(n_740),
.B2(n_672),
.Y(n_833)
);

OAI22xp5_ASAP7_75t_SL g834 ( 
.A1(n_830),
.A2(n_701),
.B1(n_755),
.B2(n_698),
.Y(n_834)
);

XNOR2xp5_ASAP7_75t_L g835 ( 
.A(n_832),
.B(n_677),
.Y(n_835)
);

OR4x1_ASAP7_75t_L g836 ( 
.A(n_833),
.B(n_735),
.C(n_649),
.D(n_625),
.Y(n_836)
);

NOR2x1_ASAP7_75t_L g837 ( 
.A(n_831),
.B(n_772),
.Y(n_837)
);

NAND2xp5_ASAP7_75t_SL g838 ( 
.A(n_834),
.B(n_772),
.Y(n_838)
);

OAI21xp5_ASAP7_75t_SL g839 ( 
.A1(n_835),
.A2(n_740),
.B(n_776),
.Y(n_839)
);

AOI22xp33_ASAP7_75t_L g840 ( 
.A1(n_838),
.A2(n_837),
.B1(n_836),
.B2(n_769),
.Y(n_840)
);

AOI22xp33_ASAP7_75t_L g841 ( 
.A1(n_839),
.A2(n_769),
.B1(n_776),
.B2(n_746),
.Y(n_841)
);

XNOR2xp5_ASAP7_75t_L g842 ( 
.A(n_840),
.B(n_749),
.Y(n_842)
);

NAND3xp33_ASAP7_75t_L g843 ( 
.A(n_842),
.B(n_841),
.C(n_733),
.Y(n_843)
);

HB1xp67_ASAP7_75t_L g844 ( 
.A(n_843),
.Y(n_844)
);

OAI221xp5_ASAP7_75t_R g845 ( 
.A1(n_844),
.A2(n_749),
.B1(n_733),
.B2(n_736),
.C(n_659),
.Y(n_845)
);

AOI211xp5_ASAP7_75t_L g846 ( 
.A1(n_845),
.A2(n_736),
.B(n_659),
.C(n_653),
.Y(n_846)
);


endmodule