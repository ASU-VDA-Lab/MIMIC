module real_aes_8458_n_103 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_102, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_101, n_63, n_1, n_53, n_36, n_103);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_102;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_101;
input n_63;
input n_1;
input n_53;
input n_36;
output n_103;
wire n_480;
wire n_113;
wire n_476;
wire n_758;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_750;
wire n_631;
wire n_287;
wire n_357;
wire n_503;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_112;
wire n_364;
wire n_421;
wire n_319;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_242;
wire n_169;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_752;
wire n_448;
wire n_545;
wire n_341;
wire n_556;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_379;
wire n_374;
wire n_453;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_519;
wire n_564;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_478;
wire n_356;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_466;
wire n_559;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_746;
wire n_755;
wire n_153;
wire n_316;
wire n_532;
wire n_284;
wire n_656;
wire n_178;
wire n_409;
wire n_748;
wire n_523;
wire n_298;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_310;
wire n_455;
wire n_725;
wire n_164;
wire n_671;
wire n_231;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_454;
wire n_122;
wire n_443;
wire n_565;
wire n_760;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_745;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_449;
wire n_182;
wire n_417;
wire n_754;
wire n_363;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_527;
wire n_505;
wire n_434;
wire n_502;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_617;
wire n_552;
wire n_402;
wire n_602;
wire n_733;
wire n_171;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_751;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_756;
wire n_288;
wire n_404;
wire n_713;
wire n_598;
wire n_728;
wire n_735;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_749;
wire n_162;
wire n_385;
wire n_275;
wire n_214;
wire n_358;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_498;
wire n_481;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_633;
wire n_679;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_741;
wire n_753;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_140;
wire n_521;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_479;
wire n_338;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_757;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_270;
wire n_507;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_168;
wire n_241;
wire n_175;
wire n_687;
wire n_729;
wire n_646;
wire n_710;
wire n_650;
wire n_105;
wire n_743;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_601;
wire n_500;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
NAND3xp33_ASAP7_75t_SL g106 ( .A(n_0), .B(n_107), .C(n_108), .Y(n_106) );
INVx1_ASAP7_75t_L g447 ( .A(n_0), .Y(n_447) );
INVx1_ASAP7_75t_L g536 ( .A(n_1), .Y(n_536) );
INVx1_ASAP7_75t_L g199 ( .A(n_2), .Y(n_199) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_3), .A2(n_39), .B1(n_161), .B2(n_478), .Y(n_495) );
AOI21xp33_ASAP7_75t_L g140 ( .A1(n_4), .A2(n_141), .B(n_148), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g527 ( .A(n_5), .B(n_134), .Y(n_527) );
AND2x6_ASAP7_75t_L g146 ( .A(n_6), .B(n_147), .Y(n_146) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_7), .A2(n_240), .B(n_241), .Y(n_239) );
NOR2xp33_ASAP7_75t_L g112 ( .A(n_8), .B(n_41), .Y(n_112) );
INVx1_ASAP7_75t_L g158 ( .A(n_9), .Y(n_158) );
NAND2xp5_ASAP7_75t_L g231 ( .A(n_10), .B(n_232), .Y(n_231) );
INVx1_ASAP7_75t_L g139 ( .A(n_11), .Y(n_139) );
NAND2xp5_ASAP7_75t_L g473 ( .A(n_12), .B(n_171), .Y(n_473) );
INVx1_ASAP7_75t_L g246 ( .A(n_13), .Y(n_246) );
INVx1_ASAP7_75t_L g531 ( .A(n_14), .Y(n_531) );
NAND2xp5_ASAP7_75t_L g512 ( .A(n_15), .B(n_135), .Y(n_512) );
AOI22xp5_ASAP7_75t_L g746 ( .A1(n_16), .A2(n_747), .B1(n_748), .B2(n_751), .Y(n_746) );
CKINVDCx20_ASAP7_75t_R g751 ( .A(n_16), .Y(n_751) );
AO32x2_ASAP7_75t_L g493 ( .A1(n_17), .A2(n_134), .A3(n_168), .B1(n_494), .B2(n_498), .Y(n_493) );
NAND2xp5_ASAP7_75t_SL g476 ( .A(n_18), .B(n_161), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g261 ( .A(n_19), .B(n_187), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g538 ( .A(n_20), .B(n_135), .Y(n_538) );
AOI22xp33_ASAP7_75t_L g497 ( .A1(n_21), .A2(n_52), .B1(n_161), .B2(n_478), .Y(n_497) );
NAND2xp5_ASAP7_75t_SL g211 ( .A(n_22), .B(n_141), .Y(n_211) );
AOI22xp33_ASAP7_75t_SL g506 ( .A1(n_23), .A2(n_79), .B1(n_161), .B2(n_171), .Y(n_506) );
NAND2xp5_ASAP7_75t_SL g489 ( .A(n_24), .B(n_161), .Y(n_489) );
NAND2xp5_ASAP7_75t_L g190 ( .A(n_25), .B(n_132), .Y(n_190) );
A2O1A1Ixp33_ASAP7_75t_L g243 ( .A1(n_26), .A2(n_244), .B(n_245), .C(n_247), .Y(n_243) );
OAI22xp5_ASAP7_75t_SL g748 ( .A1(n_27), .A2(n_77), .B1(n_749), .B2(n_750), .Y(n_748) );
CKINVDCx20_ASAP7_75t_R g750 ( .A(n_27), .Y(n_750) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_28), .Y(n_145) );
NAND2xp5_ASAP7_75t_L g550 ( .A(n_29), .B(n_164), .Y(n_550) );
NAND2xp5_ASAP7_75t_L g201 ( .A(n_30), .B(n_156), .Y(n_201) );
INVx1_ASAP7_75t_L g177 ( .A(n_31), .Y(n_177) );
NAND2xp5_ASAP7_75t_L g491 ( .A(n_32), .B(n_164), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g451 ( .A(n_33), .B(n_443), .Y(n_451) );
INVx2_ASAP7_75t_L g144 ( .A(n_34), .Y(n_144) );
NAND2xp5_ASAP7_75t_SL g545 ( .A(n_35), .B(n_161), .Y(n_545) );
NAND2xp5_ASAP7_75t_L g479 ( .A(n_36), .B(n_164), .Y(n_479) );
OAI22xp5_ASAP7_75t_SL g122 ( .A1(n_37), .A2(n_64), .B1(n_123), .B2(n_124), .Y(n_122) );
CKINVDCx20_ASAP7_75t_R g123 ( .A(n_37), .Y(n_123) );
A2O1A1Ixp33_ASAP7_75t_L g212 ( .A1(n_38), .A2(n_146), .B(n_151), .C(n_213), .Y(n_212) );
AOI222xp33_ASAP7_75t_L g453 ( .A1(n_40), .A2(n_454), .B1(n_745), .B2(n_746), .C1(n_752), .C2(n_756), .Y(n_453) );
INVx1_ASAP7_75t_L g175 ( .A(n_42), .Y(n_175) );
NAND2xp5_ASAP7_75t_SL g260 ( .A(n_43), .B(n_156), .Y(n_260) );
NAND2xp5_ASAP7_75t_SL g521 ( .A(n_44), .B(n_161), .Y(n_521) );
OAI321xp33_ASAP7_75t_L g119 ( .A1(n_45), .A2(n_120), .A3(n_443), .B1(n_448), .B2(n_449), .C(n_451), .Y(n_119) );
CKINVDCx16_ASAP7_75t_R g448 ( .A(n_45), .Y(n_448) );
AOI22xp33_ASAP7_75t_L g505 ( .A1(n_46), .A2(n_89), .B1(n_218), .B2(n_478), .Y(n_505) );
NAND2xp5_ASAP7_75t_SL g524 ( .A(n_47), .B(n_161), .Y(n_524) );
NAND2xp5_ASAP7_75t_L g532 ( .A(n_48), .B(n_161), .Y(n_532) );
CKINVDCx16_ASAP7_75t_R g178 ( .A(n_49), .Y(n_178) );
NAND2xp5_ASAP7_75t_L g525 ( .A(n_50), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g234 ( .A(n_51), .B(n_141), .Y(n_234) );
AOI22xp33_ASAP7_75t_SL g516 ( .A1(n_53), .A2(n_62), .B1(n_161), .B2(n_171), .Y(n_516) );
AOI22xp5_ASAP7_75t_L g170 ( .A1(n_54), .A2(n_151), .B1(n_171), .B2(n_173), .Y(n_170) );
CKINVDCx20_ASAP7_75t_R g221 ( .A(n_55), .Y(n_221) );
NAND2xp5_ASAP7_75t_SL g472 ( .A(n_56), .B(n_161), .Y(n_472) );
CKINVDCx16_ASAP7_75t_R g196 ( .A(n_57), .Y(n_196) );
NAND2xp5_ASAP7_75t_SL g549 ( .A(n_58), .B(n_161), .Y(n_549) );
A2O1A1Ixp33_ASAP7_75t_L g154 ( .A1(n_59), .A2(n_155), .B(n_157), .C(n_160), .Y(n_154) );
CKINVDCx20_ASAP7_75t_R g264 ( .A(n_60), .Y(n_264) );
INVx1_ASAP7_75t_L g149 ( .A(n_61), .Y(n_149) );
INVx1_ASAP7_75t_L g147 ( .A(n_63), .Y(n_147) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_64), .Y(n_124) );
AOI22xp33_ASAP7_75t_L g103 ( .A1(n_65), .A2(n_104), .B1(n_113), .B2(n_760), .Y(n_103) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_66), .B(n_161), .Y(n_537) );
INVx1_ASAP7_75t_L g138 ( .A(n_67), .Y(n_138) );
CKINVDCx20_ASAP7_75t_R g118 ( .A(n_68), .Y(n_118) );
AO32x2_ASAP7_75t_L g503 ( .A1(n_69), .A2(n_134), .A3(n_226), .B1(n_498), .B2(n_504), .Y(n_503) );
INVx1_ASAP7_75t_L g548 ( .A(n_70), .Y(n_548) );
INVx1_ASAP7_75t_L g486 ( .A(n_71), .Y(n_486) );
A2O1A1Ixp33_ASAP7_75t_SL g186 ( .A1(n_72), .A2(n_160), .B(n_187), .C(n_188), .Y(n_186) );
INVxp67_ASAP7_75t_L g189 ( .A(n_73), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_74), .B(n_171), .Y(n_487) );
INVx1_ASAP7_75t_L g110 ( .A(n_75), .Y(n_110) );
CKINVDCx20_ASAP7_75t_R g181 ( .A(n_76), .Y(n_181) );
CKINVDCx20_ASAP7_75t_R g749 ( .A(n_77), .Y(n_749) );
INVx1_ASAP7_75t_L g257 ( .A(n_78), .Y(n_257) );
A2O1A1Ixp33_ASAP7_75t_L g258 ( .A1(n_80), .A2(n_146), .B(n_151), .C(n_259), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_81), .B(n_478), .Y(n_477) );
NAND2xp5_ASAP7_75t_SL g490 ( .A(n_82), .B(n_171), .Y(n_490) );
NAND2xp5_ASAP7_75t_SL g214 ( .A(n_83), .B(n_200), .Y(n_214) );
INVx2_ASAP7_75t_L g136 ( .A(n_84), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_85), .B(n_187), .Y(n_215) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_86), .B(n_171), .Y(n_522) );
A2O1A1Ixp33_ASAP7_75t_L g197 ( .A1(n_87), .A2(n_146), .B(n_151), .C(n_198), .Y(n_197) );
INVx2_ASAP7_75t_L g107 ( .A(n_88), .Y(n_107) );
OR2x2_ASAP7_75t_L g444 ( .A(n_88), .B(n_445), .Y(n_444) );
OR2x2_ASAP7_75t_L g459 ( .A(n_88), .B(n_446), .Y(n_459) );
AOI22xp33_ASAP7_75t_L g515 ( .A1(n_90), .A2(n_102), .B1(n_171), .B2(n_172), .Y(n_515) );
NAND2xp5_ASAP7_75t_L g163 ( .A(n_91), .B(n_164), .Y(n_163) );
CKINVDCx20_ASAP7_75t_R g204 ( .A(n_92), .Y(n_204) );
A2O1A1Ixp33_ASAP7_75t_L g228 ( .A1(n_93), .A2(n_146), .B(n_151), .C(n_229), .Y(n_228) );
CKINVDCx20_ASAP7_75t_R g236 ( .A(n_94), .Y(n_236) );
INVx1_ASAP7_75t_L g185 ( .A(n_95), .Y(n_185) );
CKINVDCx16_ASAP7_75t_R g242 ( .A(n_96), .Y(n_242) );
NAND2xp5_ASAP7_75t_SL g230 ( .A(n_97), .B(n_200), .Y(n_230) );
NAND2xp5_ASAP7_75t_L g546 ( .A(n_98), .B(n_171), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_99), .B(n_134), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g109 ( .A(n_100), .B(n_110), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g183 ( .A1(n_101), .A2(n_141), .B(n_184), .Y(n_183) );
INVx1_ASAP7_75t_SL g104 ( .A(n_105), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g761 ( .A(n_105), .Y(n_761) );
OR2x2_ASAP7_75t_SL g105 ( .A(n_106), .B(n_111), .Y(n_105) );
OR2x2_ASAP7_75t_L g461 ( .A(n_107), .B(n_446), .Y(n_461) );
NOR2x2_ASAP7_75t_L g758 ( .A(n_107), .B(n_445), .Y(n_758) );
INVx1_ASAP7_75t_SL g108 ( .A(n_109), .Y(n_108) );
INVxp67_ASAP7_75t_L g111 ( .A(n_112), .Y(n_111) );
AND2x2_ASAP7_75t_L g446 ( .A(n_112), .B(n_447), .Y(n_446) );
AO21x1_ASAP7_75t_L g113 ( .A1(n_114), .A2(n_119), .B(n_452), .Y(n_113) );
INVx1_ASAP7_75t_SL g114 ( .A(n_115), .Y(n_114) );
BUFx2_ASAP7_75t_L g115 ( .A(n_116), .Y(n_115) );
BUFx2_ASAP7_75t_L g116 ( .A(n_117), .Y(n_116) );
INVx1_ASAP7_75t_SL g759 ( .A(n_117), .Y(n_759) );
INVx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
NAND2xp5_ASAP7_75t_SL g449 ( .A(n_120), .B(n_450), .Y(n_449) );
OAI22xp5_ASAP7_75t_L g120 ( .A1(n_121), .A2(n_122), .B1(n_125), .B2(n_442), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_122), .Y(n_121) );
AOI22xp5_ASAP7_75t_L g753 ( .A1(n_125), .A2(n_463), .B1(n_754), .B2(n_755), .Y(n_753) );
INVx1_ASAP7_75t_L g125 ( .A(n_126), .Y(n_125) );
BUFx2_ASAP7_75t_L g442 ( .A(n_126), .Y(n_442) );
AND3x1_ASAP7_75t_L g126 ( .A(n_127), .B(n_364), .C(n_409), .Y(n_126) );
NOR4xp25_ASAP7_75t_L g127 ( .A(n_128), .B(n_287), .C(n_328), .D(n_345), .Y(n_127) );
A2O1A1Ixp33_ASAP7_75t_L g128 ( .A1(n_129), .A2(n_191), .B(n_207), .C(n_249), .Y(n_128) );
OR2x2_ASAP7_75t_L g129 ( .A(n_130), .B(n_165), .Y(n_129) );
NAND2xp5_ASAP7_75t_L g191 ( .A(n_130), .B(n_192), .Y(n_191) );
NOR4xp25_ASAP7_75t_L g311 ( .A(n_130), .B(n_305), .C(n_312), .D(n_318), .Y(n_311) );
AND2x2_ASAP7_75t_L g384 ( .A(n_130), .B(n_273), .Y(n_384) );
AND2x2_ASAP7_75t_L g403 ( .A(n_130), .B(n_349), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g412 ( .A(n_130), .B(n_398), .Y(n_412) );
AND2x2_ASAP7_75t_L g425 ( .A(n_130), .B(n_206), .Y(n_425) );
INVx2_ASAP7_75t_L g130 ( .A(n_131), .Y(n_130) );
INVx1_ASAP7_75t_SL g270 ( .A(n_131), .Y(n_270) );
AND2x2_ASAP7_75t_L g277 ( .A(n_131), .B(n_278), .Y(n_277) );
OR2x2_ASAP7_75t_L g327 ( .A(n_131), .B(n_166), .Y(n_327) );
AND2x2_ASAP7_75t_SL g338 ( .A(n_131), .B(n_273), .Y(n_338) );
NAND2xp5_ASAP7_75t_L g342 ( .A(n_131), .B(n_166), .Y(n_342) );
AND2x2_ASAP7_75t_L g351 ( .A(n_131), .B(n_276), .Y(n_351) );
BUFx2_ASAP7_75t_L g374 ( .A(n_131), .Y(n_374) );
AND2x2_ASAP7_75t_L g378 ( .A(n_131), .B(n_182), .Y(n_378) );
OA21x2_ASAP7_75t_L g131 ( .A1(n_132), .A2(n_140), .B(n_163), .Y(n_131) );
INVx3_ASAP7_75t_L g132 ( .A(n_133), .Y(n_132) );
NOR2xp33_ASAP7_75t_SL g220 ( .A(n_133), .B(n_221), .Y(n_220) );
NAND3xp33_ASAP7_75t_L g513 ( .A(n_133), .B(n_498), .C(n_514), .Y(n_513) );
AO21x1_ASAP7_75t_L g551 ( .A1(n_133), .A2(n_514), .B(n_552), .Y(n_551) );
INVx4_ASAP7_75t_L g133 ( .A(n_134), .Y(n_133) );
OA21x2_ASAP7_75t_L g182 ( .A1(n_134), .A2(n_183), .B(n_190), .Y(n_182) );
OA21x2_ASAP7_75t_L g518 ( .A1(n_134), .A2(n_519), .B(n_527), .Y(n_518) );
BUFx6f_ASAP7_75t_L g134 ( .A(n_135), .Y(n_134) );
INVx1_ASAP7_75t_L g168 ( .A(n_135), .Y(n_168) );
AND2x2_ASAP7_75t_L g135 ( .A(n_136), .B(n_137), .Y(n_135) );
AND2x2_ASAP7_75t_SL g164 ( .A(n_136), .B(n_137), .Y(n_164) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_138), .B(n_139), .Y(n_137) );
BUFx2_ASAP7_75t_L g240 ( .A(n_141), .Y(n_240) );
AND2x4_ASAP7_75t_L g141 ( .A(n_142), .B(n_146), .Y(n_141) );
NAND2x1p5_ASAP7_75t_L g179 ( .A(n_142), .B(n_146), .Y(n_179) );
AND2x2_ASAP7_75t_L g142 ( .A(n_143), .B(n_145), .Y(n_142) );
INVx1_ASAP7_75t_L g526 ( .A(n_143), .Y(n_526) );
INVx1_ASAP7_75t_L g143 ( .A(n_144), .Y(n_143) );
INVx2_ASAP7_75t_L g152 ( .A(n_144), .Y(n_152) );
INVx1_ASAP7_75t_L g172 ( .A(n_144), .Y(n_172) );
INVx1_ASAP7_75t_L g153 ( .A(n_145), .Y(n_153) );
BUFx6f_ASAP7_75t_L g156 ( .A(n_145), .Y(n_156) );
INVx3_ASAP7_75t_L g159 ( .A(n_145), .Y(n_159) );
BUFx6f_ASAP7_75t_L g174 ( .A(n_145), .Y(n_174) );
INVx1_ASAP7_75t_L g187 ( .A(n_145), .Y(n_187) );
INVx4_ASAP7_75t_SL g162 ( .A(n_146), .Y(n_162) );
OAI21xp5_ASAP7_75t_L g470 ( .A1(n_146), .A2(n_471), .B(n_475), .Y(n_470) );
OAI21xp5_ASAP7_75t_L g484 ( .A1(n_146), .A2(n_485), .B(n_488), .Y(n_484) );
BUFx3_ASAP7_75t_L g498 ( .A(n_146), .Y(n_498) );
OAI21xp5_ASAP7_75t_L g519 ( .A1(n_146), .A2(n_520), .B(n_523), .Y(n_519) );
OAI21xp5_ASAP7_75t_L g529 ( .A1(n_146), .A2(n_530), .B(n_534), .Y(n_529) );
O2A1O1Ixp33_ASAP7_75t_L g148 ( .A1(n_149), .A2(n_150), .B(n_154), .C(n_162), .Y(n_148) );
O2A1O1Ixp33_ASAP7_75t_L g184 ( .A1(n_150), .A2(n_162), .B(n_185), .C(n_186), .Y(n_184) );
O2A1O1Ixp33_ASAP7_75t_L g241 ( .A1(n_150), .A2(n_162), .B(n_242), .C(n_243), .Y(n_241) );
INVx5_ASAP7_75t_L g150 ( .A(n_151), .Y(n_150) );
AND2x6_ASAP7_75t_L g151 ( .A(n_152), .B(n_153), .Y(n_151) );
BUFx6f_ASAP7_75t_L g161 ( .A(n_152), .Y(n_161) );
BUFx3_ASAP7_75t_L g218 ( .A(n_152), .Y(n_218) );
INVx1_ASAP7_75t_L g478 ( .A(n_152), .Y(n_478) );
AOI21xp5_ASAP7_75t_L g475 ( .A1(n_155), .A2(n_476), .B(n_477), .Y(n_475) );
O2A1O1Ixp5_ASAP7_75t_L g547 ( .A1(n_155), .A2(n_535), .B(n_548), .C(n_549), .Y(n_547) );
INVx2_ASAP7_75t_L g155 ( .A(n_156), .Y(n_155) );
INVx4_ASAP7_75t_L g232 ( .A(n_156), .Y(n_232) );
OAI22xp5_ASAP7_75t_L g494 ( .A1(n_156), .A2(n_495), .B1(n_496), .B2(n_497), .Y(n_494) );
OAI22xp5_ASAP7_75t_SL g504 ( .A1(n_156), .A2(n_159), .B1(n_505), .B2(n_506), .Y(n_504) );
OAI22xp5_ASAP7_75t_L g514 ( .A1(n_156), .A2(n_496), .B1(n_515), .B2(n_516), .Y(n_514) );
NOR2xp33_ASAP7_75t_L g157 ( .A(n_158), .B(n_159), .Y(n_157) );
NOR2xp33_ASAP7_75t_L g188 ( .A(n_159), .B(n_189), .Y(n_188) );
INVx5_ASAP7_75t_L g200 ( .A(n_159), .Y(n_200) );
O2A1O1Ixp5_ASAP7_75t_SL g485 ( .A1(n_160), .A2(n_200), .B(n_486), .C(n_487), .Y(n_485) );
INVx3_ASAP7_75t_L g160 ( .A(n_161), .Y(n_160) );
HB1xp67_ASAP7_75t_L g233 ( .A(n_161), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g169 ( .A1(n_162), .A2(n_170), .B1(n_178), .B2(n_179), .Y(n_169) );
INVx1_ASAP7_75t_L g205 ( .A(n_164), .Y(n_205) );
INVx2_ASAP7_75t_L g226 ( .A(n_164), .Y(n_226) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_164), .A2(n_239), .B(n_248), .Y(n_238) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_164), .A2(n_470), .B(n_479), .Y(n_469) );
OA21x2_ASAP7_75t_L g483 ( .A1(n_164), .A2(n_484), .B(n_491), .Y(n_483) );
OR2x2_ASAP7_75t_L g165 ( .A(n_166), .B(n_182), .Y(n_165) );
AND2x2_ASAP7_75t_L g206 ( .A(n_166), .B(n_182), .Y(n_206) );
BUFx2_ASAP7_75t_L g280 ( .A(n_166), .Y(n_280) );
AOI22xp33_ASAP7_75t_L g312 ( .A1(n_166), .A2(n_313), .B1(n_315), .B2(n_316), .Y(n_312) );
OR2x2_ASAP7_75t_L g334 ( .A(n_166), .B(n_194), .Y(n_334) );
AND2x2_ASAP7_75t_L g398 ( .A(n_166), .B(n_276), .Y(n_398) );
INVx3_ASAP7_75t_L g166 ( .A(n_167), .Y(n_166) );
AND2x2_ASAP7_75t_L g266 ( .A(n_167), .B(n_194), .Y(n_266) );
AND2x2_ASAP7_75t_L g273 ( .A(n_167), .B(n_182), .Y(n_273) );
HB1xp67_ASAP7_75t_L g315 ( .A(n_167), .Y(n_315) );
OR2x2_ASAP7_75t_L g350 ( .A(n_167), .B(n_193), .Y(n_350) );
AO21x2_ASAP7_75t_L g167 ( .A1(n_168), .A2(n_169), .B(n_180), .Y(n_167) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_168), .B(n_181), .Y(n_180) );
AO21x2_ASAP7_75t_L g194 ( .A1(n_168), .A2(n_195), .B(n_203), .Y(n_194) );
INVx2_ASAP7_75t_L g219 ( .A(n_168), .Y(n_219) );
INVx2_ASAP7_75t_L g202 ( .A(n_171), .Y(n_202) );
INVx3_ASAP7_75t_L g171 ( .A(n_172), .Y(n_171) );
OAI22xp5_ASAP7_75t_SL g173 ( .A1(n_174), .A2(n_175), .B1(n_176), .B2(n_177), .Y(n_173) );
INVx2_ASAP7_75t_L g176 ( .A(n_174), .Y(n_176) );
INVx4_ASAP7_75t_L g244 ( .A(n_174), .Y(n_244) );
OAI21xp5_ASAP7_75t_L g195 ( .A1(n_179), .A2(n_196), .B(n_197), .Y(n_195) );
OAI21xp5_ASAP7_75t_L g256 ( .A1(n_179), .A2(n_257), .B(n_258), .Y(n_256) );
INVx1_ASAP7_75t_L g269 ( .A(n_182), .Y(n_269) );
INVx3_ASAP7_75t_L g278 ( .A(n_182), .Y(n_278) );
BUFx2_ASAP7_75t_L g302 ( .A(n_182), .Y(n_302) );
AND2x2_ASAP7_75t_L g335 ( .A(n_182), .B(n_270), .Y(n_335) );
INVx1_ASAP7_75t_L g474 ( .A(n_187), .Y(n_474) );
OAI22xp5_ASAP7_75t_L g420 ( .A1(n_191), .A2(n_421), .B1(n_422), .B2(n_423), .Y(n_420) );
AND2x2_ASAP7_75t_L g192 ( .A(n_193), .B(n_206), .Y(n_192) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_193), .B(n_278), .Y(n_282) );
INVx1_ASAP7_75t_L g310 ( .A(n_193), .Y(n_310) );
INVx3_ASAP7_75t_L g193 ( .A(n_194), .Y(n_193) );
INVx3_ASAP7_75t_L g276 ( .A(n_194), .Y(n_276) );
O2A1O1Ixp33_ASAP7_75t_L g198 ( .A1(n_199), .A2(n_200), .B(n_201), .C(n_202), .Y(n_198) );
INVx2_ASAP7_75t_L g496 ( .A(n_200), .Y(n_496) );
AOI21xp5_ASAP7_75t_L g520 ( .A1(n_200), .A2(n_521), .B(n_522), .Y(n_520) );
AOI21xp5_ASAP7_75t_L g544 ( .A1(n_200), .A2(n_545), .B(n_546), .Y(n_544) );
O2A1O1Ixp33_ASAP7_75t_L g530 ( .A1(n_202), .A2(n_531), .B(n_532), .C(n_533), .Y(n_530) );
NOR2xp33_ASAP7_75t_L g203 ( .A(n_204), .B(n_205), .Y(n_203) );
NOR2xp33_ASAP7_75t_L g235 ( .A(n_205), .B(n_236), .Y(n_235) );
NOR2xp33_ASAP7_75t_L g263 ( .A(n_205), .B(n_264), .Y(n_263) );
INVx1_ASAP7_75t_L g288 ( .A(n_206), .Y(n_288) );
NAND2x1_ASAP7_75t_SL g207 ( .A(n_208), .B(n_222), .Y(n_207) );
AND2x2_ASAP7_75t_L g286 ( .A(n_208), .B(n_237), .Y(n_286) );
HB1xp67_ASAP7_75t_L g360 ( .A(n_208), .Y(n_360) );
AND2x2_ASAP7_75t_L g387 ( .A(n_208), .B(n_307), .Y(n_387) );
AND2x2_ASAP7_75t_L g395 ( .A(n_208), .B(n_357), .Y(n_395) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_208), .B(n_252), .Y(n_422) );
INVx3_ASAP7_75t_L g208 ( .A(n_209), .Y(n_208) );
AND2x2_ASAP7_75t_L g253 ( .A(n_209), .B(n_254), .Y(n_253) );
AND2x2_ASAP7_75t_L g271 ( .A(n_209), .B(n_272), .Y(n_271) );
INVx2_ASAP7_75t_L g292 ( .A(n_209), .Y(n_292) );
INVx1_ASAP7_75t_L g298 ( .A(n_209), .Y(n_298) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_209), .B(n_314), .Y(n_313) );
AND2x2_ASAP7_75t_L g331 ( .A(n_209), .B(n_255), .Y(n_331) );
OR2x2_ASAP7_75t_L g369 ( .A(n_209), .B(n_324), .Y(n_369) );
AOI32xp33_ASAP7_75t_L g381 ( .A1(n_209), .A2(n_382), .A3(n_385), .B1(n_386), .B2(n_387), .Y(n_381) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_209), .B(n_357), .Y(n_421) );
NOR2xp33_ASAP7_75t_L g432 ( .A(n_209), .B(n_317), .Y(n_432) );
OR2x6_ASAP7_75t_L g209 ( .A(n_210), .B(n_220), .Y(n_209) );
AOI21xp5_ASAP7_75t_SL g210 ( .A1(n_211), .A2(n_212), .B(n_219), .Y(n_210) );
AOI21xp5_ASAP7_75t_L g213 ( .A1(n_214), .A2(n_215), .B(n_216), .Y(n_213) );
AOI21xp5_ASAP7_75t_L g259 ( .A1(n_216), .A2(n_260), .B(n_261), .Y(n_259) );
INVx2_ASAP7_75t_L g216 ( .A(n_217), .Y(n_216) );
INVx2_ASAP7_75t_L g217 ( .A(n_218), .Y(n_217) );
INVx1_ASAP7_75t_L g247 ( .A(n_218), .Y(n_247) );
INVx1_ASAP7_75t_L g262 ( .A(n_219), .Y(n_262) );
OA21x2_ASAP7_75t_L g528 ( .A1(n_219), .A2(n_529), .B(n_538), .Y(n_528) );
OA21x2_ASAP7_75t_L g542 ( .A1(n_219), .A2(n_543), .B(n_550), .Y(n_542) );
INVx2_ASAP7_75t_L g222 ( .A(n_223), .Y(n_222) );
OR2x2_ASAP7_75t_L g343 ( .A(n_223), .B(n_344), .Y(n_343) );
OR2x2_ASAP7_75t_L g223 ( .A(n_224), .B(n_237), .Y(n_223) );
INVx1_ASAP7_75t_L g305 ( .A(n_224), .Y(n_305) );
AND2x2_ASAP7_75t_L g307 ( .A(n_224), .B(n_308), .Y(n_307) );
NAND2xp5_ASAP7_75t_L g324 ( .A(n_224), .B(n_254), .Y(n_324) );
AND2x2_ASAP7_75t_L g357 ( .A(n_224), .B(n_333), .Y(n_357) );
AND2x2_ASAP7_75t_L g394 ( .A(n_224), .B(n_255), .Y(n_394) );
INVx2_ASAP7_75t_L g224 ( .A(n_225), .Y(n_224) );
INVx1_ASAP7_75t_L g252 ( .A(n_225), .Y(n_252) );
NAND2xp5_ASAP7_75t_L g284 ( .A(n_225), .B(n_254), .Y(n_284) );
AND2x2_ASAP7_75t_L g291 ( .A(n_225), .B(n_292), .Y(n_291) );
AND2x2_ASAP7_75t_L g332 ( .A(n_225), .B(n_333), .Y(n_332) );
AO21x2_ASAP7_75t_L g225 ( .A1(n_226), .A2(n_227), .B(n_235), .Y(n_225) );
NAND2xp5_ASAP7_75t_L g227 ( .A(n_228), .B(n_234), .Y(n_227) );
AOI21xp5_ASAP7_75t_L g229 ( .A1(n_230), .A2(n_231), .B(n_233), .Y(n_229) );
INVx2_ASAP7_75t_L g308 ( .A(n_237), .Y(n_308) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_237), .B(n_254), .Y(n_317) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_237), .B(n_299), .Y(n_380) );
INVx1_ASAP7_75t_L g402 ( .A(n_237), .Y(n_402) );
INVx1_ASAP7_75t_L g419 ( .A(n_237), .Y(n_419) );
INVx2_ASAP7_75t_L g237 ( .A(n_238), .Y(n_237) );
AND2x2_ASAP7_75t_L g272 ( .A(n_238), .B(n_254), .Y(n_272) );
AND2x2_ASAP7_75t_L g294 ( .A(n_238), .B(n_255), .Y(n_294) );
INVx1_ASAP7_75t_L g333 ( .A(n_238), .Y(n_333) );
NOR2xp33_ASAP7_75t_L g245 ( .A(n_244), .B(n_246), .Y(n_245) );
AOI21xp5_ASAP7_75t_L g488 ( .A1(n_244), .A2(n_489), .B(n_490), .Y(n_488) );
INVx1_ASAP7_75t_L g533 ( .A(n_244), .Y(n_533) );
AOI221x1_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_265), .B1(n_271), .B2(n_273), .C(n_274), .Y(n_249) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_250), .A2(n_338), .B1(n_405), .B2(n_406), .Y(n_404) );
AND2x2_ASAP7_75t_L g250 ( .A(n_251), .B(n_253), .Y(n_250) );
AND2x2_ASAP7_75t_L g296 ( .A(n_251), .B(n_297), .Y(n_296) );
AND2x2_ASAP7_75t_L g391 ( .A(n_251), .B(n_271), .Y(n_391) );
INVx1_ASAP7_75t_L g251 ( .A(n_252), .Y(n_251) );
AND2x2_ASAP7_75t_L g347 ( .A(n_252), .B(n_272), .Y(n_347) );
INVx1_ASAP7_75t_L g359 ( .A(n_253), .Y(n_359) );
AND2x2_ASAP7_75t_L g370 ( .A(n_253), .B(n_357), .Y(n_370) );
AND2x2_ASAP7_75t_L g437 ( .A(n_253), .B(n_332), .Y(n_437) );
INVx2_ASAP7_75t_L g299 ( .A(n_254), .Y(n_299) );
INVx2_ASAP7_75t_L g254 ( .A(n_255), .Y(n_254) );
AO21x2_ASAP7_75t_L g255 ( .A1(n_256), .A2(n_262), .B(n_263), .Y(n_255) );
AND2x2_ASAP7_75t_L g265 ( .A(n_266), .B(n_267), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g372 ( .A(n_266), .B(n_373), .Y(n_372) );
INVx1_ASAP7_75t_L g389 ( .A(n_266), .Y(n_389) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_267), .B(n_350), .Y(n_353) );
INVx3_ASAP7_75t_SL g267 ( .A(n_268), .Y(n_267) );
AOI21xp5_ASAP7_75t_L g433 ( .A1(n_268), .A2(n_389), .B(n_434), .Y(n_433) );
AND2x4_ASAP7_75t_L g268 ( .A(n_269), .B(n_270), .Y(n_268) );
NOR2xp33_ASAP7_75t_SL g411 ( .A(n_271), .B(n_297), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_272), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g363 ( .A(n_272), .B(n_291), .Y(n_363) );
NAND2xp5_ASAP7_75t_L g440 ( .A(n_272), .B(n_298), .Y(n_440) );
AND2x2_ASAP7_75t_L g309 ( .A(n_273), .B(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g376 ( .A(n_273), .Y(n_376) );
AOI21xp33_ASAP7_75t_L g274 ( .A1(n_275), .A2(n_279), .B(n_283), .Y(n_274) );
NAND2x1_ASAP7_75t_L g275 ( .A(n_276), .B(n_277), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g301 ( .A(n_276), .B(n_302), .Y(n_301) );
AND2x2_ASAP7_75t_L g325 ( .A(n_276), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_SL g337 ( .A(n_276), .Y(n_337) );
NOR2xp33_ASAP7_75t_L g382 ( .A(n_276), .B(n_383), .Y(n_382) );
INVx1_ASAP7_75t_L g361 ( .A(n_277), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_277), .B(n_398), .Y(n_397) );
NAND2xp5_ASAP7_75t_L g414 ( .A(n_277), .B(n_280), .Y(n_414) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_280), .B(n_281), .Y(n_279) );
AOI211xp5_ASAP7_75t_L g348 ( .A1(n_280), .A2(n_319), .B(n_349), .C(n_351), .Y(n_348) );
AOI221xp5_ASAP7_75t_L g366 ( .A1(n_280), .A2(n_367), .B1(n_370), .B2(n_371), .C(n_375), .Y(n_366) );
AND2x2_ASAP7_75t_L g362 ( .A(n_281), .B(n_315), .Y(n_362) );
INVx1_ASAP7_75t_L g281 ( .A(n_282), .Y(n_281) );
OR2x2_ASAP7_75t_L g283 ( .A(n_284), .B(n_285), .Y(n_283) );
INVx1_ASAP7_75t_L g285 ( .A(n_286), .Y(n_285) );
AND2x2_ASAP7_75t_L g322 ( .A(n_286), .B(n_323), .Y(n_322) );
AND2x2_ASAP7_75t_L g393 ( .A(n_286), .B(n_394), .Y(n_393) );
OAI211xp5_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_289), .B(n_295), .C(n_320), .Y(n_287) );
NAND3xp33_ASAP7_75t_SL g406 ( .A(n_288), .B(n_407), .C(n_408), .Y(n_406) );
OR2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_293), .Y(n_289) );
OR2x2_ASAP7_75t_L g379 ( .A(n_290), .B(n_380), .Y(n_379) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
INVx1_ASAP7_75t_L g293 ( .A(n_294), .Y(n_293) );
AOI221xp5_ASAP7_75t_L g295 ( .A1(n_296), .A2(n_300), .B1(n_303), .B2(n_309), .C(n_311), .Y(n_295) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_297), .B(n_307), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g339 ( .A(n_297), .B(n_340), .Y(n_339) );
AND2x2_ASAP7_75t_L g297 ( .A(n_298), .B(n_299), .Y(n_297) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
INVx1_ASAP7_75t_L g319 ( .A(n_302), .Y(n_319) );
OAI22xp5_ASAP7_75t_L g358 ( .A1(n_302), .A2(n_359), .B1(n_360), .B2(n_361), .Y(n_358) );
OR2x2_ASAP7_75t_L g439 ( .A(n_302), .B(n_350), .Y(n_439) );
NAND2xp5_ASAP7_75t_SL g303 ( .A(n_304), .B(n_306), .Y(n_303) );
INVxp67_ASAP7_75t_L g413 ( .A(n_305), .Y(n_413) );
NAND2xp5_ASAP7_75t_L g427 ( .A(n_307), .B(n_428), .Y(n_427) );
INVxp67_ASAP7_75t_L g314 ( .A(n_308), .Y(n_314) );
NAND2xp5_ASAP7_75t_L g318 ( .A(n_310), .B(n_319), .Y(n_318) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_310), .B(n_357), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g416 ( .A(n_310), .B(n_377), .Y(n_416) );
HB1xp67_ASAP7_75t_L g340 ( .A(n_314), .Y(n_340) );
INVx1_ASAP7_75t_L g316 ( .A(n_317), .Y(n_316) );
OR2x2_ASAP7_75t_L g430 ( .A(n_319), .B(n_350), .Y(n_430) );
INVx1_ASAP7_75t_L g320 ( .A(n_321), .Y(n_320) );
AND2x2_ASAP7_75t_L g321 ( .A(n_322), .B(n_325), .Y(n_321) );
INVx1_ASAP7_75t_L g323 ( .A(n_324), .Y(n_323) );
INVx1_ASAP7_75t_SL g408 ( .A(n_325), .Y(n_408) );
INVx1_ASAP7_75t_L g326 ( .A(n_327), .Y(n_326) );
OAI322xp33_ASAP7_75t_SL g328 ( .A1(n_329), .A2(n_334), .A3(n_335), .B1(n_336), .B2(n_339), .C1(n_341), .C2(n_343), .Y(n_328) );
OAI322xp33_ASAP7_75t_L g410 ( .A1(n_329), .A2(n_411), .A3(n_412), .B1(n_413), .B2(n_414), .C1(n_415), .C2(n_417), .Y(n_410) );
CKINVDCx16_ASAP7_75t_R g329 ( .A(n_330), .Y(n_329) );
AND2x2_ASAP7_75t_L g330 ( .A(n_331), .B(n_332), .Y(n_330) );
INVx4_ASAP7_75t_L g344 ( .A(n_331), .Y(n_344) );
AND2x2_ASAP7_75t_L g405 ( .A(n_331), .B(n_357), .Y(n_405) );
AND2x2_ASAP7_75t_L g418 ( .A(n_331), .B(n_419), .Y(n_418) );
CKINVDCx16_ASAP7_75t_R g429 ( .A(n_334), .Y(n_429) );
INVx1_ASAP7_75t_L g407 ( .A(n_335), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_337), .B(n_338), .Y(n_336) );
OR2x2_ASAP7_75t_L g341 ( .A(n_337), .B(n_342), .Y(n_341) );
AND2x2_ASAP7_75t_L g424 ( .A(n_337), .B(n_425), .Y(n_424) );
NAND2xp5_ASAP7_75t_L g435 ( .A(n_337), .B(n_378), .Y(n_435) );
OR2x2_ASAP7_75t_L g368 ( .A(n_340), .B(n_369), .Y(n_368) );
INVxp33_ASAP7_75t_L g385 ( .A(n_340), .Y(n_385) );
OAI221xp5_ASAP7_75t_SL g345 ( .A1(n_344), .A2(n_346), .B1(n_348), .B2(n_352), .C(n_354), .Y(n_345) );
NOR2xp67_ASAP7_75t_L g401 ( .A(n_344), .B(n_402), .Y(n_401) );
INVx1_ASAP7_75t_L g428 ( .A(n_344), .Y(n_428) );
INVx1_ASAP7_75t_SL g346 ( .A(n_347), .Y(n_346) );
INVx3_ASAP7_75t_SL g349 ( .A(n_350), .Y(n_349) );
AOI322xp5_ASAP7_75t_L g392 ( .A1(n_351), .A2(n_376), .A3(n_393), .B1(n_395), .B2(n_396), .C1(n_399), .C2(n_403), .Y(n_392) );
INVxp67_ASAP7_75t_L g352 ( .A(n_353), .Y(n_352) );
AOI22xp5_ASAP7_75t_L g354 ( .A1(n_355), .A2(n_358), .B1(n_362), .B2(n_363), .Y(n_354) );
INVx1_ASAP7_75t_L g355 ( .A(n_356), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g364 ( .A(n_365), .B(n_388), .Y(n_364) );
NAND2xp5_ASAP7_75t_SL g365 ( .A(n_366), .B(n_381), .Y(n_365) );
INVx1_ASAP7_75t_L g367 ( .A(n_368), .Y(n_367) );
NAND2xp5_ASAP7_75t_SL g399 ( .A(n_369), .B(n_400), .Y(n_399) );
INVx1_ASAP7_75t_SL g371 ( .A(n_372), .Y(n_371) );
NAND2xp33_ASAP7_75t_SL g386 ( .A(n_372), .B(n_383), .Y(n_386) );
INVx1_ASAP7_75t_SL g373 ( .A(n_374), .Y(n_373) );
OAI322xp33_ASAP7_75t_L g426 ( .A1(n_374), .A2(n_427), .A3(n_429), .B1(n_430), .B2(n_431), .C1(n_433), .C2(n_436), .Y(n_426) );
AOI21xp33_ASAP7_75t_SL g375 ( .A1(n_376), .A2(n_377), .B(n_379), .Y(n_375) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx2_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
NAND2xp5_ASAP7_75t_L g441 ( .A(n_384), .B(n_432), .Y(n_441) );
OAI211xp5_ASAP7_75t_SL g388 ( .A1(n_389), .A2(n_390), .B(n_392), .C(n_404), .Y(n_388) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g400 ( .A(n_401), .Y(n_400) );
NOR4xp25_ASAP7_75t_L g409 ( .A(n_410), .B(n_420), .C(n_426), .D(n_438), .Y(n_409) );
INVxp67_ASAP7_75t_L g415 ( .A(n_416), .Y(n_415) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
INVx1_ASAP7_75t_SL g423 ( .A(n_424), .Y(n_423) );
INVxp67_ASAP7_75t_L g431 ( .A(n_432), .Y(n_431) );
INVx1_ASAP7_75t_L g434 ( .A(n_435), .Y(n_434) );
CKINVDCx14_ASAP7_75t_R g436 ( .A(n_437), .Y(n_436) );
OAI21xp5_ASAP7_75t_SL g438 ( .A1(n_439), .A2(n_440), .B(n_441), .Y(n_438) );
AOI22xp5_ASAP7_75t_L g455 ( .A1(n_442), .A2(n_456), .B1(n_460), .B2(n_462), .Y(n_455) );
INVx1_ASAP7_75t_L g450 ( .A(n_443), .Y(n_450) );
INVx2_ASAP7_75t_L g443 ( .A(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g445 ( .A(n_446), .Y(n_445) );
AOI21xp33_ASAP7_75t_L g452 ( .A1(n_451), .A2(n_453), .B(n_759), .Y(n_452) );
INVx1_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
INVx1_ASAP7_75t_SL g456 ( .A(n_457), .Y(n_456) );
INVx2_ASAP7_75t_L g457 ( .A(n_458), .Y(n_457) );
INVx1_ASAP7_75t_L g458 ( .A(n_459), .Y(n_458) );
INVx1_ASAP7_75t_L g754 ( .A(n_459), .Y(n_754) );
INVx1_ASAP7_75t_L g460 ( .A(n_461), .Y(n_460) );
INVx6_ASAP7_75t_L g755 ( .A(n_461), .Y(n_755) );
INVx1_ASAP7_75t_L g462 ( .A(n_463), .Y(n_462) );
OR2x2_ASAP7_75t_L g463 ( .A(n_464), .B(n_667), .Y(n_463) );
NAND5xp2_ASAP7_75t_L g464 ( .A(n_465), .B(n_586), .C(n_601), .D(n_627), .E(n_649), .Y(n_464) );
NOR2xp33_ASAP7_75t_SL g465 ( .A(n_466), .B(n_566), .Y(n_465) );
OAI221xp5_ASAP7_75t_L g466 ( .A1(n_467), .A2(n_507), .B1(n_539), .B2(n_555), .C(n_556), .Y(n_466) );
NOR2xp33_ASAP7_75t_SL g467 ( .A(n_468), .B(n_499), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g615 ( .A(n_468), .B(n_616), .Y(n_615) );
INVx1_ASAP7_75t_SL g743 ( .A(n_468), .Y(n_743) );
AND2x2_ASAP7_75t_L g468 ( .A(n_469), .B(n_480), .Y(n_468) );
INVx1_ASAP7_75t_L g583 ( .A(n_469), .Y(n_583) );
AND2x2_ASAP7_75t_L g585 ( .A(n_469), .B(n_493), .Y(n_585) );
AND2x2_ASAP7_75t_L g595 ( .A(n_469), .B(n_492), .Y(n_595) );
HB1xp67_ASAP7_75t_L g613 ( .A(n_469), .Y(n_613) );
INVx1_ASAP7_75t_L g623 ( .A(n_469), .Y(n_623) );
OR2x2_ASAP7_75t_L g661 ( .A(n_469), .B(n_560), .Y(n_661) );
INVx2_ASAP7_75t_L g711 ( .A(n_469), .Y(n_711) );
NAND2xp5_ASAP7_75t_L g728 ( .A(n_469), .B(n_559), .Y(n_728) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_472), .A2(n_473), .B(n_474), .Y(n_471) );
NOR2xp67_ASAP7_75t_L g480 ( .A(n_481), .B(n_492), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_482), .Y(n_481) );
HB1xp67_ASAP7_75t_L g577 ( .A(n_482), .Y(n_577) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_482), .B(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_SL g643 ( .A(n_482), .B(n_583), .Y(n_643) );
INVx2_ASAP7_75t_L g482 ( .A(n_483), .Y(n_482) );
HB1xp67_ASAP7_75t_L g501 ( .A(n_483), .Y(n_501) );
INVx2_ASAP7_75t_L g560 ( .A(n_483), .Y(n_560) );
OR2x2_ASAP7_75t_L g622 ( .A(n_483), .B(n_623), .Y(n_622) );
AND2x2_ASAP7_75t_L g561 ( .A(n_492), .B(n_503), .Y(n_561) );
AND2x2_ASAP7_75t_L g578 ( .A(n_492), .B(n_558), .Y(n_578) );
INVx2_ASAP7_75t_L g492 ( .A(n_493), .Y(n_492) );
AND2x2_ASAP7_75t_L g502 ( .A(n_493), .B(n_503), .Y(n_502) );
BUFx2_ASAP7_75t_L g581 ( .A(n_493), .Y(n_581) );
AND2x2_ASAP7_75t_L g710 ( .A(n_493), .B(n_711), .Y(n_710) );
AOI21xp5_ASAP7_75t_L g523 ( .A1(n_496), .A2(n_524), .B(n_525), .Y(n_523) );
O2A1O1Ixp33_ASAP7_75t_L g534 ( .A1(n_496), .A2(n_535), .B(n_536), .C(n_537), .Y(n_534) );
OAI21xp5_ASAP7_75t_L g543 ( .A1(n_498), .A2(n_544), .B(n_547), .Y(n_543) );
INVx1_ASAP7_75t_L g555 ( .A(n_499), .Y(n_555) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_502), .Y(n_499) );
AND2x2_ASAP7_75t_L g673 ( .A(n_500), .B(n_561), .Y(n_673) );
INVx1_ASAP7_75t_L g500 ( .A(n_501), .Y(n_500) );
AND2x2_ASAP7_75t_L g674 ( .A(n_501), .B(n_585), .Y(n_674) );
O2A1O1Ixp33_ASAP7_75t_L g641 ( .A1(n_502), .A2(n_642), .B(n_644), .C(n_646), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g651 ( .A(n_502), .B(n_642), .Y(n_651) );
AOI221xp5_ASAP7_75t_L g714 ( .A1(n_502), .A2(n_572), .B1(n_715), .B2(n_716), .C(n_718), .Y(n_714) );
INVx1_ASAP7_75t_L g558 ( .A(n_503), .Y(n_558) );
INVx1_ASAP7_75t_L g594 ( .A(n_503), .Y(n_594) );
BUFx6f_ASAP7_75t_L g603 ( .A(n_503), .Y(n_603) );
INVx1_ASAP7_75t_SL g507 ( .A(n_508), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_509), .B(n_517), .Y(n_508) );
AND2x2_ASAP7_75t_L g620 ( .A(n_509), .B(n_565), .Y(n_620) );
NAND2xp5_ASAP7_75t_L g639 ( .A(n_509), .B(n_640), .Y(n_639) );
INVx2_ASAP7_75t_L g509 ( .A(n_510), .Y(n_509) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_510), .B(n_589), .Y(n_588) );
OR2x2_ASAP7_75t_L g712 ( .A(n_510), .B(n_713), .Y(n_712) );
INVx1_ASAP7_75t_L g744 ( .A(n_510), .Y(n_744) );
INVx2_ASAP7_75t_L g510 ( .A(n_511), .Y(n_510) );
INVx3_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
AND2x2_ASAP7_75t_L g600 ( .A(n_511), .B(n_554), .Y(n_600) );
NOR2x1_ASAP7_75t_L g609 ( .A(n_511), .B(n_610), .Y(n_609) );
AND2x2_ASAP7_75t_L g616 ( .A(n_511), .B(n_617), .Y(n_616) );
AND2x4_ASAP7_75t_L g511 ( .A(n_512), .B(n_513), .Y(n_511) );
INVx1_ASAP7_75t_L g552 ( .A(n_512), .Y(n_552) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_517), .B(n_656), .Y(n_691) );
INVx1_ASAP7_75t_SL g695 ( .A(n_517), .Y(n_695) );
AND2x2_ASAP7_75t_L g517 ( .A(n_518), .B(n_528), .Y(n_517) );
INVx3_ASAP7_75t_L g554 ( .A(n_518), .Y(n_554) );
AND2x2_ASAP7_75t_L g565 ( .A(n_518), .B(n_542), .Y(n_565) );
AND2x2_ASAP7_75t_L g587 ( .A(n_518), .B(n_588), .Y(n_587) );
AND2x2_ASAP7_75t_L g632 ( .A(n_518), .B(n_626), .Y(n_632) );
NAND2xp5_ASAP7_75t_L g713 ( .A(n_518), .B(n_564), .Y(n_713) );
INVx2_ASAP7_75t_L g535 ( .A(n_526), .Y(n_535) );
AND2x2_ASAP7_75t_L g553 ( .A(n_528), .B(n_554), .Y(n_553) );
INVx2_ASAP7_75t_L g564 ( .A(n_528), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_528), .B(n_542), .Y(n_589) );
AND2x2_ASAP7_75t_L g625 ( .A(n_528), .B(n_626), .Y(n_625) );
INVx1_ASAP7_75t_L g539 ( .A(n_540), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_541), .B(n_553), .Y(n_540) );
INVx1_ASAP7_75t_L g605 ( .A(n_541), .Y(n_605) );
AND2x2_ASAP7_75t_L g647 ( .A(n_541), .B(n_648), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g653 ( .A(n_541), .B(n_568), .Y(n_653) );
AOI21xp5_ASAP7_75t_SL g727 ( .A1(n_541), .A2(n_559), .B(n_582), .Y(n_727) );
AND2x2_ASAP7_75t_L g541 ( .A(n_542), .B(n_551), .Y(n_541) );
OR2x2_ASAP7_75t_L g570 ( .A(n_542), .B(n_551), .Y(n_570) );
AND2x2_ASAP7_75t_L g617 ( .A(n_542), .B(n_554), .Y(n_617) );
INVx2_ASAP7_75t_L g626 ( .A(n_542), .Y(n_626) );
INVx1_ASAP7_75t_L g732 ( .A(n_542), .Y(n_732) );
AND2x2_ASAP7_75t_L g656 ( .A(n_551), .B(n_626), .Y(n_656) );
INVx1_ASAP7_75t_L g681 ( .A(n_551), .Y(n_681) );
AND2x2_ASAP7_75t_L g590 ( .A(n_553), .B(n_574), .Y(n_590) );
AND2x2_ASAP7_75t_L g602 ( .A(n_553), .B(n_603), .Y(n_602) );
INVx2_ASAP7_75t_SL g720 ( .A(n_553), .Y(n_720) );
INVx2_ASAP7_75t_L g610 ( .A(n_554), .Y(n_610) );
AND2x2_ASAP7_75t_L g648 ( .A(n_554), .B(n_564), .Y(n_648) );
NAND2xp5_ASAP7_75t_L g731 ( .A(n_554), .B(n_732), .Y(n_731) );
OAI21xp33_ASAP7_75t_L g556 ( .A1(n_557), .A2(n_561), .B(n_562), .Y(n_556) );
AND2x2_ASAP7_75t_L g663 ( .A(n_557), .B(n_664), .Y(n_663) );
INVx1_ASAP7_75t_L g717 ( .A(n_557), .Y(n_717) );
AND2x2_ASAP7_75t_L g557 ( .A(n_558), .B(n_559), .Y(n_557) );
INVx1_ASAP7_75t_L g637 ( .A(n_558), .Y(n_637) );
BUFx2_ASAP7_75t_L g736 ( .A(n_558), .Y(n_736) );
BUFx2_ASAP7_75t_L g607 ( .A(n_559), .Y(n_607) );
AND2x2_ASAP7_75t_L g709 ( .A(n_559), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_L g559 ( .A(n_560), .Y(n_559) );
INVx1_ASAP7_75t_L g692 ( .A(n_560), .Y(n_692) );
AND2x4_ASAP7_75t_L g619 ( .A(n_561), .B(n_582), .Y(n_619) );
NAND2xp5_ASAP7_75t_SL g655 ( .A(n_561), .B(n_643), .Y(n_655) );
AOI32xp33_ASAP7_75t_L g579 ( .A1(n_562), .A2(n_580), .A3(n_582), .B1(n_584), .B2(n_585), .Y(n_579) );
AND2x2_ASAP7_75t_L g562 ( .A(n_563), .B(n_565), .Y(n_562) );
INVx3_ASAP7_75t_L g568 ( .A(n_563), .Y(n_568) );
OR2x2_ASAP7_75t_L g704 ( .A(n_563), .B(n_660), .Y(n_704) );
INVx2_ASAP7_75t_L g563 ( .A(n_564), .Y(n_563) );
AND2x2_ASAP7_75t_L g573 ( .A(n_564), .B(n_574), .Y(n_573) );
AND2x2_ASAP7_75t_L g680 ( .A(n_564), .B(n_681), .Y(n_680) );
AND2x2_ASAP7_75t_L g572 ( .A(n_565), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g584 ( .A(n_565), .B(n_574), .Y(n_584) );
INVx1_ASAP7_75t_L g705 ( .A(n_565), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g738 ( .A(n_565), .B(n_680), .Y(n_738) );
A2O1A1Ixp33_ASAP7_75t_L g566 ( .A1(n_567), .A2(n_571), .B(n_575), .C(n_579), .Y(n_566) );
OAI322xp33_ASAP7_75t_L g675 ( .A1(n_567), .A2(n_612), .A3(n_676), .B1(n_678), .B2(n_682), .C1(n_683), .C2(n_687), .Y(n_675) );
NAND2xp5_ASAP7_75t_L g567 ( .A(n_568), .B(n_569), .Y(n_567) );
INVxp67_ASAP7_75t_L g640 ( .A(n_568), .Y(n_640) );
INVx1_ASAP7_75t_SL g569 ( .A(n_570), .Y(n_569) );
OR2x2_ASAP7_75t_L g694 ( .A(n_570), .B(n_695), .Y(n_694) );
NOR2xp33_ASAP7_75t_L g741 ( .A(n_570), .B(n_610), .Y(n_741) );
INVxp67_ASAP7_75t_L g571 ( .A(n_572), .Y(n_571) );
INVx1_ASAP7_75t_L g633 ( .A(n_573), .Y(n_633) );
OR2x2_ASAP7_75t_L g719 ( .A(n_574), .B(n_720), .Y(n_719) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_577), .B(n_636), .Y(n_635) );
AND2x2_ASAP7_75t_L g628 ( .A(n_578), .B(n_607), .Y(n_628) );
AND2x2_ASAP7_75t_L g699 ( .A(n_578), .B(n_612), .Y(n_699) );
NAND2xp5_ASAP7_75t_L g721 ( .A(n_578), .B(n_686), .Y(n_721) );
AOI221xp5_ASAP7_75t_L g586 ( .A1(n_580), .A2(n_587), .B1(n_590), .B2(n_591), .C(n_596), .Y(n_586) );
OR2x2_ASAP7_75t_L g597 ( .A(n_580), .B(n_593), .Y(n_597) );
AND2x2_ASAP7_75t_L g685 ( .A(n_580), .B(n_686), .Y(n_685) );
AOI32xp33_ASAP7_75t_L g724 ( .A1(n_580), .A2(n_610), .A3(n_725), .B1(n_726), .B2(n_729), .Y(n_724) );
INVx2_ASAP7_75t_L g580 ( .A(n_581), .Y(n_580) );
NAND3xp33_ASAP7_75t_L g658 ( .A(n_581), .B(n_617), .C(n_640), .Y(n_658) );
AND2x2_ASAP7_75t_L g684 ( .A(n_581), .B(n_677), .Y(n_684) );
INVxp67_ASAP7_75t_L g664 ( .A(n_582), .Y(n_664) );
BUFx3_ASAP7_75t_L g582 ( .A(n_583), .Y(n_582) );
NAND2xp5_ASAP7_75t_SL g693 ( .A(n_585), .B(n_637), .Y(n_693) );
INVx2_ASAP7_75t_L g703 ( .A(n_585), .Y(n_703) );
NOR2xp33_ASAP7_75t_L g716 ( .A(n_585), .B(n_717), .Y(n_716) );
INVx1_ASAP7_75t_L g672 ( .A(n_588), .Y(n_672) );
OR2x2_ASAP7_75t_L g598 ( .A(n_589), .B(n_599), .Y(n_598) );
NOR2xp33_ASAP7_75t_L g708 ( .A(n_591), .B(n_709), .Y(n_708) );
AND2x2_ASAP7_75t_L g591 ( .A(n_592), .B(n_595), .Y(n_591) );
INVx1_ASAP7_75t_SL g592 ( .A(n_593), .Y(n_592) );
HB1xp67_ASAP7_75t_L g677 ( .A(n_594), .Y(n_677) );
AND2x2_ASAP7_75t_L g636 ( .A(n_595), .B(n_637), .Y(n_636) );
INVx1_ASAP7_75t_L g682 ( .A(n_595), .Y(n_682) );
HB1xp67_ASAP7_75t_L g707 ( .A(n_595), .Y(n_707) );
NOR2xp33_ASAP7_75t_L g596 ( .A(n_597), .B(n_598), .Y(n_596) );
AOI21xp33_ASAP7_75t_SL g621 ( .A1(n_597), .A2(n_622), .B(n_624), .Y(n_621) );
INVx1_ASAP7_75t_L g599 ( .A(n_600), .Y(n_599) );
AND2x2_ASAP7_75t_L g715 ( .A(n_600), .B(n_625), .Y(n_715) );
AOI211xp5_ASAP7_75t_L g601 ( .A1(n_602), .A2(n_604), .B(n_614), .C(n_621), .Y(n_601) );
AND2x2_ASAP7_75t_L g645 ( .A(n_603), .B(n_613), .Y(n_645) );
INVx2_ASAP7_75t_L g660 ( .A(n_603), .Y(n_660) );
OR2x2_ASAP7_75t_L g698 ( .A(n_603), .B(n_661), .Y(n_698) );
NAND2xp5_ASAP7_75t_L g740 ( .A(n_603), .B(n_741), .Y(n_740) );
AOI211xp5_ASAP7_75t_SL g604 ( .A1(n_605), .A2(n_606), .B(n_608), .C(n_611), .Y(n_604) );
INVxp67_ASAP7_75t_L g606 ( .A(n_607), .Y(n_606) );
NAND2xp5_ASAP7_75t_L g644 ( .A(n_607), .B(n_645), .Y(n_644) );
OAI211xp5_ASAP7_75t_L g726 ( .A1(n_608), .A2(n_703), .B(n_727), .C(n_728), .Y(n_726) );
INVx1_ASAP7_75t_L g608 ( .A(n_609), .Y(n_608) );
NAND2x1p5_ASAP7_75t_L g624 ( .A(n_609), .B(n_625), .Y(n_624) );
AND2x2_ASAP7_75t_L g666 ( .A(n_610), .B(n_656), .Y(n_666) );
INVx1_ASAP7_75t_L g671 ( .A(n_610), .Y(n_671) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
INVx1_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
NAND2xp5_ASAP7_75t_SL g614 ( .A(n_615), .B(n_618), .Y(n_614) );
INVxp33_ASAP7_75t_L g722 ( .A(n_616), .Y(n_722) );
AND2x2_ASAP7_75t_L g701 ( .A(n_617), .B(n_680), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g618 ( .A(n_619), .B(n_620), .Y(n_618) );
AOI21xp5_ASAP7_75t_L g683 ( .A1(n_622), .A2(n_684), .B(n_685), .Y(n_683) );
OAI322xp33_ASAP7_75t_L g702 ( .A1(n_624), .A2(n_703), .A3(n_704), .B1(n_705), .B2(n_706), .C1(n_708), .C2(n_712), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_628), .A2(n_629), .B1(n_634), .B2(n_638), .C(n_641), .Y(n_627) );
INVx2_ASAP7_75t_L g629 ( .A(n_630), .Y(n_629) );
OR2x2_ASAP7_75t_L g630 ( .A(n_631), .B(n_633), .Y(n_630) );
INVx1_ASAP7_75t_L g631 ( .A(n_632), .Y(n_631) );
AND2x2_ASAP7_75t_L g679 ( .A(n_632), .B(n_680), .Y(n_679) );
INVx1_ASAP7_75t_L g634 ( .A(n_635), .Y(n_634) );
INVx1_ASAP7_75t_L g723 ( .A(n_636), .Y(n_723) );
INVxp67_ASAP7_75t_L g638 ( .A(n_639), .Y(n_638) );
NOR2xp33_ASAP7_75t_L g725 ( .A(n_639), .B(n_659), .Y(n_725) );
INVx2_ASAP7_75t_L g642 ( .A(n_643), .Y(n_642) );
INVx1_ASAP7_75t_SL g646 ( .A(n_647), .Y(n_646) );
AND2x2_ASAP7_75t_L g688 ( .A(n_648), .B(n_656), .Y(n_688) );
AOI221xp5_ASAP7_75t_L g649 ( .A1(n_650), .A2(n_652), .B1(n_654), .B2(n_656), .C(n_657), .Y(n_649) );
INVx1_ASAP7_75t_L g650 ( .A(n_651), .Y(n_650) );
AOI221xp5_ASAP7_75t_L g668 ( .A1(n_652), .A2(n_669), .B1(n_673), .B2(n_674), .C(n_675), .Y(n_668) );
INVx1_ASAP7_75t_L g652 ( .A(n_653), .Y(n_652) );
INVxp67_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
NAND2xp5_ASAP7_75t_L g670 ( .A(n_656), .B(n_671), .Y(n_670) );
OAI22xp5_ASAP7_75t_L g657 ( .A1(n_658), .A2(n_659), .B1(n_662), .B2(n_665), .Y(n_657) );
OR2x2_ASAP7_75t_L g659 ( .A(n_660), .B(n_661), .Y(n_659) );
INVx2_ASAP7_75t_SL g686 ( .A(n_661), .Y(n_686) );
INVxp67_ASAP7_75t_L g662 ( .A(n_663), .Y(n_662) );
INVx1_ASAP7_75t_L g665 ( .A(n_666), .Y(n_665) );
NAND5xp2_ASAP7_75t_L g667 ( .A(n_668), .B(n_689), .C(n_714), .D(n_724), .E(n_734), .Y(n_667) );
NAND2xp5_ASAP7_75t_SL g669 ( .A(n_670), .B(n_672), .Y(n_669) );
NOR4xp25_ASAP7_75t_L g742 ( .A(n_671), .B(n_677), .C(n_743), .D(n_744), .Y(n_742) );
AOI221xp5_ASAP7_75t_L g734 ( .A1(n_674), .A2(n_735), .B1(n_737), .B2(n_739), .C(n_742), .Y(n_734) );
INVx1_ASAP7_75t_L g676 ( .A(n_677), .Y(n_676) );
INVx1_ASAP7_75t_L g678 ( .A(n_679), .Y(n_678) );
INVx1_ASAP7_75t_L g733 ( .A(n_680), .Y(n_733) );
OAI322xp33_ASAP7_75t_L g690 ( .A1(n_684), .A2(n_691), .A3(n_692), .B1(n_693), .B2(n_694), .C1(n_696), .C2(n_700), .Y(n_690) );
INVx1_ASAP7_75t_SL g687 ( .A(n_688), .Y(n_687) );
NOR2xp33_ASAP7_75t_L g689 ( .A(n_690), .B(n_702), .Y(n_689) );
NOR2xp33_ASAP7_75t_L g696 ( .A(n_697), .B(n_699), .Y(n_696) );
INVx2_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_L g700 ( .A(n_701), .Y(n_700) );
INVx1_ASAP7_75t_L g706 ( .A(n_707), .Y(n_706) );
AND2x2_ASAP7_75t_L g735 ( .A(n_710), .B(n_736), .Y(n_735) );
OAI22xp33_ASAP7_75t_L g718 ( .A1(n_719), .A2(n_721), .B1(n_722), .B2(n_723), .Y(n_718) );
INVx1_ASAP7_75t_L g729 ( .A(n_730), .Y(n_729) );
OR2x2_ASAP7_75t_L g730 ( .A(n_731), .B(n_733), .Y(n_730) );
INVx1_ASAP7_75t_L g737 ( .A(n_738), .Y(n_737) );
INVxp67_ASAP7_75t_L g739 ( .A(n_740), .Y(n_739) );
INVx1_ASAP7_75t_L g745 ( .A(n_746), .Y(n_745) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
INVx1_ASAP7_75t_SL g756 ( .A(n_757), .Y(n_756) );
INVx2_ASAP7_75t_L g757 ( .A(n_758), .Y(n_757) );
INVx1_ASAP7_75t_SL g760 ( .A(n_761), .Y(n_760) );
endmodule