module fake_jpeg_16357_n_290 (n_11, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_6, n_5, n_7, n_290);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_290;

wire n_159;
wire n_117;
wire n_253;
wire n_286;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_182;
wire n_19;
wire n_84;
wire n_59;
wire n_98;
wire n_252;
wire n_251;
wire n_273;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_279;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_127;
wire n_76;
wire n_154;
wire n_278;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_281;
wire n_31;
wire n_155;
wire n_207;
wire n_277;
wire n_255;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_284;
wire n_272;
wire n_288;
wire n_280;
wire n_171;
wire n_263;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_289;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_267;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_274;
wire n_186;
wire n_24;
wire n_44;
wire n_276;
wire n_143;
wire n_202;
wire n_17;
wire n_25;
wire n_269;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_287;
wire n_121;
wire n_99;
wire n_130;
wire n_102;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_257;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_18;
wire n_20;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_259;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_266;
wire n_34;
wire n_283;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_261;
wire n_89;
wire n_146;
wire n_104;
wire n_285;
wire n_215;
wire n_262;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_271;
wire n_216;
wire n_217;
wire n_264;
wire n_184;
wire n_53;
wire n_268;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_265;
wire n_176;
wire n_199;
wire n_112;
wire n_260;
wire n_270;
wire n_222;
wire n_95;
wire n_275;
wire n_221;
wire n_151;
wire n_256;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_140;
wire n_82;
wire n_128;
wire n_118;
wire n_258;
wire n_282;
wire n_96;

BUFx3_ASAP7_75t_L g13 ( 
.A(n_5),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_10),
.Y(n_14)
);

INVx6_ASAP7_75t_L g15 ( 
.A(n_7),
.Y(n_15)
);

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

INVx1_ASAP7_75t_L g17 ( 
.A(n_9),
.Y(n_17)
);

BUFx10_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_2),
.Y(n_19)
);

INVx8_ASAP7_75t_L g20 ( 
.A(n_0),
.Y(n_20)
);

CKINVDCx14_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

BUFx5_ASAP7_75t_L g22 ( 
.A(n_9),
.Y(n_22)
);

INVx2_ASAP7_75t_L g23 ( 
.A(n_6),
.Y(n_23)
);

INVx3_ASAP7_75t_L g24 ( 
.A(n_0),
.Y(n_24)
);

INVx1_ASAP7_75t_SL g25 ( 
.A(n_9),
.Y(n_25)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_6),
.Y(n_27)
);

INVx13_ASAP7_75t_L g28 ( 
.A(n_18),
.Y(n_28)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_28),
.Y(n_40)
);

BUFx3_ASAP7_75t_L g29 ( 
.A(n_18),
.Y(n_29)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_29),
.Y(n_47)
);

INVx4_ASAP7_75t_L g30 ( 
.A(n_18),
.Y(n_30)
);

INVx4_ASAP7_75t_L g46 ( 
.A(n_30),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_31),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g43 ( 
.A(n_32),
.B(n_36),
.Y(n_43)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_18),
.Y(n_33)
);

INVx5_ASAP7_75t_L g38 ( 
.A(n_33),
.Y(n_38)
);

BUFx4f_ASAP7_75t_L g34 ( 
.A(n_16),
.Y(n_34)
);

INVx4_ASAP7_75t_L g51 ( 
.A(n_34),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g35 ( 
.A(n_16),
.Y(n_35)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_35),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_SL g36 ( 
.A(n_17),
.B(n_0),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_16),
.Y(n_37)
);

INVx3_ASAP7_75t_L g41 ( 
.A(n_37),
.Y(n_41)
);

AOI22xp33_ASAP7_75t_L g39 ( 
.A1(n_36),
.A2(n_15),
.B1(n_23),
.B2(n_25),
.Y(n_39)
);

AOI22xp5_ASAP7_75t_L g55 ( 
.A1(n_39),
.A2(n_52),
.B1(n_15),
.B2(n_24),
.Y(n_55)
);

OR2x2_ASAP7_75t_L g42 ( 
.A(n_32),
.B(n_26),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_42),
.B(n_50),
.Y(n_65)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_31),
.Y(n_44)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_31),
.Y(n_45)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_45),
.Y(n_67)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_31),
.Y(n_48)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

INVx3_ASAP7_75t_L g50 ( 
.A(n_35),
.Y(n_50)
);

OA22x2_ASAP7_75t_L g52 ( 
.A1(n_34),
.A2(n_23),
.B1(n_15),
.B2(n_18),
.Y(n_52)
);

INVx4_ASAP7_75t_L g54 ( 
.A(n_47),
.Y(n_54)
);

INVx11_ASAP7_75t_L g77 ( 
.A(n_54),
.Y(n_77)
);

AND2x2_ASAP7_75t_L g75 ( 
.A(n_55),
.B(n_28),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_38),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_L g87 ( 
.A1(n_56),
.A2(n_68),
.B(n_71),
.Y(n_87)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_43),
.B(n_32),
.Y(n_57)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_57),
.B(n_70),
.Y(n_78)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_52),
.A2(n_34),
.B1(n_28),
.B2(n_33),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_SL g92 ( 
.A1(n_58),
.A2(n_69),
.B1(n_72),
.B2(n_51),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_49),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_60),
.B(n_61),
.Y(n_96)
);

INVxp67_ASAP7_75t_L g61 ( 
.A(n_52),
.Y(n_61)
);

INVx5_ASAP7_75t_SL g62 ( 
.A(n_40),
.Y(n_62)
);

OAI22xp33_ASAP7_75t_SL g84 ( 
.A1(n_62),
.A2(n_64),
.B1(n_53),
.B2(n_51),
.Y(n_84)
);

CKINVDCx20_ASAP7_75t_R g64 ( 
.A(n_49),
.Y(n_64)
);

CKINVDCx9p33_ASAP7_75t_R g66 ( 
.A(n_40),
.Y(n_66)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_66),
.Y(n_76)
);

AOI22xp33_ASAP7_75t_SL g68 ( 
.A1(n_38),
.A2(n_25),
.B1(n_24),
.B2(n_20),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_L g69 ( 
.A1(n_52),
.A2(n_34),
.B1(n_20),
.B2(n_33),
.Y(n_69)
);

XNOR2xp5_ASAP7_75t_L g70 ( 
.A(n_42),
.B(n_34),
.Y(n_70)
);

AOI21xp5_ASAP7_75t_L g71 ( 
.A1(n_41),
.A2(n_34),
.B(n_2),
.Y(n_71)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_41),
.A2(n_33),
.B1(n_30),
.B2(n_37),
.Y(n_72)
);

INVx5_ASAP7_75t_L g73 ( 
.A(n_46),
.Y(n_73)
);

INVx3_ASAP7_75t_L g79 ( 
.A(n_73),
.Y(n_79)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_46),
.B(n_17),
.Y(n_74)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_74),
.Y(n_82)
);

AOI22xp5_ASAP7_75t_L g99 ( 
.A1(n_75),
.A2(n_58),
.B1(n_65),
.B2(n_67),
.Y(n_99)
);

OR2x2_ASAP7_75t_L g80 ( 
.A(n_70),
.B(n_26),
.Y(n_80)
);

NOR2xp33_ASAP7_75t_SL g115 ( 
.A(n_80),
.B(n_81),
.Y(n_115)
);

NAND2xp5_ASAP7_75t_L g81 ( 
.A(n_57),
.B(n_53),
.Y(n_81)
);

INVx2_ASAP7_75t_L g83 ( 
.A(n_73),
.Y(n_83)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_83),
.Y(n_107)
);

CKINVDCx14_ASAP7_75t_R g118 ( 
.A(n_84),
.Y(n_118)
);

INVx1_ASAP7_75t_L g85 ( 
.A(n_63),
.Y(n_85)
);

INVx1_ASAP7_75t_L g101 ( 
.A(n_85),
.Y(n_101)
);

BUFx2_ASAP7_75t_L g86 ( 
.A(n_66),
.Y(n_86)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_86),
.Y(n_119)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_73),
.Y(n_88)
);

INVx2_ASAP7_75t_L g110 ( 
.A(n_88),
.Y(n_110)
);

OAI22xp33_ASAP7_75t_L g89 ( 
.A1(n_69),
.A2(n_50),
.B1(n_48),
.B2(n_45),
.Y(n_89)
);

OAI22xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_94),
.B1(n_62),
.B2(n_60),
.Y(n_111)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_63),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g103 ( 
.A(n_90),
.B(n_91),
.Y(n_103)
);

INVx4_ASAP7_75t_L g91 ( 
.A(n_59),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_L g97 ( 
.A1(n_92),
.A2(n_71),
.B1(n_58),
.B2(n_72),
.Y(n_97)
);

INVx4_ASAP7_75t_L g93 ( 
.A(n_59),
.Y(n_93)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_93),
.B(n_54),
.Y(n_105)
);

OAI22xp5_ASAP7_75t_SL g94 ( 
.A1(n_55),
.A2(n_44),
.B1(n_30),
.B2(n_28),
.Y(n_94)
);

INVx2_ASAP7_75t_L g95 ( 
.A(n_67),
.Y(n_95)
);

INVx3_ASAP7_75t_L g102 ( 
.A(n_95),
.Y(n_102)
);

AOI22xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_37),
.B1(n_35),
.B2(n_14),
.Y(n_136)
);

OR2x2_ASAP7_75t_L g98 ( 
.A(n_82),
.B(n_65),
.Y(n_98)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_98),
.B(n_116),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_L g126 ( 
.A1(n_99),
.A2(n_111),
.B1(n_113),
.B2(n_79),
.Y(n_126)
);

HAxp5_ASAP7_75t_SL g100 ( 
.A(n_87),
.B(n_58),
.CON(n_100),
.SN(n_100)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_100),
.B(n_112),
.Y(n_123)
);

AND2x2_ASAP7_75t_SL g104 ( 
.A(n_81),
.B(n_58),
.Y(n_104)
);

INVx1_ASAP7_75t_L g120 ( 
.A(n_104),
.Y(n_120)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_105),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_91),
.B(n_74),
.Y(n_106)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_106),
.Y(n_124)
);

AND2x2_ASAP7_75t_SL g108 ( 
.A(n_78),
.B(n_64),
.Y(n_108)
);

MAJIxp5_ASAP7_75t_L g135 ( 
.A(n_108),
.B(n_80),
.C(n_29),
.Y(n_135)
);

CKINVDCx16_ASAP7_75t_R g109 ( 
.A(n_96),
.Y(n_109)
);

NAND2xp5_ASAP7_75t_SL g131 ( 
.A(n_109),
.B(n_85),
.Y(n_131)
);

INVx8_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

OAI22xp5_ASAP7_75t_SL g113 ( 
.A1(n_87),
.A2(n_30),
.B1(n_62),
.B2(n_37),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g114 ( 
.A(n_93),
.B(n_54),
.Y(n_114)
);

INVx1_ASAP7_75t_L g139 ( 
.A(n_114),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_95),
.B(n_18),
.Y(n_116)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_78),
.B(n_29),
.C(n_13),
.Y(n_117)
);

XNOR2xp5_ASAP7_75t_SL g137 ( 
.A(n_117),
.B(n_35),
.Y(n_137)
);

AOI22x1_ASAP7_75t_L g122 ( 
.A1(n_97),
.A2(n_92),
.B1(n_94),
.B2(n_89),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_SL g162 ( 
.A1(n_122),
.A2(n_130),
.B1(n_136),
.B2(n_112),
.Y(n_162)
);

AND2x2_ASAP7_75t_L g164 ( 
.A(n_126),
.B(n_111),
.Y(n_164)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_101),
.Y(n_127)
);

NAND2xp5_ASAP7_75t_SL g149 ( 
.A(n_127),
.B(n_128),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g128 ( 
.A(n_101),
.Y(n_128)
);

XOR2xp5_ASAP7_75t_L g129 ( 
.A(n_117),
.B(n_75),
.Y(n_129)
);

NAND2xp5_ASAP7_75t_L g160 ( 
.A(n_129),
.B(n_135),
.Y(n_160)
);

AOI22x1_ASAP7_75t_L g130 ( 
.A1(n_113),
.A2(n_75),
.B1(n_83),
.B2(n_88),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g154 ( 
.A(n_131),
.B(n_132),
.Y(n_154)
);

NOR2xp33_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_77),
.Y(n_132)
);

INVxp33_ASAP7_75t_L g133 ( 
.A(n_105),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g159 ( 
.A(n_133),
.B(n_140),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_118),
.A2(n_76),
.B1(n_77),
.B2(n_17),
.Y(n_134)
);

CKINVDCx16_ASAP7_75t_R g145 ( 
.A(n_134),
.Y(n_145)
);

OAI21xp5_ASAP7_75t_L g144 ( 
.A1(n_137),
.A2(n_115),
.B(n_98),
.Y(n_144)
);

XNOR2xp5_ASAP7_75t_SL g138 ( 
.A(n_117),
.B(n_11),
.Y(n_138)
);

OAI21xp33_ASAP7_75t_L g147 ( 
.A1(n_138),
.A2(n_109),
.B(n_98),
.Y(n_147)
);

MAJIxp5_ASAP7_75t_L g140 ( 
.A(n_108),
.B(n_29),
.C(n_13),
.Y(n_140)
);

NAND2xp5_ASAP7_75t_L g141 ( 
.A(n_108),
.B(n_27),
.Y(n_141)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_141),
.Y(n_148)
);

OAI22xp5_ASAP7_75t_L g142 ( 
.A1(n_118),
.A2(n_14),
.B1(n_27),
.B2(n_21),
.Y(n_142)
);

INVxp67_ASAP7_75t_L g158 ( 
.A(n_142),
.Y(n_158)
);

MAJIxp5_ASAP7_75t_L g143 ( 
.A(n_108),
.B(n_104),
.C(n_115),
.Y(n_143)
);

NOR2xp33_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_104),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_L g170 ( 
.A(n_144),
.B(n_163),
.Y(n_170)
);

CKINVDCx20_ASAP7_75t_R g146 ( 
.A(n_139),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_146),
.B(n_164),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_SL g190 ( 
.A(n_147),
.B(n_116),
.Y(n_190)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_125),
.Y(n_150)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_150),
.Y(n_173)
);

HB1xp67_ASAP7_75t_L g151 ( 
.A(n_125),
.Y(n_151)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_151),
.B(n_119),
.Y(n_193)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_124),
.Y(n_152)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_152),
.Y(n_180)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_121),
.Y(n_153)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_153),
.Y(n_183)
);

OR2x2_ASAP7_75t_L g155 ( 
.A(n_120),
.B(n_99),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_168),
.Y(n_175)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_121),
.Y(n_156)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_156),
.Y(n_186)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_141),
.B(n_99),
.Y(n_157)
);

NOR2xp33_ASAP7_75t_SL g192 ( 
.A(n_157),
.B(n_102),
.Y(n_192)
);

AOI21xp5_ASAP7_75t_L g161 ( 
.A1(n_123),
.A2(n_104),
.B(n_103),
.Y(n_161)
);

AOI21xp5_ASAP7_75t_L g188 ( 
.A1(n_161),
.A2(n_166),
.B(n_114),
.Y(n_188)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_162),
.A2(n_122),
.B1(n_140),
.B2(n_135),
.Y(n_179)
);

CKINVDCx20_ASAP7_75t_R g165 ( 
.A(n_120),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g176 ( 
.A(n_165),
.B(n_104),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_130),
.A2(n_107),
.B1(n_110),
.B2(n_102),
.Y(n_166)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_136),
.Y(n_167)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_167),
.Y(n_184)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_133),
.Y(n_168)
);

INVx13_ASAP7_75t_L g169 ( 
.A(n_130),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g171 ( 
.A(n_169),
.B(n_106),
.Y(n_171)
);

AOI22xp33_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_179),
.B1(n_188),
.B2(n_190),
.Y(n_210)
);

NOR2xp33_ASAP7_75t_L g174 ( 
.A(n_152),
.B(n_103),
.Y(n_174)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_174),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_176),
.Y(n_195)
);

HB1xp67_ASAP7_75t_L g177 ( 
.A(n_168),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_177),
.B(n_150),
.Y(n_197)
);

MAJIxp5_ASAP7_75t_L g178 ( 
.A(n_160),
.B(n_143),
.C(n_129),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g213 ( 
.A(n_178),
.B(n_13),
.C(n_22),
.Y(n_213)
);

XNOR2x1_ASAP7_75t_L g181 ( 
.A(n_160),
.B(n_138),
.Y(n_181)
);

XOR2xp5_ASAP7_75t_L g203 ( 
.A(n_181),
.B(n_182),
.Y(n_203)
);

XOR2xp5_ASAP7_75t_L g182 ( 
.A(n_159),
.B(n_137),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_L g185 ( 
.A(n_146),
.B(n_110),
.Y(n_185)
);

INVx1_ASAP7_75t_L g196 ( 
.A(n_185),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g187 ( 
.A1(n_169),
.A2(n_122),
.B1(n_165),
.B2(n_167),
.Y(n_187)
);

INVx1_ASAP7_75t_L g204 ( 
.A(n_187),
.Y(n_204)
);

INVxp67_ASAP7_75t_L g189 ( 
.A(n_149),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_189),
.B(n_154),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_SL g191 ( 
.A1(n_162),
.A2(n_102),
.B1(n_107),
.B2(n_119),
.Y(n_191)
);

AOI22xp5_ASAP7_75t_L g199 ( 
.A1(n_191),
.A2(n_164),
.B1(n_156),
.B2(n_153),
.Y(n_199)
);

CKINVDCx14_ASAP7_75t_R g208 ( 
.A(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_193),
.B(n_158),
.Y(n_205)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_197),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g198 ( 
.A(n_184),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g215 ( 
.A(n_198),
.B(n_205),
.Y(n_215)
);

OAI22xp5_ASAP7_75t_SL g223 ( 
.A1(n_199),
.A2(n_209),
.B1(n_212),
.B2(n_210),
.Y(n_223)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_182),
.B(n_161),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g219 ( 
.A(n_200),
.B(n_213),
.C(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g229 ( 
.A(n_201),
.B(n_202),
.Y(n_229)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_189),
.B(n_148),
.Y(n_202)
);

HB1xp67_ASAP7_75t_L g206 ( 
.A(n_180),
.Y(n_206)
);

HB1xp67_ASAP7_75t_L g227 ( 
.A(n_206),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g207 ( 
.A(n_180),
.B(n_148),
.Y(n_207)
);

NOR2xp33_ASAP7_75t_SL g216 ( 
.A(n_207),
.B(n_173),
.Y(n_216)
);

AOI22xp5_ASAP7_75t_L g209 ( 
.A1(n_172),
.A2(n_164),
.B1(n_158),
.B2(n_155),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_175),
.B(n_155),
.Y(n_211)
);

XOR2xp5_ASAP7_75t_L g214 ( 
.A(n_211),
.B(n_187),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_L g212 ( 
.A1(n_175),
.A2(n_145),
.B1(n_157),
.B2(n_144),
.Y(n_212)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_214),
.B(n_216),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_SL g217 ( 
.A(n_200),
.B(n_181),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g237 ( 
.A(n_217),
.B(n_219),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_SL g218 ( 
.A(n_201),
.B(n_183),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_218),
.B(n_1),
.Y(n_245)
);

NAND3xp33_ASAP7_75t_L g220 ( 
.A(n_211),
.B(n_190),
.C(n_170),
.Y(n_220)
);

AOI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_220),
.A2(n_195),
.B1(n_194),
.B2(n_196),
.Y(n_239)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_203),
.B(n_170),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g236 ( 
.A(n_221),
.B(n_225),
.C(n_226),
.Y(n_236)
);

AOI22xp5_ASAP7_75t_L g222 ( 
.A1(n_204),
.A2(n_173),
.B1(n_186),
.B2(n_183),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_222),
.A2(n_224),
.B1(n_21),
.B2(n_19),
.Y(n_241)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_223),
.B(n_228),
.Y(n_232)
);

AOI22xp5_ASAP7_75t_L g224 ( 
.A1(n_208),
.A2(n_186),
.B1(n_191),
.B2(n_188),
.Y(n_224)
);

AOI21xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_179),
.B(n_10),
.Y(n_225)
);

XOR2xp5_ASAP7_75t_L g226 ( 
.A(n_203),
.B(n_22),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g228 ( 
.A(n_199),
.B(n_22),
.Y(n_228)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_209),
.B(n_19),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g234 ( 
.A(n_230),
.B(n_213),
.Y(n_234)
);

BUFx12_ASAP7_75t_L g233 ( 
.A(n_215),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_L g257 ( 
.A(n_233),
.B(n_238),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_SL g251 ( 
.A(n_234),
.B(n_243),
.Y(n_251)
);

BUFx12_ASAP7_75t_L g238 ( 
.A(n_231),
.Y(n_238)
);

INVx1_ASAP7_75t_L g249 ( 
.A(n_239),
.Y(n_249)
);

BUFx12_ASAP7_75t_L g240 ( 
.A(n_220),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_240),
.B(n_242),
.Y(n_258)
);

INVx1_ASAP7_75t_L g255 ( 
.A(n_241),
.Y(n_255)
);

BUFx12_ASAP7_75t_L g242 ( 
.A(n_229),
.Y(n_242)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_230),
.A2(n_12),
.B1(n_11),
.B2(n_8),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_226),
.B(n_12),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_244),
.B(n_246),
.Y(n_253)
);

CKINVDCx20_ASAP7_75t_R g248 ( 
.A(n_245),
.Y(n_248)
);

HB1xp67_ASAP7_75t_L g246 ( 
.A(n_227),
.Y(n_246)
);

AOI21xp5_ASAP7_75t_L g247 ( 
.A1(n_240),
.A2(n_228),
.B(n_221),
.Y(n_247)
);

INVx1_ASAP7_75t_L g260 ( 
.A(n_247),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g250 ( 
.A(n_236),
.B(n_217),
.C(n_19),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g263 ( 
.A(n_250),
.B(n_252),
.C(n_254),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g252 ( 
.A(n_237),
.B(n_19),
.C(n_2),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_232),
.B(n_1),
.C(n_2),
.Y(n_254)
);

AOI21xp5_ASAP7_75t_L g256 ( 
.A1(n_235),
.A2(n_12),
.B(n_11),
.Y(n_256)
);

OAI21xp5_ASAP7_75t_L g266 ( 
.A1(n_256),
.A2(n_8),
.B(n_3),
.Y(n_266)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_257),
.B(n_235),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_SL g275 ( 
.A(n_259),
.B(n_262),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_248),
.B(n_246),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_261),
.B(n_264),
.Y(n_277)
);

NAND2xp5_ASAP7_75t_L g262 ( 
.A(n_258),
.B(n_245),
.Y(n_262)
);

AND2x2_ASAP7_75t_L g264 ( 
.A(n_249),
.B(n_242),
.Y(n_264)
);

NAND2xp5_ASAP7_75t_SL g265 ( 
.A(n_253),
.B(n_238),
.Y(n_265)
);

OAI21xp5_ASAP7_75t_L g273 ( 
.A1(n_265),
.A2(n_1),
.B(n_3),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_267),
.Y(n_276)
);

NOR2xp33_ASAP7_75t_SL g267 ( 
.A(n_251),
.B(n_233),
.Y(n_267)
);

HB1xp67_ASAP7_75t_L g268 ( 
.A(n_254),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g270 ( 
.A(n_268),
.B(n_269),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_252),
.B(n_8),
.Y(n_269)
);

OAI21xp5_ASAP7_75t_SL g271 ( 
.A1(n_261),
.A2(n_247),
.B(n_255),
.Y(n_271)
);

OAI21xp5_ASAP7_75t_SL g279 ( 
.A1(n_271),
.A2(n_1),
.B(n_4),
.Y(n_279)
);

AND3x1_ASAP7_75t_L g272 ( 
.A(n_260),
.B(n_250),
.C(n_3),
.Y(n_272)
);

AOI322xp5_ASAP7_75t_L g281 ( 
.A1(n_272),
.A2(n_4),
.A3(n_5),
.B1(n_6),
.B2(n_7),
.C1(n_276),
.C2(n_277),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g280 ( 
.A(n_273),
.B(n_4),
.Y(n_280)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_265),
.B(n_86),
.Y(n_274)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_274),
.B(n_263),
.Y(n_278)
);

NAND2xp5_ASAP7_75t_L g283 ( 
.A(n_278),
.B(n_279),
.Y(n_283)
);

AND2x2_ASAP7_75t_L g284 ( 
.A(n_280),
.B(n_281),
.Y(n_284)
);

AOI22xp5_ASAP7_75t_SL g282 ( 
.A1(n_272),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_SL g285 ( 
.A(n_284),
.B(n_275),
.Y(n_285)
);

INVx1_ASAP7_75t_L g286 ( 
.A(n_285),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g287 ( 
.A(n_286),
.B(n_270),
.Y(n_287)
);

CKINVDCx20_ASAP7_75t_R g288 ( 
.A(n_287),
.Y(n_288)
);

AO21x1_ASAP7_75t_L g289 ( 
.A1(n_288),
.A2(n_283),
.B(n_281),
.Y(n_289)
);

A2O1A1Ixp33_ASAP7_75t_L g290 ( 
.A1(n_289),
.A2(n_282),
.B(n_274),
.C(n_5),
.Y(n_290)
);


endmodule