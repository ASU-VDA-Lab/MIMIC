module fake_jpeg_16726_n_18 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_18);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_18;

wire n_13;
wire n_16;
wire n_10;
wire n_9;
wire n_14;
wire n_11;
wire n_17;
wire n_12;
wire n_15;

INVx6_ASAP7_75t_L g9 ( 
.A(n_6),
.Y(n_9)
);

AOI22xp33_ASAP7_75t_L g10 ( 
.A1(n_3),
.A2(n_7),
.B1(n_0),
.B2(n_1),
.Y(n_10)
);

NAND3xp33_ASAP7_75t_L g11 ( 
.A(n_6),
.B(n_8),
.C(n_0),
.Y(n_11)
);

INVx8_ASAP7_75t_L g12 ( 
.A(n_3),
.Y(n_12)
);

INVxp67_ASAP7_75t_L g13 ( 
.A(n_10),
.Y(n_13)
);

CKINVDCx16_ASAP7_75t_R g15 ( 
.A(n_13),
.Y(n_15)
);

OAI22xp5_ASAP7_75t_SL g14 ( 
.A1(n_9),
.A2(n_1),
.B1(n_2),
.B2(n_4),
.Y(n_14)
);

OAI22xp5_ASAP7_75t_SL g16 ( 
.A1(n_15),
.A2(n_9),
.B1(n_12),
.B2(n_14),
.Y(n_16)
);

AOI31xp67_ASAP7_75t_L g17 ( 
.A1(n_16),
.A2(n_9),
.A3(n_15),
.B(n_12),
.Y(n_17)
);

AOI322xp5_ASAP7_75t_L g18 ( 
.A1(n_17),
.A2(n_2),
.A3(n_4),
.B1(n_5),
.B2(n_11),
.C1(n_12),
.C2(n_9),
.Y(n_18)
);


endmodule