module fake_jpeg_20973_n_255 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_255);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_255;

wire n_159;
wire n_117;
wire n_253;
wire n_229;
wire n_144;
wire n_225;
wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_180;
wire n_245;
wire n_147;
wire n_158;
wire n_73;
wire n_14;
wire n_152;
wire n_19;
wire n_182;
wire n_59;
wire n_84;
wire n_98;
wire n_251;
wire n_252;
wire n_178;
wire n_228;
wire n_231;
wire n_166;
wire n_203;
wire n_65;
wire n_110;
wire n_134;
wire n_191;
wire n_193;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_127;
wire n_154;
wire n_205;
wire n_28;
wire n_38;
wire n_26;
wire n_181;
wire n_88;
wire n_116;
wire n_126;
wire n_114;
wire n_74;
wire n_137;
wire n_220;
wire n_31;
wire n_155;
wire n_207;
wire n_238;
wire n_235;
wire n_29;
wire n_103;
wire n_50;
wire n_150;
wire n_236;
wire n_160;
wire n_15;
wire n_124;
wire n_141;
wire n_194;
wire n_13;
wire n_175;
wire n_187;
wire n_57;
wire n_21;
wire n_223;
wire n_234;
wire n_171;
wire n_23;
wire n_119;
wire n_69;
wire n_27;
wire n_201;
wire n_195;
wire n_83;
wire n_179;
wire n_40;
wire n_250;
wire n_71;
wire n_80;
wire n_125;
wire n_185;
wire n_81;
wire n_204;
wire n_224;
wire n_129;
wire n_109;
wire n_113;
wire n_148;
wire n_248;
wire n_30;
wire n_168;
wire n_106;
wire n_111;
wire n_197;
wire n_186;
wire n_44;
wire n_24;
wire n_143;
wire n_202;
wire n_25;
wire n_17;
wire n_75;
wire n_122;
wire n_246;
wire n_37;
wire n_233;
wire n_102;
wire n_99;
wire n_121;
wire n_130;
wire n_70;
wire n_219;
wire n_177;
wire n_196;
wire n_66;
wire n_142;
wire n_85;
wire n_163;
wire n_77;
wire n_136;
wire n_61;
wire n_45;
wire n_139;
wire n_254;
wire n_172;
wire n_173;
wire n_244;
wire n_232;
wire n_78;
wire n_165;
wire n_20;
wire n_18;
wire n_145;
wire n_241;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_214;
wire n_58;
wire n_41;
wire n_128;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_218;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_239;
wire n_164;
wire n_243;
wire n_89;
wire n_146;
wire n_104;
wire n_215;
wire n_131;
wire n_56;
wire n_212;
wire n_240;
wire n_211;
wire n_230;
wire n_183;
wire n_79;
wire n_162;
wire n_170;
wire n_12;
wire n_132;
wire n_133;
wire n_249;
wire n_67;
wire n_216;
wire n_217;
wire n_184;
wire n_53;
wire n_33;
wire n_54;
wire n_93;
wire n_91;
wire n_227;
wire n_161;
wire n_209;
wire n_208;
wire n_22;
wire n_138;
wire n_101;
wire n_226;
wire n_210;
wire n_35;
wire n_48;
wire n_149;
wire n_157;
wire n_87;
wire n_46;
wire n_247;
wire n_200;
wire n_86;
wire n_156;
wire n_192;
wire n_115;
wire n_123;
wire n_176;
wire n_199;
wire n_112;
wire n_222;
wire n_95;
wire n_221;
wire n_151;
wire n_97;
wire n_169;
wire n_242;
wire n_153;
wire n_213;
wire n_135;
wire n_189;
wire n_237;
wire n_36;
wire n_188;
wire n_62;
wire n_167;
wire n_174;
wire n_198;
wire n_120;
wire n_190;
wire n_43;
wire n_32;
wire n_100;
wire n_118;
wire n_82;
wire n_140;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_0),
.Y(n_12)
);

CKINVDCx20_ASAP7_75t_R g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx5_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

INVx2_ASAP7_75t_L g15 ( 
.A(n_8),
.Y(n_15)
);

INVx1_ASAP7_75t_L g16 ( 
.A(n_4),
.Y(n_16)
);

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_3),
.Y(n_17)
);

CKINVDCx20_ASAP7_75t_R g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_7),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_3),
.Y(n_20)
);

BUFx3_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_11),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_3),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_1),
.Y(n_24)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_15),
.B(n_11),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_28),
.Y(n_37)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_23),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_26),
.Y(n_36)
);

INVx6_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

INVx8_ASAP7_75t_L g42 ( 
.A(n_27),
.Y(n_42)
);

INVx2_ASAP7_75t_SL g28 ( 
.A(n_23),
.Y(n_28)
);

INVx3_ASAP7_75t_L g29 ( 
.A(n_15),
.Y(n_29)
);

INVx2_ASAP7_75t_L g35 ( 
.A(n_29),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_16),
.Y(n_30)
);

NOR2xp33_ASAP7_75t_L g40 ( 
.A(n_30),
.B(n_31),
.Y(n_40)
);

INVx3_ASAP7_75t_L g31 ( 
.A(n_15),
.Y(n_31)
);

INVx2_ASAP7_75t_L g32 ( 
.A(n_23),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g38 ( 
.A(n_32),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_22),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_33),
.Y(n_34)
);

CKINVDCx5p33_ASAP7_75t_R g39 ( 
.A(n_30),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_20),
.Y(n_54)
);

INVx4_ASAP7_75t_L g41 ( 
.A(n_26),
.Y(n_41)
);

INVx3_ASAP7_75t_L g47 ( 
.A(n_41),
.Y(n_47)
);

INVx4_ASAP7_75t_L g43 ( 
.A(n_26),
.Y(n_43)
);

INVx1_ASAP7_75t_L g45 ( 
.A(n_43),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g44 ( 
.A(n_37),
.B(n_30),
.Y(n_44)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_44),
.B(n_59),
.Y(n_69)
);

HAxp5_ASAP7_75t_SL g46 ( 
.A(n_39),
.B(n_25),
.CON(n_46),
.SN(n_46)
);

AOI22xp5_ASAP7_75t_SL g74 ( 
.A1(n_46),
.A2(n_12),
.B1(n_13),
.B2(n_17),
.Y(n_74)
);

INVx3_ASAP7_75t_L g48 ( 
.A(n_35),
.Y(n_48)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_48),
.Y(n_61)
);

AND2x2_ASAP7_75t_L g49 ( 
.A(n_37),
.B(n_25),
.Y(n_49)
);

OAI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_49),
.A2(n_54),
.B(n_58),
.Y(n_70)
);

AOI22xp33_ASAP7_75t_L g50 ( 
.A1(n_39),
.A2(n_32),
.B1(n_27),
.B2(n_28),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g68 ( 
.A1(n_50),
.A2(n_56),
.B1(n_43),
.B2(n_41),
.Y(n_68)
);

HB1xp67_ASAP7_75t_L g51 ( 
.A(n_39),
.Y(n_51)
);

INVx1_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

OAI22xp5_ASAP7_75t_SL g52 ( 
.A1(n_37),
.A2(n_32),
.B1(n_27),
.B2(n_31),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g62 ( 
.A1(n_52),
.A2(n_55),
.B1(n_28),
.B2(n_34),
.Y(n_62)
);

INVx1_ASAP7_75t_L g53 ( 
.A(n_40),
.Y(n_53)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_53),
.Y(n_65)
);

OAI22xp5_ASAP7_75t_L g55 ( 
.A1(n_40),
.A2(n_27),
.B1(n_31),
.B2(n_29),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g56 ( 
.A1(n_35),
.A2(n_27),
.B1(n_28),
.B2(n_18),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_36),
.Y(n_57)
);

INVx4_ASAP7_75t_L g66 ( 
.A(n_57),
.Y(n_66)
);

OA22x2_ASAP7_75t_L g58 ( 
.A1(n_34),
.A2(n_28),
.B1(n_31),
.B2(n_29),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_40),
.B(n_26),
.Y(n_59)
);

NAND2xp5_ASAP7_75t_L g60 ( 
.A(n_35),
.B(n_26),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_60),
.B(n_42),
.Y(n_73)
);

OAI22xp5_ASAP7_75t_SL g87 ( 
.A1(n_62),
.A2(n_64),
.B1(n_43),
.B2(n_65),
.Y(n_87)
);

INVx2_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_63),
.Y(n_94)
);

OAI22xp5_ASAP7_75t_SL g67 ( 
.A1(n_53),
.A2(n_34),
.B1(n_35),
.B2(n_29),
.Y(n_67)
);

AOI22xp5_ASAP7_75t_L g80 ( 
.A1(n_67),
.A2(n_68),
.B1(n_55),
.B2(n_52),
.Y(n_80)
);

INVx2_ASAP7_75t_L g71 ( 
.A(n_48),
.Y(n_71)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_71),
.Y(n_91)
);

INVx3_ASAP7_75t_L g72 ( 
.A(n_47),
.Y(n_72)
);

CKINVDCx14_ASAP7_75t_R g81 ( 
.A(n_72),
.Y(n_81)
);

AND2x2_ASAP7_75t_L g90 ( 
.A(n_73),
.B(n_74),
.Y(n_90)
);

AOI22xp33_ASAP7_75t_SL g75 ( 
.A1(n_47),
.A2(n_43),
.B1(n_41),
.B2(n_42),
.Y(n_75)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_75),
.A2(n_76),
.B1(n_42),
.B2(n_57),
.Y(n_95)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_51),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_60),
.Y(n_77)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_77),
.Y(n_83)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_47),
.Y(n_78)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_78),
.Y(n_84)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_57),
.Y(n_79)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_79),
.Y(n_88)
);

AOI22xp5_ASAP7_75t_L g98 ( 
.A1(n_80),
.A2(n_85),
.B1(n_86),
.B2(n_87),
.Y(n_98)
);

MAJIxp5_ASAP7_75t_L g82 ( 
.A(n_69),
.B(n_49),
.C(n_44),
.Y(n_82)
);

MAJIxp5_ASAP7_75t_L g100 ( 
.A(n_82),
.B(n_93),
.C(n_85),
.Y(n_100)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_65),
.A2(n_49),
.B1(n_59),
.B2(n_54),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_L g86 ( 
.A1(n_62),
.A2(n_49),
.B1(n_58),
.B2(n_43),
.Y(n_86)
);

AOI21xp5_ASAP7_75t_L g89 ( 
.A1(n_70),
.A2(n_45),
.B(n_58),
.Y(n_89)
);

OAI21xp5_ASAP7_75t_SL g105 ( 
.A1(n_89),
.A2(n_96),
.B(n_90),
.Y(n_105)
);

AOI22xp5_ASAP7_75t_L g92 ( 
.A1(n_69),
.A2(n_58),
.B1(n_42),
.B2(n_41),
.Y(n_92)
);

NAND2xp5_ASAP7_75t_L g112 ( 
.A(n_92),
.B(n_86),
.Y(n_112)
);

MAJIxp5_ASAP7_75t_L g93 ( 
.A(n_70),
.B(n_58),
.C(n_45),
.Y(n_93)
);

OAI22xp33_ASAP7_75t_SL g99 ( 
.A1(n_95),
.A2(n_66),
.B1(n_79),
.B2(n_42),
.Y(n_99)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_67),
.Y(n_96)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_96),
.Y(n_108)
);

AOI21xp5_ASAP7_75t_L g97 ( 
.A1(n_90),
.A2(n_64),
.B(n_61),
.Y(n_97)
);

OAI21xp5_ASAP7_75t_L g136 ( 
.A1(n_97),
.A2(n_105),
.B(n_111),
.Y(n_136)
);

AOI22xp5_ASAP7_75t_L g132 ( 
.A1(n_99),
.A2(n_112),
.B1(n_91),
.B2(n_66),
.Y(n_132)
);

XNOR2xp5_ASAP7_75t_L g124 ( 
.A(n_100),
.B(n_102),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_SL g101 ( 
.A(n_83),
.B(n_92),
.Y(n_101)
);

NAND2xp5_ASAP7_75t_L g117 ( 
.A(n_101),
.B(n_109),
.Y(n_117)
);

XOR2xp5_ASAP7_75t_L g102 ( 
.A(n_82),
.B(n_74),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g103 ( 
.A(n_84),
.Y(n_103)
);

OR2x2_ASAP7_75t_L g128 ( 
.A(n_103),
.B(n_115),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g104 ( 
.A(n_83),
.B(n_72),
.Y(n_104)
);

NOR2xp33_ASAP7_75t_SL g118 ( 
.A(n_104),
.B(n_78),
.Y(n_118)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_91),
.Y(n_106)
);

INVx3_ASAP7_75t_L g133 ( 
.A(n_106),
.Y(n_133)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_81),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_L g120 ( 
.A(n_107),
.B(n_113),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_87),
.B(n_71),
.Y(n_109)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_84),
.Y(n_110)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_110),
.Y(n_116)
);

OAI21xp5_ASAP7_75t_SL g111 ( 
.A1(n_89),
.A2(n_19),
.B(n_16),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g113 ( 
.A(n_90),
.B(n_38),
.Y(n_113)
);

NAND2xp5_ASAP7_75t_SL g114 ( 
.A(n_93),
.B(n_80),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g127 ( 
.A(n_114),
.B(n_61),
.Y(n_127)
);

NOR2xp33_ASAP7_75t_L g115 ( 
.A(n_94),
.B(n_63),
.Y(n_115)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_118),
.Y(n_141)
);

INVx1_ASAP7_75t_L g119 ( 
.A(n_115),
.Y(n_119)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_119),
.Y(n_144)
);

MAJIxp5_ASAP7_75t_L g121 ( 
.A(n_100),
.B(n_94),
.C(n_88),
.Y(n_121)
);

MAJIxp5_ASAP7_75t_L g146 ( 
.A(n_121),
.B(n_38),
.C(n_33),
.Y(n_146)
);

INVx1_ASAP7_75t_L g122 ( 
.A(n_110),
.Y(n_122)
);

INVx1_ASAP7_75t_L g147 ( 
.A(n_122),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_108),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_123),
.B(n_126),
.Y(n_150)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_108),
.Y(n_125)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_125),
.Y(n_153)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_106),
.Y(n_126)
);

OAI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_127),
.A2(n_132),
.B1(n_36),
.B2(n_38),
.Y(n_152)
);

CKINVDCx20_ASAP7_75t_R g129 ( 
.A(n_103),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_129),
.B(n_130),
.Y(n_158)
);

INVx3_ASAP7_75t_SL g130 ( 
.A(n_107),
.Y(n_130)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_102),
.B(n_88),
.Y(n_131)
);

XOR2xp5_ASAP7_75t_L g154 ( 
.A(n_131),
.B(n_14),
.Y(n_154)
);

INVx2_ASAP7_75t_L g134 ( 
.A(n_107),
.Y(n_134)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_134),
.Y(n_149)
);

OAI22xp5_ASAP7_75t_SL g135 ( 
.A1(n_98),
.A2(n_38),
.B1(n_33),
.B2(n_36),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g138 ( 
.A1(n_135),
.A2(n_109),
.B1(n_101),
.B2(n_112),
.Y(n_138)
);

OAI21xp5_ASAP7_75t_L g137 ( 
.A1(n_105),
.A2(n_18),
.B(n_13),
.Y(n_137)
);

OAI21xp5_ASAP7_75t_L g143 ( 
.A1(n_137),
.A2(n_20),
.B(n_18),
.Y(n_143)
);

OAI22xp5_ASAP7_75t_SL g178 ( 
.A1(n_138),
.A2(n_139),
.B1(n_140),
.B2(n_142),
.Y(n_178)
);

AOI22xp5_ASAP7_75t_L g139 ( 
.A1(n_135),
.A2(n_114),
.B1(n_98),
.B2(n_113),
.Y(n_139)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_117),
.A2(n_119),
.B1(n_125),
.B2(n_132),
.Y(n_140)
);

AOI22xp5_ASAP7_75t_L g142 ( 
.A1(n_117),
.A2(n_111),
.B1(n_97),
.B2(n_33),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g163 ( 
.A(n_143),
.B(n_160),
.Y(n_163)
);

XOR2xp5_ASAP7_75t_SL g145 ( 
.A(n_136),
.B(n_10),
.Y(n_145)
);

AOI22xp33_ASAP7_75t_SL g162 ( 
.A1(n_145),
.A2(n_141),
.B1(n_144),
.B2(n_149),
.Y(n_162)
);

MAJIxp5_ASAP7_75t_L g166 ( 
.A(n_146),
.B(n_155),
.C(n_156),
.Y(n_166)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_136),
.A2(n_38),
.B1(n_36),
.B2(n_33),
.Y(n_148)
);

AOI22xp5_ASAP7_75t_L g164 ( 
.A1(n_148),
.A2(n_152),
.B1(n_153),
.B2(n_147),
.Y(n_164)
);

XNOR2xp5_ASAP7_75t_SL g151 ( 
.A(n_124),
.B(n_14),
.Y(n_151)
);

XNOR2xp5_ASAP7_75t_L g171 ( 
.A(n_151),
.B(n_154),
.Y(n_171)
);

XNOR2xp5_ASAP7_75t_SL g155 ( 
.A(n_124),
.B(n_14),
.Y(n_155)
);

MAJIxp5_ASAP7_75t_L g156 ( 
.A(n_121),
.B(n_131),
.C(n_116),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_SL g157 ( 
.A(n_137),
.B(n_128),
.Y(n_157)
);

NAND2xp5_ASAP7_75t_SL g173 ( 
.A(n_157),
.B(n_12),
.Y(n_173)
);

XOR2xp5_ASAP7_75t_L g159 ( 
.A(n_120),
.B(n_21),
.Y(n_159)
);

MAJIxp5_ASAP7_75t_L g172 ( 
.A(n_159),
.B(n_122),
.C(n_116),
.Y(n_172)
);

AOI22xp5_ASAP7_75t_L g160 ( 
.A1(n_130),
.A2(n_36),
.B1(n_24),
.B2(n_19),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_150),
.B(n_134),
.Y(n_161)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_161),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_L g184 ( 
.A1(n_162),
.A2(n_143),
.B1(n_154),
.B2(n_151),
.Y(n_184)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_164),
.Y(n_191)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_158),
.Y(n_165)
);

INVx1_ASAP7_75t_L g192 ( 
.A(n_165),
.Y(n_192)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_140),
.Y(n_167)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_167),
.Y(n_197)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_160),
.Y(n_168)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_168),
.B(n_169),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_138),
.B(n_128),
.Y(n_169)
);

CKINVDCx16_ASAP7_75t_R g170 ( 
.A(n_142),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_170),
.B(n_174),
.Y(n_182)
);

XOR2xp5_ASAP7_75t_L g187 ( 
.A(n_172),
.B(n_14),
.Y(n_187)
);

CKINVDCx14_ASAP7_75t_R g183 ( 
.A(n_173),
.Y(n_183)
);

NAND2xp5_ASAP7_75t_SL g174 ( 
.A(n_146),
.B(n_133),
.Y(n_174)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_148),
.Y(n_175)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_175),
.B(n_176),
.Y(n_181)
);

INVx8_ASAP7_75t_L g176 ( 
.A(n_145),
.Y(n_176)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_156),
.B(n_133),
.C(n_22),
.Y(n_177)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_177),
.B(n_22),
.C(n_24),
.Y(n_188)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_159),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_179),
.B(n_21),
.Y(n_195)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_139),
.A2(n_10),
.B1(n_1),
.B2(n_2),
.Y(n_180)
);

OAI22xp5_ASAP7_75t_SL g185 ( 
.A1(n_180),
.A2(n_24),
.B1(n_19),
.B2(n_16),
.Y(n_185)
);

XOR2xp5_ASAP7_75t_L g201 ( 
.A(n_184),
.B(n_186),
.Y(n_201)
);

INVx1_ASAP7_75t_L g210 ( 
.A(n_185),
.Y(n_210)
);

XNOR2xp5_ASAP7_75t_SL g186 ( 
.A(n_171),
.B(n_155),
.Y(n_186)
);

XOR2xp5_ASAP7_75t_L g204 ( 
.A(n_187),
.B(n_178),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g202 ( 
.A(n_188),
.B(n_193),
.C(n_196),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_177),
.B(n_22),
.C(n_20),
.Y(n_193)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_165),
.B(n_21),
.Y(n_194)
);

AOI21xp5_ASAP7_75t_L g209 ( 
.A1(n_194),
.A2(n_0),
.B(n_1),
.Y(n_209)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_195),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g196 ( 
.A(n_166),
.B(n_172),
.C(n_171),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_SL g198 ( 
.A1(n_190),
.A2(n_180),
.B1(n_169),
.B2(n_168),
.Y(n_198)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_198),
.B(n_200),
.Y(n_211)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_196),
.B(n_166),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_SL g203 ( 
.A1(n_190),
.A2(n_163),
.B1(n_164),
.B2(n_176),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g220 ( 
.A(n_203),
.B(n_208),
.Y(n_220)
);

XOR2xp5_ASAP7_75t_L g221 ( 
.A(n_204),
.B(n_205),
.Y(n_221)
);

XOR2xp5_ASAP7_75t_L g205 ( 
.A(n_186),
.B(n_178),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g206 ( 
.A(n_187),
.B(n_163),
.Y(n_206)
);

XNOR2xp5_ASAP7_75t_L g214 ( 
.A(n_206),
.B(n_209),
.Y(n_214)
);

OR2x2_ASAP7_75t_L g207 ( 
.A(n_181),
.B(n_17),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g213 ( 
.A1(n_207),
.A2(n_183),
.B1(n_192),
.B2(n_189),
.Y(n_213)
);

INVx2_ASAP7_75t_L g208 ( 
.A(n_194),
.Y(n_208)
);

MAJIxp5_ASAP7_75t_L g212 ( 
.A(n_202),
.B(n_182),
.C(n_191),
.Y(n_212)
);

OR2x2_ASAP7_75t_L g223 ( 
.A(n_212),
.B(n_215),
.Y(n_223)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_213),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_207),
.B(n_197),
.Y(n_215)
);

NOR2xp33_ASAP7_75t_L g216 ( 
.A(n_199),
.B(n_193),
.Y(n_216)
);

NOR2xp33_ASAP7_75t_L g229 ( 
.A(n_216),
.B(n_218),
.Y(n_229)
);

AOI21xp5_ASAP7_75t_L g217 ( 
.A1(n_202),
.A2(n_188),
.B(n_185),
.Y(n_217)
);

NAND2xp5_ASAP7_75t_SL g225 ( 
.A(n_217),
.B(n_219),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_210),
.B(n_204),
.Y(n_218)
);

AOI21xp5_ASAP7_75t_L g219 ( 
.A1(n_205),
.A2(n_0),
.B(n_1),
.Y(n_219)
);

XNOR2xp5_ASAP7_75t_L g222 ( 
.A(n_214),
.B(n_206),
.Y(n_222)
);

OR2x2_ASAP7_75t_L g236 ( 
.A(n_222),
.B(n_226),
.Y(n_236)
);

NOR2xp33_ASAP7_75t_L g226 ( 
.A(n_211),
.B(n_201),
.Y(n_226)
);

XOR2xp5_ASAP7_75t_L g227 ( 
.A(n_221),
.B(n_201),
.Y(n_227)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_227),
.B(n_231),
.Y(n_235)
);

XNOR2xp5_ASAP7_75t_L g228 ( 
.A(n_214),
.B(n_21),
.Y(n_228)
);

NOR2xp33_ASAP7_75t_L g233 ( 
.A(n_228),
.B(n_230),
.Y(n_233)
);

NOR2xp33_ASAP7_75t_SL g230 ( 
.A(n_212),
.B(n_17),
.Y(n_230)
);

XNOR2xp5_ASAP7_75t_L g231 ( 
.A(n_221),
.B(n_0),
.Y(n_231)
);

AO21x1_ASAP7_75t_L g232 ( 
.A1(n_229),
.A2(n_220),
.B(n_4),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g241 ( 
.A1(n_232),
.A2(n_234),
.B(n_237),
.Y(n_241)
);

NOR2xp33_ASAP7_75t_SL g234 ( 
.A(n_223),
.B(n_13),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g237 ( 
.A1(n_224),
.A2(n_12),
.B(n_4),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g238 ( 
.A(n_225),
.B(n_2),
.C(n_5),
.Y(n_238)
);

NAND2xp5_ASAP7_75t_SL g242 ( 
.A(n_238),
.B(n_2),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_SL g239 ( 
.A1(n_225),
.A2(n_2),
.B(n_5),
.Y(n_239)
);

AOI21xp5_ASAP7_75t_SL g243 ( 
.A1(n_239),
.A2(n_5),
.B(n_6),
.Y(n_243)
);

XNOR2xp5_ASAP7_75t_L g240 ( 
.A(n_235),
.B(n_229),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_240),
.B(n_242),
.Y(n_246)
);

AOI21xp33_ASAP7_75t_L g245 ( 
.A1(n_243),
.A2(n_234),
.B(n_7),
.Y(n_245)
);

XNOR2xp5_ASAP7_75t_L g244 ( 
.A(n_233),
.B(n_5),
.Y(n_244)
);

NOR2xp67_ASAP7_75t_SL g247 ( 
.A(n_244),
.B(n_6),
.Y(n_247)
);

AO21x2_ASAP7_75t_L g248 ( 
.A1(n_245),
.A2(n_247),
.B(n_241),
.Y(n_248)
);

AOI21x1_ASAP7_75t_L g250 ( 
.A1(n_248),
.A2(n_249),
.B(n_6),
.Y(n_250)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_246),
.B(n_236),
.C(n_7),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g251 ( 
.A(n_250),
.B(n_6),
.C(n_7),
.Y(n_251)
);

NAND2xp5_ASAP7_75t_SL g252 ( 
.A(n_251),
.B(n_8),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_252),
.B(n_8),
.C(n_9),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g254 ( 
.A1(n_253),
.A2(n_8),
.B(n_9),
.Y(n_254)
);

AO21x1_ASAP7_75t_L g255 ( 
.A1(n_254),
.A2(n_9),
.B(n_232),
.Y(n_255)
);


endmodule