module real_aes_6573_n_101 (n_17, n_28, n_76, n_56, n_34, n_98, n_90, n_82, n_65, n_47, n_74, n_58, n_32, n_30, n_51, n_27, n_61, n_29, n_20, n_52, n_57, n_64, n_66, n_18, n_21, n_31, n_8, n_10, n_83, n_22, n_3, n_41, n_75, n_19, n_71, n_40, n_49, n_91, n_100, n_43, n_96, n_54, n_35, n_42, n_99, n_15, n_9, n_23, n_72, n_95, n_44, n_7, n_4, n_80, n_6, n_12, n_68, n_79, n_69, n_46, n_59, n_25, n_73, n_77, n_81, n_48, n_37, n_97, n_70, n_50, n_89, n_26, n_86, n_93, n_13, n_24, n_2, n_55, n_62, n_84, n_67, n_92, n_33, n_88, n_14, n_11, n_85, n_16, n_94, n_39, n_5, n_45, n_60, n_38, n_87, n_0, n_78, n_63, n_1, n_53, n_36, n_101);
input n_17;
input n_28;
input n_76;
input n_56;
input n_34;
input n_98;
input n_90;
input n_82;
input n_65;
input n_47;
input n_74;
input n_58;
input n_32;
input n_30;
input n_51;
input n_27;
input n_61;
input n_29;
input n_20;
input n_52;
input n_57;
input n_64;
input n_66;
input n_18;
input n_21;
input n_31;
input n_8;
input n_10;
input n_83;
input n_22;
input n_3;
input n_41;
input n_75;
input n_19;
input n_71;
input n_40;
input n_49;
input n_91;
input n_100;
input n_43;
input n_96;
input n_54;
input n_35;
input n_42;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_95;
input n_44;
input n_7;
input n_4;
input n_80;
input n_6;
input n_12;
input n_68;
input n_79;
input n_69;
input n_46;
input n_59;
input n_25;
input n_73;
input n_77;
input n_81;
input n_48;
input n_37;
input n_97;
input n_70;
input n_50;
input n_89;
input n_26;
input n_86;
input n_93;
input n_13;
input n_24;
input n_2;
input n_55;
input n_62;
input n_84;
input n_67;
input n_92;
input n_33;
input n_88;
input n_14;
input n_11;
input n_85;
input n_16;
input n_94;
input n_39;
input n_5;
input n_45;
input n_60;
input n_38;
input n_87;
input n_0;
input n_78;
input n_63;
input n_1;
input n_53;
input n_36;
output n_101;
wire n_480;
wire n_113;
wire n_476;
wire n_599;
wire n_187;
wire n_436;
wire n_684;
wire n_257;
wire n_390;
wire n_185;
wire n_285;
wire n_624;
wire n_618;
wire n_522;
wire n_485;
wire n_222;
wire n_631;
wire n_503;
wire n_287;
wire n_357;
wire n_635;
wire n_386;
wire n_673;
wire n_518;
wire n_254;
wire n_207;
wire n_665;
wire n_667;
wire n_577;
wire n_580;
wire n_469;
wire n_181;
wire n_362;
wire n_124;
wire n_191;
wire n_209;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_299;
wire n_657;
wire n_322;
wire n_328;
wire n_718;
wire n_318;
wire n_355;
wire n_239;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_112;
wire n_319;
wire n_421;
wire n_364;
wire n_555;
wire n_329;
wire n_132;
wire n_131;
wire n_144;
wire n_461;
wire n_169;
wire n_242;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_429;
wire n_172;
wire n_448;
wire n_556;
wire n_341;
wire n_545;
wire n_593;
wire n_232;
wire n_460;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_537;
wire n_320;
wire n_551;
wire n_666;
wire n_560;
wire n_260;
wire n_660;
wire n_594;
wire n_186;
wire n_138;
wire n_696;
wire n_704;
wire n_453;
wire n_379;
wire n_374;
wire n_647;
wire n_235;
wire n_399;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_245;
wire n_161;
wire n_189;
wire n_271;
wire n_489;
wire n_427;
wire n_548;
wire n_678;
wire n_145;
wire n_415;
wire n_572;
wire n_227;
wire n_564;
wire n_519;
wire n_638;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_512;
wire n_395;
wire n_332;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_116;
wire n_625;
wire n_462;
wire n_289;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_716;
wire n_213;
wire n_356;
wire n_478;
wire n_584;
wire n_408;
wire n_553;
wire n_184;
wire n_372;
wire n_528;
wire n_578;
wire n_202;
wire n_495;
wire n_370;
wire n_384;
wire n_121;
wire n_352;
wire n_125;
wire n_216;
wire n_467;
wire n_327;
wire n_106;
wire n_559;
wire n_466;
wire n_636;
wire n_263;
wire n_477;
wire n_515;
wire n_230;
wire n_680;
wire n_595;
wire n_248;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_174;
wire n_570;
wire n_675;
wire n_530;
wire n_104;
wire n_535;
wire n_732;
wire n_211;
wire n_281;
wire n_496;
wire n_693;
wire n_173;
wire n_468;
wire n_234;
wire n_284;
wire n_153;
wire n_316;
wire n_532;
wire n_656;
wire n_178;
wire n_409;
wire n_298;
wire n_523;
wire n_439;
wire n_576;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_297;
wire n_383;
wire n_529;
wire n_119;
wire n_504;
wire n_725;
wire n_310;
wire n_455;
wire n_164;
wire n_671;
wire n_231;
wire n_102;
wire n_547;
wire n_659;
wire n_634;
wire n_682;
wire n_454;
wire n_122;
wire n_565;
wire n_443;
wire n_608;
wire n_534;
wire n_708;
wire n_141;
wire n_128;
wire n_111;
wire n_167;
wire n_457;
wire n_179;
wire n_129;
wire n_345;
wire n_304;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_278;
wire n_236;
wire n_664;
wire n_367;
wire n_267;
wire n_218;
wire n_737;
wire n_581;
wire n_610;
wire n_204;
wire n_620;
wire n_582;
wire n_641;
wire n_722;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_425;
wire n_609;
wire n_331;
wire n_182;
wire n_417;
wire n_363;
wire n_449;
wire n_607;
wire n_323;
wire n_690;
wire n_629;
wire n_199;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_142;
wire n_561;
wire n_437;
wire n_223;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_655;
wire n_654;
wire n_505;
wire n_502;
wire n_527;
wire n_434;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_406;
wire n_426;
wire n_244;
wire n_118;
wire n_139;
wire n_733;
wire n_402;
wire n_617;
wire n_552;
wire n_602;
wire n_171;
wire n_658;
wire n_676;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_146;
wire n_432;
wire n_226;
wire n_255;
wire n_286;
wire n_416;
wire n_410;
wire n_120;
wire n_490;
wire n_261;
wire n_238;
wire n_619;
wire n_391;
wire n_360;
wire n_695;
wire n_685;
wire n_165;
wire n_361;
wire n_632;
wire n_246;
wire n_176;
wire n_412;
wire n_163;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_488;
wire n_501;
wire n_251;
wire n_642;
wire n_613;
wire n_220;
wire n_387;
wire n_197;
wire n_296;
wire n_702;
wire n_256;
wire n_302;
wire n_464;
wire n_351;
wire n_126;
wire n_200;
wire n_604;
wire n_115;
wire n_734;
wire n_110;
wire n_392;
wire n_562;
wire n_150;
wire n_147;
wire n_404;
wire n_288;
wire n_598;
wire n_713;
wire n_735;
wire n_728;
wire n_334;
wire n_274;
wire n_160;
wire n_303;
wire n_569;
wire n_563;
wire n_188;
wire n_269;
wire n_430;
wire n_568;
wire n_201;
wire n_413;
wire n_471;
wire n_306;
wire n_579;
wire n_158;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_193;
wire n_397;
wire n_293;
wire n_162;
wire n_358;
wire n_385;
wire n_275;
wire n_214;
wire n_649;
wire n_663;
wire n_588;
wire n_109;
wire n_536;
wire n_203;
wire n_707;
wire n_622;
wire n_470;
wire n_133;
wire n_494;
wire n_711;
wire n_377;
wire n_273;
wire n_723;
wire n_114;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_154;
wire n_127;
wire n_511;
wire n_484;
wire n_326;
wire n_492;
wire n_509;
wire n_407;
wire n_217;
wire n_419;
wire n_730;
wire n_643;
wire n_486;
wire n_411;
wire n_697;
wire n_291;
wire n_148;
wire n_481;
wire n_498;
wire n_691;
wire n_159;
wire n_108;
wire n_373;
wire n_648;
wire n_589;
wire n_628;
wire n_487;
wire n_233;
wire n_290;
wire n_365;
wire n_653;
wire n_526;
wire n_637;
wire n_155;
wire n_243;
wire n_692;
wire n_544;
wire n_268;
wire n_136;
wire n_157;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_229;
wire n_107;
wire n_482;
wire n_520;
wire n_679;
wire n_633;
wire n_149;
wire n_472;
wire n_452;
wire n_190;
wire n_262;
wire n_630;
wire n_689;
wire n_715;
wire n_134;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_195;
wire n_438;
wire n_300;
wire n_252;
wire n_314;
wire n_283;
wire n_249;
wire n_623;
wire n_446;
wire n_721;
wire n_221;
wire n_681;
wire n_156;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_183;
wire n_266;
wire n_712;
wire n_205;
wire n_433;
wire n_516;
wire n_177;
wire n_335;
wire n_313;
wire n_627;
wire n_739;
wire n_521;
wire n_140;
wire n_418;
wire n_422;
wire n_219;
wire n_524;
wire n_705;
wire n_180;
wire n_212;
wire n_210;
wire n_575;
wire n_325;
wire n_338;
wire n_479;
wire n_442;
wire n_698;
wire n_371;
wire n_740;
wire n_166;
wire n_103;
wire n_541;
wire n_224;
wire n_151;
wire n_546;
wire n_587;
wire n_639;
wire n_130;
wire n_253;
wire n_459;
wire n_558;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_152;
wire n_198;
wire n_228;
wire n_272;
wire n_196;
wire n_583;
wire n_347;
wire n_315;
wire n_414;
wire n_123;
wire n_279;
wire n_686;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_450;
wire n_117;
wire n_208;
wire n_215;
wire n_441;
wire n_135;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_474;
wire n_170;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_729;
wire n_168;
wire n_175;
wire n_241;
wire n_687;
wire n_646;
wire n_650;
wire n_710;
wire n_105;
wire n_294;
wire n_393;
wire n_258;
wire n_652;
wire n_206;
wire n_703;
wire n_307;
wire n_500;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_194;
wire n_137;
wire n_225;
wire n_424;
wire n_574;
wire n_337;
wire n_247;
wire n_240;
wire n_259;
wire n_143;
wire n_192;
wire n_475;
wire n_554;
wire n_264;
wire n_237;
wire n_668;
INVx1_ASAP7_75t_L g106 ( .A(n_0), .Y(n_106) );
A2O1A1Ixp33_ASAP7_75t_L g483 ( .A1(n_1), .A2(n_141), .B(n_144), .C(n_484), .Y(n_483) );
INVx1_ASAP7_75t_L g207 ( .A(n_2), .Y(n_207) );
AOI21xp5_ASAP7_75t_L g525 ( .A1(n_3), .A2(n_136), .B(n_526), .Y(n_525) );
NAND2xp5_ASAP7_75t_L g531 ( .A(n_4), .B(n_217), .Y(n_531) );
AOI21xp33_ASAP7_75t_L g218 ( .A1(n_5), .A2(n_136), .B(n_219), .Y(n_218) );
AND2x6_ASAP7_75t_L g141 ( .A(n_6), .B(n_142), .Y(n_141) );
AOI21xp5_ASAP7_75t_L g186 ( .A1(n_7), .A2(n_187), .B(n_188), .Y(n_186) );
NAND2xp5_ASAP7_75t_L g104 ( .A(n_8), .B(n_41), .Y(n_104) );
NOR2xp33_ASAP7_75t_L g121 ( .A(n_8), .B(n_41), .Y(n_121) );
OAI22xp5_ASAP7_75t_L g124 ( .A1(n_9), .A2(n_31), .B1(n_125), .B2(n_126), .Y(n_124) );
CKINVDCx20_ASAP7_75t_R g126 ( .A(n_9), .Y(n_126) );
INVx1_ASAP7_75t_L g466 ( .A(n_10), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g175 ( .A(n_11), .B(n_176), .Y(n_175) );
INVx1_ASAP7_75t_L g224 ( .A(n_12), .Y(n_224) );
NAND2xp5_ASAP7_75t_SL g487 ( .A(n_13), .B(n_177), .Y(n_487) );
INVx1_ASAP7_75t_L g162 ( .A(n_14), .Y(n_162) );
INVx1_ASAP7_75t_L g195 ( .A(n_15), .Y(n_195) );
A2O1A1Ixp33_ASAP7_75t_L g474 ( .A1(n_16), .A2(n_150), .B(n_196), .C(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_17), .B(n_217), .Y(n_477) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_18), .B(n_152), .Y(n_269) );
NAND2xp5_ASAP7_75t_SL g135 ( .A(n_19), .B(n_136), .Y(n_135) );
NAND2xp5_ASAP7_75t_L g566 ( .A(n_20), .B(n_567), .Y(n_566) );
A2O1A1Ixp33_ASAP7_75t_L g495 ( .A1(n_21), .A2(n_176), .B(n_210), .C(n_496), .Y(n_495) );
NAND2xp5_ASAP7_75t_L g245 ( .A(n_22), .B(n_217), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g520 ( .A(n_23), .B(n_177), .Y(n_520) );
A2O1A1Ixp33_ASAP7_75t_L g191 ( .A1(n_24), .A2(n_192), .B(n_194), .C(n_196), .Y(n_191) );
NAND2xp5_ASAP7_75t_SL g506 ( .A(n_25), .B(n_177), .Y(n_506) );
CKINVDCx16_ASAP7_75t_R g516 ( .A(n_26), .Y(n_516) );
INVx1_ASAP7_75t_L g505 ( .A(n_27), .Y(n_505) );
BUFx6f_ASAP7_75t_L g140 ( .A(n_28), .Y(n_140) );
CKINVDCx20_ASAP7_75t_R g482 ( .A(n_29), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g208 ( .A(n_30), .B(n_177), .Y(n_208) );
INVx1_ASAP7_75t_L g125 ( .A(n_31), .Y(n_125) );
INVx1_ASAP7_75t_L g563 ( .A(n_32), .Y(n_563) );
INVx1_ASAP7_75t_L g234 ( .A(n_33), .Y(n_234) );
INVx2_ASAP7_75t_L g139 ( .A(n_34), .Y(n_139) );
CKINVDCx20_ASAP7_75t_R g489 ( .A(n_35), .Y(n_489) );
A2O1A1Ixp33_ASAP7_75t_L g528 ( .A1(n_36), .A2(n_176), .B(n_225), .C(n_529), .Y(n_528) );
INVxp67_ASAP7_75t_L g564 ( .A(n_37), .Y(n_564) );
A2O1A1Ixp33_ASAP7_75t_L g143 ( .A1(n_38), .A2(n_141), .B(n_144), .C(n_147), .Y(n_143) );
A2O1A1Ixp33_ASAP7_75t_L g503 ( .A1(n_39), .A2(n_144), .B(n_504), .C(n_509), .Y(n_503) );
CKINVDCx14_ASAP7_75t_R g527 ( .A(n_40), .Y(n_527) );
INVx1_ASAP7_75t_L g232 ( .A(n_42), .Y(n_232) );
A2O1A1Ixp33_ASAP7_75t_L g464 ( .A1(n_43), .A2(n_154), .B(n_222), .C(n_465), .Y(n_464) );
NAND2xp5_ASAP7_75t_SL g268 ( .A(n_44), .B(n_177), .Y(n_268) );
CKINVDCx20_ASAP7_75t_R g511 ( .A(n_45), .Y(n_511) );
CKINVDCx20_ASAP7_75t_R g560 ( .A(n_46), .Y(n_560) );
INVx1_ASAP7_75t_L g494 ( .A(n_47), .Y(n_494) );
CKINVDCx16_ASAP7_75t_R g235 ( .A(n_48), .Y(n_235) );
NAND2xp5_ASAP7_75t_L g180 ( .A(n_49), .B(n_136), .Y(n_180) );
CKINVDCx20_ASAP7_75t_R g122 ( .A(n_50), .Y(n_122) );
AOI22xp5_ASAP7_75t_L g230 ( .A1(n_51), .A2(n_144), .B1(n_210), .B2(n_231), .Y(n_230) );
CKINVDCx20_ASAP7_75t_R g164 ( .A(n_52), .Y(n_164) );
CKINVDCx16_ASAP7_75t_R g203 ( .A(n_53), .Y(n_203) );
A2O1A1Ixp33_ASAP7_75t_L g221 ( .A1(n_54), .A2(n_222), .B(n_223), .C(n_225), .Y(n_221) );
CKINVDCx14_ASAP7_75t_R g463 ( .A(n_55), .Y(n_463) );
CKINVDCx20_ASAP7_75t_R g272 ( .A(n_56), .Y(n_272) );
INVx1_ASAP7_75t_L g220 ( .A(n_57), .Y(n_220) );
INVx1_ASAP7_75t_L g142 ( .A(n_58), .Y(n_142) );
INVx1_ASAP7_75t_L g161 ( .A(n_59), .Y(n_161) );
INVx1_ASAP7_75t_SL g530 ( .A(n_60), .Y(n_530) );
CKINVDCx20_ASAP7_75t_R g115 ( .A(n_61), .Y(n_115) );
NAND2xp5_ASAP7_75t_L g498 ( .A(n_62), .B(n_217), .Y(n_498) );
INVx1_ASAP7_75t_L g519 ( .A(n_63), .Y(n_519) );
A2O1A1Ixp33_ASAP7_75t_SL g242 ( .A1(n_64), .A2(n_152), .B(n_225), .C(n_243), .Y(n_242) );
INVxp67_ASAP7_75t_L g244 ( .A(n_65), .Y(n_244) );
INVx1_ASAP7_75t_L g109 ( .A(n_66), .Y(n_109) );
AOI21xp5_ASAP7_75t_L g461 ( .A1(n_67), .A2(n_136), .B(n_462), .Y(n_461) );
CKINVDCx20_ASAP7_75t_R g523 ( .A(n_68), .Y(n_523) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_69), .Y(n_237) );
AOI21xp5_ASAP7_75t_L g471 ( .A1(n_70), .A2(n_136), .B(n_472), .Y(n_471) );
INVx1_ASAP7_75t_L g265 ( .A(n_71), .Y(n_265) );
AOI21xp5_ASAP7_75t_L g558 ( .A1(n_72), .A2(n_187), .B(n_559), .Y(n_558) );
INVx1_ASAP7_75t_L g473 ( .A(n_73), .Y(n_473) );
CKINVDCx16_ASAP7_75t_R g502 ( .A(n_74), .Y(n_502) );
OAI22xp5_ASAP7_75t_SL g735 ( .A1(n_75), .A2(n_76), .B1(n_736), .B2(n_737), .Y(n_735) );
CKINVDCx20_ASAP7_75t_R g737 ( .A(n_75), .Y(n_737) );
CKINVDCx20_ASAP7_75t_R g736 ( .A(n_76), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g266 ( .A1(n_77), .A2(n_141), .B(n_144), .C(n_267), .Y(n_266) );
AOI21xp5_ASAP7_75t_L g492 ( .A1(n_78), .A2(n_136), .B(n_493), .Y(n_492) );
INVx1_ASAP7_75t_L g476 ( .A(n_79), .Y(n_476) );
AOI222xp33_ASAP7_75t_SL g123 ( .A1(n_80), .A2(n_124), .B1(n_127), .B2(n_724), .C1(n_725), .C2(n_729), .Y(n_123) );
NAND2xp5_ASAP7_75t_SL g148 ( .A(n_81), .B(n_149), .Y(n_148) );
INVx2_ASAP7_75t_L g159 ( .A(n_82), .Y(n_159) );
INVx1_ASAP7_75t_L g485 ( .A(n_83), .Y(n_485) );
NAND2xp5_ASAP7_75t_L g151 ( .A(n_84), .B(n_152), .Y(n_151) );
A2O1A1Ixp33_ASAP7_75t_L g205 ( .A1(n_85), .A2(n_141), .B(n_144), .C(n_206), .Y(n_205) );
NAND3xp33_ASAP7_75t_SL g105 ( .A(n_86), .B(n_106), .C(n_107), .Y(n_105) );
OR2x2_ASAP7_75t_L g118 ( .A(n_86), .B(n_119), .Y(n_118) );
INVx2_ASAP7_75t_L g453 ( .A(n_86), .Y(n_453) );
OR2x2_ASAP7_75t_L g723 ( .A(n_86), .B(n_120), .Y(n_723) );
A2O1A1Ixp33_ASAP7_75t_L g517 ( .A1(n_87), .A2(n_144), .B(n_518), .C(n_521), .Y(n_517) );
NAND2xp5_ASAP7_75t_L g226 ( .A(n_88), .B(n_170), .Y(n_226) );
CKINVDCx20_ASAP7_75t_R g213 ( .A(n_89), .Y(n_213) );
AOI22xp33_ASAP7_75t_L g101 ( .A1(n_90), .A2(n_102), .B1(n_110), .B2(n_739), .Y(n_101) );
A2O1A1Ixp33_ASAP7_75t_L g172 ( .A1(n_91), .A2(n_141), .B(n_144), .C(n_173), .Y(n_172) );
CKINVDCx20_ASAP7_75t_R g182 ( .A(n_92), .Y(n_182) );
INVx1_ASAP7_75t_L g241 ( .A(n_93), .Y(n_241) );
CKINVDCx16_ASAP7_75t_R g189 ( .A(n_94), .Y(n_189) );
NAND2xp5_ASAP7_75t_SL g174 ( .A(n_95), .B(n_149), .Y(n_174) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_96), .B(n_166), .Y(n_467) );
NAND2xp5_ASAP7_75t_L g198 ( .A(n_97), .B(n_166), .Y(n_198) );
NAND2xp5_ASAP7_75t_L g108 ( .A(n_98), .B(n_109), .Y(n_108) );
AOI21xp5_ASAP7_75t_L g239 ( .A1(n_99), .A2(n_136), .B(n_240), .Y(n_239) );
INVx2_ASAP7_75t_L g497 ( .A(n_100), .Y(n_497) );
INVx1_ASAP7_75t_SL g102 ( .A(n_103), .Y(n_102) );
CKINVDCx12_ASAP7_75t_R g740 ( .A(n_103), .Y(n_740) );
OR2x2_ASAP7_75t_L g103 ( .A(n_104), .B(n_105), .Y(n_103) );
AND2x2_ASAP7_75t_L g120 ( .A(n_106), .B(n_121), .Y(n_120) );
INVx1_ASAP7_75t_SL g107 ( .A(n_108), .Y(n_107) );
AOI22x1_ASAP7_75t_L g110 ( .A1(n_111), .A2(n_123), .B1(n_732), .B2(n_733), .Y(n_110) );
NOR2xp33_ASAP7_75t_L g111 ( .A(n_112), .B(n_116), .Y(n_111) );
INVx1_ASAP7_75t_SL g112 ( .A(n_113), .Y(n_112) );
INVx1_ASAP7_75t_SL g732 ( .A(n_113), .Y(n_732) );
BUFx2_ASAP7_75t_L g113 ( .A(n_114), .Y(n_113) );
INVx2_ASAP7_75t_L g114 ( .A(n_115), .Y(n_114) );
AOI21xp5_ASAP7_75t_L g733 ( .A1(n_116), .A2(n_734), .B(n_738), .Y(n_733) );
NOR2xp33_ASAP7_75t_SL g116 ( .A(n_117), .B(n_122), .Y(n_116) );
BUFx2_ASAP7_75t_L g117 ( .A(n_118), .Y(n_117) );
HB1xp67_ASAP7_75t_L g738 ( .A(n_118), .Y(n_738) );
NOR2x2_ASAP7_75t_L g731 ( .A(n_119), .B(n_453), .Y(n_731) );
INVx2_ASAP7_75t_L g119 ( .A(n_120), .Y(n_119) );
OR2x2_ASAP7_75t_L g452 ( .A(n_120), .B(n_453), .Y(n_452) );
INVx1_ASAP7_75t_L g724 ( .A(n_124), .Y(n_724) );
OAI22xp5_ASAP7_75t_SL g127 ( .A1(n_128), .A2(n_452), .B1(n_454), .B2(n_723), .Y(n_127) );
INVx2_ASAP7_75t_L g726 ( .A(n_128), .Y(n_726) );
AND2x2_ASAP7_75t_SL g128 ( .A(n_129), .B(n_421), .Y(n_128) );
NOR3xp33_ASAP7_75t_L g129 ( .A(n_130), .B(n_314), .C(n_387), .Y(n_129) );
OAI211xp5_ASAP7_75t_SL g130 ( .A1(n_131), .A2(n_199), .B(n_246), .C(n_298), .Y(n_130) );
INVxp67_ASAP7_75t_L g131 ( .A(n_132), .Y(n_131) );
AND2x2_ASAP7_75t_L g132 ( .A(n_133), .B(n_167), .Y(n_132) );
AND2x2_ASAP7_75t_L g262 ( .A(n_133), .B(n_263), .Y(n_262) );
INVx3_ASAP7_75t_L g281 ( .A(n_133), .Y(n_281) );
INVx2_ASAP7_75t_L g296 ( .A(n_133), .Y(n_296) );
INVx1_ASAP7_75t_L g326 ( .A(n_133), .Y(n_326) );
AND2x2_ASAP7_75t_L g376 ( .A(n_133), .B(n_297), .Y(n_376) );
AOI32xp33_ASAP7_75t_L g403 ( .A1(n_133), .A2(n_331), .A3(n_404), .B1(n_406), .B2(n_407), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_133), .B(n_252), .Y(n_409) );
AND2x2_ASAP7_75t_L g436 ( .A(n_133), .B(n_279), .Y(n_436) );
NOR2xp33_ASAP7_75t_L g444 ( .A(n_133), .B(n_445), .Y(n_444) );
OR2x6_ASAP7_75t_L g133 ( .A(n_134), .B(n_163), .Y(n_133) );
AOI21xp5_ASAP7_75t_SL g134 ( .A1(n_135), .A2(n_143), .B(n_156), .Y(n_134) );
BUFx2_ASAP7_75t_L g187 ( .A(n_136), .Y(n_187) );
AND2x4_ASAP7_75t_L g136 ( .A(n_137), .B(n_141), .Y(n_136) );
NAND2x1p5_ASAP7_75t_L g204 ( .A(n_137), .B(n_141), .Y(n_204) );
AND2x2_ASAP7_75t_L g137 ( .A(n_138), .B(n_140), .Y(n_137) );
INVx1_ASAP7_75t_L g508 ( .A(n_138), .Y(n_508) );
INVx1_ASAP7_75t_L g138 ( .A(n_139), .Y(n_138) );
INVx2_ASAP7_75t_L g145 ( .A(n_139), .Y(n_145) );
INVx1_ASAP7_75t_L g211 ( .A(n_139), .Y(n_211) );
INVx1_ASAP7_75t_L g146 ( .A(n_140), .Y(n_146) );
INVx3_ASAP7_75t_L g150 ( .A(n_140), .Y(n_150) );
INVx1_ASAP7_75t_L g152 ( .A(n_140), .Y(n_152) );
BUFx6f_ASAP7_75t_L g177 ( .A(n_140), .Y(n_177) );
BUFx6f_ASAP7_75t_L g193 ( .A(n_140), .Y(n_193) );
INVx4_ASAP7_75t_SL g197 ( .A(n_141), .Y(n_197) );
BUFx3_ASAP7_75t_L g509 ( .A(n_141), .Y(n_509) );
INVx5_ASAP7_75t_L g190 ( .A(n_144), .Y(n_190) );
AND2x6_ASAP7_75t_L g144 ( .A(n_145), .B(n_146), .Y(n_144) );
BUFx3_ASAP7_75t_L g155 ( .A(n_145), .Y(n_155) );
BUFx6f_ASAP7_75t_L g179 ( .A(n_145), .Y(n_179) );
AOI21xp5_ASAP7_75t_L g147 ( .A1(n_148), .A2(n_151), .B(n_153), .Y(n_147) );
O2A1O1Ixp33_ASAP7_75t_L g206 ( .A1(n_149), .A2(n_207), .B(n_208), .C(n_209), .Y(n_206) );
O2A1O1Ixp33_ASAP7_75t_L g504 ( .A1(n_149), .A2(n_505), .B(n_506), .C(n_507), .Y(n_504) );
OAI22xp33_ASAP7_75t_L g562 ( .A1(n_149), .A2(n_192), .B1(n_563), .B2(n_564), .Y(n_562) );
INVx5_ASAP7_75t_L g149 ( .A(n_150), .Y(n_149) );
NOR2xp33_ASAP7_75t_L g223 ( .A(n_150), .B(n_224), .Y(n_223) );
NOR2xp33_ASAP7_75t_L g243 ( .A(n_150), .B(n_244), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g465 ( .A(n_150), .B(n_466), .Y(n_465) );
AOI21xp5_ASAP7_75t_L g267 ( .A1(n_153), .A2(n_268), .B(n_269), .Y(n_267) );
O2A1O1Ixp5_ASAP7_75t_L g484 ( .A1(n_153), .A2(n_485), .B(n_486), .C(n_487), .Y(n_484) );
O2A1O1Ixp33_ASAP7_75t_L g518 ( .A1(n_153), .A2(n_486), .B(n_519), .C(n_520), .Y(n_518) );
INVx2_ASAP7_75t_L g153 ( .A(n_154), .Y(n_153) );
INVx2_ASAP7_75t_L g154 ( .A(n_155), .Y(n_154) );
INVx1_ASAP7_75t_L g196 ( .A(n_155), .Y(n_196) );
INVx1_ASAP7_75t_L g270 ( .A(n_156), .Y(n_270) );
INVx2_ASAP7_75t_L g156 ( .A(n_157), .Y(n_156) );
AO21x2_ASAP7_75t_L g201 ( .A1(n_157), .A2(n_202), .B(n_212), .Y(n_201) );
AO21x2_ASAP7_75t_L g228 ( .A1(n_157), .A2(n_229), .B(n_236), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g236 ( .A(n_157), .B(n_237), .Y(n_236) );
INVx1_ASAP7_75t_L g157 ( .A(n_158), .Y(n_157) );
BUFx6f_ASAP7_75t_L g166 ( .A(n_158), .Y(n_166) );
AND2x2_ASAP7_75t_L g158 ( .A(n_159), .B(n_160), .Y(n_158) );
AND2x2_ASAP7_75t_SL g170 ( .A(n_159), .B(n_160), .Y(n_170) );
NAND2xp5_ASAP7_75t_L g160 ( .A(n_161), .B(n_162), .Y(n_160) );
NOR2xp33_ASAP7_75t_SL g163 ( .A(n_164), .B(n_165), .Y(n_163) );
INVx3_ASAP7_75t_L g217 ( .A(n_165), .Y(n_217) );
NOR2xp33_ASAP7_75t_L g488 ( .A(n_165), .B(n_489), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g510 ( .A(n_165), .B(n_511), .Y(n_510) );
AO21x2_ASAP7_75t_L g514 ( .A1(n_165), .A2(n_515), .B(n_522), .Y(n_514) );
INVx4_ASAP7_75t_L g165 ( .A(n_166), .Y(n_165) );
OA21x2_ASAP7_75t_L g238 ( .A1(n_166), .A2(n_239), .B(n_245), .Y(n_238) );
HB1xp67_ASAP7_75t_L g470 ( .A(n_166), .Y(n_470) );
AND2x2_ASAP7_75t_L g325 ( .A(n_167), .B(n_326), .Y(n_325) );
INVx1_ASAP7_75t_L g347 ( .A(n_167), .Y(n_347) );
AND2x2_ASAP7_75t_L g432 ( .A(n_167), .B(n_262), .Y(n_432) );
AND2x2_ASAP7_75t_L g435 ( .A(n_167), .B(n_436), .Y(n_435) );
AND2x2_ASAP7_75t_L g167 ( .A(n_168), .B(n_184), .Y(n_167) );
INVx2_ASAP7_75t_L g254 ( .A(n_168), .Y(n_254) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_168), .B(n_279), .Y(n_285) );
AND2x2_ASAP7_75t_L g295 ( .A(n_168), .B(n_296), .Y(n_295) );
INVx1_ASAP7_75t_L g331 ( .A(n_168), .Y(n_331) );
AO21x2_ASAP7_75t_L g168 ( .A1(n_169), .A2(n_171), .B(n_181), .Y(n_168) );
NOR2xp33_ASAP7_75t_L g522 ( .A(n_169), .B(n_523), .Y(n_522) );
INVx1_ASAP7_75t_L g567 ( .A(n_169), .Y(n_567) );
INVx2_ASAP7_75t_L g169 ( .A(n_170), .Y(n_169) );
INVx1_ASAP7_75t_L g183 ( .A(n_170), .Y(n_183) );
OA21x2_ASAP7_75t_L g185 ( .A1(n_170), .A2(n_186), .B(n_198), .Y(n_185) );
OA21x2_ASAP7_75t_L g460 ( .A1(n_170), .A2(n_461), .B(n_467), .Y(n_460) );
O2A1O1Ixp33_ASAP7_75t_L g501 ( .A1(n_170), .A2(n_204), .B(n_502), .C(n_503), .Y(n_501) );
NAND2xp5_ASAP7_75t_L g171 ( .A(n_172), .B(n_180), .Y(n_171) );
AOI21xp5_ASAP7_75t_L g173 ( .A1(n_174), .A2(n_175), .B(n_178), .Y(n_173) );
NOR2xp33_ASAP7_75t_L g529 ( .A(n_176), .B(n_530), .Y(n_529) );
INVx4_ASAP7_75t_L g176 ( .A(n_177), .Y(n_176) );
INVx2_ASAP7_75t_L g222 ( .A(n_177), .Y(n_222) );
HB1xp67_ASAP7_75t_L g178 ( .A(n_179), .Y(n_178) );
INVx3_ASAP7_75t_L g225 ( .A(n_179), .Y(n_225) );
NOR2xp33_ASAP7_75t_L g181 ( .A(n_182), .B(n_183), .Y(n_181) );
NOR2xp33_ASAP7_75t_L g212 ( .A(n_183), .B(n_213), .Y(n_212) );
NOR2xp33_ASAP7_75t_L g271 ( .A(n_183), .B(n_272), .Y(n_271) );
AO21x2_ASAP7_75t_L g480 ( .A1(n_183), .A2(n_481), .B(n_488), .Y(n_480) );
AND2x2_ASAP7_75t_L g273 ( .A(n_184), .B(n_254), .Y(n_273) );
INVx1_ASAP7_75t_L g184 ( .A(n_185), .Y(n_184) );
INVx2_ASAP7_75t_L g255 ( .A(n_185), .Y(n_255) );
AND2x2_ASAP7_75t_L g297 ( .A(n_185), .B(n_279), .Y(n_297) );
AND2x2_ASAP7_75t_L g366 ( .A(n_185), .B(n_263), .Y(n_366) );
O2A1O1Ixp33_ASAP7_75t_L g188 ( .A1(n_189), .A2(n_190), .B(n_191), .C(n_197), .Y(n_188) );
O2A1O1Ixp33_ASAP7_75t_L g219 ( .A1(n_190), .A2(n_197), .B(n_220), .C(n_221), .Y(n_219) );
O2A1O1Ixp33_ASAP7_75t_L g240 ( .A1(n_190), .A2(n_197), .B(n_241), .C(n_242), .Y(n_240) );
O2A1O1Ixp33_ASAP7_75t_SL g462 ( .A1(n_190), .A2(n_197), .B(n_463), .C(n_464), .Y(n_462) );
O2A1O1Ixp33_ASAP7_75t_SL g472 ( .A1(n_190), .A2(n_197), .B(n_473), .C(n_474), .Y(n_472) );
O2A1O1Ixp33_ASAP7_75t_SL g493 ( .A1(n_190), .A2(n_197), .B(n_494), .C(n_495), .Y(n_493) );
O2A1O1Ixp33_ASAP7_75t_L g526 ( .A1(n_190), .A2(n_197), .B(n_527), .C(n_528), .Y(n_526) );
O2A1O1Ixp33_ASAP7_75t_SL g559 ( .A1(n_190), .A2(n_197), .B(n_560), .C(n_561), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g194 ( .A(n_192), .B(n_195), .Y(n_194) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_192), .B(n_476), .Y(n_475) );
NOR2xp33_ASAP7_75t_L g496 ( .A(n_192), .B(n_497), .Y(n_496) );
INVx4_ASAP7_75t_L g192 ( .A(n_193), .Y(n_192) );
OAI22xp5_ASAP7_75t_SL g231 ( .A1(n_193), .A2(n_232), .B1(n_233), .B2(n_234), .Y(n_231) );
INVx2_ASAP7_75t_L g233 ( .A(n_193), .Y(n_233) );
OAI22xp33_ASAP7_75t_L g229 ( .A1(n_197), .A2(n_204), .B1(n_230), .B2(n_235), .Y(n_229) );
INVx1_ASAP7_75t_L g521 ( .A(n_197), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g199 ( .A(n_200), .B(n_214), .Y(n_199) );
OR2x2_ASAP7_75t_L g260 ( .A(n_200), .B(n_228), .Y(n_260) );
INVx1_ASAP7_75t_L g339 ( .A(n_200), .Y(n_339) );
AND2x2_ASAP7_75t_L g353 ( .A(n_200), .B(n_354), .Y(n_353) );
NAND2xp5_ASAP7_75t_L g385 ( .A(n_200), .B(n_227), .Y(n_385) );
NAND2xp5_ASAP7_75t_L g405 ( .A(n_200), .B(n_351), .Y(n_405) );
AND2x2_ASAP7_75t_L g413 ( .A(n_200), .B(n_414), .Y(n_413) );
INVx3_ASAP7_75t_L g200 ( .A(n_201), .Y(n_200) );
INVx3_ASAP7_75t_L g250 ( .A(n_201), .Y(n_250) );
AND2x2_ASAP7_75t_L g320 ( .A(n_201), .B(n_228), .Y(n_320) );
OAI21xp5_ASAP7_75t_L g202 ( .A1(n_203), .A2(n_204), .B(n_205), .Y(n_202) );
OAI21xp5_ASAP7_75t_L g264 ( .A1(n_204), .A2(n_265), .B(n_266), .Y(n_264) );
OAI21xp5_ASAP7_75t_L g481 ( .A1(n_204), .A2(n_482), .B(n_483), .Y(n_481) );
OAI21xp5_ASAP7_75t_L g515 ( .A1(n_204), .A2(n_516), .B(n_517), .Y(n_515) );
INVx2_ASAP7_75t_L g209 ( .A(n_210), .Y(n_209) );
INVx3_ASAP7_75t_L g210 ( .A(n_211), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g443 ( .A(n_214), .B(n_444), .Y(n_443) );
INVx2_ASAP7_75t_L g447 ( .A(n_214), .Y(n_447) );
AND2x2_ASAP7_75t_L g214 ( .A(n_215), .B(n_227), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g313 ( .A(n_215), .B(n_291), .Y(n_313) );
OR2x2_ASAP7_75t_L g342 ( .A(n_215), .B(n_343), .Y(n_342) );
AND2x2_ASAP7_75t_L g374 ( .A(n_215), .B(n_354), .Y(n_374) );
INVx1_ASAP7_75t_SL g394 ( .A(n_215), .Y(n_394) );
AND2x2_ASAP7_75t_L g398 ( .A(n_215), .B(n_259), .Y(n_398) );
INVx2_ASAP7_75t_L g215 ( .A(n_216), .Y(n_215) );
AND2x2_ASAP7_75t_SL g251 ( .A(n_216), .B(n_227), .Y(n_251) );
AND2x2_ASAP7_75t_L g258 ( .A(n_216), .B(n_238), .Y(n_258) );
NAND2xp5_ASAP7_75t_L g282 ( .A(n_216), .B(n_283), .Y(n_282) );
OR2x2_ASAP7_75t_L g301 ( .A(n_216), .B(n_283), .Y(n_301) );
INVx1_ASAP7_75t_SL g308 ( .A(n_216), .Y(n_308) );
BUFx2_ASAP7_75t_L g319 ( .A(n_216), .Y(n_319) );
AND2x2_ASAP7_75t_L g335 ( .A(n_216), .B(n_250), .Y(n_335) );
AND2x2_ASAP7_75t_L g350 ( .A(n_216), .B(n_351), .Y(n_350) );
AND2x2_ASAP7_75t_L g414 ( .A(n_216), .B(n_228), .Y(n_414) );
OA21x2_ASAP7_75t_L g216 ( .A1(n_217), .A2(n_218), .B(n_226), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g334 ( .A(n_227), .B(n_335), .Y(n_334) );
AND2x2_ASAP7_75t_L g338 ( .A(n_227), .B(n_339), .Y(n_338) );
AOI221xp5_ASAP7_75t_L g355 ( .A1(n_227), .A2(n_356), .B1(n_359), .B2(n_362), .C(n_367), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g429 ( .A(n_227), .B(n_430), .Y(n_429) );
AND2x2_ASAP7_75t_L g227 ( .A(n_228), .B(n_238), .Y(n_227) );
INVx3_ASAP7_75t_L g283 ( .A(n_228), .Y(n_283) );
INVx2_ASAP7_75t_L g486 ( .A(n_233), .Y(n_486) );
BUFx2_ASAP7_75t_L g293 ( .A(n_238), .Y(n_293) );
AND2x2_ASAP7_75t_L g307 ( .A(n_238), .B(n_308), .Y(n_307) );
INVx1_ASAP7_75t_L g324 ( .A(n_238), .Y(n_324) );
OR2x2_ASAP7_75t_L g343 ( .A(n_238), .B(n_283), .Y(n_343) );
INVx3_ASAP7_75t_L g351 ( .A(n_238), .Y(n_351) );
AND2x2_ASAP7_75t_L g354 ( .A(n_238), .B(n_283), .Y(n_354) );
AOI221xp5_ASAP7_75t_L g246 ( .A1(n_247), .A2(n_252), .B1(n_256), .B2(n_261), .C(n_274), .Y(n_246) );
INVx1_ASAP7_75t_L g247 ( .A(n_248), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_249), .B(n_251), .Y(n_248) );
NAND2xp5_ASAP7_75t_L g448 ( .A(n_249), .B(n_323), .Y(n_448) );
OR2x2_ASAP7_75t_L g451 ( .A(n_249), .B(n_282), .Y(n_451) );
INVx1_ASAP7_75t_SL g249 ( .A(n_250), .Y(n_249) );
OAI221xp5_ASAP7_75t_SL g274 ( .A1(n_250), .A2(n_275), .B1(n_282), .B2(n_284), .C(n_287), .Y(n_274) );
AND2x2_ASAP7_75t_L g291 ( .A(n_250), .B(n_283), .Y(n_291) );
AND2x2_ASAP7_75t_L g299 ( .A(n_250), .B(n_300), .Y(n_299) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_250), .B(n_307), .Y(n_306) );
NAND2x1_ASAP7_75t_L g349 ( .A(n_250), .B(n_350), .Y(n_349) );
OR2x2_ASAP7_75t_L g401 ( .A(n_250), .B(n_343), .Y(n_401) );
AOI22xp5_ASAP7_75t_L g389 ( .A1(n_252), .A2(n_361), .B1(n_390), .B2(n_392), .Y(n_389) );
INVx2_ASAP7_75t_L g252 ( .A(n_253), .Y(n_252) );
AOI322xp5_ASAP7_75t_L g298 ( .A1(n_253), .A2(n_262), .A3(n_299), .B1(n_302), .B2(n_305), .C1(n_309), .C2(n_312), .Y(n_298) );
OR2x2_ASAP7_75t_L g310 ( .A(n_253), .B(n_311), .Y(n_310) );
OR2x2_ASAP7_75t_L g253 ( .A(n_254), .B(n_255), .Y(n_253) );
NAND2xp5_ASAP7_75t_L g278 ( .A(n_254), .B(n_279), .Y(n_278) );
AND2x2_ASAP7_75t_L g289 ( .A(n_254), .B(n_263), .Y(n_289) );
INVx1_ASAP7_75t_L g304 ( .A(n_254), .Y(n_304) );
AND2x2_ASAP7_75t_L g370 ( .A(n_254), .B(n_371), .Y(n_370) );
AND2x2_ASAP7_75t_L g280 ( .A(n_255), .B(n_281), .Y(n_280) );
INVx2_ASAP7_75t_L g371 ( .A(n_255), .Y(n_371) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_255), .B(n_279), .Y(n_445) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_258), .B(n_259), .Y(n_257) );
NAND2xp5_ASAP7_75t_L g393 ( .A(n_259), .B(n_394), .Y(n_393) );
INVx3_ASAP7_75t_SL g259 ( .A(n_260), .Y(n_259) );
OR2x2_ASAP7_75t_L g345 ( .A(n_260), .B(n_292), .Y(n_345) );
OR2x2_ASAP7_75t_L g442 ( .A(n_260), .B(n_293), .Y(n_442) );
INVx1_ASAP7_75t_L g423 ( .A(n_261), .Y(n_423) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_273), .Y(n_261) );
INVx4_ASAP7_75t_L g311 ( .A(n_262), .Y(n_311) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_262), .B(n_330), .Y(n_336) );
INVx2_ASAP7_75t_L g279 ( .A(n_263), .Y(n_279) );
AO21x2_ASAP7_75t_L g263 ( .A1(n_264), .A2(n_270), .B(n_271), .Y(n_263) );
AO21x2_ASAP7_75t_L g556 ( .A1(n_270), .A2(n_557), .B(n_565), .Y(n_556) );
INVx1_ASAP7_75t_L g574 ( .A(n_270), .Y(n_574) );
INVx1_ASAP7_75t_L g361 ( .A(n_273), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g402 ( .A(n_273), .B(n_333), .Y(n_402) );
AOI21xp33_ASAP7_75t_L g348 ( .A1(n_275), .A2(n_349), .B(n_352), .Y(n_348) );
INVx2_ASAP7_75t_L g275 ( .A(n_276), .Y(n_275) );
AND2x2_ASAP7_75t_L g276 ( .A(n_277), .B(n_280), .Y(n_276) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx2_ASAP7_75t_L g333 ( .A(n_279), .Y(n_333) );
INVx1_ASAP7_75t_L g360 ( .A(n_279), .Y(n_360) );
INVx1_ASAP7_75t_L g286 ( .A(n_280), .Y(n_286) );
AND2x2_ASAP7_75t_L g288 ( .A(n_280), .B(n_289), .Y(n_288) );
AND2x2_ASAP7_75t_L g384 ( .A(n_281), .B(n_370), .Y(n_384) );
AND2x2_ASAP7_75t_L g406 ( .A(n_281), .B(n_366), .Y(n_406) );
BUFx2_ASAP7_75t_L g358 ( .A(n_283), .Y(n_358) );
OR2x2_ASAP7_75t_L g284 ( .A(n_285), .B(n_286), .Y(n_284) );
AOI32xp33_ASAP7_75t_L g287 ( .A1(n_288), .A2(n_290), .A3(n_291), .B1(n_292), .B2(n_294), .Y(n_287) );
INVx1_ASAP7_75t_L g368 ( .A(n_288), .Y(n_368) );
AOI22xp33_ASAP7_75t_L g415 ( .A1(n_288), .A2(n_416), .B1(n_417), .B2(n_419), .Y(n_415) );
INVx1_ASAP7_75t_L g290 ( .A(n_291), .Y(n_290) );
NOR2xp33_ASAP7_75t_L g321 ( .A(n_291), .B(n_322), .Y(n_321) );
NAND2xp5_ASAP7_75t_L g391 ( .A(n_291), .B(n_350), .Y(n_391) );
AND2x2_ASAP7_75t_L g438 ( .A(n_291), .B(n_323), .Y(n_438) );
NAND2xp5_ASAP7_75t_L g386 ( .A(n_292), .B(n_339), .Y(n_386) );
INVx1_ASAP7_75t_L g292 ( .A(n_293), .Y(n_292) );
INVx1_ASAP7_75t_L g439 ( .A(n_294), .Y(n_439) );
AND2x2_ASAP7_75t_L g294 ( .A(n_295), .B(n_297), .Y(n_294) );
INVx1_ASAP7_75t_L g364 ( .A(n_295), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_297), .B(n_304), .Y(n_303) );
AND2x2_ASAP7_75t_L g411 ( .A(n_297), .B(n_331), .Y(n_411) );
NAND2xp5_ASAP7_75t_L g418 ( .A(n_297), .B(n_326), .Y(n_418) );
INVx1_ASAP7_75t_SL g400 ( .A(n_299), .Y(n_400) );
NAND2xp5_ASAP7_75t_L g378 ( .A(n_300), .B(n_351), .Y(n_378) );
NOR4xp25_ASAP7_75t_L g424 ( .A(n_300), .B(n_323), .C(n_425), .D(n_428), .Y(n_424) );
INVx1_ASAP7_75t_L g300 ( .A(n_301), .Y(n_300) );
NOR2xp33_ASAP7_75t_L g404 ( .A(n_301), .B(n_405), .Y(n_404) );
INVx1_ASAP7_75t_L g302 ( .A(n_303), .Y(n_302) );
INVxp67_ASAP7_75t_L g381 ( .A(n_304), .Y(n_381) );
INVx1_ASAP7_75t_L g305 ( .A(n_306), .Y(n_305) );
OAI21xp33_ASAP7_75t_L g431 ( .A1(n_307), .A2(n_398), .B(n_432), .Y(n_431) );
AND2x4_ASAP7_75t_L g323 ( .A(n_308), .B(n_324), .Y(n_323) );
INVx1_ASAP7_75t_L g309 ( .A(n_310), .Y(n_309) );
INVx1_ASAP7_75t_L g372 ( .A(n_311), .Y(n_372) );
INVx1_ASAP7_75t_L g312 ( .A(n_313), .Y(n_312) );
NAND4xp25_ASAP7_75t_SL g314 ( .A(n_315), .B(n_340), .C(n_355), .D(n_375), .Y(n_314) );
O2A1O1Ixp33_ASAP7_75t_L g315 ( .A1(n_316), .A2(n_321), .B(n_325), .C(n_327), .Y(n_315) );
INVx1_ASAP7_75t_SL g316 ( .A(n_317), .Y(n_316) );
NAND2xp5_ASAP7_75t_L g317 ( .A(n_318), .B(n_320), .Y(n_317) );
INVx1_ASAP7_75t_SL g318 ( .A(n_319), .Y(n_318) );
AND2x2_ASAP7_75t_L g407 ( .A(n_320), .B(n_350), .Y(n_407) );
AND2x2_ASAP7_75t_L g416 ( .A(n_320), .B(n_394), .Y(n_416) );
INVx3_ASAP7_75t_SL g322 ( .A(n_323), .Y(n_322) );
NAND2xp5_ASAP7_75t_L g420 ( .A(n_323), .B(n_358), .Y(n_420) );
AND2x2_ASAP7_75t_L g332 ( .A(n_326), .B(n_333), .Y(n_332) );
OAI22xp5_ASAP7_75t_L g327 ( .A1(n_328), .A2(n_334), .B1(n_336), .B2(n_337), .Y(n_327) );
INVx1_ASAP7_75t_L g328 ( .A(n_329), .Y(n_328) );
AND2x2_ASAP7_75t_L g329 ( .A(n_330), .B(n_332), .Y(n_329) );
AND2x2_ASAP7_75t_L g430 ( .A(n_330), .B(n_376), .Y(n_430) );
INVx1_ASAP7_75t_L g330 ( .A(n_331), .Y(n_330) );
NAND2xp5_ASAP7_75t_L g397 ( .A(n_332), .B(n_381), .Y(n_397) );
NOR2xp33_ASAP7_75t_L g346 ( .A(n_333), .B(n_347), .Y(n_346) );
INVx1_ASAP7_75t_L g337 ( .A(n_338), .Y(n_337) );
O2A1O1Ixp33_ASAP7_75t_L g340 ( .A1(n_341), .A2(n_344), .B(n_346), .C(n_348), .Y(n_340) );
AOI221xp5_ASAP7_75t_L g375 ( .A1(n_341), .A2(n_376), .B1(n_377), .B2(n_379), .C(n_382), .Y(n_375) );
INVx1_ASAP7_75t_SL g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g344 ( .A(n_345), .Y(n_344) );
OAI221xp5_ASAP7_75t_L g433 ( .A1(n_349), .A2(n_434), .B1(n_437), .B2(n_439), .C(n_440), .Y(n_433) );
NAND2xp5_ASAP7_75t_L g357 ( .A(n_350), .B(n_358), .Y(n_357) );
INVx1_ASAP7_75t_SL g352 ( .A(n_353), .Y(n_352) );
INVx1_ASAP7_75t_L g356 ( .A(n_357), .Y(n_356) );
NAND2xp5_ASAP7_75t_L g426 ( .A(n_358), .B(n_427), .Y(n_426) );
NOR2xp33_ASAP7_75t_L g359 ( .A(n_360), .B(n_361), .Y(n_359) );
INVx1_ASAP7_75t_L g388 ( .A(n_360), .Y(n_388) );
INVx1_ASAP7_75t_SL g362 ( .A(n_363), .Y(n_362) );
OAI22xp5_ASAP7_75t_L g382 ( .A1(n_363), .A2(n_383), .B1(n_385), .B2(n_386), .Y(n_382) );
OR2x2_ASAP7_75t_L g363 ( .A(n_364), .B(n_365), .Y(n_363) );
INVx1_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
AOI21xp33_ASAP7_75t_L g367 ( .A1(n_368), .A2(n_369), .B(n_373), .Y(n_367) );
NAND2xp5_ASAP7_75t_L g369 ( .A(n_370), .B(n_372), .Y(n_369) );
NAND2xp5_ASAP7_75t_L g380 ( .A(n_372), .B(n_381), .Y(n_380) );
INVx1_ASAP7_75t_L g373 ( .A(n_374), .Y(n_373) );
INVx1_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
INVx1_ASAP7_75t_L g379 ( .A(n_380), .Y(n_379) );
OAI221xp5_ASAP7_75t_L g446 ( .A1(n_383), .A2(n_409), .B1(n_447), .B2(n_448), .C(n_449), .Y(n_446) );
INVx1_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
INVx1_ASAP7_75t_L g428 ( .A(n_385), .Y(n_428) );
OAI211xp5_ASAP7_75t_SL g387 ( .A1(n_388), .A2(n_389), .B(n_395), .C(n_415), .Y(n_387) );
INVx1_ASAP7_75t_L g390 ( .A(n_391), .Y(n_390) );
INVx1_ASAP7_75t_L g392 ( .A(n_393), .Y(n_392) );
AOI211xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_398), .B(n_399), .C(n_408), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
A2O1A1Ixp33_ASAP7_75t_L g399 ( .A1(n_400), .A2(n_401), .B(n_402), .C(n_403), .Y(n_399) );
INVx1_ASAP7_75t_L g427 ( .A(n_405), .Y(n_427) );
OAI21xp5_ASAP7_75t_SL g449 ( .A1(n_406), .A2(n_432), .B(n_450), .Y(n_449) );
AOI21xp33_ASAP7_75t_L g408 ( .A1(n_409), .A2(n_410), .B(n_412), .Y(n_408) );
INVx1_ASAP7_75t_SL g410 ( .A(n_411), .Y(n_410) );
INVxp67_ASAP7_75t_L g412 ( .A(n_413), .Y(n_412) );
INVx1_ASAP7_75t_L g417 ( .A(n_418), .Y(n_417) );
OAI21xp5_ASAP7_75t_SL g441 ( .A1(n_418), .A2(n_442), .B(n_443), .Y(n_441) );
INVx1_ASAP7_75t_L g419 ( .A(n_420), .Y(n_419) );
NOR3xp33_ASAP7_75t_L g421 ( .A(n_422), .B(n_433), .C(n_446), .Y(n_421) );
OAI211xp5_ASAP7_75t_L g422 ( .A1(n_423), .A2(n_424), .B(n_429), .C(n_431), .Y(n_422) );
INVx1_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
CKINVDCx14_ASAP7_75t_R g434 ( .A(n_435), .Y(n_434) );
INVx2_ASAP7_75t_L g437 ( .A(n_438), .Y(n_437) );
INVx1_ASAP7_75t_L g440 ( .A(n_441), .Y(n_440) );
INVx1_ASAP7_75t_L g450 ( .A(n_451), .Y(n_450) );
INVx1_ASAP7_75t_L g728 ( .A(n_452), .Y(n_728) );
INVx2_ASAP7_75t_L g454 ( .A(n_455), .Y(n_454) );
OAI22xp5_ASAP7_75t_SL g725 ( .A1(n_455), .A2(n_723), .B1(n_726), .B2(n_727), .Y(n_725) );
XOR2xp5_ASAP7_75t_L g734 ( .A(n_455), .B(n_735), .Y(n_734) );
OR2x2_ASAP7_75t_L g455 ( .A(n_456), .B(n_653), .Y(n_455) );
NAND5xp2_ASAP7_75t_L g456 ( .A(n_457), .B(n_568), .C(n_600), .D(n_617), .E(n_640), .Y(n_456) );
AOI221xp5_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_499), .B1(n_532), .B2(n_536), .C(n_540), .Y(n_457) );
INVx1_ASAP7_75t_L g680 ( .A(n_458), .Y(n_680) );
AND2x2_ASAP7_75t_L g458 ( .A(n_459), .B(n_478), .Y(n_458) );
AND3x2_ASAP7_75t_L g655 ( .A(n_459), .B(n_480), .C(n_656), .Y(n_655) );
AND2x2_ASAP7_75t_L g459 ( .A(n_460), .B(n_468), .Y(n_459) );
NAND2xp5_ASAP7_75t_L g537 ( .A(n_460), .B(n_538), .Y(n_537) );
BUFx3_ASAP7_75t_L g547 ( .A(n_460), .Y(n_547) );
AND2x2_ASAP7_75t_L g551 ( .A(n_460), .B(n_490), .Y(n_551) );
INVx2_ASAP7_75t_L g577 ( .A(n_460), .Y(n_577) );
OR2x2_ASAP7_75t_L g588 ( .A(n_460), .B(n_491), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g607 ( .A(n_460), .B(n_479), .Y(n_607) );
NAND2xp5_ASAP7_75t_L g625 ( .A(n_460), .B(n_626), .Y(n_625) );
AND2x2_ASAP7_75t_L g667 ( .A(n_460), .B(n_491), .Y(n_667) );
HB1xp67_ASAP7_75t_L g550 ( .A(n_468), .Y(n_550) );
AND2x2_ASAP7_75t_L g608 ( .A(n_468), .B(n_609), .Y(n_608) );
NAND2xp5_ASAP7_75t_L g627 ( .A(n_468), .B(n_479), .Y(n_627) );
INVx1_ASAP7_75t_SL g468 ( .A(n_469), .Y(n_468) );
OR2x2_ASAP7_75t_L g539 ( .A(n_469), .B(n_479), .Y(n_539) );
HB1xp67_ASAP7_75t_L g546 ( .A(n_469), .Y(n_546) );
AND2x2_ASAP7_75t_L g594 ( .A(n_469), .B(n_491), .Y(n_594) );
NAND3xp33_ASAP7_75t_L g619 ( .A(n_469), .B(n_478), .C(n_577), .Y(n_619) );
AND2x2_ASAP7_75t_L g684 ( .A(n_469), .B(n_480), .Y(n_684) );
AND2x2_ASAP7_75t_L g718 ( .A(n_469), .B(n_479), .Y(n_718) );
OA21x2_ASAP7_75t_L g469 ( .A1(n_470), .A2(n_471), .B(n_477), .Y(n_469) );
OA21x2_ASAP7_75t_L g491 ( .A1(n_470), .A2(n_492), .B(n_498), .Y(n_491) );
OA21x2_ASAP7_75t_L g524 ( .A1(n_470), .A2(n_525), .B(n_531), .Y(n_524) );
INVxp67_ASAP7_75t_L g548 ( .A(n_478), .Y(n_548) );
AND2x2_ASAP7_75t_L g478 ( .A(n_479), .B(n_490), .Y(n_478) );
NAND2xp5_ASAP7_75t_L g595 ( .A(n_479), .B(n_577), .Y(n_595) );
NAND2xp5_ASAP7_75t_L g616 ( .A(n_479), .B(n_608), .Y(n_616) );
AND2x2_ASAP7_75t_L g666 ( .A(n_479), .B(n_667), .Y(n_666) );
INVx1_ASAP7_75t_L g694 ( .A(n_479), .Y(n_694) );
INVx4_ASAP7_75t_L g479 ( .A(n_480), .Y(n_479) );
AND2x2_ASAP7_75t_L g601 ( .A(n_480), .B(n_594), .Y(n_601) );
BUFx3_ASAP7_75t_L g633 ( .A(n_480), .Y(n_633) );
INVx2_ASAP7_75t_L g609 ( .A(n_490), .Y(n_609) );
INVx2_ASAP7_75t_L g490 ( .A(n_491), .Y(n_490) );
HB1xp67_ASAP7_75t_L g578 ( .A(n_491), .Y(n_578) );
AOI22xp33_ASAP7_75t_L g668 ( .A1(n_499), .A2(n_669), .B1(n_671), .B2(n_672), .Y(n_668) );
AND2x2_ASAP7_75t_L g499 ( .A(n_500), .B(n_512), .Y(n_499) );
AND2x2_ASAP7_75t_L g532 ( .A(n_500), .B(n_533), .Y(n_532) );
INVx3_ASAP7_75t_SL g543 ( .A(n_500), .Y(n_543) );
NAND2xp5_ASAP7_75t_L g604 ( .A(n_500), .B(n_572), .Y(n_604) );
OR2x2_ASAP7_75t_L g623 ( .A(n_500), .B(n_513), .Y(n_623) );
AND2x2_ASAP7_75t_L g628 ( .A(n_500), .B(n_580), .Y(n_628) );
AND2x2_ASAP7_75t_L g631 ( .A(n_500), .B(n_573), .Y(n_631) );
AND2x2_ASAP7_75t_L g643 ( .A(n_500), .B(n_524), .Y(n_643) );
AND2x2_ASAP7_75t_L g659 ( .A(n_500), .B(n_514), .Y(n_659) );
AND2x4_ASAP7_75t_L g662 ( .A(n_500), .B(n_534), .Y(n_662) );
OR2x2_ASAP7_75t_L g679 ( .A(n_500), .B(n_615), .Y(n_679) );
OR2x2_ASAP7_75t_L g710 ( .A(n_500), .B(n_556), .Y(n_710) );
NAND2xp5_ASAP7_75t_SL g712 ( .A(n_500), .B(n_638), .Y(n_712) );
OR2x6_ASAP7_75t_L g500 ( .A(n_501), .B(n_510), .Y(n_500) );
INVx2_ASAP7_75t_L g507 ( .A(n_508), .Y(n_507) );
NAND2xp5_ASAP7_75t_SL g561 ( .A(n_508), .B(n_562), .Y(n_561) );
AND2x2_ASAP7_75t_L g586 ( .A(n_512), .B(n_554), .Y(n_586) );
NAND2xp5_ASAP7_75t_L g705 ( .A(n_512), .B(n_573), .Y(n_705) );
AND2x2_ASAP7_75t_L g512 ( .A(n_513), .B(n_524), .Y(n_512) );
AND2x2_ASAP7_75t_L g542 ( .A(n_513), .B(n_543), .Y(n_542) );
AND2x2_ASAP7_75t_L g572 ( .A(n_513), .B(n_573), .Y(n_572) );
AND2x2_ASAP7_75t_L g580 ( .A(n_513), .B(n_556), .Y(n_580) );
AND2x2_ASAP7_75t_L g598 ( .A(n_513), .B(n_534), .Y(n_598) );
OR2x2_ASAP7_75t_L g615 ( .A(n_513), .B(n_573), .Y(n_615) );
INVx2_ASAP7_75t_SL g513 ( .A(n_514), .Y(n_513) );
BUFx2_ASAP7_75t_L g535 ( .A(n_514), .Y(n_535) );
AND2x2_ASAP7_75t_L g638 ( .A(n_514), .B(n_524), .Y(n_638) );
INVx2_ASAP7_75t_L g534 ( .A(n_524), .Y(n_534) );
INVx1_ASAP7_75t_L g650 ( .A(n_524), .Y(n_650) );
AND2x2_ASAP7_75t_L g700 ( .A(n_524), .B(n_543), .Y(n_700) );
AND2x2_ASAP7_75t_L g553 ( .A(n_533), .B(n_554), .Y(n_553) );
AND2x2_ASAP7_75t_L g584 ( .A(n_533), .B(n_543), .Y(n_584) );
NAND2xp5_ASAP7_75t_L g630 ( .A(n_533), .B(n_631), .Y(n_630) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g571 ( .A(n_534), .B(n_543), .Y(n_571) );
OR2x2_ASAP7_75t_L g687 ( .A(n_535), .B(n_661), .Y(n_687) );
INVx1_ASAP7_75t_L g536 ( .A(n_537), .Y(n_536) );
NAND2xp5_ASAP7_75t_L g673 ( .A(n_538), .B(n_667), .Y(n_673) );
INVx2_ASAP7_75t_SL g538 ( .A(n_539), .Y(n_538) );
OAI32xp33_ASAP7_75t_L g629 ( .A1(n_539), .A2(n_630), .A3(n_632), .B1(n_634), .B2(n_635), .Y(n_629) );
OR2x2_ASAP7_75t_L g646 ( .A(n_539), .B(n_588), .Y(n_646) );
OAI21xp33_ASAP7_75t_SL g671 ( .A1(n_539), .A2(n_549), .B(n_576), .Y(n_671) );
OAI22xp33_ASAP7_75t_L g540 ( .A1(n_541), .A2(n_544), .B1(n_549), .B2(n_552), .Y(n_540) );
INVxp33_ASAP7_75t_L g541 ( .A(n_542), .Y(n_541) );
NAND2xp5_ASAP7_75t_L g611 ( .A(n_542), .B(n_612), .Y(n_611) );
NAND2xp5_ASAP7_75t_L g579 ( .A(n_543), .B(n_580), .Y(n_579) );
AND2x2_ASAP7_75t_L g597 ( .A(n_543), .B(n_598), .Y(n_597) );
AND2x2_ASAP7_75t_L g697 ( .A(n_543), .B(n_638), .Y(n_697) );
OR2x2_ASAP7_75t_L g721 ( .A(n_543), .B(n_615), .Y(n_721) );
AOI21xp33_ASAP7_75t_L g704 ( .A1(n_544), .A2(n_603), .B(n_705), .Y(n_704) );
OR2x2_ASAP7_75t_L g544 ( .A(n_545), .B(n_548), .Y(n_544) );
NAND2xp5_ASAP7_75t_L g545 ( .A(n_546), .B(n_547), .Y(n_545) );
INVx1_ASAP7_75t_L g581 ( .A(n_546), .Y(n_581) );
NAND2xp5_ASAP7_75t_L g599 ( .A(n_546), .B(n_551), .Y(n_599) );
AND2x2_ASAP7_75t_L g621 ( .A(n_547), .B(n_594), .Y(n_621) );
INVx1_ASAP7_75t_L g634 ( .A(n_547), .Y(n_634) );
OR2x2_ASAP7_75t_L g639 ( .A(n_547), .B(n_573), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g549 ( .A(n_550), .B(n_551), .Y(n_549) );
NOR2xp33_ASAP7_75t_L g587 ( .A(n_550), .B(n_588), .Y(n_587) );
OAI22xp33_ASAP7_75t_L g569 ( .A1(n_551), .A2(n_570), .B1(n_575), .B2(n_579), .Y(n_569) );
INVx1_ASAP7_75t_L g552 ( .A(n_553), .Y(n_552) );
OAI22xp5_ASAP7_75t_L g618 ( .A1(n_554), .A2(n_612), .B1(n_619), .B2(n_620), .Y(n_618) );
AND2x2_ASAP7_75t_L g696 ( .A(n_554), .B(n_697), .Y(n_696) );
INVx2_ASAP7_75t_L g554 ( .A(n_555), .Y(n_554) );
INVx1_ASAP7_75t_SL g555 ( .A(n_556), .Y(n_555) );
NAND2xp5_ASAP7_75t_L g649 ( .A(n_556), .B(n_650), .Y(n_649) );
AND2x2_ASAP7_75t_L g715 ( .A(n_556), .B(n_598), .Y(n_715) );
INVx1_ASAP7_75t_L g557 ( .A(n_558), .Y(n_557) );
OA21x2_ASAP7_75t_L g573 ( .A1(n_558), .A2(n_566), .B(n_574), .Y(n_573) );
INVx1_ASAP7_75t_L g565 ( .A(n_566), .Y(n_565) );
AOI221xp5_ASAP7_75t_L g568 ( .A1(n_569), .A2(n_581), .B1(n_582), .B2(n_587), .C(n_589), .Y(n_568) );
NAND2xp5_ASAP7_75t_L g570 ( .A(n_571), .B(n_572), .Y(n_570) );
NAND2xp5_ASAP7_75t_L g603 ( .A(n_571), .B(n_573), .Y(n_603) );
NAND2xp5_ASAP7_75t_L g613 ( .A(n_571), .B(n_614), .Y(n_613) );
INVx1_ASAP7_75t_L g590 ( .A(n_572), .Y(n_590) );
O2A1O1Ixp33_ASAP7_75t_L g677 ( .A1(n_572), .A2(n_678), .B(n_679), .C(n_680), .Y(n_677) );
AND2x2_ASAP7_75t_L g682 ( .A(n_572), .B(n_662), .Y(n_682) );
O2A1O1Ixp33_ASAP7_75t_SL g720 ( .A1(n_572), .A2(n_661), .B(n_721), .C(n_722), .Y(n_720) );
BUFx3_ASAP7_75t_L g612 ( .A(n_573), .Y(n_612) );
INVx1_ASAP7_75t_L g575 ( .A(n_576), .Y(n_575) );
NAND2xp5_ASAP7_75t_L g676 ( .A(n_576), .B(n_633), .Y(n_676) );
AOI211xp5_ASAP7_75t_L g695 ( .A1(n_576), .A2(n_696), .B(n_698), .C(n_704), .Y(n_695) );
AND2x2_ASAP7_75t_L g576 ( .A(n_577), .B(n_578), .Y(n_576) );
INVxp67_ASAP7_75t_L g656 ( .A(n_578), .Y(n_656) );
NAND2xp5_ASAP7_75t_L g699 ( .A(n_580), .B(n_700), .Y(n_699) );
NAND2xp5_ASAP7_75t_SL g582 ( .A(n_583), .B(n_585), .Y(n_582) );
INVx1_ASAP7_75t_SL g583 ( .A(n_584), .Y(n_583) );
AOI211xp5_ASAP7_75t_L g600 ( .A1(n_584), .A2(n_601), .B(n_602), .C(n_610), .Y(n_600) );
INVx1_ASAP7_75t_L g585 ( .A(n_586), .Y(n_585) );
INVx1_ASAP7_75t_L g685 ( .A(n_588), .Y(n_685) );
OR2x2_ASAP7_75t_L g702 ( .A(n_588), .B(n_632), .Y(n_702) );
OAI22xp5_ASAP7_75t_L g589 ( .A1(n_590), .A2(n_591), .B1(n_596), .B2(n_599), .Y(n_589) );
OAI22xp33_ASAP7_75t_L g602 ( .A1(n_591), .A2(n_603), .B1(n_604), .B2(n_605), .Y(n_602) );
INVx1_ASAP7_75t_L g591 ( .A(n_592), .Y(n_591) );
NOR2xp33_ASAP7_75t_L g592 ( .A(n_593), .B(n_595), .Y(n_592) );
OR2x2_ASAP7_75t_L g689 ( .A(n_593), .B(n_633), .Y(n_689) );
INVx1_ASAP7_75t_SL g593 ( .A(n_594), .Y(n_593) );
AND2x2_ASAP7_75t_L g644 ( .A(n_594), .B(n_634), .Y(n_644) );
INVx1_ASAP7_75t_L g652 ( .A(n_595), .Y(n_652) );
INVx1_ASAP7_75t_L g596 ( .A(n_597), .Y(n_596) );
NAND2xp5_ASAP7_75t_L g660 ( .A(n_598), .B(n_612), .Y(n_660) );
INVx1_ASAP7_75t_L g605 ( .A(n_606), .Y(n_605) );
AND2x2_ASAP7_75t_L g606 ( .A(n_607), .B(n_608), .Y(n_606) );
NAND2xp5_ASAP7_75t_SL g651 ( .A(n_608), .B(n_652), .Y(n_651) );
INVx2_ASAP7_75t_L g717 ( .A(n_609), .Y(n_717) );
AOI21xp33_ASAP7_75t_L g610 ( .A1(n_611), .A2(n_613), .B(n_616), .Y(n_610) );
INVx1_ASAP7_75t_L g647 ( .A(n_611), .Y(n_647) );
NAND2xp5_ASAP7_75t_SL g622 ( .A(n_612), .B(n_623), .Y(n_622) );
NAND2xp5_ASAP7_75t_L g642 ( .A(n_612), .B(n_643), .Y(n_642) );
NAND2x1p5_ASAP7_75t_L g663 ( .A(n_612), .B(n_638), .Y(n_663) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_612), .B(n_659), .Y(n_670) );
OAI211xp5_ASAP7_75t_L g674 ( .A1(n_612), .A2(n_622), .B(n_662), .C(n_675), .Y(n_674) );
INVx1_ASAP7_75t_SL g614 ( .A(n_615), .Y(n_614) );
AOI221xp5_ASAP7_75t_SL g617 ( .A1(n_618), .A2(n_622), .B1(n_624), .B2(n_628), .C(n_629), .Y(n_617) );
INVx1_ASAP7_75t_L g620 ( .A(n_621), .Y(n_620) );
INVxp67_ASAP7_75t_L g624 ( .A(n_625), .Y(n_624) );
NAND2xp5_ASAP7_75t_L g708 ( .A(n_626), .B(n_634), .Y(n_708) );
INVx1_ASAP7_75t_L g626 ( .A(n_627), .Y(n_626) );
O2A1O1Ixp33_ASAP7_75t_L g719 ( .A1(n_628), .A2(n_643), .B(n_645), .C(n_720), .Y(n_719) );
NAND2xp5_ASAP7_75t_L g703 ( .A(n_631), .B(n_638), .Y(n_703) );
NAND2xp5_ASAP7_75t_SL g722 ( .A(n_632), .B(n_685), .Y(n_722) );
CKINVDCx16_ASAP7_75t_R g632 ( .A(n_633), .Y(n_632) );
INVxp33_ASAP7_75t_L g635 ( .A(n_636), .Y(n_635) );
NOR2xp33_ASAP7_75t_L g636 ( .A(n_637), .B(n_639), .Y(n_636) );
AOI21xp33_ASAP7_75t_SL g648 ( .A1(n_637), .A2(n_649), .B(n_651), .Y(n_648) );
NOR2xp33_ASAP7_75t_L g709 ( .A(n_637), .B(n_710), .Y(n_709) );
INVx2_ASAP7_75t_SL g637 ( .A(n_638), .Y(n_637) );
NAND2xp5_ASAP7_75t_L g691 ( .A(n_638), .B(n_692), .Y(n_691) );
AOI221xp5_ASAP7_75t_L g640 ( .A1(n_641), .A2(n_644), .B1(n_645), .B2(n_647), .C(n_648), .Y(n_640) );
INVx1_ASAP7_75t_L g641 ( .A(n_642), .Y(n_641) );
NAND2xp5_ASAP7_75t_L g693 ( .A(n_644), .B(n_694), .Y(n_693) );
INVx1_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
INVx1_ASAP7_75t_L g678 ( .A(n_650), .Y(n_678) );
NAND5xp2_ASAP7_75t_L g653 ( .A(n_654), .B(n_681), .C(n_695), .D(n_706), .E(n_719), .Y(n_653) );
AOI211xp5_ASAP7_75t_L g654 ( .A1(n_655), .A2(n_657), .B(n_664), .C(n_677), .Y(n_654) );
INVx2_ASAP7_75t_SL g701 ( .A(n_655), .Y(n_701) );
NAND4xp25_ASAP7_75t_SL g657 ( .A(n_658), .B(n_660), .C(n_661), .D(n_663), .Y(n_657) );
INVx1_ASAP7_75t_L g658 ( .A(n_659), .Y(n_658) );
INVx3_ASAP7_75t_L g661 ( .A(n_662), .Y(n_661) );
OAI211xp5_ASAP7_75t_SL g664 ( .A1(n_663), .A2(n_665), .B(n_668), .C(n_674), .Y(n_664) );
CKINVDCx20_ASAP7_75t_R g665 ( .A(n_666), .Y(n_665) );
AOI221xp5_ASAP7_75t_L g706 ( .A1(n_666), .A2(n_707), .B1(n_709), .B2(n_711), .C(n_713), .Y(n_706) );
INVx1_ASAP7_75t_L g669 ( .A(n_670), .Y(n_669) );
INVx1_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx1_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
AOI221xp5_ASAP7_75t_SL g681 ( .A1(n_682), .A2(n_683), .B1(n_686), .B2(n_688), .C(n_690), .Y(n_681) );
AND2x2_ASAP7_75t_L g683 ( .A(n_684), .B(n_685), .Y(n_683) );
INVx1_ASAP7_75t_L g686 ( .A(n_687), .Y(n_686) );
INVx1_ASAP7_75t_L g688 ( .A(n_689), .Y(n_688) );
OAI22xp5_ASAP7_75t_L g713 ( .A1(n_689), .A2(n_712), .B1(n_714), .B2(n_716), .Y(n_713) );
INVx1_ASAP7_75t_L g690 ( .A(n_691), .Y(n_690) );
INVx1_ASAP7_75t_SL g692 ( .A(n_693), .Y(n_692) );
OAI22xp5_ASAP7_75t_L g698 ( .A1(n_699), .A2(n_701), .B1(n_702), .B2(n_703), .Y(n_698) );
INVx1_ASAP7_75t_L g707 ( .A(n_708), .Y(n_707) );
INVx1_ASAP7_75t_L g711 ( .A(n_712), .Y(n_711) );
INVx1_ASAP7_75t_SL g714 ( .A(n_715), .Y(n_714) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_718), .Y(n_716) );
INVx2_ASAP7_75t_L g727 ( .A(n_728), .Y(n_727) );
INVx1_ASAP7_75t_SL g729 ( .A(n_730), .Y(n_729) );
INVx3_ASAP7_75t_SL g730 ( .A(n_731), .Y(n_730) );
CKINVDCx20_ASAP7_75t_R g739 ( .A(n_740), .Y(n_739) );
endmodule