module fake_jpeg_17446_n_114 (n_11, n_3, n_2, n_1, n_0, n_10, n_4, n_8, n_9, n_6, n_5, n_7, n_114);

input n_11;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_4;
input n_8;
input n_9;
input n_6;
input n_5;
input n_7;

output n_114;

wire n_105;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_84;
wire n_98;
wire n_65;
wire n_110;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_88;
wire n_74;
wire n_31;
wire n_29;
wire n_103;
wire n_50;
wire n_15;
wire n_13;
wire n_57;
wire n_21;
wire n_23;
wire n_69;
wire n_27;
wire n_83;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_109;
wire n_113;
wire n_30;
wire n_106;
wire n_111;
wire n_24;
wire n_44;
wire n_25;
wire n_17;
wire n_75;
wire n_37;
wire n_102;
wire n_99;
wire n_70;
wire n_66;
wire n_85;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_20;
wire n_18;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_58;
wire n_41;
wire n_90;
wire n_60;
wire n_92;
wire n_63;
wire n_34;
wire n_39;
wire n_107;
wire n_72;
wire n_89;
wire n_104;
wire n_56;
wire n_79;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_91;
wire n_93;
wire n_22;
wire n_101;
wire n_48;
wire n_35;
wire n_87;
wire n_46;
wire n_86;
wire n_112;
wire n_95;
wire n_97;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_100;
wire n_82;
wire n_96;

CKINVDCx20_ASAP7_75t_R g12 ( 
.A(n_11),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

BUFx6f_ASAP7_75t_L g14 ( 
.A(n_11),
.Y(n_14)
);

BUFx6f_ASAP7_75t_L g15 ( 
.A(n_9),
.Y(n_15)
);

CKINVDCx5p33_ASAP7_75t_R g16 ( 
.A(n_7),
.Y(n_16)
);

BUFx5_ASAP7_75t_L g17 ( 
.A(n_5),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_7),
.Y(n_18)
);

BUFx16f_ASAP7_75t_L g19 ( 
.A(n_0),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_4),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_6),
.Y(n_22)
);

BUFx3_ASAP7_75t_L g23 ( 
.A(n_8),
.Y(n_23)
);

BUFx6f_ASAP7_75t_L g24 ( 
.A(n_9),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_6),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_13),
.Y(n_26)
);

INVx3_ASAP7_75t_L g35 ( 
.A(n_26),
.Y(n_35)
);

INVx4_ASAP7_75t_L g27 ( 
.A(n_20),
.Y(n_27)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_27),
.B(n_34),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g28 ( 
.A(n_20),
.Y(n_28)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_28),
.Y(n_39)
);

INVx11_ASAP7_75t_L g29 ( 
.A(n_19),
.Y(n_29)
);

INVx6_ASAP7_75t_L g36 ( 
.A(n_29),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g30 ( 
.A(n_25),
.B(n_0),
.Y(n_30)
);

INVx1_ASAP7_75t_L g41 ( 
.A(n_30),
.Y(n_41)
);

INVx2_ASAP7_75t_L g31 ( 
.A(n_13),
.Y(n_31)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_31),
.Y(n_42)
);

NOR2xp33_ASAP7_75t_L g32 ( 
.A(n_23),
.B(n_0),
.Y(n_32)
);

INVx1_ASAP7_75t_L g46 ( 
.A(n_32),
.Y(n_46)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_33),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_23),
.B(n_1),
.Y(n_34)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_32),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_37),
.B(n_40),
.Y(n_55)
);

INVxp67_ASAP7_75t_L g40 ( 
.A(n_34),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_L g43 ( 
.A1(n_31),
.A2(n_19),
.B1(n_12),
.B2(n_24),
.Y(n_43)
);

AOI22xp33_ASAP7_75t_SL g59 ( 
.A1(n_43),
.A2(n_29),
.B1(n_15),
.B2(n_24),
.Y(n_59)
);

AOI22xp5_ASAP7_75t_SL g45 ( 
.A1(n_27),
.A2(n_16),
.B1(n_22),
.B2(n_18),
.Y(n_45)
);

OR2x2_ASAP7_75t_L g50 ( 
.A(n_45),
.B(n_17),
.Y(n_50)
);

NAND2xp5_ASAP7_75t_L g47 ( 
.A(n_40),
.B(n_30),
.Y(n_47)
);

MAJIxp5_ASAP7_75t_L g66 ( 
.A(n_47),
.B(n_49),
.C(n_54),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_SL g48 ( 
.A(n_41),
.B(n_5),
.Y(n_48)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_48),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g49 ( 
.A(n_41),
.B(n_28),
.Y(n_49)
);

OAI22xp33_ASAP7_75t_SL g71 ( 
.A1(n_50),
.A2(n_60),
.B1(n_36),
.B2(n_55),
.Y(n_71)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_42),
.Y(n_51)
);

INVx1_ASAP7_75t_L g68 ( 
.A(n_51),
.Y(n_68)
);

INVxp67_ASAP7_75t_L g52 ( 
.A(n_45),
.Y(n_52)
);

CKINVDCx16_ASAP7_75t_R g73 ( 
.A(n_52),
.Y(n_73)
);

NOR2xp67_ASAP7_75t_SL g53 ( 
.A(n_46),
.B(n_20),
.Y(n_53)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_53),
.A2(n_61),
.B(n_49),
.Y(n_74)
);

XOR2xp5_ASAP7_75t_L g54 ( 
.A(n_38),
.B(n_27),
.Y(n_54)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_56),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g57 ( 
.A(n_35),
.B(n_28),
.Y(n_57)
);

INVx1_ASAP7_75t_L g65 ( 
.A(n_57),
.Y(n_65)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_44),
.Y(n_58)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_58),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g62 ( 
.A1(n_59),
.A2(n_29),
.B1(n_36),
.B2(n_33),
.Y(n_62)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_44),
.Y(n_60)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_39),
.B(n_28),
.Y(n_61)
);

AOI22xp33_ASAP7_75t_L g75 ( 
.A1(n_62),
.A2(n_58),
.B1(n_51),
.B2(n_33),
.Y(n_75)
);

XOR2xp5_ASAP7_75t_L g64 ( 
.A(n_54),
.B(n_28),
.Y(n_64)
);

XOR2xp5_ASAP7_75t_L g82 ( 
.A(n_64),
.B(n_69),
.Y(n_82)
);

AND2x6_ASAP7_75t_L g67 ( 
.A(n_52),
.B(n_1),
.Y(n_67)
);

BUFx12_ASAP7_75t_L g80 ( 
.A(n_67),
.Y(n_80)
);

XOR2xp5_ASAP7_75t_L g69 ( 
.A(n_47),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_71),
.B(n_21),
.Y(n_84)
);

NAND2xp5_ASAP7_75t_L g85 ( 
.A(n_74),
.B(n_21),
.Y(n_85)
);

OAI22xp5_ASAP7_75t_SL g89 ( 
.A1(n_75),
.A2(n_77),
.B1(n_85),
.B2(n_73),
.Y(n_89)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_76),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g77 ( 
.A1(n_65),
.A2(n_50),
.B1(n_57),
.B2(n_61),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g78 ( 
.A(n_70),
.B(n_14),
.Y(n_78)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_78),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g79 ( 
.A(n_63),
.B(n_15),
.Y(n_79)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_79),
.Y(n_92)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_65),
.B(n_10),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g88 ( 
.A(n_81),
.B(n_84),
.Y(n_88)
);

XNOR2xp5_ASAP7_75t_L g83 ( 
.A(n_64),
.B(n_39),
.Y(n_83)
);

MAJIxp5_ASAP7_75t_L g86 ( 
.A(n_83),
.B(n_66),
.C(n_69),
.Y(n_86)
);

XNOR2xp5_ASAP7_75t_L g95 ( 
.A(n_86),
.B(n_91),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g97 ( 
.A(n_89),
.B(n_93),
.Y(n_97)
);

AOI21xp5_ASAP7_75t_L g91 ( 
.A1(n_83),
.A2(n_74),
.B(n_67),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_SL g93 ( 
.A1(n_77),
.A2(n_66),
.B1(n_68),
.B2(n_26),
.Y(n_93)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_87),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_94),
.B(n_96),
.Y(n_100)
);

XOR2xp5_ASAP7_75t_L g96 ( 
.A(n_86),
.B(n_82),
.Y(n_96)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_90),
.Y(n_98)
);

NOR2xp33_ASAP7_75t_L g102 ( 
.A(n_98),
.B(n_76),
.Y(n_102)
);

OAI221xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_88),
.B1(n_93),
.B2(n_82),
.C(n_89),
.Y(n_99)
);

OAI21xp5_ASAP7_75t_L g101 ( 
.A1(n_99),
.A2(n_97),
.B(n_95),
.Y(n_101)
);

MAJIxp5_ASAP7_75t_L g106 ( 
.A(n_101),
.B(n_96),
.C(n_80),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_102),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_L g103 ( 
.A1(n_95),
.A2(n_80),
.B1(n_92),
.B2(n_26),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_103),
.A2(n_80),
.B1(n_2),
.B2(n_3),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g105 ( 
.A(n_100),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g109 ( 
.A(n_105),
.B(n_8),
.Y(n_109)
);

XNOR2xp5_ASAP7_75t_L g108 ( 
.A(n_106),
.B(n_104),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g110 ( 
.A(n_107),
.B(n_1),
.Y(n_110)
);

OAI22xp5_ASAP7_75t_L g111 ( 
.A1(n_108),
.A2(n_109),
.B1(n_110),
.B2(n_106),
.Y(n_111)
);

OAI21xp5_ASAP7_75t_SL g113 ( 
.A1(n_111),
.A2(n_112),
.B(n_2),
.Y(n_113)
);

OAI21xp5_ASAP7_75t_SL g112 ( 
.A1(n_109),
.A2(n_2),
.B(n_3),
.Y(n_112)
);

HAxp5_ASAP7_75t_SL g114 ( 
.A(n_113),
.B(n_3),
.CON(n_114),
.SN(n_114)
);


endmodule