module fake_jpeg_23516_n_34 (n_3, n_2, n_1, n_0, n_4, n_5, n_34);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_5;

output n_34;

wire n_13;
wire n_21;
wire n_33;
wire n_10;
wire n_23;
wire n_27;
wire n_6;
wire n_22;
wire n_14;
wire n_19;
wire n_18;
wire n_20;
wire n_30;
wire n_16;
wire n_24;
wire n_28;
wire n_26;
wire n_9;
wire n_11;
wire n_17;
wire n_25;
wire n_31;
wire n_29;
wire n_12;
wire n_32;
wire n_8;
wire n_15;
wire n_7;

BUFx4f_ASAP7_75t_SL g6 ( 
.A(n_1),
.Y(n_6)
);

INVx4_ASAP7_75t_L g7 ( 
.A(n_0),
.Y(n_7)
);

INVx3_ASAP7_75t_L g8 ( 
.A(n_5),
.Y(n_8)
);

INVx2_ASAP7_75t_L g9 ( 
.A(n_2),
.Y(n_9)
);

BUFx6f_ASAP7_75t_L g10 ( 
.A(n_3),
.Y(n_10)
);

INVx8_ASAP7_75t_L g11 ( 
.A(n_1),
.Y(n_11)
);

INVx6_ASAP7_75t_L g12 ( 
.A(n_5),
.Y(n_12)
);

BUFx6f_ASAP7_75t_L g13 ( 
.A(n_6),
.Y(n_13)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_13),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g14 ( 
.A(n_6),
.Y(n_14)
);

NAND2xp5_ASAP7_75t_L g22 ( 
.A(n_14),
.B(n_15),
.Y(n_22)
);

CKINVDCx14_ASAP7_75t_R g15 ( 
.A(n_6),
.Y(n_15)
);

INVxp67_ASAP7_75t_L g16 ( 
.A(n_8),
.Y(n_16)
);

A2O1A1Ixp33_ASAP7_75t_L g20 ( 
.A1(n_16),
.A2(n_10),
.B(n_9),
.C(n_8),
.Y(n_20)
);

AOI22xp33_ASAP7_75t_L g17 ( 
.A1(n_12),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_17)
);

OAI22xp5_ASAP7_75t_L g23 ( 
.A1(n_17),
.A2(n_12),
.B1(n_11),
.B2(n_7),
.Y(n_23)
);

MAJIxp5_ASAP7_75t_L g18 ( 
.A(n_9),
.B(n_0),
.C(n_2),
.Y(n_18)
);

MAJIxp5_ASAP7_75t_L g21 ( 
.A(n_18),
.B(n_10),
.C(n_4),
.Y(n_21)
);

INVxp67_ASAP7_75t_L g24 ( 
.A(n_20),
.Y(n_24)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_23),
.C(n_18),
.Y(n_25)
);

NAND2xp5_ASAP7_75t_L g28 ( 
.A(n_25),
.B(n_21),
.Y(n_28)
);

NOR2xp33_ASAP7_75t_SL g26 ( 
.A(n_22),
.B(n_3),
.Y(n_26)
);

NOR2xp33_ASAP7_75t_SL g27 ( 
.A(n_26),
.B(n_4),
.Y(n_27)
);

NAND2xp5_ASAP7_75t_SL g30 ( 
.A(n_27),
.B(n_28),
.Y(n_30)
);

AOI22xp5_ASAP7_75t_SL g29 ( 
.A1(n_28),
.A2(n_24),
.B1(n_7),
.B2(n_16),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_SL g31 ( 
.A(n_29),
.B(n_20),
.Y(n_31)
);

OAI21xp5_ASAP7_75t_L g32 ( 
.A1(n_31),
.A2(n_30),
.B(n_29),
.Y(n_32)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_32),
.B(n_13),
.Y(n_33)
);

XNOR2xp5_ASAP7_75t_L g34 ( 
.A(n_33),
.B(n_19),
.Y(n_34)
);


endmodule