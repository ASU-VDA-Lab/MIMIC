module fake_aes_8019_n_716 (n_44, n_69, n_22, n_57, n_52, n_26, n_50, n_33, n_73, n_49, n_60, n_41, n_35, n_65, n_9, n_10, n_19, n_74, n_7, n_29, n_45, n_62, n_36, n_47, n_37, n_34, n_5, n_23, n_8, n_16, n_13, n_70, n_17, n_63, n_14, n_71, n_56, n_42, n_24, n_78, n_6, n_4, n_40, n_38, n_64, n_46, n_31, n_58, n_32, n_0, n_55, n_12, n_75, n_72, n_43, n_76, n_68, n_27, n_53, n_67, n_77, n_20, n_2, n_54, n_28, n_48, n_11, n_25, n_30, n_59, n_3, n_18, n_66, n_1, n_15, n_61, n_21, n_51, n_39, n_716);
input n_44;
input n_69;
input n_22;
input n_57;
input n_52;
input n_26;
input n_50;
input n_33;
input n_73;
input n_49;
input n_60;
input n_41;
input n_35;
input n_65;
input n_9;
input n_10;
input n_19;
input n_74;
input n_7;
input n_29;
input n_45;
input n_62;
input n_36;
input n_47;
input n_37;
input n_34;
input n_5;
input n_23;
input n_8;
input n_16;
input n_13;
input n_70;
input n_17;
input n_63;
input n_14;
input n_71;
input n_56;
input n_42;
input n_24;
input n_78;
input n_6;
input n_4;
input n_40;
input n_38;
input n_64;
input n_46;
input n_31;
input n_58;
input n_32;
input n_0;
input n_55;
input n_12;
input n_75;
input n_72;
input n_43;
input n_76;
input n_68;
input n_27;
input n_53;
input n_67;
input n_77;
input n_20;
input n_2;
input n_54;
input n_28;
input n_48;
input n_11;
input n_25;
input n_30;
input n_59;
input n_3;
input n_18;
input n_66;
input n_1;
input n_15;
input n_61;
input n_21;
input n_51;
input n_39;
output n_716;
wire n_117;
wire n_663;
wire n_707;
wire n_361;
wire n_513;
wire n_185;
wire n_705;
wire n_603;
wire n_604;
wire n_590;
wire n_407;
wire n_646;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_607;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_667;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_701;
wire n_612;
wire n_154;
wire n_328;
wire n_655;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_645;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_637;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_288;
wire n_383;
wire n_661;
wire n_672;
wire n_532;
wire n_627;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_659;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_588;
wire n_275;
wire n_715;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_587;
wire n_662;
wire n_162;
wire n_678;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_617;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_628;
wire n_411;
wire n_598;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_599;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_694;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_609;
wire n_636;
wire n_366;
wire n_596;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_702;
wire n_572;
wire n_324;
wire n_392;
wire n_668;
wire n_652;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_680;
wire n_642;
wire n_586;
wire n_671;
wire n_244;
wire n_540;
wire n_638;
wire n_563;
wire n_119;
wire n_141;
wire n_560;
wire n_517;
wire n_479;
wire n_97;
wire n_167;
wire n_623;
wire n_593;
wire n_697;
wire n_554;
wire n_712;
wire n_447;
wire n_608;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_630;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_692;
wire n_647;
wire n_367;
wire n_644;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_624;
wire n_108;
wire n_91;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_711;
wire n_318;
wire n_471;
wire n_632;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_613;
wire n_648;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_665;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_708;
wire n_191;
wire n_307;
wire n_634;
wire n_610;
wire n_696;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_676;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_235;
wire n_243;
wire n_415;
wire n_394;
wire n_482;
wire n_442;
wire n_331;
wire n_485;
wire n_703;
wire n_352;
wire n_619;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_699;
wire n_693;
wire n_256;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_651;
wire n_674;
wire n_172;
wire n_329;
wire n_251;
wire n_635;
wire n_689;
wire n_525;
wire n_218;
wire n_507;
wire n_605;
wire n_611;
wire n_704;
wire n_633;
wire n_271;
wire n_626;
wire n_302;
wire n_466;
wire n_710;
wire n_270;
wire n_685;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_664;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_660;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_622;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_601;
wire n_87;
wire n_379;
wire n_641;
wire n_614;
wire n_527;
wire n_98;
wire n_649;
wire n_276;
wire n_526;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_420;
wire n_423;
wire n_342;
wire n_446;
wire n_666;
wire n_621;
wire n_370;
wire n_589;
wire n_643;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_687;
wire n_193;
wire n_273;
wire n_505;
wire n_706;
wire n_390;
wire n_682;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_90;
wire n_357;
wire n_653;
wire n_260;
wire n_539;
wire n_201;
wire n_197;
wire n_591;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_673;
wire n_669;
wire n_178;
wire n_616;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_654;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_376;
wire n_639;
wire n_552;
wire n_677;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_520;
wire n_681;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_615;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_656;
wire n_438;
wire n_134;
wire n_640;
wire n_429;
wire n_488;
wire n_233;
wire n_686;
wire n_684;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_679;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_597;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_584;
wire n_497;
wire n_339;
wire n_657;
wire n_583;
wire n_620;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_561;
wire n_335;
wire n_272;
wire n_700;
wire n_594;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_602;
wire n_198;
wire n_169;
wire n_424;
wire n_714;
wire n_629;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_675;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_698;
wire n_380;
wire n_618;
wire n_690;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_600;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_451;
wire n_487;
wire n_371;
wire n_688;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_670;
wire n_84;
wire n_266;
wire n_683;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_592;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_658;
wire n_691;
wire n_444;
wire n_176;
wire n_650;
wire n_625;
wire n_695;
wire n_521;
wire n_469;
wire n_585;
wire n_713;
wire n_123;
wire n_457;
wire n_595;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_631;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_606;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_709;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_132;
wire n_109;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
INVx1_ASAP7_75t_L g79 ( .A(n_14), .Y(n_79) );
CKINVDCx5p33_ASAP7_75t_R g80 ( .A(n_13), .Y(n_80) );
CKINVDCx5p33_ASAP7_75t_R g81 ( .A(n_47), .Y(n_81) );
INVx1_ASAP7_75t_L g82 ( .A(n_28), .Y(n_82) );
NOR2xp67_ASAP7_75t_L g83 ( .A(n_68), .B(n_53), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_2), .Y(n_84) );
CKINVDCx5p33_ASAP7_75t_R g85 ( .A(n_69), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_73), .Y(n_86) );
CKINVDCx5p33_ASAP7_75t_R g87 ( .A(n_54), .Y(n_87) );
INVx2_ASAP7_75t_L g88 ( .A(n_30), .Y(n_88) );
CKINVDCx14_ASAP7_75t_R g89 ( .A(n_1), .Y(n_89) );
INVx2_ASAP7_75t_L g90 ( .A(n_64), .Y(n_90) );
CKINVDCx5p33_ASAP7_75t_R g91 ( .A(n_67), .Y(n_91) );
INVxp33_ASAP7_75t_L g92 ( .A(n_43), .Y(n_92) );
INVx1_ASAP7_75t_L g93 ( .A(n_74), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_63), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_17), .Y(n_95) );
CKINVDCx5p33_ASAP7_75t_R g96 ( .A(n_65), .Y(n_96) );
BUFx6f_ASAP7_75t_L g97 ( .A(n_18), .Y(n_97) );
INVx1_ASAP7_75t_SL g98 ( .A(n_70), .Y(n_98) );
CKINVDCx16_ASAP7_75t_R g99 ( .A(n_44), .Y(n_99) );
HB1xp67_ASAP7_75t_L g100 ( .A(n_75), .Y(n_100) );
INVx1_ASAP7_75t_L g101 ( .A(n_14), .Y(n_101) );
INVx2_ASAP7_75t_L g102 ( .A(n_60), .Y(n_102) );
INVxp67_ASAP7_75t_L g103 ( .A(n_9), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_26), .Y(n_104) );
CKINVDCx20_ASAP7_75t_R g105 ( .A(n_15), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_25), .Y(n_106) );
CKINVDCx5p33_ASAP7_75t_R g107 ( .A(n_27), .Y(n_107) );
BUFx3_ASAP7_75t_L g108 ( .A(n_51), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_12), .Y(n_109) );
INVx2_ASAP7_75t_L g110 ( .A(n_3), .Y(n_110) );
INVx1_ASAP7_75t_SL g111 ( .A(n_62), .Y(n_111) );
INVx1_ASAP7_75t_L g112 ( .A(n_61), .Y(n_112) );
BUFx5_ASAP7_75t_L g113 ( .A(n_32), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_4), .Y(n_114) );
INVx2_ASAP7_75t_L g115 ( .A(n_49), .Y(n_115) );
INVx1_ASAP7_75t_L g116 ( .A(n_10), .Y(n_116) );
INVx1_ASAP7_75t_L g117 ( .A(n_58), .Y(n_117) );
OR2x2_ASAP7_75t_L g118 ( .A(n_66), .B(n_22), .Y(n_118) );
BUFx2_ASAP7_75t_L g119 ( .A(n_56), .Y(n_119) );
BUFx10_ASAP7_75t_L g120 ( .A(n_78), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_48), .Y(n_121) );
CKINVDCx5p33_ASAP7_75t_R g122 ( .A(n_20), .Y(n_122) );
INVx1_ASAP7_75t_L g123 ( .A(n_71), .Y(n_123) );
CKINVDCx20_ASAP7_75t_R g124 ( .A(n_76), .Y(n_124) );
INVx1_ASAP7_75t_L g125 ( .A(n_12), .Y(n_125) );
INVx1_ASAP7_75t_L g126 ( .A(n_6), .Y(n_126) );
CKINVDCx5p33_ASAP7_75t_R g127 ( .A(n_72), .Y(n_127) );
AND2x4_ASAP7_75t_L g128 ( .A(n_110), .B(n_0), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_110), .Y(n_129) );
INVx2_ASAP7_75t_L g130 ( .A(n_113), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_82), .Y(n_131) );
BUFx3_ASAP7_75t_L g132 ( .A(n_108), .Y(n_132) );
INVx3_ASAP7_75t_L g133 ( .A(n_120), .Y(n_133) );
CKINVDCx5p33_ASAP7_75t_R g134 ( .A(n_89), .Y(n_134) );
INVx3_ASAP7_75t_L g135 ( .A(n_120), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_89), .Y(n_136) );
NAND2xp5_ASAP7_75t_L g137 ( .A(n_119), .B(n_0), .Y(n_137) );
AOI22xp5_ASAP7_75t_L g138 ( .A1(n_99), .A2(n_1), .B1(n_2), .B2(n_3), .Y(n_138) );
INVx2_ASAP7_75t_L g139 ( .A(n_113), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_86), .Y(n_140) );
INVx3_ASAP7_75t_L g141 ( .A(n_120), .Y(n_141) );
INVx2_ASAP7_75t_L g142 ( .A(n_113), .Y(n_142) );
NOR2xp33_ASAP7_75t_L g143 ( .A(n_100), .B(n_4), .Y(n_143) );
CKINVDCx5p33_ASAP7_75t_R g144 ( .A(n_124), .Y(n_144) );
BUFx6f_ASAP7_75t_L g145 ( .A(n_97), .Y(n_145) );
OAI22xp5_ASAP7_75t_SL g146 ( .A1(n_105), .A2(n_5), .B1(n_6), .B2(n_7), .Y(n_146) );
INVxp67_ASAP7_75t_L g147 ( .A(n_79), .Y(n_147) );
INVx3_ASAP7_75t_L g148 ( .A(n_84), .Y(n_148) );
INVx1_ASAP7_75t_L g149 ( .A(n_93), .Y(n_149) );
INVx1_ASAP7_75t_L g150 ( .A(n_94), .Y(n_150) );
INVx2_ASAP7_75t_L g151 ( .A(n_113), .Y(n_151) );
INVx6_ASAP7_75t_L g152 ( .A(n_113), .Y(n_152) );
AOI22xp5_ASAP7_75t_L g153 ( .A1(n_124), .A2(n_5), .B1(n_7), .B2(n_8), .Y(n_153) );
NAND2xp5_ASAP7_75t_L g154 ( .A(n_103), .B(n_8), .Y(n_154) );
BUFx2_ASAP7_75t_L g155 ( .A(n_80), .Y(n_155) );
OAI22xp5_ASAP7_75t_L g156 ( .A1(n_92), .A2(n_9), .B1(n_10), .B2(n_11), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_81), .Y(n_157) );
INVx2_ASAP7_75t_L g158 ( .A(n_113), .Y(n_158) );
AOI22xp5_ASAP7_75t_L g159 ( .A1(n_101), .A2(n_11), .B1(n_13), .B2(n_15), .Y(n_159) );
HB1xp67_ASAP7_75t_L g160 ( .A(n_109), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_95), .Y(n_161) );
INVx2_ASAP7_75t_L g162 ( .A(n_113), .Y(n_162) );
INVx1_ASAP7_75t_L g163 ( .A(n_104), .Y(n_163) );
INVx1_ASAP7_75t_L g164 ( .A(n_112), .Y(n_164) );
BUFx6f_ASAP7_75t_L g165 ( .A(n_97), .Y(n_165) );
NOR2x1_ASAP7_75t_L g166 ( .A(n_114), .B(n_16), .Y(n_166) );
INVx1_ASAP7_75t_L g167 ( .A(n_117), .Y(n_167) );
INVx1_ASAP7_75t_L g168 ( .A(n_121), .Y(n_168) );
BUFx6f_ASAP7_75t_L g169 ( .A(n_97), .Y(n_169) );
BUFx6f_ASAP7_75t_L g170 ( .A(n_97), .Y(n_170) );
INVx2_ASAP7_75t_L g171 ( .A(n_88), .Y(n_171) );
BUFx6f_ASAP7_75t_L g172 ( .A(n_145), .Y(n_172) );
INVx1_ASAP7_75t_L g173 ( .A(n_128), .Y(n_173) );
INVx4_ASAP7_75t_L g174 ( .A(n_152), .Y(n_174) );
INVx1_ASAP7_75t_L g175 ( .A(n_128), .Y(n_175) );
INVx6_ASAP7_75t_L g176 ( .A(n_128), .Y(n_176) );
NAND2xp5_ASAP7_75t_SL g177 ( .A(n_131), .B(n_106), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_148), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_133), .B(n_92), .Y(n_179) );
NOR2xp33_ASAP7_75t_L g180 ( .A(n_133), .B(n_106), .Y(n_180) );
OR2x2_ASAP7_75t_L g181 ( .A(n_155), .B(n_116), .Y(n_181) );
INVx2_ASAP7_75t_L g182 ( .A(n_130), .Y(n_182) );
INVx2_ASAP7_75t_L g183 ( .A(n_130), .Y(n_183) );
AND3x2_ASAP7_75t_L g184 ( .A(n_136), .B(n_126), .C(n_125), .Y(n_184) );
BUFx4f_ASAP7_75t_L g185 ( .A(n_133), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_148), .Y(n_186) );
INVx2_ASAP7_75t_L g187 ( .A(n_139), .Y(n_187) );
INVxp33_ASAP7_75t_L g188 ( .A(n_155), .Y(n_188) );
BUFx3_ASAP7_75t_L g189 ( .A(n_132), .Y(n_189) );
AOI22xp33_ASAP7_75t_L g190 ( .A1(n_131), .A2(n_123), .B1(n_102), .B2(n_88), .Y(n_190) );
NAND2xp33_ASAP7_75t_L g191 ( .A(n_134), .B(n_91), .Y(n_191) );
NAND2xp5_ASAP7_75t_L g192 ( .A(n_135), .B(n_127), .Y(n_192) );
INVxp67_ASAP7_75t_SL g193 ( .A(n_160), .Y(n_193) );
BUFx6f_ASAP7_75t_L g194 ( .A(n_145), .Y(n_194) );
NAND2xp5_ASAP7_75t_L g195 ( .A(n_135), .B(n_127), .Y(n_195) );
INVx2_ASAP7_75t_SL g196 ( .A(n_157), .Y(n_196) );
AND2x2_ASAP7_75t_L g197 ( .A(n_135), .B(n_81), .Y(n_197) );
BUFx6f_ASAP7_75t_L g198 ( .A(n_145), .Y(n_198) );
INVx2_ASAP7_75t_L g199 ( .A(n_139), .Y(n_199) );
NAND2xp5_ASAP7_75t_SL g200 ( .A(n_140), .B(n_102), .Y(n_200) );
INVx2_ASAP7_75t_L g201 ( .A(n_132), .Y(n_201) );
INVx2_ASAP7_75t_L g202 ( .A(n_152), .Y(n_202) );
AND2x6_ASAP7_75t_L g203 ( .A(n_166), .B(n_108), .Y(n_203) );
NAND2xp33_ASAP7_75t_L g204 ( .A(n_134), .B(n_107), .Y(n_204) );
NAND2xp5_ASAP7_75t_L g205 ( .A(n_141), .B(n_85), .Y(n_205) );
INVx2_ASAP7_75t_L g206 ( .A(n_152), .Y(n_206) );
INVx1_ASAP7_75t_L g207 ( .A(n_148), .Y(n_207) );
AND2x2_ASAP7_75t_L g208 ( .A(n_141), .B(n_85), .Y(n_208) );
INVx3_ASAP7_75t_L g209 ( .A(n_141), .Y(n_209) );
INVx2_ASAP7_75t_SL g210 ( .A(n_157), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_140), .B(n_122), .Y(n_211) );
OR2x2_ASAP7_75t_L g212 ( .A(n_147), .B(n_122), .Y(n_212) );
BUFx4f_ASAP7_75t_L g213 ( .A(n_152), .Y(n_213) );
NAND2xp33_ASAP7_75t_L g214 ( .A(n_149), .B(n_96), .Y(n_214) );
NAND2xp5_ASAP7_75t_L g215 ( .A(n_149), .B(n_87), .Y(n_215) );
INVxp67_ASAP7_75t_L g216 ( .A(n_137), .Y(n_216) );
INVx4_ASAP7_75t_L g217 ( .A(n_142), .Y(n_217) );
INVx2_ASAP7_75t_L g218 ( .A(n_171), .Y(n_218) );
INVx4_ASAP7_75t_L g219 ( .A(n_142), .Y(n_219) );
BUFx6f_ASAP7_75t_L g220 ( .A(n_145), .Y(n_220) );
INVx2_ASAP7_75t_L g221 ( .A(n_151), .Y(n_221) );
NOR2xp33_ASAP7_75t_L g222 ( .A(n_150), .B(n_115), .Y(n_222) );
AND2x4_ASAP7_75t_L g223 ( .A(n_150), .B(n_115), .Y(n_223) );
BUFx6f_ASAP7_75t_L g224 ( .A(n_145), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_165), .Y(n_225) );
AOI22xp33_ASAP7_75t_L g226 ( .A1(n_161), .A2(n_90), .B1(n_118), .B2(n_98), .Y(n_226) );
INVx1_ASAP7_75t_L g227 ( .A(n_171), .Y(n_227) );
INVx4_ASAP7_75t_SL g228 ( .A(n_165), .Y(n_228) );
NOR2xp33_ASAP7_75t_L g229 ( .A(n_161), .B(n_90), .Y(n_229) );
CKINVDCx20_ASAP7_75t_R g230 ( .A(n_144), .Y(n_230) );
INVx1_ASAP7_75t_L g231 ( .A(n_129), .Y(n_231) );
NAND2xp5_ASAP7_75t_L g232 ( .A(n_163), .B(n_87), .Y(n_232) );
INVx1_ASAP7_75t_L g233 ( .A(n_129), .Y(n_233) );
OR2x2_ASAP7_75t_L g234 ( .A(n_163), .B(n_111), .Y(n_234) );
BUFx2_ASAP7_75t_L g235 ( .A(n_144), .Y(n_235) );
NAND2xp5_ASAP7_75t_SL g236 ( .A(n_164), .B(n_83), .Y(n_236) );
CKINVDCx20_ASAP7_75t_R g237 ( .A(n_146), .Y(n_237) );
OR2x2_ASAP7_75t_L g238 ( .A(n_193), .B(n_154), .Y(n_238) );
NAND2xp5_ASAP7_75t_SL g239 ( .A(n_216), .B(n_143), .Y(n_239) );
INVx4_ASAP7_75t_L g240 ( .A(n_174), .Y(n_240) );
INVx2_ASAP7_75t_L g241 ( .A(n_189), .Y(n_241) );
OAI21xp5_ASAP7_75t_L g242 ( .A1(n_182), .A2(n_158), .B(n_151), .Y(n_242) );
INVx1_ASAP7_75t_L g243 ( .A(n_186), .Y(n_243) );
NOR2xp33_ASAP7_75t_L g244 ( .A(n_216), .B(n_168), .Y(n_244) );
AOI21xp5_ASAP7_75t_L g245 ( .A1(n_192), .A2(n_162), .B(n_158), .Y(n_245) );
NAND2xp5_ASAP7_75t_SL g246 ( .A(n_217), .B(n_162), .Y(n_246) );
NOR2xp33_ASAP7_75t_L g247 ( .A(n_195), .B(n_164), .Y(n_247) );
NAND2xp5_ASAP7_75t_L g248 ( .A(n_179), .B(n_168), .Y(n_248) );
INVx1_ASAP7_75t_L g249 ( .A(n_186), .Y(n_249) );
BUFx8_ASAP7_75t_L g250 ( .A(n_235), .Y(n_250) );
INVx2_ASAP7_75t_L g251 ( .A(n_189), .Y(n_251) );
AOI22xp5_ASAP7_75t_L g252 ( .A1(n_193), .A2(n_156), .B1(n_138), .B2(n_153), .Y(n_252) );
INVx1_ASAP7_75t_L g253 ( .A(n_178), .Y(n_253) );
CKINVDCx5p33_ASAP7_75t_R g254 ( .A(n_230), .Y(n_254) );
NOR2xp33_ASAP7_75t_L g255 ( .A(n_205), .B(n_167), .Y(n_255) );
INVx3_ASAP7_75t_L g256 ( .A(n_209), .Y(n_256) );
NAND2xp5_ASAP7_75t_L g257 ( .A(n_179), .B(n_167), .Y(n_257) );
INVxp67_ASAP7_75t_L g258 ( .A(n_212), .Y(n_258) );
BUFx3_ASAP7_75t_L g259 ( .A(n_201), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_207), .Y(n_260) );
INVx1_ASAP7_75t_SL g261 ( .A(n_188), .Y(n_261) );
AOI22xp33_ASAP7_75t_L g262 ( .A1(n_173), .A2(n_159), .B1(n_170), .B2(n_165), .Y(n_262) );
BUFx6f_ASAP7_75t_L g263 ( .A(n_218), .Y(n_263) );
NAND2xp5_ASAP7_75t_L g264 ( .A(n_211), .B(n_215), .Y(n_264) );
AOI22xp5_ASAP7_75t_L g265 ( .A1(n_226), .A2(n_105), .B1(n_169), .B2(n_165), .Y(n_265) );
NAND2xp5_ASAP7_75t_SL g266 ( .A(n_217), .B(n_169), .Y(n_266) );
HB1xp67_ASAP7_75t_L g267 ( .A(n_188), .Y(n_267) );
INVx1_ASAP7_75t_L g268 ( .A(n_176), .Y(n_268) );
NOR2x2_ASAP7_75t_L g269 ( .A(n_237), .B(n_19), .Y(n_269) );
AOI22xp33_ASAP7_75t_L g270 ( .A1(n_175), .A2(n_170), .B1(n_169), .B2(n_165), .Y(n_270) );
NAND2xp5_ASAP7_75t_L g271 ( .A(n_232), .B(n_169), .Y(n_271) );
NAND2xp5_ASAP7_75t_SL g272 ( .A(n_219), .B(n_169), .Y(n_272) );
NAND2xp5_ASAP7_75t_L g273 ( .A(n_197), .B(n_170), .Y(n_273) );
INVx1_ASAP7_75t_L g274 ( .A(n_176), .Y(n_274) );
A2O1A1Ixp33_ASAP7_75t_L g275 ( .A1(n_222), .A2(n_170), .B(n_23), .C(n_24), .Y(n_275) );
INVx2_ASAP7_75t_L g276 ( .A(n_209), .Y(n_276) );
AND2x2_ASAP7_75t_L g277 ( .A(n_181), .B(n_170), .Y(n_277) );
INVx2_ASAP7_75t_SL g278 ( .A(n_208), .Y(n_278) );
INVx2_ASAP7_75t_L g279 ( .A(n_231), .Y(n_279) );
NAND2xp5_ASAP7_75t_SL g280 ( .A(n_219), .B(n_21), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_233), .Y(n_281) );
NAND2xp5_ASAP7_75t_SL g282 ( .A(n_182), .B(n_29), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g283 ( .A(n_234), .B(n_31), .Y(n_283) );
INVx1_ASAP7_75t_SL g284 ( .A(n_196), .Y(n_284) );
BUFx4f_ASAP7_75t_L g285 ( .A(n_210), .Y(n_285) );
OAI22xp5_ASAP7_75t_L g286 ( .A1(n_176), .A2(n_33), .B1(n_34), .B2(n_35), .Y(n_286) );
NOR2xp33_ASAP7_75t_L g287 ( .A(n_185), .B(n_36), .Y(n_287) );
INVx1_ASAP7_75t_L g288 ( .A(n_227), .Y(n_288) );
AOI22xp33_ASAP7_75t_L g289 ( .A1(n_223), .A2(n_37), .B1(n_38), .B2(n_39), .Y(n_289) );
INVx2_ASAP7_75t_L g290 ( .A(n_183), .Y(n_290) );
AOI22xp5_ASAP7_75t_L g291 ( .A1(n_226), .A2(n_40), .B1(n_41), .B2(n_42), .Y(n_291) );
AND3x1_ASAP7_75t_L g292 ( .A(n_190), .B(n_45), .C(n_46), .Y(n_292) );
OAI22xp5_ASAP7_75t_L g293 ( .A1(n_190), .A2(n_50), .B1(n_52), .B2(n_55), .Y(n_293) );
AO22x1_ASAP7_75t_L g294 ( .A1(n_203), .A2(n_57), .B1(n_59), .B2(n_77), .Y(n_294) );
BUFx3_ASAP7_75t_L g295 ( .A(n_185), .Y(n_295) );
INVx1_ASAP7_75t_L g296 ( .A(n_223), .Y(n_296) );
NOR2xp33_ASAP7_75t_L g297 ( .A(n_214), .B(n_180), .Y(n_297) );
NAND2xp5_ASAP7_75t_L g298 ( .A(n_180), .B(n_229), .Y(n_298) );
INVx1_ASAP7_75t_SL g299 ( .A(n_184), .Y(n_299) );
NAND2xp5_ASAP7_75t_SL g300 ( .A(n_183), .B(n_221), .Y(n_300) );
INVx1_ASAP7_75t_L g301 ( .A(n_177), .Y(n_301) );
AOI22xp33_ASAP7_75t_L g302 ( .A1(n_222), .A2(n_229), .B1(n_203), .B2(n_177), .Y(n_302) );
NAND2xp5_ASAP7_75t_L g303 ( .A(n_203), .B(n_174), .Y(n_303) );
NAND2xp5_ASAP7_75t_L g304 ( .A(n_203), .B(n_236), .Y(n_304) );
INVx2_ASAP7_75t_SL g305 ( .A(n_184), .Y(n_305) );
INVx1_ASAP7_75t_L g306 ( .A(n_200), .Y(n_306) );
O2A1O1Ixp33_ASAP7_75t_L g307 ( .A1(n_200), .A2(n_204), .B(n_191), .C(n_236), .Y(n_307) );
OAI22xp5_ASAP7_75t_L g308 ( .A1(n_248), .A2(n_187), .B1(n_221), .B2(n_199), .Y(n_308) );
NOR2xp33_ASAP7_75t_R g309 ( .A(n_254), .B(n_203), .Y(n_309) );
NAND2x1p5_ASAP7_75t_L g310 ( .A(n_240), .B(n_213), .Y(n_310) );
INVx3_ASAP7_75t_SL g311 ( .A(n_261), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_264), .A2(n_213), .B(n_206), .Y(n_312) );
OAI22xp5_ASAP7_75t_L g313 ( .A1(n_257), .A2(n_252), .B1(n_265), .B2(n_298), .Y(n_313) );
HB1xp67_ASAP7_75t_L g314 ( .A(n_267), .Y(n_314) );
NOR2xp33_ASAP7_75t_R g315 ( .A(n_250), .B(n_187), .Y(n_315) );
AND2x4_ASAP7_75t_L g316 ( .A(n_278), .B(n_202), .Y(n_316) );
OAI21xp5_ASAP7_75t_L g317 ( .A1(n_245), .A2(n_199), .B(n_228), .Y(n_317) );
NOR2xp33_ASAP7_75t_L g318 ( .A(n_258), .B(n_172), .Y(n_318) );
INVx1_ASAP7_75t_SL g319 ( .A(n_267), .Y(n_319) );
AOI21xp5_ASAP7_75t_L g320 ( .A1(n_300), .A2(n_172), .B(n_194), .Y(n_320) );
BUFx12f_ASAP7_75t_L g321 ( .A(n_250), .Y(n_321) );
BUFx2_ASAP7_75t_L g322 ( .A(n_284), .Y(n_322) );
AOI22xp33_ASAP7_75t_L g323 ( .A1(n_244), .A2(n_172), .B1(n_194), .B2(n_198), .Y(n_323) );
INVx2_ASAP7_75t_L g324 ( .A(n_263), .Y(n_324) );
NAND2xp5_ASAP7_75t_SL g325 ( .A(n_238), .B(n_228), .Y(n_325) );
BUFx2_ASAP7_75t_L g326 ( .A(n_285), .Y(n_326) );
AOI21xp5_ASAP7_75t_L g327 ( .A1(n_300), .A2(n_172), .B(n_194), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_244), .B(n_228), .Y(n_328) );
O2A1O1Ixp33_ASAP7_75t_L g329 ( .A1(n_239), .A2(n_194), .B(n_198), .C(n_220), .Y(n_329) );
NAND2xp5_ASAP7_75t_L g330 ( .A(n_247), .B(n_198), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_277), .Y(n_331) );
O2A1O1Ixp33_ASAP7_75t_L g332 ( .A1(n_296), .A2(n_198), .B(n_220), .C(n_224), .Y(n_332) );
INVx1_ASAP7_75t_L g333 ( .A(n_253), .Y(n_333) );
AOI21xp5_ASAP7_75t_L g334 ( .A1(n_273), .A2(n_225), .B(n_220), .Y(n_334) );
INVx3_ASAP7_75t_SL g335 ( .A(n_269), .Y(n_335) );
NAND2xp5_ASAP7_75t_L g336 ( .A(n_247), .B(n_220), .Y(n_336) );
AOI21xp5_ASAP7_75t_L g337 ( .A1(n_246), .A2(n_224), .B(n_225), .Y(n_337) );
A2O1A1Ixp33_ASAP7_75t_SL g338 ( .A1(n_287), .A2(n_224), .B(n_225), .C(n_297), .Y(n_338) );
AND2x4_ASAP7_75t_L g339 ( .A(n_295), .B(n_224), .Y(n_339) );
A2O1A1Ixp33_ASAP7_75t_L g340 ( .A1(n_255), .A2(n_225), .B(n_297), .C(n_281), .Y(n_340) );
INVx2_ASAP7_75t_L g341 ( .A(n_263), .Y(n_341) );
AOI21xp5_ASAP7_75t_L g342 ( .A1(n_246), .A2(n_255), .B(n_271), .Y(n_342) );
BUFx12f_ASAP7_75t_L g343 ( .A(n_305), .Y(n_343) );
AND2x2_ASAP7_75t_L g344 ( .A(n_285), .B(n_299), .Y(n_344) );
OR2x2_ASAP7_75t_L g345 ( .A(n_262), .B(n_304), .Y(n_345) );
AO32x1_ASAP7_75t_L g346 ( .A1(n_293), .A2(n_286), .A3(n_292), .B1(n_241), .B2(n_251), .Y(n_346) );
INVx2_ASAP7_75t_L g347 ( .A(n_263), .Y(n_347) );
INVx3_ASAP7_75t_SL g348 ( .A(n_240), .Y(n_348) );
AOI21xp5_ASAP7_75t_L g349 ( .A1(n_303), .A2(n_260), .B(n_242), .Y(n_349) );
BUFx2_ASAP7_75t_L g350 ( .A(n_256), .Y(n_350) );
AOI21xp5_ASAP7_75t_L g351 ( .A1(n_301), .A2(n_306), .B(n_272), .Y(n_351) );
AO22x1_ASAP7_75t_L g352 ( .A1(n_287), .A2(n_283), .B1(n_256), .B2(n_274), .Y(n_352) );
NOR2xp33_ASAP7_75t_R g353 ( .A(n_268), .B(n_262), .Y(n_353) );
NOR3xp33_ASAP7_75t_L g354 ( .A(n_307), .B(n_294), .C(n_249), .Y(n_354) );
BUFx2_ASAP7_75t_L g355 ( .A(n_288), .Y(n_355) );
NAND2xp5_ASAP7_75t_L g356 ( .A(n_279), .B(n_302), .Y(n_356) );
NOR2xp33_ASAP7_75t_L g357 ( .A(n_243), .B(n_276), .Y(n_357) );
NAND2xp5_ASAP7_75t_SL g358 ( .A(n_302), .B(n_291), .Y(n_358) );
NAND2xp5_ASAP7_75t_L g359 ( .A(n_259), .B(n_290), .Y(n_359) );
NAND2xp5_ASAP7_75t_L g360 ( .A(n_263), .B(n_289), .Y(n_360) );
OAI22xp5_ASAP7_75t_L g361 ( .A1(n_289), .A2(n_280), .B1(n_270), .B2(n_275), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_313), .A2(n_280), .B1(n_272), .B2(n_266), .Y(n_362) );
INVx4_ASAP7_75t_L g363 ( .A(n_311), .Y(n_363) );
AOI21xp33_ASAP7_75t_L g364 ( .A1(n_313), .A2(n_266), .B(n_282), .Y(n_364) );
NAND2xp5_ASAP7_75t_L g365 ( .A(n_319), .B(n_282), .Y(n_365) );
INVx1_ASAP7_75t_L g366 ( .A(n_314), .Y(n_366) );
INVx1_ASAP7_75t_L g367 ( .A(n_333), .Y(n_367) );
OAI21xp5_ASAP7_75t_L g368 ( .A1(n_342), .A2(n_270), .B(n_349), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_358), .A2(n_351), .B(n_360), .Y(n_369) );
INVx1_ASAP7_75t_L g370 ( .A(n_355), .Y(n_370) );
INVx1_ASAP7_75t_L g371 ( .A(n_319), .Y(n_371) );
OAI21x1_ASAP7_75t_L g372 ( .A1(n_320), .A2(n_327), .B(n_317), .Y(n_372) );
OAI21xp5_ASAP7_75t_L g373 ( .A1(n_340), .A2(n_308), .B(n_330), .Y(n_373) );
INVx1_ASAP7_75t_L g374 ( .A(n_331), .Y(n_374) );
INVx2_ASAP7_75t_SL g375 ( .A(n_315), .Y(n_375) );
AO32x2_ASAP7_75t_L g376 ( .A1(n_361), .A2(n_308), .A3(n_346), .B1(n_338), .B2(n_354), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_322), .A2(n_316), .B1(n_335), .B2(n_356), .C(n_344), .Y(n_377) );
AOI22xp5_ASAP7_75t_L g378 ( .A1(n_326), .A2(n_343), .B1(n_348), .B2(n_316), .Y(n_378) );
INVx1_ASAP7_75t_L g379 ( .A(n_318), .Y(n_379) );
A2O1A1Ixp33_ASAP7_75t_L g380 ( .A1(n_345), .A2(n_360), .B(n_312), .C(n_330), .Y(n_380) );
NOR2xp33_ASAP7_75t_L g381 ( .A(n_350), .B(n_357), .Y(n_381) );
AOI22xp5_ASAP7_75t_L g382 ( .A1(n_359), .A2(n_321), .B1(n_325), .B2(n_361), .Y(n_382) );
INVx1_ASAP7_75t_SL g383 ( .A(n_309), .Y(n_383) );
AOI31xp67_ASAP7_75t_L g384 ( .A1(n_324), .A2(n_347), .A3(n_341), .B(n_336), .Y(n_384) );
NOR2xp33_ASAP7_75t_SL g385 ( .A(n_310), .B(n_328), .Y(n_385) );
CKINVDCx20_ASAP7_75t_R g386 ( .A(n_353), .Y(n_386) );
INVx1_ASAP7_75t_SL g387 ( .A(n_328), .Y(n_387) );
A2O1A1Ixp33_ASAP7_75t_L g388 ( .A1(n_329), .A2(n_317), .B(n_334), .C(n_332), .Y(n_388) );
BUFx3_ASAP7_75t_L g389 ( .A(n_339), .Y(n_389) );
BUFx12f_ASAP7_75t_L g390 ( .A(n_310), .Y(n_390) );
BUFx3_ASAP7_75t_L g391 ( .A(n_339), .Y(n_391) );
INVx1_ASAP7_75t_L g392 ( .A(n_346), .Y(n_392) );
OAI21x1_ASAP7_75t_L g393 ( .A1(n_337), .A2(n_323), .B(n_352), .Y(n_393) );
OAI21x1_ASAP7_75t_L g394 ( .A1(n_346), .A2(n_327), .B(n_320), .Y(n_394) );
INVx2_ASAP7_75t_L g395 ( .A(n_384), .Y(n_395) );
AOI21xp5_ASAP7_75t_L g396 ( .A1(n_369), .A2(n_364), .B(n_388), .Y(n_396) );
OA21x2_ASAP7_75t_L g397 ( .A1(n_394), .A2(n_392), .B(n_380), .Y(n_397) );
OA21x2_ASAP7_75t_L g398 ( .A1(n_380), .A2(n_372), .B(n_373), .Y(n_398) );
NAND2xp5_ASAP7_75t_L g399 ( .A(n_367), .B(n_374), .Y(n_399) );
INVx1_ASAP7_75t_L g400 ( .A(n_371), .Y(n_400) );
INVx1_ASAP7_75t_L g401 ( .A(n_379), .Y(n_401) );
AOI222xp33_ASAP7_75t_L g402 ( .A1(n_377), .A2(n_370), .B1(n_366), .B2(n_381), .C1(n_375), .C2(n_386), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_381), .B(n_387), .Y(n_403) );
AND2x2_ASAP7_75t_L g404 ( .A(n_382), .B(n_389), .Y(n_404) );
A2O1A1Ixp33_ASAP7_75t_L g405 ( .A1(n_365), .A2(n_362), .B(n_388), .C(n_368), .Y(n_405) );
INVx2_ASAP7_75t_L g406 ( .A(n_376), .Y(n_406) );
AOI22xp5_ASAP7_75t_L g407 ( .A1(n_386), .A2(n_385), .B1(n_363), .B2(n_390), .Y(n_407) );
NAND2xp5_ASAP7_75t_L g408 ( .A(n_378), .B(n_389), .Y(n_408) );
NAND2xp5_ASAP7_75t_L g409 ( .A(n_391), .B(n_383), .Y(n_409) );
OA21x2_ASAP7_75t_L g410 ( .A1(n_393), .A2(n_362), .B(n_376), .Y(n_410) );
OAI21x1_ASAP7_75t_L g411 ( .A1(n_376), .A2(n_391), .B(n_363), .Y(n_411) );
AOI21xp5_ASAP7_75t_L g412 ( .A1(n_376), .A2(n_369), .B(n_364), .Y(n_412) );
AOI21xp5_ASAP7_75t_L g413 ( .A1(n_369), .A2(n_364), .B(n_388), .Y(n_413) );
OA21x2_ASAP7_75t_L g414 ( .A1(n_394), .A2(n_392), .B(n_369), .Y(n_414) );
INVx2_ASAP7_75t_L g415 ( .A(n_384), .Y(n_415) );
AOI21xp5_ASAP7_75t_L g416 ( .A1(n_369), .A2(n_364), .B(n_388), .Y(n_416) );
AOI221xp5_ASAP7_75t_L g417 ( .A1(n_377), .A2(n_258), .B1(n_193), .B2(n_244), .C(n_313), .Y(n_417) );
OR2x6_ASAP7_75t_L g418 ( .A(n_390), .B(n_389), .Y(n_418) );
NAND2xp5_ASAP7_75t_SL g419 ( .A(n_363), .B(n_322), .Y(n_419) );
AO31x2_ASAP7_75t_L g420 ( .A1(n_380), .A2(n_392), .A3(n_369), .B(n_388), .Y(n_420) );
NAND2xp5_ASAP7_75t_L g421 ( .A(n_367), .B(n_193), .Y(n_421) );
OAI221xp5_ASAP7_75t_L g422 ( .A1(n_377), .A2(n_252), .B1(n_258), .B2(n_235), .C(n_261), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_367), .Y(n_423) );
INVx2_ASAP7_75t_L g424 ( .A(n_395), .Y(n_424) );
AOI322xp5_ASAP7_75t_L g425 ( .A1(n_417), .A2(n_407), .A3(n_401), .B1(n_423), .B2(n_403), .C1(n_399), .C2(n_419), .Y(n_425) );
OR2x2_ASAP7_75t_L g426 ( .A(n_401), .B(n_423), .Y(n_426) );
INVx2_ASAP7_75t_L g427 ( .A(n_395), .Y(n_427) );
INVx3_ASAP7_75t_L g428 ( .A(n_398), .Y(n_428) );
OA21x2_ASAP7_75t_L g429 ( .A1(n_396), .A2(n_413), .B(n_416), .Y(n_429) );
INVx2_ASAP7_75t_L g430 ( .A(n_415), .Y(n_430) );
INVx2_ASAP7_75t_L g431 ( .A(n_415), .Y(n_431) );
INVx2_ASAP7_75t_L g432 ( .A(n_414), .Y(n_432) );
INVx1_ASAP7_75t_L g433 ( .A(n_400), .Y(n_433) );
INVx1_ASAP7_75t_L g434 ( .A(n_400), .Y(n_434) );
INVx1_ASAP7_75t_L g435 ( .A(n_420), .Y(n_435) );
INVx1_ASAP7_75t_L g436 ( .A(n_420), .Y(n_436) );
AND2x2_ASAP7_75t_L g437 ( .A(n_404), .B(n_406), .Y(n_437) );
INVx4_ASAP7_75t_L g438 ( .A(n_418), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_414), .Y(n_439) );
AOI22xp33_ASAP7_75t_SL g440 ( .A1(n_403), .A2(n_422), .B1(n_404), .B2(n_408), .Y(n_440) );
AND2x2_ASAP7_75t_L g441 ( .A(n_406), .B(n_398), .Y(n_441) );
INVx1_ASAP7_75t_L g442 ( .A(n_420), .Y(n_442) );
AND2x2_ASAP7_75t_L g443 ( .A(n_398), .B(n_420), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_398), .B(n_420), .Y(n_444) );
OR2x2_ASAP7_75t_L g445 ( .A(n_405), .B(n_411), .Y(n_445) );
INVx2_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
OR2x2_ASAP7_75t_L g447 ( .A(n_411), .B(n_397), .Y(n_447) );
OAI21x1_ASAP7_75t_L g448 ( .A1(n_412), .A2(n_397), .B(n_414), .Y(n_448) );
INVx1_ASAP7_75t_L g449 ( .A(n_397), .Y(n_449) );
OR2x2_ASAP7_75t_L g450 ( .A(n_397), .B(n_410), .Y(n_450) );
INVx1_ASAP7_75t_L g451 ( .A(n_410), .Y(n_451) );
AND2x4_ASAP7_75t_L g452 ( .A(n_407), .B(n_418), .Y(n_452) );
INVx3_ASAP7_75t_L g453 ( .A(n_410), .Y(n_453) );
BUFx2_ASAP7_75t_L g454 ( .A(n_418), .Y(n_454) );
INVx1_ASAP7_75t_L g455 ( .A(n_410), .Y(n_455) );
AND2x4_ASAP7_75t_L g456 ( .A(n_418), .B(n_409), .Y(n_456) );
OA21x2_ASAP7_75t_L g457 ( .A1(n_421), .A2(n_402), .B(n_418), .Y(n_457) );
AO21x2_ASAP7_75t_L g458 ( .A1(n_402), .A2(n_412), .B(n_396), .Y(n_458) );
INVx2_ASAP7_75t_L g459 ( .A(n_395), .Y(n_459) );
INVx1_ASAP7_75t_L g460 ( .A(n_424), .Y(n_460) );
AND2x2_ASAP7_75t_L g461 ( .A(n_437), .B(n_443), .Y(n_461) );
INVxp67_ASAP7_75t_SL g462 ( .A(n_426), .Y(n_462) );
AND2x2_ASAP7_75t_L g463 ( .A(n_437), .B(n_443), .Y(n_463) );
INVx1_ASAP7_75t_L g464 ( .A(n_424), .Y(n_464) );
OR2x2_ASAP7_75t_L g465 ( .A(n_437), .B(n_458), .Y(n_465) );
INVxp67_ASAP7_75t_SL g466 ( .A(n_426), .Y(n_466) );
INVx1_ASAP7_75t_L g467 ( .A(n_424), .Y(n_467) );
AND2x2_ASAP7_75t_L g468 ( .A(n_443), .B(n_444), .Y(n_468) );
INVx1_ASAP7_75t_L g469 ( .A(n_426), .Y(n_469) );
BUFx6f_ASAP7_75t_L g470 ( .A(n_432), .Y(n_470) );
AND2x4_ASAP7_75t_L g471 ( .A(n_452), .B(n_438), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_433), .Y(n_472) );
INVx1_ASAP7_75t_L g473 ( .A(n_427), .Y(n_473) );
AND2x2_ASAP7_75t_L g474 ( .A(n_444), .B(n_458), .Y(n_474) );
AND2x4_ASAP7_75t_L g475 ( .A(n_452), .B(n_438), .Y(n_475) );
BUFx6f_ASAP7_75t_L g476 ( .A(n_432), .Y(n_476) );
INVx1_ASAP7_75t_L g477 ( .A(n_427), .Y(n_477) );
INVx1_ASAP7_75t_L g478 ( .A(n_430), .Y(n_478) );
AND2x2_ASAP7_75t_L g479 ( .A(n_444), .B(n_458), .Y(n_479) );
OAI22xp5_ASAP7_75t_L g480 ( .A1(n_440), .A2(n_457), .B1(n_438), .B2(n_452), .Y(n_480) );
AND2x4_ASAP7_75t_L g481 ( .A(n_452), .B(n_438), .Y(n_481) );
NOR2xp33_ASAP7_75t_L g482 ( .A(n_452), .B(n_456), .Y(n_482) );
INVx1_ASAP7_75t_SL g483 ( .A(n_454), .Y(n_483) );
AND2x2_ASAP7_75t_L g484 ( .A(n_458), .B(n_434), .Y(n_484) );
AND2x2_ASAP7_75t_L g485 ( .A(n_433), .B(n_434), .Y(n_485) );
INVx1_ASAP7_75t_L g486 ( .A(n_454), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_441), .B(n_436), .Y(n_487) );
NAND2xp5_ASAP7_75t_L g488 ( .A(n_425), .B(n_440), .Y(n_488) );
INVxp67_ASAP7_75t_SL g489 ( .A(n_457), .Y(n_489) );
AND2x2_ASAP7_75t_L g490 ( .A(n_441), .B(n_442), .Y(n_490) );
INVx3_ASAP7_75t_L g491 ( .A(n_428), .Y(n_491) );
INVx1_ASAP7_75t_L g492 ( .A(n_431), .Y(n_492) );
AND2x2_ASAP7_75t_L g493 ( .A(n_441), .B(n_442), .Y(n_493) );
AND2x2_ASAP7_75t_L g494 ( .A(n_435), .B(n_436), .Y(n_494) );
NAND2xp5_ASAP7_75t_L g495 ( .A(n_425), .B(n_457), .Y(n_495) );
INVx1_ASAP7_75t_SL g496 ( .A(n_456), .Y(n_496) );
OR2x2_ASAP7_75t_L g497 ( .A(n_457), .B(n_435), .Y(n_497) );
BUFx3_ASAP7_75t_L g498 ( .A(n_456), .Y(n_498) );
INVx1_ASAP7_75t_L g499 ( .A(n_431), .Y(n_499) );
HB1xp67_ASAP7_75t_L g500 ( .A(n_456), .Y(n_500) );
BUFx2_ASAP7_75t_L g501 ( .A(n_456), .Y(n_501) );
AND2x4_ASAP7_75t_L g502 ( .A(n_428), .B(n_453), .Y(n_502) );
AND2x4_ASAP7_75t_L g503 ( .A(n_428), .B(n_453), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_431), .Y(n_504) );
AOI221xp5_ASAP7_75t_L g505 ( .A1(n_428), .A2(n_455), .B1(n_451), .B2(n_453), .C(n_449), .Y(n_505) );
INVx5_ASAP7_75t_SL g506 ( .A(n_459), .Y(n_506) );
AND2x2_ASAP7_75t_L g507 ( .A(n_468), .B(n_453), .Y(n_507) );
AND2x2_ASAP7_75t_L g508 ( .A(n_468), .B(n_455), .Y(n_508) );
AND2x2_ASAP7_75t_L g509 ( .A(n_461), .B(n_451), .Y(n_509) );
NAND2xp5_ASAP7_75t_L g510 ( .A(n_462), .B(n_457), .Y(n_510) );
INVx1_ASAP7_75t_L g511 ( .A(n_472), .Y(n_511) );
AND2x2_ASAP7_75t_L g512 ( .A(n_474), .B(n_449), .Y(n_512) );
INVx1_ASAP7_75t_L g513 ( .A(n_485), .Y(n_513) );
INVx1_ASAP7_75t_L g514 ( .A(n_485), .Y(n_514) );
INVx1_ASAP7_75t_L g515 ( .A(n_460), .Y(n_515) );
AND2x2_ASAP7_75t_L g516 ( .A(n_461), .B(n_445), .Y(n_516) );
AND2x2_ASAP7_75t_L g517 ( .A(n_463), .B(n_445), .Y(n_517) );
AND2x2_ASAP7_75t_L g518 ( .A(n_474), .B(n_445), .Y(n_518) );
OR2x2_ASAP7_75t_L g519 ( .A(n_465), .B(n_450), .Y(n_519) );
INVx1_ASAP7_75t_L g520 ( .A(n_460), .Y(n_520) );
INVx2_ASAP7_75t_L g521 ( .A(n_470), .Y(n_521) );
AND2x2_ASAP7_75t_L g522 ( .A(n_463), .B(n_450), .Y(n_522) );
AND2x2_ASAP7_75t_L g523 ( .A(n_479), .B(n_450), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_464), .Y(n_524) );
INVx1_ASAP7_75t_L g525 ( .A(n_464), .Y(n_525) );
INVx2_ASAP7_75t_L g526 ( .A(n_470), .Y(n_526) );
AND2x2_ASAP7_75t_L g527 ( .A(n_479), .B(n_459), .Y(n_527) );
AND2x2_ASAP7_75t_L g528 ( .A(n_487), .B(n_429), .Y(n_528) );
INVxp67_ASAP7_75t_SL g529 ( .A(n_470), .Y(n_529) );
INVx1_ASAP7_75t_L g530 ( .A(n_467), .Y(n_530) );
INVxp67_ASAP7_75t_L g531 ( .A(n_484), .Y(n_531) );
AND2x2_ASAP7_75t_L g532 ( .A(n_487), .B(n_429), .Y(n_532) );
OAI22xp33_ASAP7_75t_L g533 ( .A1(n_488), .A2(n_447), .B1(n_439), .B2(n_446), .Y(n_533) );
INVx1_ASAP7_75t_L g534 ( .A(n_467), .Y(n_534) );
INVx1_ASAP7_75t_L g535 ( .A(n_473), .Y(n_535) );
NAND2xp5_ASAP7_75t_L g536 ( .A(n_466), .B(n_429), .Y(n_536) );
INVx1_ASAP7_75t_L g537 ( .A(n_473), .Y(n_537) );
INVx2_ASAP7_75t_L g538 ( .A(n_470), .Y(n_538) );
OR2x2_ASAP7_75t_L g539 ( .A(n_465), .B(n_429), .Y(n_539) );
AND2x2_ASAP7_75t_L g540 ( .A(n_490), .B(n_429), .Y(n_540) );
AND2x2_ASAP7_75t_L g541 ( .A(n_490), .B(n_439), .Y(n_541) );
AND2x2_ASAP7_75t_L g542 ( .A(n_493), .B(n_439), .Y(n_542) );
INVx1_ASAP7_75t_L g543 ( .A(n_477), .Y(n_543) );
INVxp67_ASAP7_75t_L g544 ( .A(n_484), .Y(n_544) );
AND2x2_ASAP7_75t_L g545 ( .A(n_493), .B(n_446), .Y(n_545) );
AND2x4_ASAP7_75t_L g546 ( .A(n_502), .B(n_446), .Y(n_546) );
INVx1_ASAP7_75t_L g547 ( .A(n_477), .Y(n_547) );
NAND2xp5_ASAP7_75t_SL g548 ( .A(n_506), .B(n_447), .Y(n_548) );
AND2x2_ASAP7_75t_L g549 ( .A(n_494), .B(n_447), .Y(n_549) );
AND2x2_ASAP7_75t_L g550 ( .A(n_494), .B(n_448), .Y(n_550) );
INVx1_ASAP7_75t_L g551 ( .A(n_478), .Y(n_551) );
AND2x2_ASAP7_75t_L g552 ( .A(n_501), .B(n_448), .Y(n_552) );
AND2x2_ASAP7_75t_L g553 ( .A(n_501), .B(n_448), .Y(n_553) );
AND2x2_ASAP7_75t_L g554 ( .A(n_482), .B(n_502), .Y(n_554) );
NAND2xp5_ASAP7_75t_L g555 ( .A(n_469), .B(n_495), .Y(n_555) );
INVxp67_ASAP7_75t_L g556 ( .A(n_497), .Y(n_556) );
AND2x2_ASAP7_75t_L g557 ( .A(n_502), .B(n_503), .Y(n_557) );
AND2x4_ASAP7_75t_L g558 ( .A(n_503), .B(n_471), .Y(n_558) );
AND2x2_ASAP7_75t_L g559 ( .A(n_503), .B(n_498), .Y(n_559) );
AND2x2_ASAP7_75t_SL g560 ( .A(n_471), .B(n_481), .Y(n_560) );
HB1xp67_ASAP7_75t_L g561 ( .A(n_478), .Y(n_561) );
INVx2_ASAP7_75t_L g562 ( .A(n_476), .Y(n_562) );
AND2x2_ASAP7_75t_L g563 ( .A(n_498), .B(n_500), .Y(n_563) );
BUFx3_ASAP7_75t_L g564 ( .A(n_476), .Y(n_564) );
NAND2xp5_ASAP7_75t_L g565 ( .A(n_513), .B(n_497), .Y(n_565) );
AND2x2_ASAP7_75t_L g566 ( .A(n_518), .B(n_481), .Y(n_566) );
INVx3_ASAP7_75t_L g567 ( .A(n_560), .Y(n_567) );
INVx1_ASAP7_75t_SL g568 ( .A(n_541), .Y(n_568) );
AND2x2_ASAP7_75t_L g569 ( .A(n_518), .B(n_481), .Y(n_569) );
NAND2x1_ASAP7_75t_SL g570 ( .A(n_524), .B(n_471), .Y(n_570) );
INVx1_ASAP7_75t_L g571 ( .A(n_511), .Y(n_571) );
INVxp67_ASAP7_75t_L g572 ( .A(n_555), .Y(n_572) );
INVx2_ASAP7_75t_L g573 ( .A(n_545), .Y(n_573) );
INVx1_ASAP7_75t_L g574 ( .A(n_511), .Y(n_574) );
INVx2_ASAP7_75t_SL g575 ( .A(n_560), .Y(n_575) );
INVx1_ASAP7_75t_L g576 ( .A(n_515), .Y(n_576) );
INVx1_ASAP7_75t_L g577 ( .A(n_515), .Y(n_577) );
AND2x2_ASAP7_75t_L g578 ( .A(n_518), .B(n_475), .Y(n_578) );
OR2x2_ASAP7_75t_L g579 ( .A(n_519), .B(n_496), .Y(n_579) );
OR2x2_ASAP7_75t_L g580 ( .A(n_519), .B(n_480), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_520), .Y(n_581) );
OR2x2_ASAP7_75t_L g582 ( .A(n_531), .B(n_489), .Y(n_582) );
INVx2_ASAP7_75t_L g583 ( .A(n_545), .Y(n_583) );
BUFx3_ASAP7_75t_L g584 ( .A(n_564), .Y(n_584) );
AND2x2_ASAP7_75t_L g585 ( .A(n_523), .B(n_475), .Y(n_585) );
INVx1_ASAP7_75t_L g586 ( .A(n_513), .Y(n_586) );
INVx1_ASAP7_75t_L g587 ( .A(n_514), .Y(n_587) );
INVx2_ASAP7_75t_L g588 ( .A(n_545), .Y(n_588) );
NAND2xp5_ASAP7_75t_L g589 ( .A(n_514), .B(n_486), .Y(n_589) );
INVx2_ASAP7_75t_L g590 ( .A(n_520), .Y(n_590) );
AND2x2_ASAP7_75t_SL g591 ( .A(n_560), .B(n_475), .Y(n_591) );
NAND2xp5_ASAP7_75t_L g592 ( .A(n_555), .B(n_505), .Y(n_592) );
NAND2xp5_ASAP7_75t_L g593 ( .A(n_512), .B(n_483), .Y(n_593) );
AND2x2_ASAP7_75t_L g594 ( .A(n_523), .B(n_491), .Y(n_594) );
HB1xp67_ASAP7_75t_L g595 ( .A(n_524), .Y(n_595) );
INVx1_ASAP7_75t_L g596 ( .A(n_525), .Y(n_596) );
HB1xp67_ASAP7_75t_L g597 ( .A(n_561), .Y(n_597) );
NAND2xp5_ASAP7_75t_L g598 ( .A(n_512), .B(n_492), .Y(n_598) );
INVx1_ASAP7_75t_L g599 ( .A(n_525), .Y(n_599) );
OR2x2_ASAP7_75t_L g600 ( .A(n_531), .B(n_492), .Y(n_600) );
INVx1_ASAP7_75t_L g601 ( .A(n_530), .Y(n_601) );
INVx1_ASAP7_75t_L g602 ( .A(n_530), .Y(n_602) );
OR2x2_ASAP7_75t_L g603 ( .A(n_544), .B(n_504), .Y(n_603) );
INVx1_ASAP7_75t_L g604 ( .A(n_534), .Y(n_604) );
INVx1_ASAP7_75t_L g605 ( .A(n_534), .Y(n_605) );
INVx2_ASAP7_75t_L g606 ( .A(n_535), .Y(n_606) );
CKINVDCx16_ASAP7_75t_R g607 ( .A(n_508), .Y(n_607) );
AND2x2_ASAP7_75t_L g608 ( .A(n_507), .B(n_512), .Y(n_608) );
INVx1_ASAP7_75t_L g609 ( .A(n_535), .Y(n_609) );
NAND2xp5_ASAP7_75t_L g610 ( .A(n_509), .B(n_504), .Y(n_610) );
INVx1_ASAP7_75t_L g611 ( .A(n_537), .Y(n_611) );
INVx2_ASAP7_75t_L g612 ( .A(n_537), .Y(n_612) );
INVx1_ASAP7_75t_L g613 ( .A(n_543), .Y(n_613) );
NOR2xp33_ASAP7_75t_SL g614 ( .A(n_561), .B(n_499), .Y(n_614) );
INVx1_ASAP7_75t_L g615 ( .A(n_543), .Y(n_615) );
INVx3_ASAP7_75t_L g616 ( .A(n_546), .Y(n_616) );
HB1xp67_ASAP7_75t_L g617 ( .A(n_556), .Y(n_617) );
HB1xp67_ASAP7_75t_L g618 ( .A(n_595), .Y(n_618) );
AND2x2_ASAP7_75t_L g619 ( .A(n_607), .B(n_557), .Y(n_619) );
INVx1_ASAP7_75t_L g620 ( .A(n_617), .Y(n_620) );
AND2x2_ASAP7_75t_L g621 ( .A(n_608), .B(n_557), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g622 ( .A(n_572), .B(n_544), .Y(n_622) );
AND2x2_ASAP7_75t_L g623 ( .A(n_608), .B(n_554), .Y(n_623) );
NAND2xp5_ASAP7_75t_L g624 ( .A(n_592), .B(n_556), .Y(n_624) );
AND2x4_ASAP7_75t_L g625 ( .A(n_567), .B(n_558), .Y(n_625) );
INVx1_ASAP7_75t_SL g626 ( .A(n_568), .Y(n_626) );
NOR2xp33_ASAP7_75t_SL g627 ( .A(n_591), .B(n_522), .Y(n_627) );
INVx1_ASAP7_75t_L g628 ( .A(n_571), .Y(n_628) );
INVx2_ASAP7_75t_L g629 ( .A(n_590), .Y(n_629) );
O2A1O1Ixp33_ASAP7_75t_L g630 ( .A1(n_580), .A2(n_533), .B(n_510), .C(n_539), .Y(n_630) );
NAND2xp5_ASAP7_75t_L g631 ( .A(n_586), .B(n_528), .Y(n_631) );
AOI22xp33_ASAP7_75t_L g632 ( .A1(n_591), .A2(n_533), .B1(n_510), .B2(n_532), .Y(n_632) );
NOR2xp33_ASAP7_75t_L g633 ( .A(n_587), .B(n_554), .Y(n_633) );
AND2x2_ASAP7_75t_L g634 ( .A(n_585), .B(n_559), .Y(n_634) );
NAND2xp5_ASAP7_75t_L g635 ( .A(n_580), .B(n_540), .Y(n_635) );
OR2x2_ASAP7_75t_L g636 ( .A(n_610), .B(n_522), .Y(n_636) );
AND2x4_ASAP7_75t_L g637 ( .A(n_567), .B(n_558), .Y(n_637) );
NOR2xp33_ASAP7_75t_L g638 ( .A(n_585), .B(n_517), .Y(n_638) );
OAI21xp5_ASAP7_75t_SL g639 ( .A1(n_567), .A2(n_548), .B(n_558), .Y(n_639) );
NAND2xp5_ASAP7_75t_L g640 ( .A(n_565), .B(n_540), .Y(n_640) );
AND2x2_ASAP7_75t_L g641 ( .A(n_566), .B(n_559), .Y(n_641) );
NAND2xp33_ASAP7_75t_L g642 ( .A(n_575), .B(n_527), .Y(n_642) );
NAND2x1_ASAP7_75t_L g643 ( .A(n_575), .B(n_558), .Y(n_643) );
INVx1_ASAP7_75t_L g644 ( .A(n_574), .Y(n_644) );
NAND3xp33_ASAP7_75t_SL g645 ( .A(n_614), .B(n_539), .C(n_536), .Y(n_645) );
NOR3xp33_ASAP7_75t_L g646 ( .A(n_589), .B(n_536), .C(n_532), .Y(n_646) );
INVx2_ASAP7_75t_L g647 ( .A(n_590), .Y(n_647) );
OR2x2_ASAP7_75t_L g648 ( .A(n_573), .B(n_549), .Y(n_648) );
OR2x2_ASAP7_75t_L g649 ( .A(n_573), .B(n_583), .Y(n_649) );
NOR2xp33_ASAP7_75t_L g650 ( .A(n_566), .B(n_517), .Y(n_650) );
AND2x2_ASAP7_75t_L g651 ( .A(n_569), .B(n_549), .Y(n_651) );
INVx1_ASAP7_75t_L g652 ( .A(n_576), .Y(n_652) );
OAI21xp33_ASAP7_75t_L g653 ( .A1(n_570), .A2(n_528), .B(n_516), .Y(n_653) );
NAND2x1_ASAP7_75t_L g654 ( .A(n_616), .B(n_546), .Y(n_654) );
AND2x2_ASAP7_75t_L g655 ( .A(n_569), .B(n_508), .Y(n_655) );
NAND2xp5_ASAP7_75t_L g656 ( .A(n_646), .B(n_597), .Y(n_656) );
AND2x2_ASAP7_75t_L g657 ( .A(n_619), .B(n_578), .Y(n_657) );
INVx2_ASAP7_75t_L g658 ( .A(n_618), .Y(n_658) );
NAND4xp25_ASAP7_75t_SL g659 ( .A(n_632), .B(n_578), .C(n_593), .D(n_594), .Y(n_659) );
OAI22xp5_ASAP7_75t_SL g660 ( .A1(n_643), .A2(n_582), .B1(n_570), .B2(n_584), .Y(n_660) );
OAI22xp33_ASAP7_75t_L g661 ( .A1(n_627), .A2(n_582), .B1(n_616), .B2(n_579), .Y(n_661) );
OAI322xp33_ASAP7_75t_L g662 ( .A1(n_624), .A2(n_579), .A3(n_603), .B1(n_600), .B2(n_598), .C1(n_583), .C2(n_588), .Y(n_662) );
AOI22xp5_ASAP7_75t_L g663 ( .A1(n_646), .A2(n_594), .B1(n_616), .B2(n_509), .Y(n_663) );
O2A1O1Ixp5_ASAP7_75t_L g664 ( .A1(n_654), .A2(n_615), .B(n_596), .C(n_599), .Y(n_664) );
INVx1_ASAP7_75t_L g665 ( .A(n_618), .Y(n_665) );
O2A1O1Ixp5_ASAP7_75t_L g666 ( .A1(n_620), .A2(n_622), .B(n_637), .C(n_625), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_632), .A2(n_600), .B1(n_603), .B2(n_588), .Y(n_667) );
NAND2xp5_ASAP7_75t_L g668 ( .A(n_635), .B(n_516), .Y(n_668) );
O2A1O1Ixp33_ASAP7_75t_SL g669 ( .A1(n_639), .A2(n_602), .B(n_611), .C(n_609), .Y(n_669) );
NAND2xp5_ASAP7_75t_SL g670 ( .A(n_653), .B(n_584), .Y(n_670) );
OAI21xp33_ASAP7_75t_L g671 ( .A1(n_631), .A2(n_550), .B(n_507), .Y(n_671) );
AOI22xp5_ASAP7_75t_L g672 ( .A1(n_642), .A2(n_550), .B1(n_507), .B2(n_527), .Y(n_672) );
INVxp67_ASAP7_75t_L g673 ( .A(n_626), .Y(n_673) );
INVx2_ASAP7_75t_SL g674 ( .A(n_634), .Y(n_674) );
HB1xp67_ASAP7_75t_L g675 ( .A(n_649), .Y(n_675) );
OR2x2_ASAP7_75t_L g676 ( .A(n_640), .B(n_541), .Y(n_676) );
NAND2xp5_ASAP7_75t_L g677 ( .A(n_630), .B(n_613), .Y(n_677) );
NAND2xp5_ASAP7_75t_L g678 ( .A(n_655), .B(n_613), .Y(n_678) );
NAND2xp5_ASAP7_75t_L g679 ( .A(n_677), .B(n_633), .Y(n_679) );
INVx1_ASAP7_75t_L g680 ( .A(n_665), .Y(n_680) );
AOI21xp33_ASAP7_75t_L g681 ( .A1(n_656), .A2(n_642), .B(n_644), .Y(n_681) );
INVx1_ASAP7_75t_L g682 ( .A(n_675), .Y(n_682) );
AOI221xp5_ASAP7_75t_L g683 ( .A1(n_667), .A2(n_633), .B1(n_645), .B2(n_638), .C(n_650), .Y(n_683) );
INVx1_ASAP7_75t_L g684 ( .A(n_678), .Y(n_684) );
INVxp67_ASAP7_75t_L g685 ( .A(n_656), .Y(n_685) );
OAI21xp33_ASAP7_75t_L g686 ( .A1(n_659), .A2(n_650), .B(n_638), .Y(n_686) );
INVx1_ASAP7_75t_L g687 ( .A(n_664), .Y(n_687) );
NAND3xp33_ASAP7_75t_L g688 ( .A(n_666), .B(n_628), .C(n_652), .Y(n_688) );
INVx1_ASAP7_75t_L g689 ( .A(n_658), .Y(n_689) );
OAI322xp33_ASAP7_75t_SL g690 ( .A1(n_668), .A2(n_576), .A3(n_601), .B1(n_577), .B2(n_581), .C1(n_605), .C2(n_604), .Y(n_690) );
AOI22xp5_ASAP7_75t_L g691 ( .A1(n_667), .A2(n_637), .B1(n_625), .B2(n_623), .Y(n_691) );
CKINVDCx20_ASAP7_75t_R g692 ( .A(n_673), .Y(n_692) );
AOI322xp5_ASAP7_75t_L g693 ( .A1(n_686), .A2(n_661), .A3(n_671), .B1(n_663), .B2(n_670), .C1(n_674), .C2(n_657), .Y(n_693) );
A2O1A1Ixp33_ASAP7_75t_SL g694 ( .A1(n_687), .A2(n_672), .B(n_629), .C(n_647), .Y(n_694) );
AOI221xp5_ASAP7_75t_L g695 ( .A1(n_690), .A2(n_662), .B1(n_669), .B2(n_660), .C(n_637), .Y(n_695) );
OAI21xp33_ASAP7_75t_L g696 ( .A1(n_683), .A2(n_676), .B(n_636), .Y(n_696) );
OAI211xp5_ASAP7_75t_SL g697 ( .A1(n_685), .A2(n_648), .B(n_577), .C(n_601), .Y(n_697) );
OAI211xp5_ASAP7_75t_SL g698 ( .A1(n_685), .A2(n_581), .B(n_647), .C(n_629), .Y(n_698) );
OAI221xp5_ASAP7_75t_SL g699 ( .A1(n_691), .A2(n_621), .B1(n_641), .B2(n_651), .C(n_553), .Y(n_699) );
AOI21xp33_ASAP7_75t_L g700 ( .A1(n_679), .A2(n_612), .B(n_606), .Y(n_700) );
NAND3xp33_ASAP7_75t_SL g701 ( .A(n_693), .B(n_692), .C(n_688), .Y(n_701) );
AOI211xp5_ASAP7_75t_L g702 ( .A1(n_699), .A2(n_681), .B(n_682), .C(n_680), .Y(n_702) );
NOR3xp33_ASAP7_75t_L g703 ( .A(n_695), .B(n_684), .C(n_689), .Y(n_703) );
OAI221xp5_ASAP7_75t_L g704 ( .A1(n_694), .A2(n_612), .B1(n_606), .B2(n_529), .C(n_551), .Y(n_704) );
AOI221xp5_ASAP7_75t_L g705 ( .A1(n_696), .A2(n_552), .B1(n_553), .B2(n_563), .C(n_551), .Y(n_705) );
INVxp33_ASAP7_75t_L g706 ( .A(n_703), .Y(n_706) );
NOR2x1_ASAP7_75t_L g707 ( .A(n_701), .B(n_698), .Y(n_707) );
NAND5xp2_ASAP7_75t_L g708 ( .A(n_702), .B(n_700), .C(n_552), .D(n_563), .E(n_529), .Y(n_708) );
INVx2_ASAP7_75t_L g709 ( .A(n_707), .Y(n_709) );
OAI22x1_ASAP7_75t_L g710 ( .A1(n_706), .A2(n_705), .B1(n_704), .B2(n_697), .Y(n_710) );
INVx4_ASAP7_75t_L g711 ( .A(n_709), .Y(n_711) );
XOR2xp5_ASAP7_75t_L g712 ( .A(n_711), .B(n_710), .Y(n_712) );
XNOR2xp5_ASAP7_75t_L g713 ( .A(n_712), .B(n_708), .Y(n_713) );
OAI21xp5_ASAP7_75t_SL g714 ( .A1(n_713), .A2(n_546), .B(n_547), .Y(n_714) );
AO221x2_ASAP7_75t_L g715 ( .A1(n_714), .A2(n_521), .B1(n_562), .B2(n_526), .C(n_538), .Y(n_715) );
AOI22xp5_ASAP7_75t_L g716 ( .A1(n_715), .A2(n_546), .B1(n_542), .B2(n_491), .Y(n_716) );
endmodule