module real_jpeg_26524_n_29 (n_17, n_8, n_0, n_21, n_141, n_2, n_139, n_142, n_143, n_10, n_137, n_9, n_12, n_135, n_24, n_6, n_136, n_28, n_23, n_11, n_14, n_138, n_25, n_7, n_22, n_18, n_3, n_144, n_5, n_4, n_1, n_26, n_27, n_20, n_19, n_140, n_16, n_15, n_13, n_29);

input n_17;
input n_8;
input n_0;
input n_21;
input n_141;
input n_2;
input n_139;
input n_142;
input n_143;
input n_10;
input n_137;
input n_9;
input n_12;
input n_135;
input n_24;
input n_6;
input n_136;
input n_28;
input n_23;
input n_11;
input n_14;
input n_138;
input n_25;
input n_7;
input n_22;
input n_18;
input n_3;
input n_144;
input n_5;
input n_4;
input n_1;
input n_26;
input n_27;
input n_20;
input n_19;
input n_140;
input n_16;
input n_15;
input n_13;

output n_29;

wire n_108;
wire n_54;
wire n_37;
wire n_73;
wire n_35;
wire n_38;
wire n_91;
wire n_49;
wire n_114;
wire n_68;
wire n_78;
wire n_83;
wire n_104;
wire n_64;
wire n_131;
wire n_47;
wire n_87;
wire n_40;
wire n_105;
wire n_115;
wire n_98;
wire n_56;
wire n_48;
wire n_126;
wire n_120;
wire n_113;
wire n_93;
wire n_95;
wire n_65;
wire n_33;
wire n_76;
wire n_67;
wire n_79;
wire n_107;
wire n_66;
wire n_44;
wire n_62;
wire n_121;
wire n_106;
wire n_45;
wire n_112;
wire n_42;
wire n_77;
wire n_109;
wire n_39;
wire n_122;
wire n_94;
wire n_118;
wire n_123;
wire n_116;
wire n_50;
wire n_69;
wire n_31;
wire n_129;
wire n_72;
wire n_100;
wire n_51;
wire n_71;
wire n_90;
wire n_61;
wire n_110;
wire n_117;
wire n_99;
wire n_86;
wire n_70;
wire n_41;
wire n_74;
wire n_80;
wire n_32;
wire n_30;
wire n_130;
wire n_103;
wire n_43;
wire n_57;
wire n_84;
wire n_82;
wire n_111;
wire n_132;
wire n_125;
wire n_55;
wire n_58;
wire n_52;
wire n_63;
wire n_124;
wire n_92;
wire n_75;
wire n_97;
wire n_34;
wire n_60;
wire n_46;
wire n_88;
wire n_59;
wire n_128;
wire n_133;
wire n_53;
wire n_127;
wire n_119;
wire n_36;
wire n_81;
wire n_102;
wire n_85;
wire n_101;
wire n_96;
wire n_89;

CKINVDCx20_ASAP7_75t_R g44 ( 
.A(n_0),
.Y(n_44)
);

NOR2xp33_ASAP7_75t_L g65 ( 
.A(n_1),
.B(n_66),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_1),
.B(n_66),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_2),
.B(n_109),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_L g111 ( 
.A(n_2),
.B(n_109),
.Y(n_111)
);

NOR2xp33_ASAP7_75t_L g117 ( 
.A(n_3),
.B(n_118),
.Y(n_117)
);

NAND2xp5_ASAP7_75t_L g120 ( 
.A(n_3),
.B(n_118),
.Y(n_120)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_4),
.B(n_56),
.C(n_121),
.Y(n_55)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_5),
.Y(n_34)
);

BUFx12_ASAP7_75t_L g61 ( 
.A(n_5),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_SL g78 ( 
.A(n_5),
.B(n_79),
.Y(n_78)
);

NOR2xp33_ASAP7_75t_SL g81 ( 
.A(n_5),
.B(n_82),
.Y(n_81)
);

BUFx12_ASAP7_75t_L g92 ( 
.A(n_5),
.Y(n_92)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_6),
.Y(n_114)
);

NAND2xp5_ASAP7_75t_SL g80 ( 
.A(n_7),
.B(n_81),
.Y(n_80)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_8),
.Y(n_54)
);

NAND2xp5_ASAP7_75t_SL g59 ( 
.A(n_9),
.B(n_60),
.Y(n_59)
);

OR2x2_ASAP7_75t_L g107 ( 
.A(n_9),
.B(n_60),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_10),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_11),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g52 ( 
.A(n_12),
.B(n_53),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g123 ( 
.A(n_12),
.B(n_53),
.Y(n_123)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g131 ( 
.A(n_14),
.Y(n_131)
);

OAI21xp5_ASAP7_75t_SL g30 ( 
.A1(n_15),
.A2(n_31),
.B(n_35),
.Y(n_30)
);

NAND2xp5_ASAP7_75t_L g35 ( 
.A(n_15),
.B(n_31),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g37 ( 
.A(n_15),
.B(n_38),
.Y(n_37)
);

NOR2xp33_ASAP7_75t_SL g42 ( 
.A(n_15),
.B(n_43),
.Y(n_42)
);

NAND2xp5_ASAP7_75t_L g132 ( 
.A(n_15),
.B(n_43),
.Y(n_132)
);

NAND2xp5_ASAP7_75t_L g133 ( 
.A(n_15),
.B(n_38),
.Y(n_133)
);

CKINVDCx20_ASAP7_75t_R g39 ( 
.A(n_16),
.Y(n_39)
);

CKINVDCx20_ASAP7_75t_R g122 ( 
.A(n_17),
.Y(n_122)
);

NOR2xp33_ASAP7_75t_L g70 ( 
.A(n_18),
.B(n_71),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_SL g100 ( 
.A(n_18),
.B(n_71),
.Y(n_100)
);

NOR2xp33_ASAP7_75t_L g77 ( 
.A(n_19),
.B(n_78),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_SL g83 ( 
.A(n_19),
.B(n_78),
.Y(n_83)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_20),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g94 ( 
.A(n_20),
.B(n_91),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_SL g47 ( 
.A(n_21),
.B(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g129 ( 
.A(n_21),
.B(n_48),
.Y(n_129)
);

CKINVDCx20_ASAP7_75t_R g102 ( 
.A(n_22),
.Y(n_102)
);

CKINVDCx20_ASAP7_75t_R g126 ( 
.A(n_23),
.Y(n_126)
);

MAJIxp5_ASAP7_75t_L g45 ( 
.A(n_24),
.B(n_46),
.C(n_130),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g85 ( 
.A(n_25),
.Y(n_85)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_26),
.Y(n_96)
);

CKINVDCx20_ASAP7_75t_R g127 ( 
.A(n_27),
.Y(n_127)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_28),
.Y(n_32)
);

XOR2xp5_ASAP7_75t_L g29 ( 
.A(n_30),
.B(n_36),
.Y(n_29)
);

NOR2xp33_ASAP7_75t_L g31 ( 
.A(n_32),
.B(n_33),
.Y(n_31)
);

NOR2xp33_ASAP7_75t_L g38 ( 
.A(n_33),
.B(n_39),
.Y(n_38)
);

NOR2xp33_ASAP7_75t_L g43 ( 
.A(n_33),
.B(n_44),
.Y(n_43)
);

NOR2xp33_ASAP7_75t_L g48 ( 
.A(n_33),
.B(n_49),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g53 ( 
.A(n_33),
.B(n_54),
.Y(n_53)
);

NOR2xp33_ASAP7_75t_SL g66 ( 
.A(n_33),
.B(n_67),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_33),
.B(n_122),
.Y(n_121)
);

OR2x2_ASAP7_75t_L g125 ( 
.A(n_33),
.B(n_126),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_33),
.B(n_131),
.Y(n_130)
);

INVx11_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx4_ASAP7_75t_L g88 ( 
.A(n_34),
.Y(n_88)
);

OAI21xp5_ASAP7_75t_L g36 ( 
.A1(n_37),
.A2(n_40),
.B(n_133),
.Y(n_36)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_41),
.Y(n_40)
);

OAI21xp5_ASAP7_75t_L g41 ( 
.A1(n_42),
.A2(n_45),
.B(n_132),
.Y(n_41)
);

OAI21xp5_ASAP7_75t_L g46 ( 
.A1(n_47),
.A2(n_50),
.B(n_129),
.Y(n_46)
);

AOI21xp5_ASAP7_75t_SL g50 ( 
.A1(n_51),
.A2(n_124),
.B(n_128),
.Y(n_50)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_55),
.B(n_123),
.Y(n_51)
);

OAI21xp5_ASAP7_75t_SL g56 ( 
.A1(n_57),
.A2(n_117),
.B(n_120),
.Y(n_56)
);

AOI21xp5_ASAP7_75t_SL g57 ( 
.A1(n_58),
.A2(n_112),
.B(n_116),
.Y(n_57)
);

A2O1A1Ixp33_ASAP7_75t_SL g58 ( 
.A1(n_59),
.A2(n_63),
.B(n_108),
.C(n_111),
.Y(n_58)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_61),
.B(n_62),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_SL g71 ( 
.A(n_61),
.B(n_72),
.Y(n_71)
);

OR2x2_ASAP7_75t_L g103 ( 
.A(n_61),
.B(n_104),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_SL g109 ( 
.A(n_61),
.B(n_110),
.Y(n_109)
);

OR2x2_ASAP7_75t_L g113 ( 
.A(n_61),
.B(n_114),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g118 ( 
.A(n_61),
.B(n_119),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_64),
.B(n_107),
.Y(n_63)
);

OAI21xp5_ASAP7_75t_L g64 ( 
.A1(n_65),
.A2(n_68),
.B(n_106),
.Y(n_64)
);

AOI21xp5_ASAP7_75t_L g68 ( 
.A1(n_69),
.A2(n_101),
.B(n_105),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g69 ( 
.A1(n_70),
.A2(n_73),
.B(n_100),
.Y(n_69)
);

AOI21xp5_ASAP7_75t_L g73 ( 
.A1(n_74),
.A2(n_95),
.B(n_99),
.Y(n_73)
);

OAI21xp5_ASAP7_75t_SL g74 ( 
.A1(n_75),
.A2(n_90),
.B(n_94),
.Y(n_74)
);

AOI21xp5_ASAP7_75t_L g75 ( 
.A1(n_76),
.A2(n_84),
.B(n_89),
.Y(n_75)
);

OAI21xp5_ASAP7_75t_SL g76 ( 
.A1(n_77),
.A2(n_80),
.B(n_83),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g84 ( 
.A(n_85),
.B(n_86),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g89 ( 
.A(n_85),
.B(n_86),
.Y(n_89)
);

OR2x2_ASAP7_75t_L g86 ( 
.A(n_87),
.B(n_88),
.Y(n_86)
);

NOR2xp33_ASAP7_75t_SL g91 ( 
.A(n_92),
.B(n_93),
.Y(n_91)
);

OR2x2_ASAP7_75t_L g97 ( 
.A(n_92),
.B(n_98),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g95 ( 
.A(n_96),
.B(n_97),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_SL g99 ( 
.A(n_96),
.B(n_97),
.Y(n_99)
);

NAND2xp5_ASAP7_75t_L g101 ( 
.A(n_102),
.B(n_103),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g105 ( 
.A(n_102),
.B(n_103),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_113),
.B(n_115),
.Y(n_112)
);

NOR2xp33_ASAP7_75t_L g116 ( 
.A(n_113),
.B(n_115),
.Y(n_116)
);

NAND2xp5_ASAP7_75t_SL g124 ( 
.A(n_125),
.B(n_127),
.Y(n_124)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_125),
.B(n_127),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g62 ( 
.A(n_135),
.Y(n_62)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_136),
.Y(n_67)
);

CKINVDCx20_ASAP7_75t_R g72 ( 
.A(n_137),
.Y(n_72)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_138),
.Y(n_79)
);

CKINVDCx20_ASAP7_75t_R g82 ( 
.A(n_139),
.Y(n_82)
);

CKINVDCx20_ASAP7_75t_R g87 ( 
.A(n_140),
.Y(n_87)
);

CKINVDCx20_ASAP7_75t_R g93 ( 
.A(n_141),
.Y(n_93)
);

CKINVDCx20_ASAP7_75t_R g98 ( 
.A(n_142),
.Y(n_98)
);

CKINVDCx20_ASAP7_75t_R g104 ( 
.A(n_143),
.Y(n_104)
);

CKINVDCx20_ASAP7_75t_R g110 ( 
.A(n_144),
.Y(n_110)
);


endmodule