module fake_jpeg_7500_n_342 (n_13, n_11, n_14, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_342);

input n_13;
input n_11;
input n_14;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_342;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_16;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_172;
wire n_78;
wire n_241;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_26;
wire n_88;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_18;
wire n_20;
wire n_145;
wire n_303;
wire n_259;
wire n_90;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_55;
wire n_312;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g16 ( 
.A(n_1),
.Y(n_16)
);

BUFx6f_ASAP7_75t_L g17 ( 
.A(n_15),
.Y(n_17)
);

BUFx3_ASAP7_75t_L g18 ( 
.A(n_1),
.Y(n_18)
);

CKINVDCx20_ASAP7_75t_R g19 ( 
.A(n_0),
.Y(n_19)
);

INVx2_ASAP7_75t_L g20 ( 
.A(n_9),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_3),
.Y(n_21)
);

INVx2_ASAP7_75t_L g22 ( 
.A(n_3),
.Y(n_22)
);

INVx1_ASAP7_75t_L g23 ( 
.A(n_7),
.Y(n_23)
);

BUFx24_ASAP7_75t_L g24 ( 
.A(n_13),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_1),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

BUFx6f_ASAP7_75t_L g27 ( 
.A(n_7),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

CKINVDCx20_ASAP7_75t_R g30 ( 
.A(n_4),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx4f_ASAP7_75t_L g32 ( 
.A(n_7),
.Y(n_32)
);

BUFx6f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_11),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

INVx2_ASAP7_75t_SL g36 ( 
.A(n_18),
.Y(n_36)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_36),
.B(n_37),
.Y(n_69)
);

INVx2_ASAP7_75t_L g37 ( 
.A(n_32),
.Y(n_37)
);

INVx8_ASAP7_75t_L g38 ( 
.A(n_24),
.Y(n_38)
);

INVx6_ASAP7_75t_L g56 ( 
.A(n_38),
.Y(n_56)
);

INVx2_ASAP7_75t_L g39 ( 
.A(n_32),
.Y(n_39)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_39),
.B(n_41),
.Y(n_71)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g57 ( 
.A(n_40),
.Y(n_57)
);

INVx2_ASAP7_75t_L g41 ( 
.A(n_32),
.Y(n_41)
);

BUFx6f_ASAP7_75t_L g42 ( 
.A(n_32),
.Y(n_42)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_SL g43 ( 
.A(n_18),
.Y(n_43)
);

INVx1_ASAP7_75t_L g60 ( 
.A(n_43),
.Y(n_60)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_17),
.Y(n_44)
);

INVx3_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx3_ASAP7_75t_L g45 ( 
.A(n_17),
.Y(n_45)
);

INVx4_ASAP7_75t_L g50 ( 
.A(n_45),
.Y(n_50)
);

BUFx12f_ASAP7_75t_L g46 ( 
.A(n_24),
.Y(n_46)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_46),
.Y(n_53)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_24),
.Y(n_47)
);

INVx5_ASAP7_75t_L g49 ( 
.A(n_47),
.Y(n_49)
);

INVx4_ASAP7_75t_L g48 ( 
.A(n_24),
.Y(n_48)
);

HB1xp67_ASAP7_75t_L g65 ( 
.A(n_48),
.Y(n_65)
);

AOI22xp5_ASAP7_75t_L g51 ( 
.A1(n_40),
.A2(n_29),
.B1(n_20),
.B2(n_22),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_SL g73 ( 
.A1(n_51),
.A2(n_45),
.B1(n_23),
.B2(n_31),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_SL g52 ( 
.A(n_37),
.B(n_35),
.Y(n_52)
);

AND2x2_ASAP7_75t_L g95 ( 
.A(n_52),
.B(n_31),
.Y(n_95)
);

BUFx5_ASAP7_75t_L g55 ( 
.A(n_36),
.Y(n_55)
);

INVx3_ASAP7_75t_SL g91 ( 
.A(n_55),
.Y(n_91)
);

AOI22xp33_ASAP7_75t_SL g58 ( 
.A1(n_40),
.A2(n_29),
.B1(n_20),
.B2(n_22),
.Y(n_58)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_58),
.A2(n_64),
.B1(n_26),
.B2(n_19),
.Y(n_99)
);

INVx2_ASAP7_75t_L g61 ( 
.A(n_37),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g93 ( 
.A(n_61),
.B(n_62),
.Y(n_93)
);

INVx2_ASAP7_75t_L g62 ( 
.A(n_39),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g63 ( 
.A(n_46),
.B(n_35),
.Y(n_63)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_63),
.B(n_23),
.Y(n_87)
);

AOI22xp33_ASAP7_75t_L g64 ( 
.A1(n_45),
.A2(n_34),
.B1(n_25),
.B2(n_21),
.Y(n_64)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_39),
.Y(n_66)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_66),
.Y(n_82)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_41),
.Y(n_67)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_67),
.Y(n_88)
);

INVx3_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

INVx2_ASAP7_75t_L g70 ( 
.A(n_41),
.Y(n_70)
);

HB1xp67_ASAP7_75t_L g77 ( 
.A(n_70),
.Y(n_77)
);

OR2x4_ASAP7_75t_L g72 ( 
.A(n_52),
.B(n_42),
.Y(n_72)
);

OAI21xp5_ASAP7_75t_L g103 ( 
.A1(n_72),
.A2(n_98),
.B(n_95),
.Y(n_103)
);

AOI22xp5_ASAP7_75t_L g107 ( 
.A1(n_73),
.A2(n_98),
.B1(n_68),
.B2(n_54),
.Y(n_107)
);

XNOR2xp5_ASAP7_75t_L g74 ( 
.A(n_63),
.B(n_42),
.Y(n_74)
);

XNOR2xp5_ASAP7_75t_L g125 ( 
.A(n_74),
.B(n_24),
.Y(n_125)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_65),
.Y(n_75)
);

NOR2xp33_ASAP7_75t_L g119 ( 
.A(n_75),
.B(n_76),
.Y(n_119)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_69),
.Y(n_76)
);

AOI22xp5_ASAP7_75t_L g78 ( 
.A1(n_57),
.A2(n_48),
.B1(n_47),
.B2(n_38),
.Y(n_78)
);

OAI22xp5_ASAP7_75t_SL g110 ( 
.A1(n_78),
.A2(n_84),
.B1(n_96),
.B2(n_59),
.Y(n_110)
);

BUFx3_ASAP7_75t_L g79 ( 
.A(n_55),
.Y(n_79)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

NAND3xp33_ASAP7_75t_L g80 ( 
.A(n_50),
.B(n_48),
.C(n_15),
.Y(n_80)
);

NAND2xp5_ASAP7_75t_SL g106 ( 
.A(n_80),
.B(n_87),
.Y(n_106)
);

HB1xp67_ASAP7_75t_L g81 ( 
.A(n_61),
.Y(n_81)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_81),
.Y(n_104)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_62),
.Y(n_83)
);

INVx4_ASAP7_75t_L g114 ( 
.A(n_83),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_L g84 ( 
.A1(n_50),
.A2(n_43),
.B1(n_36),
.B2(n_34),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_49),
.Y(n_85)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_85),
.B(n_86),
.Y(n_122)
);

CKINVDCx16_ASAP7_75t_R g86 ( 
.A(n_71),
.Y(n_86)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_49),
.Y(n_89)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_89),
.B(n_94),
.Y(n_129)
);

HB1xp67_ASAP7_75t_L g90 ( 
.A(n_70),
.Y(n_90)
);

INVx2_ASAP7_75t_L g111 ( 
.A(n_90),
.Y(n_111)
);

INVx3_ASAP7_75t_L g92 ( 
.A(n_66),
.Y(n_92)
);

INVx4_ASAP7_75t_L g121 ( 
.A(n_92),
.Y(n_121)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

NAND2xp5_ASAP7_75t_SL g123 ( 
.A(n_95),
.B(n_99),
.Y(n_123)
);

AOI22xp33_ASAP7_75t_SL g96 ( 
.A1(n_56),
.A2(n_47),
.B1(n_38),
.B2(n_43),
.Y(n_96)
);

INVx2_ASAP7_75t_L g97 ( 
.A(n_51),
.Y(n_97)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_97),
.Y(n_130)
);

AO22x1_ASAP7_75t_SL g98 ( 
.A1(n_57),
.A2(n_44),
.B1(n_43),
.B2(n_36),
.Y(n_98)
);

INVx5_ASAP7_75t_L g100 ( 
.A(n_56),
.Y(n_100)
);

INVx8_ASAP7_75t_L g109 ( 
.A(n_100),
.Y(n_109)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_54),
.Y(n_101)
);

INVx1_ASAP7_75t_SL g120 ( 
.A(n_101),
.Y(n_120)
);

OAI21xp5_ASAP7_75t_SL g142 ( 
.A1(n_103),
.A2(n_102),
.B(n_88),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_74),
.B(n_60),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_118),
.Y(n_144)
);

AOI22xp33_ASAP7_75t_L g163 ( 
.A1(n_107),
.A2(n_33),
.B1(n_46),
.B2(n_28),
.Y(n_163)
);

INVx1_ASAP7_75t_L g108 ( 
.A(n_93),
.Y(n_108)
);

NAND2xp5_ASAP7_75t_SL g135 ( 
.A(n_108),
.B(n_115),
.Y(n_135)
);

AOI22xp5_ASAP7_75t_L g151 ( 
.A1(n_110),
.A2(n_127),
.B1(n_128),
.B2(n_30),
.Y(n_151)
);

INVx3_ASAP7_75t_L g113 ( 
.A(n_79),
.Y(n_113)
);

INVx4_ASAP7_75t_L g148 ( 
.A(n_113),
.Y(n_148)
);

INVx1_ASAP7_75t_L g115 ( 
.A(n_98),
.Y(n_115)
);

INVx1_ASAP7_75t_L g116 ( 
.A(n_78),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_131),
.Y(n_147)
);

MAJx2_ASAP7_75t_L g117 ( 
.A(n_72),
.B(n_60),
.C(n_46),
.Y(n_117)
);

MAJIxp5_ASAP7_75t_L g155 ( 
.A(n_117),
.B(n_46),
.C(n_18),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_L g118 ( 
.A(n_95),
.B(n_44),
.Y(n_118)
);

BUFx5_ASAP7_75t_L g124 ( 
.A(n_91),
.Y(n_124)
);

CKINVDCx14_ASAP7_75t_R g136 ( 
.A(n_124),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g139 ( 
.A(n_125),
.B(n_46),
.Y(n_139)
);

NAND2xp5_ASAP7_75t_SL g126 ( 
.A(n_75),
.B(n_19),
.Y(n_126)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_126),
.Y(n_138)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_97),
.A2(n_59),
.B1(n_44),
.B2(n_53),
.Y(n_127)
);

OAI22xp5_ASAP7_75t_SL g128 ( 
.A1(n_73),
.A2(n_53),
.B1(n_26),
.B2(n_25),
.Y(n_128)
);

INVx1_ASAP7_75t_L g131 ( 
.A(n_91),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g132 ( 
.A1(n_115),
.A2(n_100),
.B1(n_92),
.B2(n_83),
.Y(n_132)
);

AOI22xp5_ASAP7_75t_L g182 ( 
.A1(n_132),
.A2(n_111),
.B1(n_104),
.B2(n_121),
.Y(n_182)
);

INVx1_ASAP7_75t_L g133 ( 
.A(n_129),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_133),
.B(n_134),
.Y(n_164)
);

INVx1_ASAP7_75t_L g134 ( 
.A(n_119),
.Y(n_134)
);

INVx2_ASAP7_75t_L g137 ( 
.A(n_124),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_137),
.B(n_140),
.Y(n_169)
);

XNOR2xp5_ASAP7_75t_L g166 ( 
.A(n_139),
.B(n_155),
.Y(n_166)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_114),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_122),
.Y(n_141)
);

NOR2xp33_ASAP7_75t_L g187 ( 
.A(n_141),
.B(n_143),
.Y(n_187)
);

XOR2xp5_ASAP7_75t_L g183 ( 
.A(n_142),
.B(n_33),
.Y(n_183)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_127),
.Y(n_143)
);

INVx2_ASAP7_75t_L g145 ( 
.A(n_120),
.Y(n_145)
);

NOR2xp33_ASAP7_75t_L g192 ( 
.A(n_145),
.B(n_149),
.Y(n_192)
);

AOI22xp33_ASAP7_75t_SL g146 ( 
.A1(n_109),
.A2(n_85),
.B1(n_101),
.B2(n_94),
.Y(n_146)
);

OAI22xp5_ASAP7_75t_L g167 ( 
.A1(n_146),
.A2(n_151),
.B1(n_163),
.B2(n_109),
.Y(n_167)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_120),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g150 ( 
.A1(n_116),
.A2(n_30),
.B1(n_21),
.B2(n_82),
.Y(n_150)
);

INVxp67_ASAP7_75t_L g174 ( 
.A(n_150),
.Y(n_174)
);

INVx1_ASAP7_75t_L g152 ( 
.A(n_107),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_152),
.B(n_160),
.Y(n_172)
);

XOR2xp5_ASAP7_75t_L g153 ( 
.A(n_105),
.B(n_77),
.Y(n_153)
);

MAJIxp5_ASAP7_75t_L g188 ( 
.A(n_153),
.B(n_159),
.C(n_14),
.Y(n_188)
);

AOI22xp5_ASAP7_75t_L g154 ( 
.A1(n_110),
.A2(n_33),
.B1(n_17),
.B2(n_28),
.Y(n_154)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_154),
.A2(n_121),
.B1(n_114),
.B2(n_33),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g156 ( 
.A(n_112),
.B(n_10),
.Y(n_156)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_156),
.Y(n_180)
);

INVxp67_ASAP7_75t_L g157 ( 
.A(n_128),
.Y(n_157)
);

HB1xp67_ASAP7_75t_L g173 ( 
.A(n_157),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g158 ( 
.A(n_112),
.B(n_10),
.Y(n_158)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_158),
.Y(n_190)
);

XNOR2xp5_ASAP7_75t_L g159 ( 
.A(n_125),
.B(n_103),
.Y(n_159)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_118),
.Y(n_160)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_113),
.B(n_11),
.Y(n_161)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_161),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_123),
.B(n_16),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g178 ( 
.A(n_162),
.B(n_104),
.Y(n_178)
);

INVx2_ASAP7_75t_L g165 ( 
.A(n_140),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g202 ( 
.A(n_165),
.B(n_168),
.Y(n_202)
);

CKINVDCx14_ASAP7_75t_R g203 ( 
.A(n_167),
.Y(n_203)
);

INVx1_ASAP7_75t_L g168 ( 
.A(n_147),
.Y(n_168)
);

OA22x2_ASAP7_75t_L g170 ( 
.A1(n_132),
.A2(n_117),
.B1(n_130),
.B2(n_131),
.Y(n_170)
);

AOI22xp5_ASAP7_75t_L g221 ( 
.A1(n_170),
.A2(n_179),
.B1(n_184),
.B2(n_198),
.Y(n_221)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_135),
.Y(n_171)
);

NAND2xp5_ASAP7_75t_SL g209 ( 
.A(n_171),
.B(n_175),
.Y(n_209)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_152),
.A2(n_106),
.B1(n_108),
.B2(n_111),
.Y(n_175)
);

CKINVDCx20_ASAP7_75t_R g176 ( 
.A(n_140),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g224 ( 
.A(n_176),
.B(n_181),
.Y(n_224)
);

BUFx2_ASAP7_75t_L g177 ( 
.A(n_145),
.Y(n_177)
);

INVxp67_ASAP7_75t_SL g204 ( 
.A(n_177),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_SL g215 ( 
.A(n_178),
.B(n_186),
.Y(n_215)
);

CKINVDCx20_ASAP7_75t_R g181 ( 
.A(n_150),
.Y(n_181)
);

OAI22xp5_ASAP7_75t_L g205 ( 
.A1(n_182),
.A2(n_189),
.B1(n_172),
.B2(n_178),
.Y(n_205)
);

XOR2xp5_ASAP7_75t_L g199 ( 
.A(n_183),
.B(n_137),
.Y(n_199)
);

OAI22xp5_ASAP7_75t_SL g184 ( 
.A1(n_143),
.A2(n_28),
.B1(n_27),
.B2(n_16),
.Y(n_184)
);

NAND2xp5_ASAP7_75t_L g185 ( 
.A(n_144),
.B(n_27),
.Y(n_185)
);

INVx1_ASAP7_75t_L g200 ( 
.A(n_185),
.Y(n_200)
);

OAI22xp5_ASAP7_75t_L g186 ( 
.A1(n_157),
.A2(n_27),
.B1(n_16),
.B2(n_15),
.Y(n_186)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_188),
.B(n_197),
.C(n_138),
.Y(n_217)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_142),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g207 ( 
.A(n_189),
.B(n_194),
.Y(n_207)
);

NAND2xp5_ASAP7_75t_L g191 ( 
.A(n_144),
.B(n_153),
.Y(n_191)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_191),
.Y(n_201)
);

INVx1_ASAP7_75t_L g194 ( 
.A(n_149),
.Y(n_194)
);

INVx1_ASAP7_75t_L g195 ( 
.A(n_151),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g210 ( 
.A(n_195),
.B(n_196),
.Y(n_210)
);

CKINVDCx14_ASAP7_75t_R g196 ( 
.A(n_162),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g197 ( 
.A(n_159),
.B(n_0),
.C(n_1),
.Y(n_197)
);

AO22x1_ASAP7_75t_SL g198 ( 
.A1(n_154),
.A2(n_160),
.B1(n_155),
.B2(n_139),
.Y(n_198)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_199),
.B(n_226),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g230 ( 
.A(n_205),
.Y(n_230)
);

OAI22xp5_ASAP7_75t_SL g206 ( 
.A1(n_172),
.A2(n_195),
.B1(n_174),
.B2(n_198),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_206),
.A2(n_220),
.B1(n_184),
.B2(n_179),
.Y(n_236)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_192),
.Y(n_208)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_208),
.B(n_211),
.Y(n_233)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_169),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_164),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g235 ( 
.A(n_212),
.B(n_216),
.Y(n_235)
);

XOR2x1_ASAP7_75t_SL g213 ( 
.A(n_198),
.B(n_134),
.Y(n_213)
);

OAI21xp5_ASAP7_75t_L g234 ( 
.A1(n_213),
.A2(n_218),
.B(n_222),
.Y(n_234)
);

NAND2x1_ASAP7_75t_L g214 ( 
.A(n_183),
.B(n_133),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g231 ( 
.A1(n_214),
.A2(n_168),
.B1(n_171),
.B2(n_194),
.Y(n_231)
);

OR2x2_ASAP7_75t_L g216 ( 
.A(n_187),
.B(n_148),
.Y(n_216)
);

XNOR2xp5_ASAP7_75t_L g232 ( 
.A(n_217),
.B(n_166),
.Y(n_232)
);

AOI21xp5_ASAP7_75t_L g218 ( 
.A1(n_174),
.A2(n_148),
.B(n_136),
.Y(n_218)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_182),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_205),
.Y(n_245)
);

OAI22xp5_ASAP7_75t_SL g220 ( 
.A1(n_173),
.A2(n_0),
.B1(n_2),
.B2(n_3),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g222 ( 
.A1(n_170),
.A2(n_2),
.B(n_4),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g223 ( 
.A1(n_170),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_223)
);

INVx1_ASAP7_75t_L g240 ( 
.A(n_223),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_185),
.B(n_2),
.Y(n_225)
);

INVx1_ASAP7_75t_L g238 ( 
.A(n_225),
.Y(n_238)
);

OAI21xp5_ASAP7_75t_SL g226 ( 
.A1(n_170),
.A2(n_4),
.B(n_5),
.Y(n_226)
);

NAND2xp5_ASAP7_75t_L g227 ( 
.A(n_191),
.B(n_5),
.Y(n_227)
);

INVx1_ASAP7_75t_L g244 ( 
.A(n_227),
.Y(n_244)
);

MAJIxp5_ASAP7_75t_L g228 ( 
.A(n_201),
.B(n_166),
.C(n_188),
.Y(n_228)
);

MAJIxp5_ASAP7_75t_L g260 ( 
.A(n_228),
.B(n_232),
.C(n_239),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g229 ( 
.A(n_202),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g274 ( 
.A(n_229),
.B(n_237),
.Y(n_274)
);

XNOR2xp5_ASAP7_75t_L g254 ( 
.A(n_231),
.B(n_223),
.Y(n_254)
);

OAI21xp33_ASAP7_75t_SL g256 ( 
.A1(n_236),
.A2(n_222),
.B(n_221),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_216),
.B(n_193),
.Y(n_237)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_201),
.B(n_197),
.C(n_190),
.Y(n_239)
);

NAND2xp5_ASAP7_75t_SL g241 ( 
.A(n_216),
.B(n_180),
.Y(n_241)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_241),
.Y(n_258)
);

MAJIxp5_ASAP7_75t_L g242 ( 
.A(n_199),
.B(n_177),
.C(n_165),
.Y(n_242)
);

MAJIxp5_ASAP7_75t_L g264 ( 
.A(n_242),
.B(n_246),
.C(n_225),
.Y(n_264)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_245),
.Y(n_263)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_214),
.B(n_5),
.C(n_6),
.Y(n_246)
);

INVxp67_ASAP7_75t_L g247 ( 
.A(n_202),
.Y(n_247)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_247),
.B(n_248),
.Y(n_257)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_207),
.Y(n_248)
);

OAI22xp5_ASAP7_75t_L g249 ( 
.A1(n_203),
.A2(n_6),
.B1(n_7),
.B2(n_8),
.Y(n_249)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_249),
.Y(n_267)
);

NAND3xp33_ASAP7_75t_SL g250 ( 
.A(n_224),
.B(n_9),
.C(n_11),
.Y(n_250)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_250),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g251 ( 
.A(n_207),
.Y(n_251)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_251),
.Y(n_270)
);

XOR2xp5_ASAP7_75t_L g252 ( 
.A(n_213),
.B(n_9),
.Y(n_252)
);

XOR2xp5_ASAP7_75t_L g255 ( 
.A(n_252),
.B(n_226),
.Y(n_255)
);

NAND2xp5_ASAP7_75t_L g253 ( 
.A(n_227),
.B(n_6),
.Y(n_253)
);

INVx1_ASAP7_75t_L g272 ( 
.A(n_253),
.Y(n_272)
);

XNOR2xp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_246),
.Y(n_282)
);

XOR2xp5_ASAP7_75t_L g277 ( 
.A(n_255),
.B(n_261),
.Y(n_277)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_256),
.Y(n_279)
);

XNOR2xp5_ASAP7_75t_L g259 ( 
.A(n_242),
.B(n_218),
.Y(n_259)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_259),
.B(n_264),
.C(n_268),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g261 ( 
.A(n_234),
.B(n_214),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_240),
.A2(n_219),
.B1(n_209),
.B2(n_221),
.Y(n_262)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_262),
.Y(n_280)
);

OA22x2_ASAP7_75t_L g265 ( 
.A1(n_234),
.A2(n_206),
.B1(n_210),
.B2(n_209),
.Y(n_265)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_265),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g266 ( 
.A(n_232),
.B(n_217),
.C(n_200),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g276 ( 
.A(n_266),
.B(n_271),
.C(n_243),
.Y(n_276)
);

XNOR2xp5_ASAP7_75t_L g268 ( 
.A(n_233),
.B(n_210),
.Y(n_268)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_228),
.B(n_200),
.C(n_211),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_247),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g283 ( 
.A(n_273),
.B(n_204),
.Y(n_283)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_274),
.B(n_251),
.Y(n_275)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_275),
.Y(n_304)
);

MAJIxp5_ASAP7_75t_L g293 ( 
.A(n_276),
.B(n_287),
.C(n_291),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g278 ( 
.A(n_261),
.B(n_243),
.Y(n_278)
);

XOR2xp5_ASAP7_75t_L g302 ( 
.A(n_278),
.B(n_253),
.Y(n_302)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_257),
.Y(n_281)
);

NAND2xp5_ASAP7_75t_L g295 ( 
.A(n_281),
.B(n_282),
.Y(n_295)
);

CKINVDCx20_ASAP7_75t_R g299 ( 
.A(n_283),
.Y(n_299)
);

INVxp67_ASAP7_75t_L g284 ( 
.A(n_270),
.Y(n_284)
);

NAND2xp5_ASAP7_75t_L g300 ( 
.A(n_284),
.B(n_289),
.Y(n_300)
);

XNOR2xp5_ASAP7_75t_L g286 ( 
.A(n_260),
.B(n_233),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g303 ( 
.A(n_286),
.B(n_288),
.Y(n_303)
);

MAJIxp5_ASAP7_75t_L g287 ( 
.A(n_271),
.B(n_239),
.C(n_235),
.Y(n_287)
);

INVxp67_ASAP7_75t_L g289 ( 
.A(n_256),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_265),
.Y(n_290)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_290),
.B(n_252),
.Y(n_301)
);

MAJIxp5_ASAP7_75t_L g291 ( 
.A(n_266),
.B(n_235),
.C(n_230),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_SL g292 ( 
.A1(n_285),
.A2(n_263),
.B(n_245),
.Y(n_292)
);

OAI21xp5_ASAP7_75t_L g313 ( 
.A1(n_292),
.A2(n_12),
.B(n_13),
.Y(n_313)
);

MAJIxp5_ASAP7_75t_L g294 ( 
.A(n_287),
.B(n_260),
.C(n_264),
.Y(n_294)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_294),
.B(n_296),
.C(n_298),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_291),
.B(n_244),
.C(n_272),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_SL g297 ( 
.A1(n_289),
.A2(n_265),
.B1(n_236),
.B2(n_231),
.Y(n_297)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_297),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g298 ( 
.A(n_276),
.B(n_244),
.C(n_255),
.Y(n_298)
);

INVxp67_ASAP7_75t_L g318 ( 
.A(n_301),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_302),
.B(n_8),
.Y(n_317)
);

NAND2xp5_ASAP7_75t_L g309 ( 
.A(n_303),
.B(n_277),
.Y(n_309)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_279),
.A2(n_258),
.B1(n_267),
.B2(n_269),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g311 ( 
.A(n_305),
.B(n_306),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g306 ( 
.A1(n_280),
.A2(n_238),
.B1(n_215),
.B2(n_208),
.Y(n_306)
);

AOI21xp5_ASAP7_75t_L g307 ( 
.A1(n_296),
.A2(n_284),
.B(n_212),
.Y(n_307)
);

OAI21xp5_ASAP7_75t_SL g325 ( 
.A1(n_307),
.A2(n_318),
.B(n_292),
.Y(n_325)
);

AOI21xp5_ASAP7_75t_L g320 ( 
.A1(n_309),
.A2(n_314),
.B(n_295),
.Y(n_320)
);

AOI22xp5_ASAP7_75t_SL g310 ( 
.A1(n_304),
.A2(n_277),
.B1(n_278),
.B2(n_238),
.Y(n_310)
);

INVxp67_ASAP7_75t_L g322 ( 
.A(n_310),
.Y(n_322)
);

AOI31xp33_ASAP7_75t_L g312 ( 
.A1(n_305),
.A2(n_215),
.A3(n_220),
.B(n_13),
.Y(n_312)
);

FAx1_ASAP7_75t_SL g326 ( 
.A(n_312),
.B(n_313),
.CI(n_302),
.CON(n_326),
.SN(n_326)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_293),
.A2(n_14),
.B(n_12),
.Y(n_314)
);

OR2x2_ASAP7_75t_L g315 ( 
.A(n_300),
.B(n_8),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g323 ( 
.A(n_315),
.B(n_8),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_317),
.B(n_311),
.Y(n_327)
);

AOI22xp5_ASAP7_75t_L g319 ( 
.A1(n_316),
.A2(n_297),
.B1(n_306),
.B2(n_299),
.Y(n_319)
);

NOR2xp33_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_320),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g321 ( 
.A(n_308),
.B(n_298),
.Y(n_321)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_321),
.A2(n_318),
.B(n_310),
.Y(n_332)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_323),
.B(n_324),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_308),
.B(n_293),
.C(n_294),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g330 ( 
.A(n_325),
.B(n_326),
.Y(n_330)
);

NOR2xp33_ASAP7_75t_L g333 ( 
.A(n_327),
.B(n_326),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_327),
.B(n_315),
.Y(n_331)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_331),
.Y(n_336)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_332),
.B(n_333),
.Y(n_334)
);

NAND2xp5_ASAP7_75t_L g335 ( 
.A(n_328),
.B(n_321),
.Y(n_335)
);

INVxp33_ASAP7_75t_SL g337 ( 
.A(n_335),
.Y(n_337)
);

NOR3xp33_ASAP7_75t_L g338 ( 
.A(n_337),
.B(n_334),
.C(n_330),
.Y(n_338)
);

BUFx24_ASAP7_75t_SL g339 ( 
.A(n_338),
.Y(n_339)
);

BUFx24_ASAP7_75t_SL g340 ( 
.A(n_339),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g341 ( 
.A1(n_340),
.A2(n_336),
.B1(n_329),
.B2(n_322),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_341),
.B(n_332),
.C(n_322),
.Y(n_342)
);


endmodule