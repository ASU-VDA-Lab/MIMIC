module fake_netlist_1_6638_n_16 (n_1, n_2, n_0, n_16);
input n_1;
input n_2;
input n_0;
output n_16;
wire n_11;
wire n_13;
wire n_12;
wire n_6;
wire n_4;
wire n_3;
wire n_9;
wire n_5;
wire n_14;
wire n_7;
wire n_15;
wire n_10;
wire n_8;
CKINVDCx5p33_ASAP7_75t_R g3 ( .A(n_0), .Y(n_3) );
AND2x2_ASAP7_75t_L g4 ( .A(n_2), .B(n_1), .Y(n_4) );
OR2x2_ASAP7_75t_L g5 ( .A(n_1), .B(n_0), .Y(n_5) );
OAI21x1_ASAP7_75t_L g6 ( .A1(n_5), .A2(n_0), .B(n_1), .Y(n_6) );
INVx5_ASAP7_75t_L g7 ( .A(n_4), .Y(n_7) );
NAND3x1_ASAP7_75t_L g8 ( .A(n_4), .B(n_0), .C(n_1), .Y(n_8) );
AND2x2_ASAP7_75t_L g9 ( .A(n_7), .B(n_4), .Y(n_9) );
AND2x2_ASAP7_75t_L g10 ( .A(n_7), .B(n_3), .Y(n_10) );
INVxp67_ASAP7_75t_L g11 ( .A(n_10), .Y(n_11) );
OAI211xp5_ASAP7_75t_L g12 ( .A1(n_9), .A2(n_5), .B(n_7), .C(n_6), .Y(n_12) );
AOI211xp5_ASAP7_75t_L g13 ( .A1(n_11), .A2(n_9), .B(n_6), .C(n_8), .Y(n_13) );
NAND4xp25_ASAP7_75t_L g14 ( .A(n_12), .B(n_8), .C(n_2), .D(n_7), .Y(n_14) );
AOI22xp5_ASAP7_75t_L g15 ( .A1(n_14), .A2(n_12), .B1(n_7), .B2(n_2), .Y(n_15) );
OA21x2_ASAP7_75t_L g16 ( .A1(n_15), .A2(n_13), .B(n_2), .Y(n_16) );
endmodule