module fake_jpeg_31548_n_83 (n_13, n_21, n_1, n_10, n_23, n_27, n_6, n_22, n_14, n_19, n_18, n_20, n_4, n_30, n_16, n_3, n_0, n_24, n_28, n_26, n_9, n_5, n_11, n_17, n_25, n_31, n_2, n_29, n_12, n_8, n_15, n_7, n_83);

input n_13;
input n_21;
input n_1;
input n_10;
input n_23;
input n_27;
input n_6;
input n_22;
input n_14;
input n_19;
input n_18;
input n_20;
input n_4;
input n_30;
input n_16;
input n_3;
input n_0;
input n_24;
input n_28;
input n_26;
input n_9;
input n_5;
input n_11;
input n_17;
input n_25;
input n_31;
input n_2;
input n_29;
input n_12;
input n_8;
input n_15;
input n_7;

output n_83;

wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_73;
wire n_59;
wire n_65;
wire n_42;
wire n_49;
wire n_76;
wire n_38;
wire n_74;
wire n_50;
wire n_57;
wire n_69;
wire n_40;
wire n_71;
wire n_80;
wire n_81;
wire n_44;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_56;
wire n_79;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_35;
wire n_48;
wire n_46;
wire n_36;
wire n_62;
wire n_43;
wire n_32;
wire n_82;

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_22),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx4_ASAP7_75t_L g34 ( 
.A(n_8),
.Y(n_34)
);

INVx6_ASAP7_75t_L g35 ( 
.A(n_23),
.Y(n_35)
);

BUFx6f_ASAP7_75t_L g36 ( 
.A(n_30),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_2),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g38 ( 
.A(n_5),
.B(n_15),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_2),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_17),
.Y(n_40)
);

INVx1_ASAP7_75t_SL g41 ( 
.A(n_7),
.Y(n_41)
);

INVx3_ASAP7_75t_L g42 ( 
.A(n_34),
.Y(n_42)
);

INVx3_ASAP7_75t_L g53 ( 
.A(n_42),
.Y(n_53)
);

INVx11_ASAP7_75t_L g43 ( 
.A(n_36),
.Y(n_43)
);

INVx2_ASAP7_75t_L g54 ( 
.A(n_43),
.Y(n_54)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

INVx1_ASAP7_75t_SL g49 ( 
.A(n_44),
.Y(n_49)
);

INVx4_ASAP7_75t_SL g45 ( 
.A(n_41),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_38),
.B(n_0),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_L g47 ( 
.A(n_46),
.B(n_37),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_47),
.B(n_48),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g48 ( 
.A1(n_44),
.A2(n_40),
.B1(n_41),
.B2(n_33),
.Y(n_48)
);

OAI22xp5_ASAP7_75t_L g50 ( 
.A1(n_46),
.A2(n_32),
.B1(n_39),
.B2(n_6),
.Y(n_50)
);

O2A1O1Ixp33_ASAP7_75t_L g59 ( 
.A1(n_50),
.A2(n_11),
.B(n_12),
.C(n_13),
.Y(n_59)
);

CKINVDCx20_ASAP7_75t_R g51 ( 
.A(n_45),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g60 ( 
.A(n_51),
.B(n_52),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g52 ( 
.A(n_46),
.B(n_18),
.C(n_4),
.Y(n_52)
);

MAJIxp5_ASAP7_75t_L g55 ( 
.A(n_46),
.B(n_19),
.C(n_9),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_SL g56 ( 
.A(n_55),
.B(n_1),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g67 ( 
.A(n_56),
.B(n_57),
.Y(n_67)
);

INVx6_ASAP7_75t_L g57 ( 
.A(n_54),
.Y(n_57)
);

OR2x2_ASAP7_75t_SL g58 ( 
.A(n_53),
.B(n_10),
.Y(n_58)
);

MAJIxp5_ASAP7_75t_L g68 ( 
.A(n_58),
.B(n_65),
.C(n_20),
.Y(n_68)
);

OAI21xp5_ASAP7_75t_L g66 ( 
.A1(n_59),
.A2(n_62),
.B(n_63),
.Y(n_66)
);

NOR2xp33_ASAP7_75t_L g62 ( 
.A(n_48),
.B(n_14),
.Y(n_62)
);

INVx1_ASAP7_75t_L g63 ( 
.A(n_49),
.Y(n_63)
);

BUFx12f_ASAP7_75t_L g64 ( 
.A(n_51),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_L g69 ( 
.A(n_64),
.B(n_21),
.Y(n_69)
);

NAND2xp5_ASAP7_75t_SL g65 ( 
.A(n_47),
.B(n_16),
.Y(n_65)
);

NAND2xp5_ASAP7_75t_L g74 ( 
.A(n_68),
.B(n_69),
.Y(n_74)
);

AO21x2_ASAP7_75t_L g70 ( 
.A1(n_61),
.A2(n_24),
.B(n_25),
.Y(n_70)
);

NAND2xp5_ASAP7_75t_L g72 ( 
.A(n_70),
.B(n_71),
.Y(n_72)
);

OAI22xp5_ASAP7_75t_L g71 ( 
.A1(n_60),
.A2(n_26),
.B1(n_27),
.B2(n_28),
.Y(n_71)
);

CKINVDCx20_ASAP7_75t_R g73 ( 
.A(n_69),
.Y(n_73)
);

NAND2xp5_ASAP7_75t_L g75 ( 
.A(n_73),
.B(n_67),
.Y(n_75)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_75),
.Y(n_77)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_72),
.Y(n_76)
);

NAND2xp5_ASAP7_75t_L g78 ( 
.A(n_77),
.B(n_76),
.Y(n_78)
);

CKINVDCx20_ASAP7_75t_R g79 ( 
.A(n_78),
.Y(n_79)
);

AND2x2_ASAP7_75t_L g80 ( 
.A(n_79),
.B(n_66),
.Y(n_80)
);

NOR4xp25_ASAP7_75t_L g81 ( 
.A(n_80),
.B(n_74),
.C(n_70),
.D(n_29),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_L g82 ( 
.A(n_81),
.B(n_31),
.Y(n_82)
);

NOR2xp33_ASAP7_75t_L g83 ( 
.A(n_82),
.B(n_56),
.Y(n_83)
);


endmodule