module fake_ibex_1620_n_3555 (n_151, n_85, n_599, n_507, n_540, n_395, n_84, n_64, n_171, n_103, n_529, n_389, n_204, n_626, n_274, n_387, n_688, n_130, n_177, n_76, n_273, n_309, n_330, n_9, n_328, n_293, n_341, n_372, n_124, n_37, n_256, n_418, n_193, n_510, n_446, n_108, n_350, n_601, n_621, n_610, n_165, n_452, n_86, n_70, n_664, n_255, n_175, n_586, n_638, n_398, n_59, n_28, n_125, n_304, n_191, n_593, n_5, n_62, n_71, n_153, n_545, n_583, n_678, n_663, n_194, n_249, n_334, n_634, n_312, n_622, n_578, n_478, n_239, n_94, n_134, n_432, n_371, n_403, n_423, n_608, n_357, n_88, n_412, n_457, n_494, n_142, n_226, n_336, n_258, n_40, n_90, n_17, n_74, n_449, n_547, n_176, n_58, n_43, n_216, n_33, n_652, n_421, n_475, n_166, n_163, n_645, n_500, n_542, n_114, n_236, n_34, n_376, n_377, n_584, n_531, n_647, n_15, n_556, n_24, n_189, n_498, n_698, n_280, n_317, n_340, n_375, n_105, n_187, n_667, n_1, n_154, n_682, n_182, n_196, n_326, n_327, n_89, n_50, n_144, n_170, n_270, n_346, n_383, n_113, n_561, n_117, n_417, n_471, n_265, n_504, n_158, n_259, n_276, n_339, n_470, n_210, n_348, n_220, n_674, n_91, n_481, n_287, n_54, n_243, n_19, n_497, n_671, n_228, n_147, n_552, n_251, n_384, n_632, n_373, n_458, n_244, n_73, n_343, n_310, n_426, n_323, n_469, n_598, n_143, n_106, n_386, n_549, n_8, n_224, n_183, n_533, n_508, n_67, n_453, n_591, n_655, n_333, n_110, n_306, n_400, n_47, n_550, n_169, n_10, n_673, n_21, n_242, n_278, n_316, n_16, n_404, n_60, n_557, n_641, n_7, n_109, n_127, n_121, n_527, n_590, n_465, n_48, n_325, n_57, n_301, n_496, n_617, n_434, n_296, n_690, n_120, n_168, n_526, n_155, n_315, n_441, n_604, n_13, n_637, n_122, n_523, n_116, n_694, n_614, n_370, n_431, n_574, n_0, n_289, n_12, n_515, n_642, n_150, n_286, n_321, n_133, n_569, n_600, n_51, n_215, n_279, n_49, n_374, n_235, n_464, n_538, n_669, n_22, n_136, n_261, n_521, n_665, n_459, n_30, n_518, n_367, n_221, n_654, n_656, n_437, n_602, n_355, n_474, n_594, n_636, n_407, n_102, n_490, n_568, n_52, n_448, n_646, n_595, n_99, n_466, n_269, n_156, n_570, n_126, n_623, n_585, n_530, n_356, n_25, n_104, n_45, n_420, n_483, n_543, n_580, n_141, n_487, n_222, n_660, n_186, n_524, n_349, n_454, n_295, n_331, n_576, n_230, n_96, n_185, n_388, n_625, n_619, n_536, n_611, n_352, n_290, n_558, n_666, n_174, n_467, n_427, n_607, n_157, n_219, n_246, n_31, n_442, n_146, n_207, n_438, n_689, n_167, n_676, n_128, n_253, n_208, n_234, n_3, n_152, n_300, n_145, n_65, n_358, n_205, n_618, n_488, n_139, n_514, n_429, n_560, n_275, n_541, n_98, n_129, n_613, n_659, n_267, n_662, n_635, n_245, n_589, n_571, n_229, n_209, n_472, n_648, n_347, n_473, n_445, n_629, n_335, n_413, n_82, n_263, n_27, n_573, n_353, n_359, n_299, n_87, n_262, n_433, n_75, n_439, n_643, n_137, n_679, n_338, n_173, n_696, n_477, n_640, n_363, n_402, n_180, n_369, n_596, n_201, n_699, n_14, n_351, n_368, n_456, n_257, n_77, n_44, n_672, n_401, n_553, n_554, n_66, n_305, n_307, n_192, n_140, n_484, n_566, n_480, n_416, n_581, n_651, n_365, n_4, n_6, n_605, n_539, n_100, n_179, n_354, n_206, n_392, n_630, n_516, n_548, n_567, n_329, n_447, n_26, n_188, n_200, n_444, n_506, n_562, n_564, n_546, n_199, n_592, n_495, n_410, n_308, n_675, n_463, n_624, n_411, n_135, n_520, n_684, n_658, n_512, n_615, n_685, n_283, n_366, n_397, n_111, n_692, n_36, n_627, n_18, n_322, n_53, n_227, n_499, n_115, n_11, n_248, n_92, n_702, n_451, n_101, n_190, n_138, n_650, n_409, n_582, n_653, n_214, n_238, n_579, n_332, n_517, n_211, n_218, n_314, n_691, n_563, n_132, n_277, n_555, n_337, n_522, n_700, n_479, n_534, n_225, n_360, n_272, n_511, n_23, n_468, n_223, n_381, n_525, n_535, n_382, n_502, n_681, n_633, n_532, n_95, n_405, n_415, n_597, n_285, n_288, n_247, n_320, n_379, n_551, n_55, n_612, n_291, n_318, n_63, n_161, n_237, n_29, n_203, n_268, n_440, n_148, n_2, n_342, n_233, n_385, n_414, n_430, n_118, n_603, n_378, n_486, n_422, n_164, n_38, n_198, n_264, n_616, n_217, n_324, n_391, n_537, n_78, n_670, n_20, n_69, n_390, n_544, n_39, n_178, n_509, n_695, n_639, n_303, n_362, n_93, n_505, n_162, n_482, n_240, n_282, n_61, n_680, n_501, n_668, n_266, n_42, n_294, n_112, n_485, n_46, n_284, n_80, n_172, n_250, n_493, n_460, n_609, n_476, n_461, n_575, n_313, n_519, n_345, n_408, n_119, n_361, n_455, n_419, n_72, n_319, n_195, n_513, n_212, n_588, n_693, n_311, n_661, n_406, n_606, n_97, n_197, n_528, n_181, n_131, n_123, n_631, n_683, n_260, n_620, n_462, n_302, n_450, n_443, n_686, n_572, n_644, n_577, n_344, n_393, n_436, n_428, n_491, n_297, n_435, n_628, n_41, n_252, n_396, n_697, n_83, n_32, n_107, n_149, n_489, n_677, n_399, n_254, n_213, n_424, n_565, n_701, n_271, n_241, n_68, n_503, n_292, n_394, n_79, n_81, n_35, n_364, n_687, n_159, n_202, n_231, n_298, n_587, n_160, n_657, n_184, n_56, n_492, n_649, n_232, n_380, n_281, n_559, n_425, n_3555);

input n_151;
input n_85;
input n_599;
input n_507;
input n_540;
input n_395;
input n_84;
input n_64;
input n_171;
input n_103;
input n_529;
input n_389;
input n_204;
input n_626;
input n_274;
input n_387;
input n_688;
input n_130;
input n_177;
input n_76;
input n_273;
input n_309;
input n_330;
input n_9;
input n_328;
input n_293;
input n_341;
input n_372;
input n_124;
input n_37;
input n_256;
input n_418;
input n_193;
input n_510;
input n_446;
input n_108;
input n_350;
input n_601;
input n_621;
input n_610;
input n_165;
input n_452;
input n_86;
input n_70;
input n_664;
input n_255;
input n_175;
input n_586;
input n_638;
input n_398;
input n_59;
input n_28;
input n_125;
input n_304;
input n_191;
input n_593;
input n_5;
input n_62;
input n_71;
input n_153;
input n_545;
input n_583;
input n_678;
input n_663;
input n_194;
input n_249;
input n_334;
input n_634;
input n_312;
input n_622;
input n_578;
input n_478;
input n_239;
input n_94;
input n_134;
input n_432;
input n_371;
input n_403;
input n_423;
input n_608;
input n_357;
input n_88;
input n_412;
input n_457;
input n_494;
input n_142;
input n_226;
input n_336;
input n_258;
input n_40;
input n_90;
input n_17;
input n_74;
input n_449;
input n_547;
input n_176;
input n_58;
input n_43;
input n_216;
input n_33;
input n_652;
input n_421;
input n_475;
input n_166;
input n_163;
input n_645;
input n_500;
input n_542;
input n_114;
input n_236;
input n_34;
input n_376;
input n_377;
input n_584;
input n_531;
input n_647;
input n_15;
input n_556;
input n_24;
input n_189;
input n_498;
input n_698;
input n_280;
input n_317;
input n_340;
input n_375;
input n_105;
input n_187;
input n_667;
input n_1;
input n_154;
input n_682;
input n_182;
input n_196;
input n_326;
input n_327;
input n_89;
input n_50;
input n_144;
input n_170;
input n_270;
input n_346;
input n_383;
input n_113;
input n_561;
input n_117;
input n_417;
input n_471;
input n_265;
input n_504;
input n_158;
input n_259;
input n_276;
input n_339;
input n_470;
input n_210;
input n_348;
input n_220;
input n_674;
input n_91;
input n_481;
input n_287;
input n_54;
input n_243;
input n_19;
input n_497;
input n_671;
input n_228;
input n_147;
input n_552;
input n_251;
input n_384;
input n_632;
input n_373;
input n_458;
input n_244;
input n_73;
input n_343;
input n_310;
input n_426;
input n_323;
input n_469;
input n_598;
input n_143;
input n_106;
input n_386;
input n_549;
input n_8;
input n_224;
input n_183;
input n_533;
input n_508;
input n_67;
input n_453;
input n_591;
input n_655;
input n_333;
input n_110;
input n_306;
input n_400;
input n_47;
input n_550;
input n_169;
input n_10;
input n_673;
input n_21;
input n_242;
input n_278;
input n_316;
input n_16;
input n_404;
input n_60;
input n_557;
input n_641;
input n_7;
input n_109;
input n_127;
input n_121;
input n_527;
input n_590;
input n_465;
input n_48;
input n_325;
input n_57;
input n_301;
input n_496;
input n_617;
input n_434;
input n_296;
input n_690;
input n_120;
input n_168;
input n_526;
input n_155;
input n_315;
input n_441;
input n_604;
input n_13;
input n_637;
input n_122;
input n_523;
input n_116;
input n_694;
input n_614;
input n_370;
input n_431;
input n_574;
input n_0;
input n_289;
input n_12;
input n_515;
input n_642;
input n_150;
input n_286;
input n_321;
input n_133;
input n_569;
input n_600;
input n_51;
input n_215;
input n_279;
input n_49;
input n_374;
input n_235;
input n_464;
input n_538;
input n_669;
input n_22;
input n_136;
input n_261;
input n_521;
input n_665;
input n_459;
input n_30;
input n_518;
input n_367;
input n_221;
input n_654;
input n_656;
input n_437;
input n_602;
input n_355;
input n_474;
input n_594;
input n_636;
input n_407;
input n_102;
input n_490;
input n_568;
input n_52;
input n_448;
input n_646;
input n_595;
input n_99;
input n_466;
input n_269;
input n_156;
input n_570;
input n_126;
input n_623;
input n_585;
input n_530;
input n_356;
input n_25;
input n_104;
input n_45;
input n_420;
input n_483;
input n_543;
input n_580;
input n_141;
input n_487;
input n_222;
input n_660;
input n_186;
input n_524;
input n_349;
input n_454;
input n_295;
input n_331;
input n_576;
input n_230;
input n_96;
input n_185;
input n_388;
input n_625;
input n_619;
input n_536;
input n_611;
input n_352;
input n_290;
input n_558;
input n_666;
input n_174;
input n_467;
input n_427;
input n_607;
input n_157;
input n_219;
input n_246;
input n_31;
input n_442;
input n_146;
input n_207;
input n_438;
input n_689;
input n_167;
input n_676;
input n_128;
input n_253;
input n_208;
input n_234;
input n_3;
input n_152;
input n_300;
input n_145;
input n_65;
input n_358;
input n_205;
input n_618;
input n_488;
input n_139;
input n_514;
input n_429;
input n_560;
input n_275;
input n_541;
input n_98;
input n_129;
input n_613;
input n_659;
input n_267;
input n_662;
input n_635;
input n_245;
input n_589;
input n_571;
input n_229;
input n_209;
input n_472;
input n_648;
input n_347;
input n_473;
input n_445;
input n_629;
input n_335;
input n_413;
input n_82;
input n_263;
input n_27;
input n_573;
input n_353;
input n_359;
input n_299;
input n_87;
input n_262;
input n_433;
input n_75;
input n_439;
input n_643;
input n_137;
input n_679;
input n_338;
input n_173;
input n_696;
input n_477;
input n_640;
input n_363;
input n_402;
input n_180;
input n_369;
input n_596;
input n_201;
input n_699;
input n_14;
input n_351;
input n_368;
input n_456;
input n_257;
input n_77;
input n_44;
input n_672;
input n_401;
input n_553;
input n_554;
input n_66;
input n_305;
input n_307;
input n_192;
input n_140;
input n_484;
input n_566;
input n_480;
input n_416;
input n_581;
input n_651;
input n_365;
input n_4;
input n_6;
input n_605;
input n_539;
input n_100;
input n_179;
input n_354;
input n_206;
input n_392;
input n_630;
input n_516;
input n_548;
input n_567;
input n_329;
input n_447;
input n_26;
input n_188;
input n_200;
input n_444;
input n_506;
input n_562;
input n_564;
input n_546;
input n_199;
input n_592;
input n_495;
input n_410;
input n_308;
input n_675;
input n_463;
input n_624;
input n_411;
input n_135;
input n_520;
input n_684;
input n_658;
input n_512;
input n_615;
input n_685;
input n_283;
input n_366;
input n_397;
input n_111;
input n_692;
input n_36;
input n_627;
input n_18;
input n_322;
input n_53;
input n_227;
input n_499;
input n_115;
input n_11;
input n_248;
input n_92;
input n_702;
input n_451;
input n_101;
input n_190;
input n_138;
input n_650;
input n_409;
input n_582;
input n_653;
input n_214;
input n_238;
input n_579;
input n_332;
input n_517;
input n_211;
input n_218;
input n_314;
input n_691;
input n_563;
input n_132;
input n_277;
input n_555;
input n_337;
input n_522;
input n_700;
input n_479;
input n_534;
input n_225;
input n_360;
input n_272;
input n_511;
input n_23;
input n_468;
input n_223;
input n_381;
input n_525;
input n_535;
input n_382;
input n_502;
input n_681;
input n_633;
input n_532;
input n_95;
input n_405;
input n_415;
input n_597;
input n_285;
input n_288;
input n_247;
input n_320;
input n_379;
input n_551;
input n_55;
input n_612;
input n_291;
input n_318;
input n_63;
input n_161;
input n_237;
input n_29;
input n_203;
input n_268;
input n_440;
input n_148;
input n_2;
input n_342;
input n_233;
input n_385;
input n_414;
input n_430;
input n_118;
input n_603;
input n_378;
input n_486;
input n_422;
input n_164;
input n_38;
input n_198;
input n_264;
input n_616;
input n_217;
input n_324;
input n_391;
input n_537;
input n_78;
input n_670;
input n_20;
input n_69;
input n_390;
input n_544;
input n_39;
input n_178;
input n_509;
input n_695;
input n_639;
input n_303;
input n_362;
input n_93;
input n_505;
input n_162;
input n_482;
input n_240;
input n_282;
input n_61;
input n_680;
input n_501;
input n_668;
input n_266;
input n_42;
input n_294;
input n_112;
input n_485;
input n_46;
input n_284;
input n_80;
input n_172;
input n_250;
input n_493;
input n_460;
input n_609;
input n_476;
input n_461;
input n_575;
input n_313;
input n_519;
input n_345;
input n_408;
input n_119;
input n_361;
input n_455;
input n_419;
input n_72;
input n_319;
input n_195;
input n_513;
input n_212;
input n_588;
input n_693;
input n_311;
input n_661;
input n_406;
input n_606;
input n_97;
input n_197;
input n_528;
input n_181;
input n_131;
input n_123;
input n_631;
input n_683;
input n_260;
input n_620;
input n_462;
input n_302;
input n_450;
input n_443;
input n_686;
input n_572;
input n_644;
input n_577;
input n_344;
input n_393;
input n_436;
input n_428;
input n_491;
input n_297;
input n_435;
input n_628;
input n_41;
input n_252;
input n_396;
input n_697;
input n_83;
input n_32;
input n_107;
input n_149;
input n_489;
input n_677;
input n_399;
input n_254;
input n_213;
input n_424;
input n_565;
input n_701;
input n_271;
input n_241;
input n_68;
input n_503;
input n_292;
input n_394;
input n_79;
input n_81;
input n_35;
input n_364;
input n_687;
input n_159;
input n_202;
input n_231;
input n_298;
input n_587;
input n_160;
input n_657;
input n_184;
input n_56;
input n_492;
input n_649;
input n_232;
input n_380;
input n_281;
input n_559;
input n_425;

output n_3555;

wire n_1084;
wire n_2594;
wire n_1474;
wire n_1295;
wire n_1983;
wire n_2804;
wire n_3150;
wire n_992;
wire n_1582;
wire n_2201;
wire n_2512;
wire n_766;
wire n_2960;
wire n_2175;
wire n_2071;
wire n_2796;
wire n_1110;
wire n_3548;
wire n_2607;
wire n_1382;
wire n_3144;
wire n_2569;
wire n_2949;
wire n_1998;
wire n_2840;
wire n_1596;
wire n_926;
wire n_3319;
wire n_1079;
wire n_3077;
wire n_2835;
wire n_1100;
wire n_845;
wire n_2177;
wire n_2123;
wire n_1930;
wire n_1234;
wire n_3019;
wire n_2047;
wire n_1594;
wire n_1944;
wire n_2498;
wire n_1802;
wire n_2235;
wire n_773;
wire n_2038;
wire n_2504;
wire n_1469;
wire n_821;
wire n_2017;
wire n_873;
wire n_1227;
wire n_962;
wire n_1080;
wire n_862;
wire n_909;
wire n_2290;
wire n_957;
wire n_3272;
wire n_3255;
wire n_1652;
wire n_969;
wire n_1859;
wire n_2183;
wire n_1954;
wire n_2074;
wire n_2897;
wire n_1883;
wire n_1125;
wire n_733;
wire n_2687;
wire n_3456;
wire n_2037;
wire n_1226;
wire n_1034;
wire n_2383;
wire n_3132;
wire n_1765;
wire n_872;
wire n_2392;
wire n_1873;
wire n_1619;
wire n_1666;
wire n_2640;
wire n_2682;
wire n_930;
wire n_1044;
wire n_3280;
wire n_3105;
wire n_3146;
wire n_1492;
wire n_1134;
wire n_1478;
wire n_1684;
wire n_1796;
wire n_1614;
wire n_2374;
wire n_3334;
wire n_2598;
wire n_1722;
wire n_911;
wire n_2023;
wire n_781;
wire n_2720;
wire n_802;
wire n_3340;
wire n_2322;
wire n_1233;
wire n_2335;
wire n_3025;
wire n_3411;
wire n_2955;
wire n_3458;
wire n_3519;
wire n_2276;
wire n_1045;
wire n_3235;
wire n_2989;
wire n_1856;
wire n_963;
wire n_1782;
wire n_2230;
wire n_2889;
wire n_2139;
wire n_2847;
wire n_3033;
wire n_1308;
wire n_1138;
wire n_2943;
wire n_708;
wire n_1096;
wire n_2151;
wire n_2391;
wire n_1391;
wire n_3338;
wire n_3168;
wire n_884;
wire n_2396;
wire n_3135;
wire n_3440;
wire n_850;
wire n_3175;
wire n_3484;
wire n_1971;
wire n_2485;
wire n_2479;
wire n_879;
wire n_2179;
wire n_1957;
wire n_2188;
wire n_723;
wire n_1144;
wire n_2360;
wire n_2359;
wire n_2506;
wire n_1392;
wire n_2158;
wire n_1268;
wire n_2571;
wire n_3187;
wire n_739;
wire n_2724;
wire n_3086;
wire n_2475;
wire n_853;
wire n_948;
wire n_2799;
wire n_1752;
wire n_1829;
wire n_1338;
wire n_1730;
wire n_875;
wire n_1307;
wire n_1327;
wire n_2644;
wire n_876;
wire n_3211;
wire n_711;
wire n_1840;
wire n_2837;
wire n_3479;
wire n_989;
wire n_3262;
wire n_3407;
wire n_1908;
wire n_3315;
wire n_3537;
wire n_1668;
wire n_2343;
wire n_2605;
wire n_2887;
wire n_1641;
wire n_829;
wire n_2565;
wire n_825;
wire n_1480;
wire n_1463;
wire n_1823;
wire n_3251;
wire n_1681;
wire n_2921;
wire n_939;
wire n_1636;
wire n_1687;
wire n_3192;
wire n_3533;
wire n_2192;
wire n_1766;
wire n_3184;
wire n_3469;
wire n_3170;
wire n_1922;
wire n_2032;
wire n_2820;
wire n_3323;
wire n_1937;
wire n_2311;
wire n_3392;
wire n_3347;
wire n_893;
wire n_3242;
wire n_3395;
wire n_1654;
wire n_2995;
wire n_3330;
wire n_1258;
wire n_1344;
wire n_2208;
wire n_2198;
wire n_1929;
wire n_2707;
wire n_3472;
wire n_3509;
wire n_1749;
wire n_1680;
wire n_835;
wire n_1981;
wire n_1195;
wire n_2918;
wire n_3353;
wire n_824;
wire n_1945;
wire n_2638;
wire n_787;
wire n_2860;
wire n_2448;
wire n_2015;
wire n_2537;
wire n_1130;
wire n_2643;
wire n_1228;
wire n_2998;
wire n_2336;
wire n_2163;
wire n_1081;
wire n_2354;
wire n_1155;
wire n_1292;
wire n_2432;
wire n_3043;
wire n_2873;
wire n_1576;
wire n_1664;
wire n_2273;
wire n_3298;
wire n_852;
wire n_1427;
wire n_1133;
wire n_3049;
wire n_2421;
wire n_1926;
wire n_3208;
wire n_904;
wire n_2363;
wire n_2814;
wire n_3237;
wire n_3264;
wire n_3204;
wire n_2003;
wire n_1970;
wire n_2621;
wire n_1778;
wire n_2558;
wire n_2953;
wire n_2922;
wire n_2347;
wire n_3507;
wire n_3103;
wire n_2839;
wire n_1030;
wire n_1698;
wire n_1094;
wire n_2462;
wire n_1496;
wire n_1910;
wire n_715;
wire n_2436;
wire n_1663;
wire n_2333;
wire n_1214;
wire n_1274;
wire n_2705;
wire n_2527;
wire n_1606;
wire n_769;
wire n_1595;
wire n_2164;
wire n_1509;
wire n_1648;
wire n_1618;
wire n_2944;
wire n_1886;
wire n_2269;
wire n_857;
wire n_765;
wire n_1070;
wire n_1841;
wire n_2472;
wire n_777;
wire n_2685;
wire n_2846;
wire n_3197;
wire n_1955;
wire n_917;
wire n_2249;
wire n_3148;
wire n_2362;
wire n_968;
wire n_3022;
wire n_2413;
wire n_2822;
wire n_1253;
wire n_1306;
wire n_1484;
wire n_2686;
wire n_1493;
wire n_2597;
wire n_1313;
wire n_2774;
wire n_3151;
wire n_2090;
wire n_2260;
wire n_3125;
wire n_2812;
wire n_2753;
wire n_1638;
wire n_2215;
wire n_1071;
wire n_1449;
wire n_1723;
wire n_1960;
wire n_2663;
wire n_793;
wire n_3129;
wire n_937;
wire n_2595;
wire n_2116;
wire n_1645;
wire n_3186;
wire n_973;
wire n_1038;
wire n_2280;
wire n_1943;
wire n_3541;
wire n_1863;
wire n_2844;
wire n_1269;
wire n_2393;
wire n_2773;
wire n_2906;
wire n_3030;
wire n_3097;
wire n_979;
wire n_1309;
wire n_1999;
wire n_1316;
wire n_1562;
wire n_1215;
wire n_2777;
wire n_2480;
wire n_1445;
wire n_2283;
wire n_2806;
wire n_2813;
wire n_2147;
wire n_1716;
wire n_1466;
wire n_1412;
wire n_3210;
wire n_3221;
wire n_1672;
wire n_1007;
wire n_2253;
wire n_1276;
wire n_1637;
wire n_3310;
wire n_841;
wire n_2900;
wire n_772;
wire n_810;
wire n_1401;
wire n_1817;
wire n_2951;
wire n_2145;
wire n_2122;
wire n_1588;
wire n_2216;
wire n_1301;
wire n_2579;
wire n_2876;
wire n_2242;
wire n_869;
wire n_1620;
wire n_1561;
wire n_718;
wire n_3301;
wire n_2370;
wire n_2025;
wire n_1078;
wire n_2247;
wire n_3451;
wire n_1219;
wire n_713;
wire n_1865;
wire n_3177;
wire n_3518;
wire n_3399;
wire n_1252;
wire n_2022;
wire n_2730;
wire n_1170;
wire n_1927;
wire n_2373;
wire n_1869;
wire n_1853;
wire n_2275;
wire n_2980;
wire n_2189;
wire n_2482;
wire n_745;
wire n_2767;
wire n_2826;
wire n_2899;
wire n_2112;
wire n_1753;
wire n_3351;
wire n_1322;
wire n_2008;
wire n_1305;
wire n_2088;
wire n_795;
wire n_1248;
wire n_2762;
wire n_2171;
wire n_3307;
wire n_762;
wire n_1388;
wire n_2859;
wire n_800;
wire n_2564;
wire n_706;
wire n_3023;
wire n_784;
wire n_1653;
wire n_1375;
wire n_3224;
wire n_1356;
wire n_894;
wire n_1118;
wire n_2591;
wire n_1881;
wire n_1969;
wire n_709;
wire n_1296;
wire n_3060;
wire n_1326;
wire n_971;
wire n_1350;
wire n_906;
wire n_2957;
wire n_2586;
wire n_1093;
wire n_1764;
wire n_2412;
wire n_2783;
wire n_978;
wire n_899;
wire n_1799;
wire n_3293;
wire n_1019;
wire n_902;
wire n_1689;
wire n_1250;
wire n_2550;
wire n_1190;
wire n_1304;
wire n_744;
wire n_2541;
wire n_2987;
wire n_881;
wire n_3259;
wire n_1702;
wire n_3381;
wire n_734;
wire n_1558;
wire n_2750;
wire n_1650;
wire n_1520;
wire n_1073;
wire n_1453;
wire n_1108;
wire n_2722;
wire n_2509;
wire n_2727;
wire n_1794;
wire n_1423;
wire n_1239;
wire n_2399;
wire n_1370;
wire n_2719;
wire n_1209;
wire n_1708;
wire n_2213;
wire n_3038;
wire n_3521;
wire n_3203;
wire n_3295;
wire n_2723;
wire n_1616;
wire n_3199;
wire n_3093;
wire n_729;
wire n_1569;
wire n_2664;
wire n_1434;
wire n_1649;
wire n_2389;
wire n_3450;
wire n_1936;
wire n_2114;
wire n_1717;
wire n_2107;
wire n_1609;
wire n_2257;
wire n_3435;
wire n_3530;
wire n_1613;
wire n_820;
wire n_805;
wire n_1988;
wire n_1132;
wire n_892;
wire n_1467;
wire n_1803;
wire n_2401;
wire n_1787;
wire n_2782;
wire n_2511;
wire n_3217;
wire n_1281;
wire n_3094;
wire n_1447;
wire n_2166;
wire n_2451;
wire n_2150;
wire n_1549;
wire n_2631;
wire n_1867;
wire n_1531;
wire n_2919;
wire n_1332;
wire n_2660;
wire n_2661;
wire n_2292;
wire n_3510;
wire n_2334;
wire n_1424;
wire n_3467;
wire n_2444;
wire n_2350;
wire n_1742;
wire n_2625;
wire n_1818;
wire n_870;
wire n_2199;
wire n_1709;
wire n_1610;
wire n_2219;
wire n_1298;
wire n_1844;
wire n_1387;
wire n_2649;
wire n_1040;
wire n_2203;
wire n_2693;
wire n_3194;
wire n_3371;
wire n_1159;
wire n_1368;
wire n_2281;
wire n_1154;
wire n_3202;
wire n_2539;
wire n_2431;
wire n_1701;
wire n_2084;
wire n_1243;
wire n_2387;
wire n_2646;
wire n_3375;
wire n_2397;
wire n_1121;
wire n_2746;
wire n_3241;
wire n_2256;
wire n_3317;
wire n_737;
wire n_2445;
wire n_3461;
wire n_2729;
wire n_1571;
wire n_1980;
wire n_3355;
wire n_2529;
wire n_2019;
wire n_1407;
wire n_3282;
wire n_1235;
wire n_1821;
wire n_3508;
wire n_1003;
wire n_889;
wire n_2708;
wire n_3156;
wire n_3457;
wire n_2748;
wire n_816;
wire n_1058;
wire n_1835;
wire n_1862;
wire n_2224;
wire n_2697;
wire n_3531;
wire n_3415;
wire n_2470;
wire n_2355;
wire n_2890;
wire n_2731;
wire n_1543;
wire n_3466;
wire n_3386;
wire n_823;
wire n_2233;
wire n_2499;
wire n_3370;
wire n_1504;
wire n_1519;
wire n_1425;
wire n_1781;
wire n_2069;
wire n_2602;
wire n_1441;
wire n_2028;
wire n_3309;
wire n_1924;
wire n_2856;
wire n_1921;
wire n_3024;
wire n_1156;
wire n_2857;
wire n_1293;
wire n_1360;
wire n_749;
wire n_1555;
wire n_1394;
wire n_1347;
wire n_819;
wire n_2070;
wire n_1042;
wire n_822;
wire n_1888;
wire n_3471;
wire n_743;
wire n_3117;
wire n_3320;
wire n_754;
wire n_1786;
wire n_2033;
wire n_3039;
wire n_1319;
wire n_1553;
wire n_3478;
wire n_3542;
wire n_1041;
wire n_2766;
wire n_2828;
wire n_1964;
wire n_1090;
wire n_3374;
wire n_1196;
wire n_1182;
wire n_1271;
wire n_2416;
wire n_2786;
wire n_1731;
wire n_1905;
wire n_2962;
wire n_1031;
wire n_3416;
wire n_2879;
wire n_2958;
wire n_3147;
wire n_2052;
wire n_981;
wire n_2425;
wire n_2800;
wire n_3514;
wire n_3091;
wire n_3006;
wire n_3348;
wire n_2118;
wire n_2259;
wire n_2162;
wire n_2236;
wire n_3455;
wire n_2377;
wire n_2718;
wire n_2577;
wire n_1591;
wire n_3426;
wire n_3165;
wire n_2289;
wire n_2288;
wire n_2841;
wire n_3075;
wire n_1671;
wire n_1795;
wire n_1409;
wire n_1015;
wire n_3448;
wire n_2744;
wire n_2101;
wire n_2795;
wire n_3524;
wire n_1377;
wire n_2473;
wire n_1583;
wire n_3520;
wire n_1521;
wire n_2632;
wire n_1152;
wire n_2456;
wire n_2924;
wire n_3054;
wire n_2264;
wire n_2076;
wire n_1036;
wire n_974;
wire n_2599;
wire n_1831;
wire n_864;
wire n_1987;
wire n_959;
wire n_1106;
wire n_1312;
wire n_1129;
wire n_1244;
wire n_3171;
wire n_1733;
wire n_3365;
wire n_1634;
wire n_2853;
wire n_1932;
wire n_1552;
wire n_1452;
wire n_1318;
wire n_1508;
wire n_2217;
wire n_738;
wire n_1217;
wire n_2866;
wire n_3153;
wire n_3291;
wire n_2655;
wire n_3487;
wire n_2454;
wire n_1715;
wire n_1189;
wire n_3300;
wire n_761;
wire n_748;
wire n_1713;
wire n_901;
wire n_1577;
wire n_2036;
wire n_1255;
wire n_2829;
wire n_2968;
wire n_2740;
wire n_3473;
wire n_1700;
wire n_2623;
wire n_2622;
wire n_3232;
wire n_2819;
wire n_1218;
wire n_2178;
wire n_1181;
wire n_3263;
wire n_1140;
wire n_1985;
wire n_1772;
wire n_2858;
wire n_1056;
wire n_2626;
wire n_1283;
wire n_3007;
wire n_1446;
wire n_2404;
wire n_1487;
wire n_3078;
wire n_2789;
wire n_2603;
wire n_840;
wire n_1203;
wire n_1421;
wire n_3218;
wire n_2821;
wire n_2424;
wire n_846;
wire n_1793;
wire n_1237;
wire n_2573;
wire n_2390;
wire n_2880;
wire n_2423;
wire n_859;
wire n_1109;
wire n_965;
wire n_2741;
wire n_2793;
wire n_3098;
wire n_3490;
wire n_3055;
wire n_1633;
wire n_3299;
wire n_2580;
wire n_3222;
wire n_1711;
wire n_3529;
wire n_3069;
wire n_3107;
wire n_3352;
wire n_3436;
wire n_1051;
wire n_1008;
wire n_3065;
wire n_2964;
wire n_2375;
wire n_1498;
wire n_2312;
wire n_2572;
wire n_2946;
wire n_1053;
wire n_1656;
wire n_1207;
wire n_1076;
wire n_1735;
wire n_2063;
wire n_1032;
wire n_936;
wire n_3082;
wire n_2176;
wire n_1884;
wire n_1825;
wire n_2805;
wire n_1589;
wire n_2717;
wire n_2204;
wire n_2863;
wire n_2575;
wire n_1210;
wire n_2319;
wire n_2877;
wire n_1933;
wire n_2522;
wire n_3357;
wire n_1996;
wire n_1510;
wire n_1201;
wire n_1842;
wire n_2852;
wire n_2132;
wire n_3110;
wire n_1246;
wire n_1677;
wire n_732;
wire n_1236;
wire n_3364;
wire n_832;
wire n_2297;
wire n_3429;
wire n_3306;
wire n_3412;
wire n_3037;
wire n_3188;
wire n_2780;
wire n_1792;
wire n_1712;
wire n_3250;
wire n_1984;
wire n_1568;
wire n_2885;
wire n_1877;
wire n_3445;
wire n_1184;
wire n_1477;
wire n_2080;
wire n_2220;
wire n_2585;
wire n_1724;
wire n_2554;
wire n_3155;
wire n_2838;
wire n_1364;
wire n_3183;
wire n_1540;
wire n_1676;
wire n_1013;
wire n_3243;
wire n_2468;
wire n_929;
wire n_3248;
wire n_3214;
wire n_1136;
wire n_1890;
wire n_1075;
wire n_1249;
wire n_3128;
wire n_1918;
wire n_2606;
wire n_2549;
wire n_2461;
wire n_3468;
wire n_2006;
wire n_2440;
wire n_1229;
wire n_1440;
wire n_1490;
wire n_2152;
wire n_907;
wire n_1179;
wire n_1990;
wire n_1153;
wire n_1751;
wire n_2787;
wire n_2467;
wire n_2146;
wire n_2341;
wire n_3525;
wire n_1737;
wire n_3145;
wire n_2779;
wire n_1117;
wire n_1273;
wire n_2547;
wire n_2930;
wire n_2616;
wire n_1748;
wire n_2662;
wire n_1083;
wire n_3205;
wire n_1014;
wire n_724;
wire n_2883;
wire n_938;
wire n_1178;
wire n_2935;
wire n_878;
wire n_2441;
wire n_3503;
wire n_2358;
wire n_2490;
wire n_3127;
wire n_3496;
wire n_2361;
wire n_1566;
wire n_1464;
wire n_944;
wire n_3312;
wire n_3003;
wire n_1848;
wire n_2062;
wire n_2277;
wire n_2650;
wire n_1982;
wire n_2252;
wire n_2888;
wire n_2339;
wire n_1334;
wire n_1963;
wire n_3394;
wire n_1695;
wire n_1418;
wire n_3331;
wire n_2402;
wire n_1137;
wire n_2552;
wire n_2910;
wire n_2999;
wire n_2590;
wire n_3119;
wire n_1977;
wire n_2294;
wire n_1200;
wire n_2295;
wire n_2530;
wire n_3345;
wire n_2379;
wire n_1120;
wire n_2300;
wire n_2792;
wire n_1602;
wire n_2965;
wire n_1776;
wire n_2372;
wire n_3341;
wire n_2382;
wire n_1852;
wire n_1522;
wire n_2523;
wire n_2557;
wire n_3544;
wire n_1279;
wire n_2505;
wire n_931;
wire n_3488;
wire n_827;
wire n_3554;
wire n_2481;
wire n_1064;
wire n_1408;
wire n_2832;
wire n_1028;
wire n_1264;
wire n_3535;
wire n_2808;
wire n_2287;
wire n_3396;
wire n_2954;
wire n_3526;
wire n_2102;
wire n_1935;
wire n_2046;
wire n_3367;
wire n_3492;
wire n_1146;
wire n_2785;
wire n_2751;
wire n_705;
wire n_2142;
wire n_1548;
wire n_2977;
wire n_1682;
wire n_1608;
wire n_1009;
wire n_1260;
wire n_1896;
wire n_1704;
wire n_2160;
wire n_2699;
wire n_2234;
wire n_847;
wire n_2991;
wire n_1436;
wire n_3239;
wire n_2600;
wire n_1069;
wire n_1485;
wire n_2239;
wire n_1465;
wire n_1352;
wire n_1171;
wire n_1126;
wire n_1232;
wire n_1979;
wire n_2328;
wire n_2715;
wire n_1345;
wire n_2434;
wire n_837;
wire n_1590;
wire n_2332;
wire n_2971;
wire n_954;
wire n_1628;
wire n_725;
wire n_1773;
wire n_2133;
wire n_3553;
wire n_3072;
wire n_1545;
wire n_3249;
wire n_2369;
wire n_3470;
wire n_1471;
wire n_1738;
wire n_3441;
wire n_1115;
wire n_998;
wire n_1395;
wire n_1729;
wire n_2551;
wire n_3281;
wire n_801;
wire n_2823;
wire n_3274;
wire n_2094;
wire n_2613;
wire n_1479;
wire n_3505;
wire n_2306;
wire n_1046;
wire n_2419;
wire n_3397;
wire n_2934;
wire n_2807;
wire n_882;
wire n_942;
wire n_1627;
wire n_1431;
wire n_721;
wire n_2525;
wire n_814;
wire n_1864;
wire n_943;
wire n_2568;
wire n_3087;
wire n_2629;
wire n_1086;
wire n_1523;
wire n_2197;
wire n_1756;
wire n_2010;
wire n_2097;
wire n_2733;
wire n_2241;
wire n_1470;
wire n_2098;
wire n_2109;
wire n_1761;
wire n_2648;
wire n_2458;
wire n_1836;
wire n_2398;
wire n_3032;
wire n_3401;
wire n_1593;
wire n_986;
wire n_1420;
wire n_2651;
wire n_1750;
wire n_1775;
wire n_2833;
wire n_1699;
wire n_3179;
wire n_927;
wire n_1563;
wire n_2905;
wire n_3460;
wire n_803;
wire n_2570;
wire n_3123;
wire n_1875;
wire n_3379;
wire n_1615;
wire n_2184;
wire n_2418;
wire n_1087;
wire n_3390;
wire n_757;
wire n_1400;
wire n_712;
wire n_1539;
wire n_1806;
wire n_1599;
wire n_2842;
wire n_2711;
wire n_3070;
wire n_3477;
wire n_2635;
wire n_2469;
wire n_1575;
wire n_2209;
wire n_3074;
wire n_3020;
wire n_3142;
wire n_3164;
wire n_3475;
wire n_1448;
wire n_2077;
wire n_3136;
wire n_2520;
wire n_817;
wire n_2193;
wire n_2612;
wire n_3034;
wire n_2095;
wire n_3108;
wire n_2486;
wire n_2628;
wire n_2395;
wire n_951;
wire n_2521;
wire n_2908;
wire n_2053;
wire n_2752;
wire n_1580;
wire n_2124;
wire n_1574;
wire n_780;
wire n_2200;
wire n_1705;
wire n_2304;
wire n_1746;
wire n_726;
wire n_1439;
wire n_2263;
wire n_2212;
wire n_2716;
wire n_2352;
wire n_3495;
wire n_863;
wire n_2185;
wire n_3169;
wire n_1832;
wire n_1128;
wire n_2476;
wire n_2376;
wire n_2979;
wire n_3398;
wire n_1266;
wire n_1300;
wire n_2781;
wire n_3419;
wire n_807;
wire n_741;
wire n_2460;
wire n_2170;
wire n_1785;
wire n_1870;
wire n_2484;
wire n_2721;
wire n_1405;
wire n_2884;
wire n_3383;
wire n_3167;
wire n_997;
wire n_2308;
wire n_3459;
wire n_3238;
wire n_2986;
wire n_3498;
wire n_1428;
wire n_2691;
wire n_2243;
wire n_2400;
wire n_3092;
wire n_2903;
wire n_891;
wire n_3254;
wire n_2507;
wire n_2759;
wire n_3434;
wire n_1528;
wire n_1495;
wire n_3131;
wire n_2463;
wire n_2654;
wire n_717;
wire n_2975;
wire n_1357;
wire n_2503;
wire n_2478;
wire n_3178;
wire n_2794;
wire n_1512;
wire n_2496;
wire n_3378;
wire n_3481;
wire n_2974;
wire n_871;
wire n_2990;
wire n_2923;
wire n_1339;
wire n_1544;
wire n_1426;
wire n_2365;
wire n_3449;
wire n_3517;
wire n_3350;
wire n_2245;
wire n_1315;
wire n_1413;
wire n_2464;
wire n_811;
wire n_808;
wire n_945;
wire n_2925;
wire n_2270;
wire n_3260;
wire n_1706;
wire n_1560;
wire n_1592;
wire n_2776;
wire n_1461;
wire n_3166;
wire n_2695;
wire n_2630;
wire n_903;
wire n_1967;
wire n_2340;
wire n_3385;
wire n_2117;
wire n_1095;
wire n_1328;
wire n_1265;
wire n_2488;
wire n_1378;
wire n_2042;
wire n_3257;
wire n_1048;
wire n_774;
wire n_2459;
wire n_3137;
wire n_3116;
wire n_1925;
wire n_2439;
wire n_2106;
wire n_1430;
wire n_2414;
wire n_1251;
wire n_3090;
wire n_1247;
wire n_2450;
wire n_836;
wire n_1475;
wire n_3337;
wire n_2465;
wire n_1263;
wire n_3316;
wire n_1185;
wire n_1683;
wire n_1122;
wire n_2765;
wire n_3387;
wire n_890;
wire n_874;
wire n_1505;
wire n_3010;
wire n_2941;
wire n_1163;
wire n_1514;
wire n_964;
wire n_2728;
wire n_2948;
wire n_916;
wire n_3428;
wire n_2298;
wire n_2771;
wire n_3219;
wire n_2936;
wire n_895;
wire n_1035;
wire n_2427;
wire n_2045;
wire n_2985;
wire n_1535;
wire n_3158;
wire n_3106;
wire n_751;
wire n_2190;
wire n_1127;
wire n_932;
wire n_1972;
wire n_3080;
wire n_2772;
wire n_2778;
wire n_1004;
wire n_947;
wire n_831;
wire n_778;
wire n_1898;
wire n_1254;
wire n_1148;
wire n_1667;
wire n_1104;
wire n_1845;
wire n_1011;
wire n_2205;
wire n_2684;
wire n_2875;
wire n_2524;
wire n_3284;
wire n_1437;
wire n_2747;
wire n_3389;
wire n_1707;
wire n_1941;
wire n_2422;
wire n_2064;
wire n_3088;
wire n_1679;
wire n_2342;
wire n_2755;
wire n_2301;
wire n_1497;
wire n_2002;
wire n_2055;
wire n_2385;
wire n_3095;
wire n_3026;
wire n_2545;
wire n_1578;
wire n_3294;
wire n_2050;
wire n_1143;
wire n_1783;
wire n_2712;
wire n_3279;
wire n_2584;
wire n_972;
wire n_1815;
wire n_2500;
wire n_3344;
wire n_1917;
wire n_1444;
wire n_920;
wire n_2442;
wire n_1067;
wire n_3328;
wire n_2763;
wire n_2788;
wire n_994;
wire n_2000;
wire n_2089;
wire n_1857;
wire n_2761;
wire n_1920;
wire n_2696;
wire n_3252;
wire n_887;
wire n_1162;
wire n_1997;
wire n_2578;
wire n_2745;
wire n_1894;
wire n_2110;
wire n_2904;
wire n_3064;
wire n_2896;
wire n_2997;
wire n_3314;
wire n_1349;
wire n_1331;
wire n_1223;
wire n_991;
wire n_961;
wire n_2127;
wire n_1323;
wire n_1739;
wire n_3130;
wire n_1777;
wire n_3028;
wire n_3228;
wire n_1353;
wire n_3409;
wire n_2386;
wire n_3324;
wire n_1429;
wire n_3073;
wire n_2029;
wire n_3209;
wire n_2026;
wire n_1546;
wire n_3420;
wire n_1432;
wire n_2103;
wire n_3322;
wire n_1950;
wire n_1320;
wire n_996;
wire n_915;
wire n_2238;
wire n_2619;
wire n_3289;
wire n_1174;
wire n_1874;
wire n_1834;
wire n_3372;
wire n_3499;
wire n_3552;
wire n_2862;
wire n_3100;
wire n_3405;
wire n_1727;
wire n_3377;
wire n_1286;
wire n_1657;
wire n_1741;
wire n_1294;
wire n_1601;
wire n_900;
wire n_3414;
wire n_1351;
wire n_2933;
wire n_2138;
wire n_1380;
wire n_1367;
wire n_3336;
wire n_3240;
wire n_1291;
wire n_2895;
wire n_1914;
wire n_1458;
wire n_1694;
wire n_1460;
wire n_2041;
wire n_3201;
wire n_2271;
wire n_2356;
wire n_3339;
wire n_1830;
wire n_2261;
wire n_3016;
wire n_1629;
wire n_3476;
wire n_2994;
wire n_2011;
wire n_2620;
wire n_1826;
wire n_1855;
wire n_1662;
wire n_2105;
wire n_2187;
wire n_1340;
wire n_2694;
wire n_3443;
wire n_2562;
wire n_2642;
wire n_3029;
wire n_3269;
wire n_3447;
wire n_2647;
wire n_1626;
wire n_2223;
wire n_1660;
wire n_1850;
wire n_1643;
wire n_1670;
wire n_1789;
wire n_2415;
wire n_3152;
wire n_3154;
wire n_2344;
wire n_2317;
wire n_2556;
wire n_1112;
wire n_1267;
wire n_2384;
wire n_2683;
wire n_1384;
wire n_1376;
wire n_1537;
wire n_1858;
wire n_3432;
wire n_3523;
wire n_2815;
wire n_1816;
wire n_2446;
wire n_3388;
wire n_1612;
wire n_703;
wire n_2318;
wire n_1172;
wire n_2659;
wire n_1099;
wire n_2141;
wire n_3113;
wire n_2902;
wire n_2909;
wire n_1422;
wire n_1527;
wire n_3174;
wire n_3190;
wire n_1055;
wire n_1524;
wire n_798;
wire n_2849;
wire n_2947;
wire n_1754;
wire n_3048;
wire n_1177;
wire n_1025;
wire n_1991;
wire n_2566;
wire n_2679;
wire n_3292;
wire n_2210;
wire n_1517;
wire n_2502;
wire n_1225;
wire n_1962;
wire n_2346;
wire n_982;
wire n_1624;
wire n_785;
wire n_2180;
wire n_1952;
wire n_3376;
wire n_3002;
wire n_2087;
wire n_2920;
wire n_3290;
wire n_1598;
wire n_2952;
wire n_2617;
wire n_977;
wire n_2878;
wire n_1895;
wire n_2250;
wire n_719;
wire n_1491;
wire n_1860;
wire n_2831;
wire n_716;
wire n_1810;
wire n_1763;
wire n_923;
wire n_1607;
wire n_2865;
wire n_2075;
wire n_3047;
wire n_1625;
wire n_2959;
wire n_2610;
wire n_2420;
wire n_2380;
wire n_3335;
wire n_3265;
wire n_2240;
wire n_933;
wire n_2221;
wire n_1774;
wire n_1797;
wire n_2516;
wire n_2120;
wire n_1037;
wire n_2031;
wire n_1899;
wire n_3427;
wire n_1348;
wire n_1289;
wire n_838;
wire n_2892;
wire n_1021;
wire n_746;
wire n_1557;
wire n_1188;
wire n_1567;
wire n_2007;
wire n_742;
wire n_1191;
wire n_2004;
wire n_3356;
wire n_3431;
wire n_3220;
wire n_2024;
wire n_2086;
wire n_1503;
wire n_3422;
wire n_1052;
wire n_789;
wire n_1942;
wire n_3141;
wire n_2309;
wire n_842;
wire n_2274;
wire n_2698;
wire n_767;
wire n_1617;
wire n_1839;
wire n_1587;
wire n_2330;
wire n_2555;
wire n_2639;
wire n_1259;
wire n_2108;
wire n_3099;
wire n_2535;
wire n_1001;
wire n_2945;
wire n_3057;
wire n_2143;
wire n_2410;
wire n_1396;
wire n_2916;
wire n_1224;
wire n_1923;
wire n_3206;
wire n_2196;
wire n_2739;
wire n_2611;
wire n_1538;
wire n_2528;
wire n_2548;
wire n_3216;
wire n_2709;
wire n_3061;
wire n_2633;
wire n_1017;
wire n_2244;
wire n_730;
wire n_2604;
wire n_3424;
wire n_3462;
wire n_2351;
wire n_2437;
wire n_2049;
wire n_1456;
wire n_3245;
wire n_1889;
wire n_2113;
wire n_2665;
wire n_1124;
wire n_1690;
wire n_3063;
wire n_2688;
wire n_2881;
wire n_3302;
wire n_1673;
wire n_3361;
wire n_2018;
wire n_3134;
wire n_922;
wire n_2817;
wire n_1790;
wire n_993;
wire n_851;
wire n_3196;
wire n_2085;
wire n_3304;
wire n_2581;
wire n_1725;
wire n_2809;
wire n_2149;
wire n_2268;
wire n_2237;
wire n_2320;
wire n_1135;
wire n_2255;
wire n_2001;
wire n_1820;
wire n_1800;
wire n_3277;
wire n_3480;
wire n_2758;
wire n_1494;
wire n_1550;
wire n_2060;
wire n_1066;
wire n_2214;
wire n_3474;
wire n_1169;
wire n_1726;
wire n_1946;
wire n_3111;
wire n_1938;
wire n_830;
wire n_3452;
wire n_1241;
wire n_2589;
wire n_1072;
wire n_2194;
wire n_1231;
wire n_1173;
wire n_2736;
wire n_1208;
wire n_1639;
wire n_1604;
wire n_2735;
wire n_2845;
wire n_3506;
wire n_826;
wire n_1976;
wire n_2154;
wire n_2035;
wire n_1337;
wire n_2732;
wire n_3162;
wire n_2984;
wire n_1906;
wire n_3004;
wire n_1647;
wire n_1901;
wire n_3096;
wire n_3333;
wire n_839;
wire n_768;
wire n_3031;
wire n_1278;
wire n_2059;
wire n_796;
wire n_797;
wire n_3276;
wire n_1006;
wire n_2956;
wire n_1238;
wire n_1415;
wire n_976;
wire n_1710;
wire n_3021;
wire n_1063;
wire n_2153;
wire n_2452;
wire n_1270;
wire n_2891;
wire n_834;
wire n_2457;
wire n_2144;
wire n_1476;
wire n_935;
wire n_1603;
wire n_925;
wire n_2592;
wire n_1054;
wire n_2027;
wire n_3404;
wire n_2072;
wire n_2737;
wire n_2012;
wire n_722;
wire n_2251;
wire n_2963;
wire n_3512;
wire n_1644;
wire n_1406;
wire n_1489;
wire n_1880;
wire n_1993;
wire n_2137;
wire n_804;
wire n_1455;
wire n_1642;
wire n_1871;
wire n_2182;
wire n_2868;
wire n_3044;
wire n_2447;
wire n_3493;
wire n_2818;
wire n_3358;
wire n_3115;
wire n_1057;
wire n_1473;
wire n_3140;
wire n_3486;
wire n_2125;
wire n_2426;
wire n_2894;
wire n_1403;
wire n_2181;
wire n_3253;
wire n_2587;
wire n_1149;
wire n_1176;
wire n_1502;
wire n_1605;
wire n_868;
wire n_2099;
wire n_1202;
wire n_1065;
wire n_1897;
wire n_2477;
wire n_1457;
wire n_3172;
wire n_905;
wire n_2159;
wire n_3410;
wire n_975;
wire n_934;
wire n_775;
wire n_3273;
wire n_950;
wire n_2700;
wire n_1222;
wire n_3139;
wire n_1630;
wire n_3408;
wire n_2286;
wire n_3182;
wire n_1879;
wire n_1959;
wire n_2563;
wire n_1198;
wire n_2206;
wire n_1311;
wire n_3393;
wire n_1261;
wire n_2299;
wire n_3538;
wire n_2078;
wire n_3327;
wire n_2265;
wire n_776;
wire n_1114;
wire n_3513;
wire n_3011;
wire n_1167;
wire n_818;
wire n_3231;
wire n_2677;
wire n_2531;
wire n_2315;
wire n_3138;
wire n_2157;
wire n_3212;
wire n_1282;
wire n_2067;
wire n_2517;
wire n_1321;
wire n_1779;
wire n_3446;
wire n_3349;
wire n_2489;
wire n_1770;
wire n_1107;
wire n_3058;
wire n_3454;
wire n_1846;
wire n_2211;
wire n_1573;
wire n_2950;
wire n_815;
wire n_919;
wire n_2272;
wire n_1956;
wire n_2608;
wire n_3384;
wire n_2983;
wire n_1718;
wire n_2225;
wire n_3229;
wire n_2546;
wire n_1411;
wire n_2825;
wire n_1139;
wire n_1018;
wire n_858;
wire n_2345;
wire n_1324;
wire n_1669;
wire n_1501;
wire n_2742;
wire n_782;
wire n_1885;
wire n_1740;
wire n_1989;
wire n_3540;
wire n_1838;
wire n_833;
wire n_2680;
wire n_1343;
wire n_1801;
wire n_3439;
wire n_1371;
wire n_1513;
wire n_728;
wire n_3001;
wire n_2861;
wire n_2976;
wire n_2161;
wire n_2191;
wire n_2329;
wire n_1788;
wire n_2093;
wire n_2576;
wire n_786;
wire n_2348;
wire n_2417;
wire n_2675;
wire n_2043;
wire n_2366;
wire n_1621;
wire n_2338;
wire n_1919;
wire n_1342;
wire n_752;
wire n_2756;
wire n_2893;
wire n_2009;
wire n_2248;
wire n_958;
wire n_1175;
wire n_3500;
wire n_1416;
wire n_1659;
wire n_2850;
wire n_3465;
wire n_1221;
wire n_1047;
wire n_1878;
wire n_1515;
wire n_1374;
wire n_2851;
wire n_2438;
wire n_1435;
wire n_1688;
wire n_792;
wire n_2973;
wire n_1314;
wire n_1433;
wire n_2567;
wire n_3085;
wire n_3059;
wire n_1242;
wire n_1119;
wire n_2810;
wire n_2867;
wire n_2229;
wire n_1085;
wire n_3027;
wire n_2388;
wire n_2981;
wire n_3438;
wire n_2222;
wire n_3112;
wire n_1907;
wire n_3464;
wire n_885;
wire n_1530;
wire n_3215;
wire n_3413;
wire n_877;
wire n_2871;
wire n_2135;
wire n_1088;
wire n_896;
wire n_2764;
wire n_2624;
wire n_1813;
wire n_1451;
wire n_1005;
wire n_1102;
wire n_3234;
wire n_794;
wire n_2471;
wire n_1288;
wire n_1275;
wire n_985;
wire n_1165;
wire n_897;
wire n_1622;
wire n_2757;
wire n_2714;
wire n_3066;
wire n_2669;
wire n_2869;
wire n_1105;
wire n_1459;
wire n_912;
wire n_3121;
wire n_2232;
wire n_2898;
wire n_2455;
wire n_2121;
wire n_1893;
wire n_2519;
wire n_1570;
wire n_2231;
wire n_2874;
wire n_995;
wire n_2278;
wire n_1000;
wire n_2284;
wire n_1931;
wire n_2433;
wire n_2803;
wire n_2816;
wire n_3402;
wire n_1256;
wire n_2798;
wire n_3425;
wire n_1303;
wire n_1994;
wire n_1771;
wire n_3308;
wire n_1526;
wire n_764;
wire n_1507;
wire n_1206;
wire n_1809;
wire n_855;
wire n_2367;
wire n_812;
wire n_2658;
wire n_3236;
wire n_3491;
wire n_3109;
wire n_1961;
wire n_3271;
wire n_3013;
wire n_2553;
wire n_1050;
wire n_2218;
wire n_2667;
wire n_3062;
wire n_1769;
wire n_2130;
wire n_3256;
wire n_1060;
wire n_3126;
wire n_1372;
wire n_1847;
wire n_756;
wire n_1565;
wire n_1257;
wire n_2325;
wire n_2406;
wire n_1632;
wire n_2864;
wire n_3346;
wire n_3104;
wire n_3391;
wire n_1542;
wire n_946;
wire n_1547;
wire n_707;
wire n_1362;
wire n_1586;
wire n_3497;
wire n_1097;
wire n_3354;
wire n_3288;
wire n_3373;
wire n_3382;
wire n_3122;
wire n_2518;
wire n_2784;
wire n_3012;
wire n_3045;
wire n_1909;
wire n_2543;
wire n_3368;
wire n_2381;
wire n_2313;
wire n_956;
wire n_790;
wire n_2495;
wire n_2992;
wire n_1541;
wire n_2703;
wire n_1812;
wire n_3014;
wire n_1951;
wire n_1330;
wire n_1697;
wire n_2128;
wire n_2574;
wire n_1872;
wire n_1940;
wire n_2690;
wire n_1747;
wire n_1212;
wire n_1887;
wire n_1199;
wire n_3400;
wire n_2020;
wire n_3504;
wire n_1978;
wire n_2508;
wire n_3511;
wire n_2540;
wire n_1767;
wire n_1939;
wire n_2428;
wire n_3159;
wire n_1768;
wire n_1443;
wire n_2068;
wire n_2636;
wire n_2672;
wire n_3360;
wire n_1585;
wire n_1861;
wire n_2316;
wire n_3101;
wire n_1564;
wire n_1995;
wire n_1631;
wire n_2593;
wire n_1623;
wire n_2911;
wire n_861;
wire n_1828;
wire n_2364;
wire n_1389;
wire n_3303;
wire n_1131;
wire n_2641;
wire n_1798;
wire n_727;
wire n_1077;
wire n_3120;
wire n_1554;
wire n_3549;
wire n_1481;
wire n_1584;
wire n_2021;
wire n_1928;
wire n_2713;
wire n_828;
wire n_2938;
wire n_3227;
wire n_1438;
wire n_3342;
wire n_1973;
wire n_2314;
wire n_2939;
wire n_2156;
wire n_2494;
wire n_753;
wire n_2126;
wire n_1147;
wire n_747;
wire n_3403;
wire n_1363;
wire n_2228;
wire n_1691;
wire n_1098;
wire n_1366;
wire n_1518;
wire n_1187;
wire n_1361;
wire n_2034;
wire n_1693;
wire n_2790;
wire n_2872;
wire n_3102;
wire n_3173;
wire n_2411;
wire n_2081;
wire n_1892;
wire n_1061;
wire n_3539;
wire n_2266;
wire n_2993;
wire n_3433;
wire n_2061;
wire n_3018;
wire n_1373;
wire n_2449;
wire n_1686;
wire n_2131;
wire n_2526;
wire n_2830;
wire n_1302;
wire n_3017;
wire n_3083;
wire n_2083;
wire n_886;
wire n_2119;
wire n_1010;
wire n_883;
wire n_2207;
wire n_2044;
wire n_2542;
wire n_755;
wire n_2091;
wire n_2843;
wire n_3362;
wire n_3035;
wire n_3191;
wire n_1029;
wire n_3485;
wire n_2394;
wire n_3051;
wire n_770;
wire n_1572;
wire n_1635;
wire n_3305;
wire n_3149;
wire n_2827;
wire n_941;
wire n_1245;
wire n_1317;
wire n_2615;
wire n_3278;
wire n_3343;
wire n_2701;
wire n_2929;
wire n_3163;
wire n_2487;
wire n_1329;
wire n_2409;
wire n_2637;
wire n_2337;
wire n_854;
wire n_2405;
wire n_2601;
wire n_2513;
wire n_3118;
wire n_714;
wire n_1297;
wire n_1369;
wire n_1912;
wire n_3143;
wire n_1734;
wire n_3543;
wire n_1876;
wire n_2666;
wire n_3050;
wire n_2323;
wire n_3532;
wire n_740;
wire n_1811;
wire n_928;
wire n_898;
wire n_1285;
wire n_3042;
wire n_967;
wire n_2561;
wire n_736;
wire n_2913;
wire n_2491;
wire n_1529;
wire n_1381;
wire n_1824;
wire n_2254;
wire n_1597;
wire n_1161;
wire n_1103;
wire n_3522;
wire n_1486;
wire n_1068;
wire n_1833;
wire n_2914;
wire n_3551;
wire n_2371;
wire n_914;
wire n_3444;
wire n_1986;
wire n_3366;
wire n_2882;
wire n_1024;
wire n_3009;
wire n_1141;
wire n_3453;
wire n_3297;
wire n_3176;
wire n_1949;
wire n_1197;
wire n_2493;
wire n_2408;
wire n_2429;
wire n_3326;
wire n_1168;
wire n_865;
wire n_3000;
wire n_2115;
wire n_2013;
wire n_2140;
wire n_2134;
wire n_2483;
wire n_2305;
wire n_1556;
wire n_3423;
wire n_3547;
wire n_1192;
wire n_1646;
wire n_1290;
wire n_2514;
wire n_2466;
wire n_1759;
wire n_2048;
wire n_2760;
wire n_987;
wire n_750;
wire n_1299;
wire n_2942;
wire n_2096;
wire n_2129;
wire n_3230;
wire n_3545;
wire n_1101;
wire n_2532;
wire n_2079;
wire n_2296;
wire n_1720;
wire n_880;
wire n_2671;
wire n_1911;
wire n_2293;
wire n_3296;
wire n_731;
wire n_1336;
wire n_3068;
wire n_3071;
wire n_2734;
wire n_2870;
wire n_1166;
wire n_758;
wire n_720;
wire n_710;
wire n_1390;
wire n_2775;
wire n_1023;
wire n_1358;
wire n_813;
wire n_2310;
wire n_3223;
wire n_3318;
wire n_1211;
wire n_1397;
wire n_2674;
wire n_1284;
wire n_2005;
wire n_1359;
wire n_1116;
wire n_2811;
wire n_1758;
wire n_3226;
wire n_791;
wire n_1532;
wire n_2848;
wire n_1419;
wire n_2689;
wire n_1784;
wire n_1685;
wire n_1992;
wire n_1082;
wire n_3200;
wire n_3430;
wire n_1213;
wire n_2596;
wire n_2801;
wire n_1193;
wire n_1488;
wire n_849;
wire n_980;
wire n_2928;
wire n_3225;
wire n_2227;
wire n_2652;
wire n_3067;
wire n_1074;
wire n_3380;
wire n_3207;
wire n_759;
wire n_1379;
wire n_1721;
wire n_2972;
wire n_2627;
wire n_1827;
wire n_953;
wire n_1180;
wire n_1462;
wire n_3369;
wire n_3185;
wire n_2326;
wire n_1866;
wire n_1220;
wire n_1398;
wire n_2169;
wire n_2111;
wire n_1262;
wire n_1904;
wire n_2966;
wire n_3084;
wire n_3036;
wire n_1692;
wire n_2501;
wire n_2051;
wire n_1012;
wire n_1805;
wire n_960;
wire n_1022;
wire n_1760;
wire n_1240;
wire n_2173;
wire n_1183;
wire n_3285;
wire n_3160;
wire n_3483;
wire n_1204;
wire n_1151;
wire n_2824;
wire n_1814;
wire n_771;
wire n_3124;
wire n_999;
wire n_2634;
wire n_3286;
wire n_2982;
wire n_1092;
wire n_1808;
wire n_2768;
wire n_2668;
wire n_1658;
wire n_1386;
wire n_2588;
wire n_3015;
wire n_2931;
wire n_3321;
wire n_2492;
wire n_3081;
wire n_910;
wire n_2291;
wire n_3046;
wire n_844;
wire n_2172;
wire n_1728;
wire n_1020;
wire n_3076;
wire n_1142;
wire n_783;
wire n_1385;
wire n_2927;
wire n_1062;
wire n_1230;
wire n_1027;
wire n_1516;
wire n_2533;
wire n_1499;
wire n_1500;
wire n_2155;
wire n_2706;
wire n_1868;
wire n_966;
wire n_2148;
wire n_2104;
wire n_949;
wire n_704;
wire n_2303;
wire n_2618;
wire n_2653;
wire n_2855;
wire n_2357;
wire n_924;
wire n_2937;
wire n_3359;
wire n_3114;
wire n_2331;
wire n_3332;
wire n_1600;
wire n_1661;
wire n_2967;
wire n_1965;
wire n_3005;
wire n_1757;
wire n_2136;
wire n_2403;
wire n_918;
wire n_3053;
wire n_2056;
wire n_1913;
wire n_2702;
wire n_2054;
wire n_1039;
wire n_2226;
wire n_2407;
wire n_2791;
wire n_1043;
wire n_1402;
wire n_2267;
wire n_735;
wire n_1450;
wire n_2082;
wire n_2302;
wire n_2453;
wire n_2560;
wire n_3056;
wire n_3267;
wire n_2092;
wire n_3008;
wire n_1472;
wire n_1365;
wire n_2443;
wire n_3189;
wire n_3052;
wire n_2802;
wire n_2797;
wire n_2279;
wire n_1089;
wire n_1536;
wire n_1049;
wire n_1719;
wire n_2066;
wire n_1158;
wire n_1974;
wire n_2988;
wire n_763;
wire n_1882;
wire n_2770;
wire n_2961;
wire n_2704;
wire n_2996;
wire n_1915;
wire n_2836;
wire n_940;
wire n_1762;
wire n_2534;
wire n_1404;
wire n_788;
wire n_3283;
wire n_1736;
wire n_3421;
wire n_2907;
wire n_3311;
wire n_1160;
wire n_1442;
wire n_1948;
wire n_2168;
wire n_1216;
wire n_2681;
wire n_1891;
wire n_1026;
wire n_3247;
wire n_2886;
wire n_1454;
wire n_1033;
wire n_990;
wire n_1383;
wire n_1968;
wire n_2057;
wire n_2609;
wire n_2378;
wire n_888;
wire n_2749;
wire n_1325;
wire n_3133;
wire n_2754;
wire n_3527;
wire n_2014;
wire n_3041;
wire n_1483;
wire n_1703;
wire n_1205;
wire n_1822;
wire n_843;
wire n_1953;
wire n_1059;
wire n_2969;
wire n_799;
wire n_2692;
wire n_3261;
wire n_3550;
wire n_1804;
wire n_1581;
wire n_3287;
wire n_3534;
wire n_1837;
wire n_3325;
wire n_1744;
wire n_1975;
wire n_3437;
wire n_1414;
wire n_2324;
wire n_2246;
wire n_2738;
wire n_3161;
wire n_1002;
wire n_1851;
wire n_1755;
wire n_2195;
wire n_2940;
wire n_1111;
wire n_1819;
wire n_3313;
wire n_1341;
wire n_1807;
wire n_2670;
wire n_2645;
wire n_2202;
wire n_1310;
wire n_3275;
wire n_1745;
wire n_1714;
wire n_3198;
wire n_3463;
wire n_1958;
wire n_1611;
wire n_2559;
wire n_3516;
wire n_2262;
wire n_955;
wire n_1333;
wire n_1916;
wire n_2726;
wire n_2917;
wire n_2073;
wire n_952;
wire n_1675;
wire n_1947;
wire n_2165;
wire n_1640;
wire n_2016;
wire n_3157;
wire n_1551;
wire n_1145;
wire n_1533;
wire n_2307;
wire n_2515;
wire n_3546;
wire n_1511;
wire n_1791;
wire n_1113;
wire n_3089;
wire n_1651;
wire n_1966;
wire n_2058;
wire n_2678;
wire n_3406;
wire n_1468;
wire n_3442;
wire n_2327;
wire n_2656;
wire n_913;
wire n_2353;
wire n_1164;
wire n_2258;
wire n_1732;
wire n_2167;
wire n_3079;
wire n_1354;
wire n_3329;
wire n_2039;
wire n_1277;
wire n_1696;
wire n_1016;
wire n_3233;
wire n_1355;
wire n_809;
wire n_2544;
wire n_856;
wire n_779;
wire n_3193;
wire n_3501;
wire n_866;
wire n_2538;
wire n_3270;
wire n_2582;
wire n_1559;
wire n_2321;
wire n_2915;
wire n_1579;
wire n_1280;
wire n_2854;
wire n_2932;
wire n_3258;
wire n_1335;
wire n_3266;
wire n_2285;
wire n_3213;
wire n_1934;
wire n_2040;
wire n_1900;
wire n_2174;
wire n_3246;
wire n_1843;
wire n_2186;
wire n_2510;
wire n_2030;
wire n_2614;
wire n_3418;
wire n_2435;
wire n_1665;
wire n_2583;
wire n_3417;
wire n_1091;
wire n_1678;
wire n_1780;
wire n_2725;
wire n_1287;
wire n_2769;
wire n_1482;
wire n_860;
wire n_1525;
wire n_848;
wire n_3244;
wire n_3195;
wire n_2100;
wire n_2349;
wire n_1902;
wire n_2536;
wire n_2474;
wire n_1194;
wire n_1150;
wire n_1399;
wire n_1903;
wire n_1674;
wire n_1849;
wire n_867;
wire n_983;
wire n_1417;
wire n_3482;
wire n_2282;
wire n_970;
wire n_2430;
wire n_2676;
wire n_921;
wire n_2673;
wire n_3515;
wire n_3489;
wire n_2926;
wire n_1534;
wire n_2912;
wire n_3181;
wire n_908;
wire n_3536;
wire n_1346;
wire n_2834;
wire n_3268;
wire n_1123;
wire n_2710;
wire n_1272;
wire n_2497;
wire n_1393;
wire n_2970;
wire n_984;
wire n_1655;
wire n_3040;
wire n_3494;
wire n_2978;
wire n_1410;
wire n_988;
wire n_2368;
wire n_3363;
wire n_760;
wire n_3528;
wire n_1157;
wire n_3502;
wire n_806;
wire n_2657;
wire n_1186;
wire n_2065;
wire n_3180;
wire n_2901;
wire n_1743;
wire n_2743;
wire n_1854;
wire n_1506;

CKINVDCx5p33_ASAP7_75t_R g703 ( 
.A(n_455),
.Y(n_703)
);

CKINVDCx5p33_ASAP7_75t_R g704 ( 
.A(n_221),
.Y(n_704)
);

CKINVDCx16_ASAP7_75t_R g705 ( 
.A(n_59),
.Y(n_705)
);

CKINVDCx20_ASAP7_75t_R g706 ( 
.A(n_398),
.Y(n_706)
);

INVx1_ASAP7_75t_L g707 ( 
.A(n_562),
.Y(n_707)
);

BUFx5_ASAP7_75t_L g708 ( 
.A(n_291),
.Y(n_708)
);

CKINVDCx5p33_ASAP7_75t_R g709 ( 
.A(n_62),
.Y(n_709)
);

INVx1_ASAP7_75t_L g710 ( 
.A(n_376),
.Y(n_710)
);

CKINVDCx5p33_ASAP7_75t_R g711 ( 
.A(n_181),
.Y(n_711)
);

BUFx10_ASAP7_75t_L g712 ( 
.A(n_506),
.Y(n_712)
);

INVx1_ASAP7_75t_SL g713 ( 
.A(n_99),
.Y(n_713)
);

CKINVDCx5p33_ASAP7_75t_R g714 ( 
.A(n_244),
.Y(n_714)
);

CKINVDCx5p33_ASAP7_75t_R g715 ( 
.A(n_517),
.Y(n_715)
);

CKINVDCx5p33_ASAP7_75t_R g716 ( 
.A(n_393),
.Y(n_716)
);

INVx2_ASAP7_75t_SL g717 ( 
.A(n_75),
.Y(n_717)
);

INVx1_ASAP7_75t_L g718 ( 
.A(n_468),
.Y(n_718)
);

CKINVDCx5p33_ASAP7_75t_R g719 ( 
.A(n_383),
.Y(n_719)
);

INVx1_ASAP7_75t_L g720 ( 
.A(n_196),
.Y(n_720)
);

CKINVDCx20_ASAP7_75t_R g721 ( 
.A(n_135),
.Y(n_721)
);

CKINVDCx5p33_ASAP7_75t_R g722 ( 
.A(n_674),
.Y(n_722)
);

CKINVDCx5p33_ASAP7_75t_R g723 ( 
.A(n_30),
.Y(n_723)
);

OR2x2_ASAP7_75t_L g724 ( 
.A(n_561),
.B(n_50),
.Y(n_724)
);

INVx1_ASAP7_75t_L g725 ( 
.A(n_641),
.Y(n_725)
);

CKINVDCx5p33_ASAP7_75t_R g726 ( 
.A(n_680),
.Y(n_726)
);

INVx1_ASAP7_75t_L g727 ( 
.A(n_373),
.Y(n_727)
);

CKINVDCx5p33_ASAP7_75t_R g728 ( 
.A(n_628),
.Y(n_728)
);

CKINVDCx20_ASAP7_75t_R g729 ( 
.A(n_229),
.Y(n_729)
);

INVx1_ASAP7_75t_L g730 ( 
.A(n_266),
.Y(n_730)
);

INVx1_ASAP7_75t_L g731 ( 
.A(n_175),
.Y(n_731)
);

CKINVDCx5p33_ASAP7_75t_R g732 ( 
.A(n_195),
.Y(n_732)
);

INVx1_ASAP7_75t_L g733 ( 
.A(n_477),
.Y(n_733)
);

BUFx2_ASAP7_75t_L g734 ( 
.A(n_89),
.Y(n_734)
);

CKINVDCx5p33_ASAP7_75t_R g735 ( 
.A(n_274),
.Y(n_735)
);

INVx1_ASAP7_75t_L g736 ( 
.A(n_697),
.Y(n_736)
);

INVx1_ASAP7_75t_L g737 ( 
.A(n_297),
.Y(n_737)
);

CKINVDCx5p33_ASAP7_75t_R g738 ( 
.A(n_468),
.Y(n_738)
);

XOR2xp5_ASAP7_75t_L g739 ( 
.A(n_505),
.B(n_209),
.Y(n_739)
);

CKINVDCx5p33_ASAP7_75t_R g740 ( 
.A(n_363),
.Y(n_740)
);

CKINVDCx5p33_ASAP7_75t_R g741 ( 
.A(n_77),
.Y(n_741)
);

CKINVDCx5p33_ASAP7_75t_R g742 ( 
.A(n_669),
.Y(n_742)
);

INVx2_ASAP7_75t_L g743 ( 
.A(n_259),
.Y(n_743)
);

CKINVDCx5p33_ASAP7_75t_R g744 ( 
.A(n_498),
.Y(n_744)
);

CKINVDCx5p33_ASAP7_75t_R g745 ( 
.A(n_369),
.Y(n_745)
);

INVx1_ASAP7_75t_L g746 ( 
.A(n_251),
.Y(n_746)
);

CKINVDCx5p33_ASAP7_75t_R g747 ( 
.A(n_682),
.Y(n_747)
);

CKINVDCx20_ASAP7_75t_R g748 ( 
.A(n_438),
.Y(n_748)
);

NOR2xp67_ASAP7_75t_L g749 ( 
.A(n_260),
.B(n_596),
.Y(n_749)
);

CKINVDCx20_ASAP7_75t_R g750 ( 
.A(n_387),
.Y(n_750)
);

INVx1_ASAP7_75t_L g751 ( 
.A(n_224),
.Y(n_751)
);

CKINVDCx5p33_ASAP7_75t_R g752 ( 
.A(n_160),
.Y(n_752)
);

CKINVDCx5p33_ASAP7_75t_R g753 ( 
.A(n_558),
.Y(n_753)
);

INVx1_ASAP7_75t_L g754 ( 
.A(n_65),
.Y(n_754)
);

CKINVDCx16_ASAP7_75t_R g755 ( 
.A(n_13),
.Y(n_755)
);

OR2x2_ASAP7_75t_L g756 ( 
.A(n_661),
.B(n_53),
.Y(n_756)
);

CKINVDCx5p33_ASAP7_75t_R g757 ( 
.A(n_378),
.Y(n_757)
);

CKINVDCx5p33_ASAP7_75t_R g758 ( 
.A(n_307),
.Y(n_758)
);

CKINVDCx14_ASAP7_75t_R g759 ( 
.A(n_491),
.Y(n_759)
);

BUFx10_ASAP7_75t_L g760 ( 
.A(n_177),
.Y(n_760)
);

CKINVDCx5p33_ASAP7_75t_R g761 ( 
.A(n_164),
.Y(n_761)
);

INVxp67_ASAP7_75t_L g762 ( 
.A(n_593),
.Y(n_762)
);

CKINVDCx5p33_ASAP7_75t_R g763 ( 
.A(n_85),
.Y(n_763)
);

CKINVDCx5p33_ASAP7_75t_R g764 ( 
.A(n_259),
.Y(n_764)
);

NOR2xp67_ASAP7_75t_L g765 ( 
.A(n_276),
.B(n_19),
.Y(n_765)
);

BUFx6f_ASAP7_75t_L g766 ( 
.A(n_5),
.Y(n_766)
);

INVx2_ASAP7_75t_L g767 ( 
.A(n_638),
.Y(n_767)
);

INVxp67_ASAP7_75t_L g768 ( 
.A(n_325),
.Y(n_768)
);

CKINVDCx5p33_ASAP7_75t_R g769 ( 
.A(n_19),
.Y(n_769)
);

INVx2_ASAP7_75t_L g770 ( 
.A(n_544),
.Y(n_770)
);

INVx1_ASAP7_75t_L g771 ( 
.A(n_360),
.Y(n_771)
);

CKINVDCx5p33_ASAP7_75t_R g772 ( 
.A(n_535),
.Y(n_772)
);

INVx1_ASAP7_75t_L g773 ( 
.A(n_687),
.Y(n_773)
);

INVx1_ASAP7_75t_L g774 ( 
.A(n_9),
.Y(n_774)
);

INVx2_ASAP7_75t_L g775 ( 
.A(n_673),
.Y(n_775)
);

INVx1_ASAP7_75t_L g776 ( 
.A(n_679),
.Y(n_776)
);

CKINVDCx5p33_ASAP7_75t_R g777 ( 
.A(n_388),
.Y(n_777)
);

CKINVDCx5p33_ASAP7_75t_R g778 ( 
.A(n_288),
.Y(n_778)
);

CKINVDCx5p33_ASAP7_75t_R g779 ( 
.A(n_228),
.Y(n_779)
);

BUFx6f_ASAP7_75t_L g780 ( 
.A(n_453),
.Y(n_780)
);

INVx1_ASAP7_75t_L g781 ( 
.A(n_675),
.Y(n_781)
);

INVxp67_ASAP7_75t_SL g782 ( 
.A(n_632),
.Y(n_782)
);

CKINVDCx5p33_ASAP7_75t_R g783 ( 
.A(n_522),
.Y(n_783)
);

CKINVDCx5p33_ASAP7_75t_R g784 ( 
.A(n_297),
.Y(n_784)
);

INVx2_ASAP7_75t_L g785 ( 
.A(n_61),
.Y(n_785)
);

CKINVDCx20_ASAP7_75t_R g786 ( 
.A(n_542),
.Y(n_786)
);

INVx1_ASAP7_75t_L g787 ( 
.A(n_179),
.Y(n_787)
);

CKINVDCx5p33_ASAP7_75t_R g788 ( 
.A(n_179),
.Y(n_788)
);

INVx1_ASAP7_75t_L g789 ( 
.A(n_560),
.Y(n_789)
);

INVx2_ASAP7_75t_L g790 ( 
.A(n_20),
.Y(n_790)
);

CKINVDCx5p33_ASAP7_75t_R g791 ( 
.A(n_168),
.Y(n_791)
);

INVx1_ASAP7_75t_L g792 ( 
.A(n_659),
.Y(n_792)
);

CKINVDCx5p33_ASAP7_75t_R g793 ( 
.A(n_548),
.Y(n_793)
);

INVx1_ASAP7_75t_L g794 ( 
.A(n_371),
.Y(n_794)
);

CKINVDCx5p33_ASAP7_75t_R g795 ( 
.A(n_202),
.Y(n_795)
);

CKINVDCx5p33_ASAP7_75t_R g796 ( 
.A(n_152),
.Y(n_796)
);

BUFx10_ASAP7_75t_L g797 ( 
.A(n_549),
.Y(n_797)
);

CKINVDCx20_ASAP7_75t_R g798 ( 
.A(n_15),
.Y(n_798)
);

BUFx3_ASAP7_75t_L g799 ( 
.A(n_263),
.Y(n_799)
);

HB1xp67_ASAP7_75t_L g800 ( 
.A(n_632),
.Y(n_800)
);

INVx1_ASAP7_75t_L g801 ( 
.A(n_558),
.Y(n_801)
);

CKINVDCx5p33_ASAP7_75t_R g802 ( 
.A(n_99),
.Y(n_802)
);

CKINVDCx20_ASAP7_75t_R g803 ( 
.A(n_402),
.Y(n_803)
);

CKINVDCx5p33_ASAP7_75t_R g804 ( 
.A(n_275),
.Y(n_804)
);

CKINVDCx5p33_ASAP7_75t_R g805 ( 
.A(n_548),
.Y(n_805)
);

INVx1_ASAP7_75t_L g806 ( 
.A(n_488),
.Y(n_806)
);

INVx1_ASAP7_75t_L g807 ( 
.A(n_690),
.Y(n_807)
);

CKINVDCx5p33_ASAP7_75t_R g808 ( 
.A(n_613),
.Y(n_808)
);

INVx1_ASAP7_75t_L g809 ( 
.A(n_136),
.Y(n_809)
);

BUFx10_ASAP7_75t_L g810 ( 
.A(n_435),
.Y(n_810)
);

INVx1_ASAP7_75t_L g811 ( 
.A(n_51),
.Y(n_811)
);

BUFx2_ASAP7_75t_L g812 ( 
.A(n_540),
.Y(n_812)
);

CKINVDCx5p33_ASAP7_75t_R g813 ( 
.A(n_272),
.Y(n_813)
);

CKINVDCx5p33_ASAP7_75t_R g814 ( 
.A(n_317),
.Y(n_814)
);

CKINVDCx5p33_ASAP7_75t_R g815 ( 
.A(n_702),
.Y(n_815)
);

CKINVDCx20_ASAP7_75t_R g816 ( 
.A(n_157),
.Y(n_816)
);

BUFx2_ASAP7_75t_L g817 ( 
.A(n_177),
.Y(n_817)
);

INVx1_ASAP7_75t_L g818 ( 
.A(n_46),
.Y(n_818)
);

CKINVDCx5p33_ASAP7_75t_R g819 ( 
.A(n_89),
.Y(n_819)
);

INVx2_ASAP7_75t_SL g820 ( 
.A(n_492),
.Y(n_820)
);

INVx1_ASAP7_75t_L g821 ( 
.A(n_688),
.Y(n_821)
);

CKINVDCx5p33_ASAP7_75t_R g822 ( 
.A(n_149),
.Y(n_822)
);

CKINVDCx5p33_ASAP7_75t_R g823 ( 
.A(n_403),
.Y(n_823)
);

HB1xp67_ASAP7_75t_L g824 ( 
.A(n_153),
.Y(n_824)
);

INVx1_ASAP7_75t_L g825 ( 
.A(n_308),
.Y(n_825)
);

INVx1_ASAP7_75t_L g826 ( 
.A(n_511),
.Y(n_826)
);

CKINVDCx5p33_ASAP7_75t_R g827 ( 
.A(n_544),
.Y(n_827)
);

INVx1_ASAP7_75t_L g828 ( 
.A(n_75),
.Y(n_828)
);

CKINVDCx5p33_ASAP7_75t_R g829 ( 
.A(n_228),
.Y(n_829)
);

CKINVDCx20_ASAP7_75t_R g830 ( 
.A(n_154),
.Y(n_830)
);

CKINVDCx5p33_ASAP7_75t_R g831 ( 
.A(n_656),
.Y(n_831)
);

CKINVDCx16_ASAP7_75t_R g832 ( 
.A(n_651),
.Y(n_832)
);

CKINVDCx5p33_ASAP7_75t_R g833 ( 
.A(n_474),
.Y(n_833)
);

INVx1_ASAP7_75t_L g834 ( 
.A(n_169),
.Y(n_834)
);

INVx1_ASAP7_75t_L g835 ( 
.A(n_541),
.Y(n_835)
);

INVx1_ASAP7_75t_L g836 ( 
.A(n_106),
.Y(n_836)
);

INVx1_ASAP7_75t_L g837 ( 
.A(n_644),
.Y(n_837)
);

CKINVDCx5p33_ASAP7_75t_R g838 ( 
.A(n_464),
.Y(n_838)
);

HB1xp67_ASAP7_75t_L g839 ( 
.A(n_154),
.Y(n_839)
);

CKINVDCx5p33_ASAP7_75t_R g840 ( 
.A(n_278),
.Y(n_840)
);

INVx1_ASAP7_75t_L g841 ( 
.A(n_592),
.Y(n_841)
);

CKINVDCx5p33_ASAP7_75t_R g842 ( 
.A(n_234),
.Y(n_842)
);

CKINVDCx5p33_ASAP7_75t_R g843 ( 
.A(n_232),
.Y(n_843)
);

INVx1_ASAP7_75t_L g844 ( 
.A(n_458),
.Y(n_844)
);

INVx1_ASAP7_75t_L g845 ( 
.A(n_650),
.Y(n_845)
);

INVxp67_ASAP7_75t_L g846 ( 
.A(n_88),
.Y(n_846)
);

NOR2xp67_ASAP7_75t_L g847 ( 
.A(n_655),
.B(n_596),
.Y(n_847)
);

INVx1_ASAP7_75t_L g848 ( 
.A(n_72),
.Y(n_848)
);

INVx2_ASAP7_75t_L g849 ( 
.A(n_444),
.Y(n_849)
);

INVx1_ASAP7_75t_L g850 ( 
.A(n_590),
.Y(n_850)
);

INVx1_ASAP7_75t_L g851 ( 
.A(n_233),
.Y(n_851)
);

INVx1_ASAP7_75t_L g852 ( 
.A(n_140),
.Y(n_852)
);

CKINVDCx5p33_ASAP7_75t_R g853 ( 
.A(n_598),
.Y(n_853)
);

CKINVDCx5p33_ASAP7_75t_R g854 ( 
.A(n_264),
.Y(n_854)
);

CKINVDCx5p33_ASAP7_75t_R g855 ( 
.A(n_115),
.Y(n_855)
);

INVx1_ASAP7_75t_L g856 ( 
.A(n_111),
.Y(n_856)
);

CKINVDCx5p33_ASAP7_75t_R g857 ( 
.A(n_97),
.Y(n_857)
);

CKINVDCx5p33_ASAP7_75t_R g858 ( 
.A(n_584),
.Y(n_858)
);

CKINVDCx5p33_ASAP7_75t_R g859 ( 
.A(n_541),
.Y(n_859)
);

CKINVDCx5p33_ASAP7_75t_R g860 ( 
.A(n_590),
.Y(n_860)
);

INVx1_ASAP7_75t_SL g861 ( 
.A(n_580),
.Y(n_861)
);

INVx2_ASAP7_75t_L g862 ( 
.A(n_66),
.Y(n_862)
);

INVx1_ASAP7_75t_L g863 ( 
.A(n_274),
.Y(n_863)
);

CKINVDCx5p33_ASAP7_75t_R g864 ( 
.A(n_595),
.Y(n_864)
);

INVx1_ASAP7_75t_L g865 ( 
.A(n_398),
.Y(n_865)
);

INVx1_ASAP7_75t_L g866 ( 
.A(n_275),
.Y(n_866)
);

BUFx10_ASAP7_75t_L g867 ( 
.A(n_353),
.Y(n_867)
);

CKINVDCx5p33_ASAP7_75t_R g868 ( 
.A(n_249),
.Y(n_868)
);

CKINVDCx5p33_ASAP7_75t_R g869 ( 
.A(n_59),
.Y(n_869)
);

INVx2_ASAP7_75t_L g870 ( 
.A(n_560),
.Y(n_870)
);

CKINVDCx20_ASAP7_75t_R g871 ( 
.A(n_328),
.Y(n_871)
);

INVx1_ASAP7_75t_L g872 ( 
.A(n_306),
.Y(n_872)
);

CKINVDCx16_ASAP7_75t_R g873 ( 
.A(n_420),
.Y(n_873)
);

INVx2_ASAP7_75t_L g874 ( 
.A(n_686),
.Y(n_874)
);

INVx2_ASAP7_75t_SL g875 ( 
.A(n_203),
.Y(n_875)
);

INVx1_ASAP7_75t_L g876 ( 
.A(n_294),
.Y(n_876)
);

BUFx3_ASAP7_75t_L g877 ( 
.A(n_657),
.Y(n_877)
);

INVx1_ASAP7_75t_L g878 ( 
.A(n_162),
.Y(n_878)
);

INVx1_ASAP7_75t_L g879 ( 
.A(n_445),
.Y(n_879)
);

INVx1_ASAP7_75t_L g880 ( 
.A(n_492),
.Y(n_880)
);

BUFx2_ASAP7_75t_L g881 ( 
.A(n_660),
.Y(n_881)
);

INVx1_ASAP7_75t_L g882 ( 
.A(n_639),
.Y(n_882)
);

BUFx6f_ASAP7_75t_L g883 ( 
.A(n_633),
.Y(n_883)
);

INVx1_ASAP7_75t_L g884 ( 
.A(n_430),
.Y(n_884)
);

CKINVDCx5p33_ASAP7_75t_R g885 ( 
.A(n_136),
.Y(n_885)
);

INVx2_ASAP7_75t_L g886 ( 
.A(n_699),
.Y(n_886)
);

BUFx3_ASAP7_75t_L g887 ( 
.A(n_300),
.Y(n_887)
);

CKINVDCx5p33_ASAP7_75t_R g888 ( 
.A(n_670),
.Y(n_888)
);

INVx2_ASAP7_75t_L g889 ( 
.A(n_507),
.Y(n_889)
);

CKINVDCx20_ASAP7_75t_R g890 ( 
.A(n_479),
.Y(n_890)
);

INVx1_ASAP7_75t_L g891 ( 
.A(n_148),
.Y(n_891)
);

CKINVDCx5p33_ASAP7_75t_R g892 ( 
.A(n_5),
.Y(n_892)
);

CKINVDCx5p33_ASAP7_75t_R g893 ( 
.A(n_214),
.Y(n_893)
);

CKINVDCx5p33_ASAP7_75t_R g894 ( 
.A(n_533),
.Y(n_894)
);

INVx1_ASAP7_75t_L g895 ( 
.A(n_112),
.Y(n_895)
);

INVx2_ASAP7_75t_L g896 ( 
.A(n_35),
.Y(n_896)
);

INVxp33_ASAP7_75t_L g897 ( 
.A(n_138),
.Y(n_897)
);

CKINVDCx5p33_ASAP7_75t_R g898 ( 
.A(n_531),
.Y(n_898)
);

CKINVDCx5p33_ASAP7_75t_R g899 ( 
.A(n_524),
.Y(n_899)
);

CKINVDCx20_ASAP7_75t_R g900 ( 
.A(n_380),
.Y(n_900)
);

CKINVDCx5p33_ASAP7_75t_R g901 ( 
.A(n_68),
.Y(n_901)
);

INVx2_ASAP7_75t_SL g902 ( 
.A(n_369),
.Y(n_902)
);

INVx2_ASAP7_75t_L g903 ( 
.A(n_423),
.Y(n_903)
);

INVx1_ASAP7_75t_L g904 ( 
.A(n_586),
.Y(n_904)
);

INVx1_ASAP7_75t_L g905 ( 
.A(n_355),
.Y(n_905)
);

INVx1_ASAP7_75t_L g906 ( 
.A(n_441),
.Y(n_906)
);

HB1xp67_ASAP7_75t_L g907 ( 
.A(n_471),
.Y(n_907)
);

CKINVDCx5p33_ASAP7_75t_R g908 ( 
.A(n_583),
.Y(n_908)
);

INVx1_ASAP7_75t_L g909 ( 
.A(n_476),
.Y(n_909)
);

INVx2_ASAP7_75t_L g910 ( 
.A(n_240),
.Y(n_910)
);

BUFx3_ASAP7_75t_L g911 ( 
.A(n_312),
.Y(n_911)
);

CKINVDCx16_ASAP7_75t_R g912 ( 
.A(n_183),
.Y(n_912)
);

CKINVDCx5p33_ASAP7_75t_R g913 ( 
.A(n_108),
.Y(n_913)
);

INVx1_ASAP7_75t_L g914 ( 
.A(n_342),
.Y(n_914)
);

BUFx3_ASAP7_75t_L g915 ( 
.A(n_158),
.Y(n_915)
);

CKINVDCx5p33_ASAP7_75t_R g916 ( 
.A(n_479),
.Y(n_916)
);

INVx1_ASAP7_75t_L g917 ( 
.A(n_2),
.Y(n_917)
);

CKINVDCx20_ASAP7_75t_R g918 ( 
.A(n_701),
.Y(n_918)
);

CKINVDCx5p33_ASAP7_75t_R g919 ( 
.A(n_106),
.Y(n_919)
);

CKINVDCx20_ASAP7_75t_R g920 ( 
.A(n_51),
.Y(n_920)
);

CKINVDCx5p33_ASAP7_75t_R g921 ( 
.A(n_477),
.Y(n_921)
);

INVx1_ASAP7_75t_L g922 ( 
.A(n_667),
.Y(n_922)
);

INVx1_ASAP7_75t_L g923 ( 
.A(n_425),
.Y(n_923)
);

INVx1_ASAP7_75t_L g924 ( 
.A(n_138),
.Y(n_924)
);

INVx1_ASAP7_75t_L g925 ( 
.A(n_242),
.Y(n_925)
);

CKINVDCx20_ASAP7_75t_R g926 ( 
.A(n_599),
.Y(n_926)
);

INVx1_ASAP7_75t_L g927 ( 
.A(n_35),
.Y(n_927)
);

BUFx3_ASAP7_75t_L g928 ( 
.A(n_629),
.Y(n_928)
);

INVx1_ASAP7_75t_SL g929 ( 
.A(n_283),
.Y(n_929)
);

CKINVDCx5p33_ASAP7_75t_R g930 ( 
.A(n_258),
.Y(n_930)
);

CKINVDCx5p33_ASAP7_75t_R g931 ( 
.A(n_296),
.Y(n_931)
);

INVx1_ASAP7_75t_L g932 ( 
.A(n_295),
.Y(n_932)
);

INVx1_ASAP7_75t_L g933 ( 
.A(n_407),
.Y(n_933)
);

CKINVDCx5p33_ASAP7_75t_R g934 ( 
.A(n_366),
.Y(n_934)
);

INVx2_ASAP7_75t_SL g935 ( 
.A(n_426),
.Y(n_935)
);

INVx1_ASAP7_75t_L g936 ( 
.A(n_312),
.Y(n_936)
);

CKINVDCx5p33_ASAP7_75t_R g937 ( 
.A(n_329),
.Y(n_937)
);

BUFx3_ASAP7_75t_L g938 ( 
.A(n_505),
.Y(n_938)
);

CKINVDCx5p33_ASAP7_75t_R g939 ( 
.A(n_132),
.Y(n_939)
);

INVx1_ASAP7_75t_L g940 ( 
.A(n_634),
.Y(n_940)
);

INVx1_ASAP7_75t_L g941 ( 
.A(n_264),
.Y(n_941)
);

CKINVDCx5p33_ASAP7_75t_R g942 ( 
.A(n_581),
.Y(n_942)
);

INVx1_ASAP7_75t_L g943 ( 
.A(n_629),
.Y(n_943)
);

INVx1_ASAP7_75t_L g944 ( 
.A(n_48),
.Y(n_944)
);

CKINVDCx5p33_ASAP7_75t_R g945 ( 
.A(n_530),
.Y(n_945)
);

CKINVDCx12_ASAP7_75t_R g946 ( 
.A(n_636),
.Y(n_946)
);

INVxp67_ASAP7_75t_L g947 ( 
.A(n_627),
.Y(n_947)
);

INVx1_ASAP7_75t_L g948 ( 
.A(n_619),
.Y(n_948)
);

CKINVDCx5p33_ASAP7_75t_R g949 ( 
.A(n_283),
.Y(n_949)
);

CKINVDCx5p33_ASAP7_75t_R g950 ( 
.A(n_526),
.Y(n_950)
);

CKINVDCx5p33_ASAP7_75t_R g951 ( 
.A(n_422),
.Y(n_951)
);

CKINVDCx5p33_ASAP7_75t_R g952 ( 
.A(n_192),
.Y(n_952)
);

CKINVDCx5p33_ASAP7_75t_R g953 ( 
.A(n_132),
.Y(n_953)
);

INVx1_ASAP7_75t_L g954 ( 
.A(n_555),
.Y(n_954)
);

INVx1_ASAP7_75t_L g955 ( 
.A(n_461),
.Y(n_955)
);

CKINVDCx5p33_ASAP7_75t_R g956 ( 
.A(n_614),
.Y(n_956)
);

INVx2_ASAP7_75t_SL g957 ( 
.A(n_340),
.Y(n_957)
);

CKINVDCx5p33_ASAP7_75t_R g958 ( 
.A(n_609),
.Y(n_958)
);

INVx1_ASAP7_75t_L g959 ( 
.A(n_537),
.Y(n_959)
);

INVx1_ASAP7_75t_L g960 ( 
.A(n_443),
.Y(n_960)
);

CKINVDCx5p33_ASAP7_75t_R g961 ( 
.A(n_302),
.Y(n_961)
);

CKINVDCx16_ASAP7_75t_R g962 ( 
.A(n_337),
.Y(n_962)
);

INVx1_ASAP7_75t_L g963 ( 
.A(n_332),
.Y(n_963)
);

CKINVDCx5p33_ASAP7_75t_R g964 ( 
.A(n_535),
.Y(n_964)
);

INVx1_ASAP7_75t_L g965 ( 
.A(n_439),
.Y(n_965)
);

NOR2xp67_ASAP7_75t_L g966 ( 
.A(n_528),
.B(n_181),
.Y(n_966)
);

INVx2_ASAP7_75t_L g967 ( 
.A(n_176),
.Y(n_967)
);

INVx1_ASAP7_75t_L g968 ( 
.A(n_87),
.Y(n_968)
);

BUFx6f_ASAP7_75t_L g969 ( 
.A(n_455),
.Y(n_969)
);

CKINVDCx5p33_ASAP7_75t_R g970 ( 
.A(n_7),
.Y(n_970)
);

CKINVDCx5p33_ASAP7_75t_R g971 ( 
.A(n_304),
.Y(n_971)
);

CKINVDCx5p33_ASAP7_75t_R g972 ( 
.A(n_12),
.Y(n_972)
);

INVx1_ASAP7_75t_L g973 ( 
.A(n_577),
.Y(n_973)
);

CKINVDCx5p33_ASAP7_75t_R g974 ( 
.A(n_563),
.Y(n_974)
);

INVx1_ASAP7_75t_L g975 ( 
.A(n_435),
.Y(n_975)
);

BUFx3_ASAP7_75t_L g976 ( 
.A(n_131),
.Y(n_976)
);

INVx1_ASAP7_75t_L g977 ( 
.A(n_671),
.Y(n_977)
);

CKINVDCx5p33_ASAP7_75t_R g978 ( 
.A(n_631),
.Y(n_978)
);

CKINVDCx5p33_ASAP7_75t_R g979 ( 
.A(n_419),
.Y(n_979)
);

INVx2_ASAP7_75t_L g980 ( 
.A(n_43),
.Y(n_980)
);

CKINVDCx5p33_ASAP7_75t_R g981 ( 
.A(n_171),
.Y(n_981)
);

INVxp33_ASAP7_75t_L g982 ( 
.A(n_529),
.Y(n_982)
);

CKINVDCx20_ASAP7_75t_R g983 ( 
.A(n_482),
.Y(n_983)
);

CKINVDCx5p33_ASAP7_75t_R g984 ( 
.A(n_528),
.Y(n_984)
);

INVx1_ASAP7_75t_L g985 ( 
.A(n_303),
.Y(n_985)
);

INVx1_ASAP7_75t_L g986 ( 
.A(n_140),
.Y(n_986)
);

HB1xp67_ASAP7_75t_L g987 ( 
.A(n_653),
.Y(n_987)
);

CKINVDCx5p33_ASAP7_75t_R g988 ( 
.A(n_563),
.Y(n_988)
);

INVx1_ASAP7_75t_L g989 ( 
.A(n_186),
.Y(n_989)
);

CKINVDCx5p33_ASAP7_75t_R g990 ( 
.A(n_391),
.Y(n_990)
);

INVx1_ASAP7_75t_SL g991 ( 
.A(n_24),
.Y(n_991)
);

CKINVDCx5p33_ASAP7_75t_R g992 ( 
.A(n_120),
.Y(n_992)
);

BUFx2_ASAP7_75t_L g993 ( 
.A(n_252),
.Y(n_993)
);

CKINVDCx16_ASAP7_75t_R g994 ( 
.A(n_209),
.Y(n_994)
);

INVx1_ASAP7_75t_L g995 ( 
.A(n_437),
.Y(n_995)
);

CKINVDCx5p33_ASAP7_75t_R g996 ( 
.A(n_54),
.Y(n_996)
);

INVx1_ASAP7_75t_L g997 ( 
.A(n_343),
.Y(n_997)
);

INVx1_ASAP7_75t_L g998 ( 
.A(n_223),
.Y(n_998)
);

CKINVDCx5p33_ASAP7_75t_R g999 ( 
.A(n_4),
.Y(n_999)
);

CKINVDCx5p33_ASAP7_75t_R g1000 ( 
.A(n_373),
.Y(n_1000)
);

CKINVDCx5p33_ASAP7_75t_R g1001 ( 
.A(n_611),
.Y(n_1001)
);

INVxp67_ASAP7_75t_SL g1002 ( 
.A(n_555),
.Y(n_1002)
);

INVx1_ASAP7_75t_L g1003 ( 
.A(n_681),
.Y(n_1003)
);

INVx1_ASAP7_75t_L g1004 ( 
.A(n_155),
.Y(n_1004)
);

CKINVDCx20_ASAP7_75t_R g1005 ( 
.A(n_412),
.Y(n_1005)
);

CKINVDCx5p33_ASAP7_75t_R g1006 ( 
.A(n_124),
.Y(n_1006)
);

BUFx3_ASAP7_75t_L g1007 ( 
.A(n_233),
.Y(n_1007)
);

CKINVDCx5p33_ASAP7_75t_R g1008 ( 
.A(n_546),
.Y(n_1008)
);

CKINVDCx5p33_ASAP7_75t_R g1009 ( 
.A(n_265),
.Y(n_1009)
);

CKINVDCx5p33_ASAP7_75t_R g1010 ( 
.A(n_234),
.Y(n_1010)
);

INVx1_ASAP7_75t_L g1011 ( 
.A(n_232),
.Y(n_1011)
);

INVx1_ASAP7_75t_L g1012 ( 
.A(n_418),
.Y(n_1012)
);

CKINVDCx5p33_ASAP7_75t_R g1013 ( 
.A(n_71),
.Y(n_1013)
);

CKINVDCx16_ASAP7_75t_R g1014 ( 
.A(n_487),
.Y(n_1014)
);

INVx1_ASAP7_75t_L g1015 ( 
.A(n_589),
.Y(n_1015)
);

CKINVDCx5p33_ASAP7_75t_R g1016 ( 
.A(n_126),
.Y(n_1016)
);

INVx1_ASAP7_75t_L g1017 ( 
.A(n_105),
.Y(n_1017)
);

INVx2_ASAP7_75t_L g1018 ( 
.A(n_3),
.Y(n_1018)
);

CKINVDCx5p33_ASAP7_75t_R g1019 ( 
.A(n_239),
.Y(n_1019)
);

INVx1_ASAP7_75t_L g1020 ( 
.A(n_95),
.Y(n_1020)
);

INVxp67_ASAP7_75t_L g1021 ( 
.A(n_319),
.Y(n_1021)
);

CKINVDCx5p33_ASAP7_75t_R g1022 ( 
.A(n_98),
.Y(n_1022)
);

CKINVDCx5p33_ASAP7_75t_R g1023 ( 
.A(n_45),
.Y(n_1023)
);

BUFx2_ASAP7_75t_L g1024 ( 
.A(n_101),
.Y(n_1024)
);

CKINVDCx5p33_ASAP7_75t_R g1025 ( 
.A(n_349),
.Y(n_1025)
);

INVx3_ASAP7_75t_L g1026 ( 
.A(n_250),
.Y(n_1026)
);

CKINVDCx5p33_ASAP7_75t_R g1027 ( 
.A(n_227),
.Y(n_1027)
);

CKINVDCx5p33_ASAP7_75t_R g1028 ( 
.A(n_519),
.Y(n_1028)
);

BUFx2_ASAP7_75t_SL g1029 ( 
.A(n_523),
.Y(n_1029)
);

CKINVDCx5p33_ASAP7_75t_R g1030 ( 
.A(n_184),
.Y(n_1030)
);

BUFx10_ASAP7_75t_L g1031 ( 
.A(n_694),
.Y(n_1031)
);

CKINVDCx14_ASAP7_75t_R g1032 ( 
.A(n_305),
.Y(n_1032)
);

CKINVDCx5p33_ASAP7_75t_R g1033 ( 
.A(n_141),
.Y(n_1033)
);

BUFx3_ASAP7_75t_L g1034 ( 
.A(n_198),
.Y(n_1034)
);

INVx1_ASAP7_75t_L g1035 ( 
.A(n_536),
.Y(n_1035)
);

INVx1_ASAP7_75t_L g1036 ( 
.A(n_288),
.Y(n_1036)
);

BUFx3_ASAP7_75t_L g1037 ( 
.A(n_277),
.Y(n_1037)
);

INVx1_ASAP7_75t_L g1038 ( 
.A(n_188),
.Y(n_1038)
);

BUFx3_ASAP7_75t_L g1039 ( 
.A(n_252),
.Y(n_1039)
);

BUFx5_ASAP7_75t_L g1040 ( 
.A(n_331),
.Y(n_1040)
);

INVx1_ASAP7_75t_L g1041 ( 
.A(n_80),
.Y(n_1041)
);

INVxp33_ASAP7_75t_L g1042 ( 
.A(n_443),
.Y(n_1042)
);

CKINVDCx5p33_ASAP7_75t_R g1043 ( 
.A(n_621),
.Y(n_1043)
);

INVx1_ASAP7_75t_SL g1044 ( 
.A(n_302),
.Y(n_1044)
);

CKINVDCx5p33_ASAP7_75t_R g1045 ( 
.A(n_620),
.Y(n_1045)
);

CKINVDCx5p33_ASAP7_75t_R g1046 ( 
.A(n_97),
.Y(n_1046)
);

INVx1_ASAP7_75t_L g1047 ( 
.A(n_46),
.Y(n_1047)
);

INVx1_ASAP7_75t_L g1048 ( 
.A(n_70),
.Y(n_1048)
);

BUFx5_ASAP7_75t_L g1049 ( 
.A(n_88),
.Y(n_1049)
);

CKINVDCx20_ASAP7_75t_R g1050 ( 
.A(n_355),
.Y(n_1050)
);

INVx1_ASAP7_75t_L g1051 ( 
.A(n_418),
.Y(n_1051)
);

INVx1_ASAP7_75t_L g1052 ( 
.A(n_301),
.Y(n_1052)
);

CKINVDCx16_ASAP7_75t_R g1053 ( 
.A(n_103),
.Y(n_1053)
);

CKINVDCx5p33_ASAP7_75t_R g1054 ( 
.A(n_490),
.Y(n_1054)
);

INVx2_ASAP7_75t_L g1055 ( 
.A(n_22),
.Y(n_1055)
);

CKINVDCx5p33_ASAP7_75t_R g1056 ( 
.A(n_84),
.Y(n_1056)
);

INVx1_ASAP7_75t_SL g1057 ( 
.A(n_482),
.Y(n_1057)
);

INVx1_ASAP7_75t_L g1058 ( 
.A(n_395),
.Y(n_1058)
);

INVx1_ASAP7_75t_L g1059 ( 
.A(n_285),
.Y(n_1059)
);

CKINVDCx5p33_ASAP7_75t_R g1060 ( 
.A(n_463),
.Y(n_1060)
);

CKINVDCx5p33_ASAP7_75t_R g1061 ( 
.A(n_597),
.Y(n_1061)
);

CKINVDCx5p33_ASAP7_75t_R g1062 ( 
.A(n_13),
.Y(n_1062)
);

BUFx2_ASAP7_75t_L g1063 ( 
.A(n_303),
.Y(n_1063)
);

CKINVDCx5p33_ASAP7_75t_R g1064 ( 
.A(n_551),
.Y(n_1064)
);

CKINVDCx5p33_ASAP7_75t_R g1065 ( 
.A(n_183),
.Y(n_1065)
);

CKINVDCx5p33_ASAP7_75t_R g1066 ( 
.A(n_83),
.Y(n_1066)
);

BUFx3_ASAP7_75t_L g1067 ( 
.A(n_78),
.Y(n_1067)
);

BUFx2_ASAP7_75t_L g1068 ( 
.A(n_503),
.Y(n_1068)
);

CKINVDCx5p33_ASAP7_75t_R g1069 ( 
.A(n_326),
.Y(n_1069)
);

CKINVDCx5p33_ASAP7_75t_R g1070 ( 
.A(n_176),
.Y(n_1070)
);

CKINVDCx5p33_ASAP7_75t_R g1071 ( 
.A(n_224),
.Y(n_1071)
);

CKINVDCx5p33_ASAP7_75t_R g1072 ( 
.A(n_672),
.Y(n_1072)
);

CKINVDCx5p33_ASAP7_75t_R g1073 ( 
.A(n_215),
.Y(n_1073)
);

CKINVDCx5p33_ASAP7_75t_R g1074 ( 
.A(n_116),
.Y(n_1074)
);

INVx1_ASAP7_75t_L g1075 ( 
.A(n_273),
.Y(n_1075)
);

INVx1_ASAP7_75t_L g1076 ( 
.A(n_481),
.Y(n_1076)
);

INVx1_ASAP7_75t_L g1077 ( 
.A(n_386),
.Y(n_1077)
);

CKINVDCx5p33_ASAP7_75t_R g1078 ( 
.A(n_434),
.Y(n_1078)
);

CKINVDCx5p33_ASAP7_75t_R g1079 ( 
.A(n_376),
.Y(n_1079)
);

INVx1_ASAP7_75t_L g1080 ( 
.A(n_235),
.Y(n_1080)
);

CKINVDCx5p33_ASAP7_75t_R g1081 ( 
.A(n_206),
.Y(n_1081)
);

CKINVDCx20_ASAP7_75t_R g1082 ( 
.A(n_642),
.Y(n_1082)
);

BUFx2_ASAP7_75t_L g1083 ( 
.A(n_71),
.Y(n_1083)
);

INVxp33_ASAP7_75t_SL g1084 ( 
.A(n_216),
.Y(n_1084)
);

INVx1_ASAP7_75t_L g1085 ( 
.A(n_108),
.Y(n_1085)
);

CKINVDCx5p33_ASAP7_75t_R g1086 ( 
.A(n_168),
.Y(n_1086)
);

INVx1_ASAP7_75t_L g1087 ( 
.A(n_551),
.Y(n_1087)
);

INVx1_ASAP7_75t_SL g1088 ( 
.A(n_664),
.Y(n_1088)
);

CKINVDCx5p33_ASAP7_75t_R g1089 ( 
.A(n_649),
.Y(n_1089)
);

CKINVDCx5p33_ASAP7_75t_R g1090 ( 
.A(n_478),
.Y(n_1090)
);

CKINVDCx16_ASAP7_75t_R g1091 ( 
.A(n_223),
.Y(n_1091)
);

CKINVDCx5p33_ASAP7_75t_R g1092 ( 
.A(n_676),
.Y(n_1092)
);

CKINVDCx20_ASAP7_75t_R g1093 ( 
.A(n_362),
.Y(n_1093)
);

CKINVDCx5p33_ASAP7_75t_R g1094 ( 
.A(n_469),
.Y(n_1094)
);

INVx2_ASAP7_75t_L g1095 ( 
.A(n_359),
.Y(n_1095)
);

CKINVDCx5p33_ASAP7_75t_R g1096 ( 
.A(n_598),
.Y(n_1096)
);

CKINVDCx5p33_ASAP7_75t_R g1097 ( 
.A(n_689),
.Y(n_1097)
);

CKINVDCx16_ASAP7_75t_R g1098 ( 
.A(n_193),
.Y(n_1098)
);

CKINVDCx5p33_ASAP7_75t_R g1099 ( 
.A(n_405),
.Y(n_1099)
);

CKINVDCx5p33_ASAP7_75t_R g1100 ( 
.A(n_759),
.Y(n_1100)
);

AND2x4_ASAP7_75t_L g1101 ( 
.A(n_1026),
.B(n_717),
.Y(n_1101)
);

OAI21x1_ASAP7_75t_L g1102 ( 
.A1(n_767),
.A2(n_637),
.B(n_635),
.Y(n_1102)
);

HB1xp67_ASAP7_75t_L g1103 ( 
.A(n_1032),
.Y(n_1103)
);

BUFx2_ASAP7_75t_L g1104 ( 
.A(n_734),
.Y(n_1104)
);

BUFx6f_ASAP7_75t_L g1105 ( 
.A(n_883),
.Y(n_1105)
);

OA21x2_ASAP7_75t_L g1106 ( 
.A1(n_767),
.A2(n_643),
.B(n_640),
.Y(n_1106)
);

BUFx8_ASAP7_75t_SL g1107 ( 
.A(n_706),
.Y(n_1107)
);

INVx3_ASAP7_75t_L g1108 ( 
.A(n_1026),
.Y(n_1108)
);

AOI22xp5_ASAP7_75t_L g1109 ( 
.A1(n_717),
.A2(n_2),
.B1(n_0),
.B2(n_1),
.Y(n_1109)
);

BUFx6f_ASAP7_75t_L g1110 ( 
.A(n_883),
.Y(n_1110)
);

INVx3_ASAP7_75t_L g1111 ( 
.A(n_712),
.Y(n_1111)
);

INVx1_ASAP7_75t_L g1112 ( 
.A(n_987),
.Y(n_1112)
);

AND2x4_ASAP7_75t_L g1113 ( 
.A(n_820),
.B(n_0),
.Y(n_1113)
);

OAI22x1_ASAP7_75t_R g1114 ( 
.A1(n_706),
.A2(n_4),
.B1(n_1),
.B2(n_3),
.Y(n_1114)
);

INVx1_ASAP7_75t_L g1115 ( 
.A(n_820),
.Y(n_1115)
);

INVx2_ASAP7_75t_SL g1116 ( 
.A(n_712),
.Y(n_1116)
);

HB1xp67_ASAP7_75t_L g1117 ( 
.A(n_800),
.Y(n_1117)
);

BUFx6f_ASAP7_75t_L g1118 ( 
.A(n_883),
.Y(n_1118)
);

INVx1_ASAP7_75t_L g1119 ( 
.A(n_875),
.Y(n_1119)
);

INVx5_ASAP7_75t_L g1120 ( 
.A(n_1031),
.Y(n_1120)
);

HB1xp67_ASAP7_75t_L g1121 ( 
.A(n_824),
.Y(n_1121)
);

BUFx6f_ASAP7_75t_L g1122 ( 
.A(n_883),
.Y(n_1122)
);

BUFx8_ASAP7_75t_L g1123 ( 
.A(n_881),
.Y(n_1123)
);

NAND2xp5_ASAP7_75t_L g1124 ( 
.A(n_875),
.B(n_6),
.Y(n_1124)
);

AND2x4_ASAP7_75t_L g1125 ( 
.A(n_902),
.B(n_7),
.Y(n_1125)
);

AOI22xp5_ASAP7_75t_L g1126 ( 
.A1(n_902),
.A2(n_10),
.B1(n_8),
.B2(n_9),
.Y(n_1126)
);

NAND2xp33_ASAP7_75t_L g1127 ( 
.A(n_708),
.B(n_645),
.Y(n_1127)
);

INVx1_ASAP7_75t_L g1128 ( 
.A(n_935),
.Y(n_1128)
);

NAND2xp5_ASAP7_75t_L g1129 ( 
.A(n_957),
.B(n_8),
.Y(n_1129)
);

BUFx6f_ASAP7_75t_L g1130 ( 
.A(n_766),
.Y(n_1130)
);

OAI22xp5_ASAP7_75t_L g1131 ( 
.A1(n_705),
.A2(n_12),
.B1(n_10),
.B2(n_11),
.Y(n_1131)
);

HB1xp67_ASAP7_75t_L g1132 ( 
.A(n_839),
.Y(n_1132)
);

AOI22xp5_ASAP7_75t_L g1133 ( 
.A1(n_1084),
.A2(n_15),
.B1(n_11),
.B2(n_14),
.Y(n_1133)
);

BUFx12f_ASAP7_75t_L g1134 ( 
.A(n_712),
.Y(n_1134)
);

INVx5_ASAP7_75t_L g1135 ( 
.A(n_1031),
.Y(n_1135)
);

INVx2_ASAP7_75t_L g1136 ( 
.A(n_708),
.Y(n_1136)
);

OA21x2_ASAP7_75t_L g1137 ( 
.A1(n_775),
.A2(n_647),
.B(n_646),
.Y(n_1137)
);

OAI21x1_ASAP7_75t_L g1138 ( 
.A1(n_775),
.A2(n_652),
.B(n_648),
.Y(n_1138)
);

INVx3_ASAP7_75t_L g1139 ( 
.A(n_760),
.Y(n_1139)
);

AND2x6_ASAP7_75t_L g1140 ( 
.A(n_877),
.B(n_654),
.Y(n_1140)
);

INVx4_ASAP7_75t_L g1141 ( 
.A(n_1031),
.Y(n_1141)
);

HB1xp67_ASAP7_75t_L g1142 ( 
.A(n_907),
.Y(n_1142)
);

INVx1_ASAP7_75t_L g1143 ( 
.A(n_799),
.Y(n_1143)
);

INVx5_ASAP7_75t_L g1144 ( 
.A(n_877),
.Y(n_1144)
);

AND2x2_ASAP7_75t_L g1145 ( 
.A(n_897),
.B(n_14),
.Y(n_1145)
);

NOR2xp33_ASAP7_75t_L g1146 ( 
.A(n_982),
.B(n_16),
.Y(n_1146)
);

INVx3_ASAP7_75t_L g1147 ( 
.A(n_760),
.Y(n_1147)
);

AOI22xp5_ASAP7_75t_L g1148 ( 
.A1(n_1084),
.A2(n_18),
.B1(n_16),
.B2(n_17),
.Y(n_1148)
);

HB1xp67_ASAP7_75t_L g1149 ( 
.A(n_799),
.Y(n_1149)
);

INVx2_ASAP7_75t_L g1150 ( 
.A(n_708),
.Y(n_1150)
);

CKINVDCx5p33_ASAP7_75t_R g1151 ( 
.A(n_832),
.Y(n_1151)
);

AND2x2_ASAP7_75t_L g1152 ( 
.A(n_1042),
.B(n_17),
.Y(n_1152)
);

INVx1_ASAP7_75t_L g1153 ( 
.A(n_887),
.Y(n_1153)
);

BUFx6f_ASAP7_75t_L g1154 ( 
.A(n_766),
.Y(n_1154)
);

CKINVDCx5p33_ASAP7_75t_R g1155 ( 
.A(n_918),
.Y(n_1155)
);

NOR2xp33_ASAP7_75t_SL g1156 ( 
.A(n_726),
.B(n_658),
.Y(n_1156)
);

BUFx6f_ASAP7_75t_L g1157 ( 
.A(n_766),
.Y(n_1157)
);

INVxp67_ASAP7_75t_L g1158 ( 
.A(n_812),
.Y(n_1158)
);

INVx2_ASAP7_75t_L g1159 ( 
.A(n_708),
.Y(n_1159)
);

AOI22xp5_ASAP7_75t_SL g1160 ( 
.A1(n_721),
.A2(n_748),
.B1(n_750),
.B2(n_729),
.Y(n_1160)
);

AND2x4_ASAP7_75t_L g1161 ( 
.A(n_887),
.B(n_18),
.Y(n_1161)
);

HB1xp67_ASAP7_75t_L g1162 ( 
.A(n_911),
.Y(n_1162)
);

NAND2xp5_ASAP7_75t_L g1163 ( 
.A(n_817),
.B(n_20),
.Y(n_1163)
);

INVx4_ASAP7_75t_L g1164 ( 
.A(n_722),
.Y(n_1164)
);

BUFx6f_ASAP7_75t_L g1165 ( 
.A(n_766),
.Y(n_1165)
);

INVx3_ASAP7_75t_L g1166 ( 
.A(n_760),
.Y(n_1166)
);

AND2x2_ASAP7_75t_L g1167 ( 
.A(n_993),
.B(n_21),
.Y(n_1167)
);

INVx3_ASAP7_75t_L g1168 ( 
.A(n_797),
.Y(n_1168)
);

INVx1_ASAP7_75t_L g1169 ( 
.A(n_911),
.Y(n_1169)
);

AND2x6_ASAP7_75t_L g1170 ( 
.A(n_874),
.B(n_662),
.Y(n_1170)
);

NAND2xp5_ASAP7_75t_L g1171 ( 
.A(n_1024),
.B(n_21),
.Y(n_1171)
);

NOR2xp33_ASAP7_75t_L g1172 ( 
.A(n_1063),
.B(n_22),
.Y(n_1172)
);

INVx2_ASAP7_75t_L g1173 ( 
.A(n_1040),
.Y(n_1173)
);

AOI22x1_ASAP7_75t_SL g1174 ( 
.A1(n_721),
.A2(n_25),
.B1(n_23),
.B2(n_24),
.Y(n_1174)
);

BUFx3_ASAP7_75t_L g1175 ( 
.A(n_886),
.Y(n_1175)
);

NAND2xp5_ASAP7_75t_L g1176 ( 
.A(n_1068),
.B(n_1083),
.Y(n_1176)
);

OAI22x1_ASAP7_75t_R g1177 ( 
.A1(n_729),
.A2(n_26),
.B1(n_23),
.B2(n_25),
.Y(n_1177)
);

INVx2_ASAP7_75t_L g1178 ( 
.A(n_1040),
.Y(n_1178)
);

AOI22x1_ASAP7_75t_SL g1179 ( 
.A1(n_748),
.A2(n_28),
.B1(n_26),
.B2(n_27),
.Y(n_1179)
);

INVx2_ASAP7_75t_SL g1180 ( 
.A(n_797),
.Y(n_1180)
);

INVx2_ASAP7_75t_L g1181 ( 
.A(n_1040),
.Y(n_1181)
);

INVx3_ASAP7_75t_L g1182 ( 
.A(n_797),
.Y(n_1182)
);

OR2x6_ASAP7_75t_L g1183 ( 
.A(n_1029),
.B(n_27),
.Y(n_1183)
);

BUFx6f_ASAP7_75t_L g1184 ( 
.A(n_780),
.Y(n_1184)
);

AND2x4_ASAP7_75t_L g1185 ( 
.A(n_915),
.B(n_928),
.Y(n_1185)
);

INVx2_ASAP7_75t_SL g1186 ( 
.A(n_810),
.Y(n_1186)
);

CKINVDCx5p33_ASAP7_75t_R g1187 ( 
.A(n_918),
.Y(n_1187)
);

BUFx12f_ASAP7_75t_L g1188 ( 
.A(n_810),
.Y(n_1188)
);

INVx2_ASAP7_75t_L g1189 ( 
.A(n_1040),
.Y(n_1189)
);

OR2x2_ASAP7_75t_L g1190 ( 
.A(n_755),
.B(n_29),
.Y(n_1190)
);

INVx2_ASAP7_75t_L g1191 ( 
.A(n_1040),
.Y(n_1191)
);

INVx1_ASAP7_75t_L g1192 ( 
.A(n_915),
.Y(n_1192)
);

AND2x4_ASAP7_75t_L g1193 ( 
.A(n_928),
.B(n_29),
.Y(n_1193)
);

BUFx12f_ASAP7_75t_L g1194 ( 
.A(n_810),
.Y(n_1194)
);

CKINVDCx5p33_ASAP7_75t_R g1195 ( 
.A(n_1082),
.Y(n_1195)
);

INVx1_ASAP7_75t_L g1196 ( 
.A(n_938),
.Y(n_1196)
);

INVx2_ASAP7_75t_L g1197 ( 
.A(n_1108),
.Y(n_1197)
);

INVx11_ASAP7_75t_L g1198 ( 
.A(n_1123),
.Y(n_1198)
);

INVx1_ASAP7_75t_L g1199 ( 
.A(n_1113),
.Y(n_1199)
);

INVx2_ASAP7_75t_L g1200 ( 
.A(n_1108),
.Y(n_1200)
);

INVx2_ASAP7_75t_L g1201 ( 
.A(n_1185),
.Y(n_1201)
);

INVx1_ASAP7_75t_L g1202 ( 
.A(n_1125),
.Y(n_1202)
);

INVx2_ASAP7_75t_L g1203 ( 
.A(n_1185),
.Y(n_1203)
);

OAI22xp33_ASAP7_75t_L g1204 ( 
.A1(n_1133),
.A2(n_912),
.B1(n_962),
.B2(n_873),
.Y(n_1204)
);

BUFx3_ASAP7_75t_L g1205 ( 
.A(n_1101),
.Y(n_1205)
);

BUFx3_ASAP7_75t_L g1206 ( 
.A(n_1101),
.Y(n_1206)
);

AND2x2_ASAP7_75t_L g1207 ( 
.A(n_1117),
.B(n_1091),
.Y(n_1207)
);

INVx2_ASAP7_75t_L g1208 ( 
.A(n_1136),
.Y(n_1208)
);

NAND2xp33_ASAP7_75t_L g1209 ( 
.A(n_1140),
.B(n_1049),
.Y(n_1209)
);

AND2x2_ASAP7_75t_L g1210 ( 
.A(n_1117),
.B(n_1098),
.Y(n_1210)
);

BUFx6f_ASAP7_75t_L g1211 ( 
.A(n_1105),
.Y(n_1211)
);

INVx2_ASAP7_75t_L g1212 ( 
.A(n_1150),
.Y(n_1212)
);

INVx2_ASAP7_75t_L g1213 ( 
.A(n_1159),
.Y(n_1213)
);

INVx1_ASAP7_75t_L g1214 ( 
.A(n_1125),
.Y(n_1214)
);

NAND2xp5_ASAP7_75t_SL g1215 ( 
.A(n_1173),
.B(n_1178),
.Y(n_1215)
);

NAND2xp5_ASAP7_75t_L g1216 ( 
.A(n_1149),
.B(n_725),
.Y(n_1216)
);

AND2x6_ASAP7_75t_L g1217 ( 
.A(n_1161),
.B(n_1193),
.Y(n_1217)
);

OAI22xp33_ASAP7_75t_L g1218 ( 
.A1(n_1148),
.A2(n_1014),
.B1(n_1053),
.B2(n_994),
.Y(n_1218)
);

INVxp33_ASAP7_75t_SL g1219 ( 
.A(n_1103),
.Y(n_1219)
);

INVx1_ASAP7_75t_L g1220 ( 
.A(n_1149),
.Y(n_1220)
);

BUFx6f_ASAP7_75t_SL g1221 ( 
.A(n_1183),
.Y(n_1221)
);

INVx1_ASAP7_75t_L g1222 ( 
.A(n_1162),
.Y(n_1222)
);

INVx2_ASAP7_75t_L g1223 ( 
.A(n_1181),
.Y(n_1223)
);

NAND2xp5_ASAP7_75t_L g1224 ( 
.A(n_1115),
.B(n_776),
.Y(n_1224)
);

AOI21x1_ASAP7_75t_L g1225 ( 
.A1(n_1189),
.A2(n_773),
.B(n_736),
.Y(n_1225)
);

OR2x6_ASAP7_75t_L g1226 ( 
.A(n_1134),
.B(n_749),
.Y(n_1226)
);

INVx3_ASAP7_75t_L g1227 ( 
.A(n_1161),
.Y(n_1227)
);

NAND2xp5_ASAP7_75t_L g1228 ( 
.A(n_1119),
.B(n_922),
.Y(n_1228)
);

INVx2_ASAP7_75t_L g1229 ( 
.A(n_1191),
.Y(n_1229)
);

INVx2_ASAP7_75t_L g1230 ( 
.A(n_1128),
.Y(n_1230)
);

OR2x6_ASAP7_75t_L g1231 ( 
.A(n_1188),
.B(n_765),
.Y(n_1231)
);

INVx3_ASAP7_75t_L g1232 ( 
.A(n_1111),
.Y(n_1232)
);

NAND2xp33_ASAP7_75t_L g1233 ( 
.A(n_1140),
.B(n_1049),
.Y(n_1233)
);

NAND3xp33_ASAP7_75t_L g1234 ( 
.A(n_1112),
.B(n_768),
.C(n_762),
.Y(n_1234)
);

AND3x2_ASAP7_75t_L g1235 ( 
.A(n_1104),
.B(n_1132),
.C(n_1121),
.Y(n_1235)
);

INVx2_ASAP7_75t_L g1236 ( 
.A(n_1175),
.Y(n_1236)
);

INVx3_ASAP7_75t_L g1237 ( 
.A(n_1111),
.Y(n_1237)
);

INVx2_ASAP7_75t_L g1238 ( 
.A(n_1175),
.Y(n_1238)
);

INVx1_ASAP7_75t_L g1239 ( 
.A(n_1124),
.Y(n_1239)
);

BUFx6f_ASAP7_75t_L g1240 ( 
.A(n_1105),
.Y(n_1240)
);

BUFx6f_ASAP7_75t_L g1241 ( 
.A(n_1105),
.Y(n_1241)
);

AND2x2_ASAP7_75t_L g1242 ( 
.A(n_1121),
.B(n_867),
.Y(n_1242)
);

INVx3_ASAP7_75t_L g1243 ( 
.A(n_1139),
.Y(n_1243)
);

OR2x6_ASAP7_75t_L g1244 ( 
.A(n_1194),
.B(n_1183),
.Y(n_1244)
);

INVxp67_ASAP7_75t_L g1245 ( 
.A(n_1132),
.Y(n_1245)
);

AND2x2_ASAP7_75t_L g1246 ( 
.A(n_1142),
.B(n_867),
.Y(n_1246)
);

INVxp33_ASAP7_75t_SL g1247 ( 
.A(n_1151),
.Y(n_1247)
);

INVx1_ASAP7_75t_L g1248 ( 
.A(n_1129),
.Y(n_1248)
);

INVxp33_ASAP7_75t_L g1249 ( 
.A(n_1142),
.Y(n_1249)
);

INVx2_ASAP7_75t_L g1250 ( 
.A(n_1143),
.Y(n_1250)
);

INVx1_ASAP7_75t_L g1251 ( 
.A(n_1129),
.Y(n_1251)
);

INVx1_ASAP7_75t_L g1252 ( 
.A(n_1153),
.Y(n_1252)
);

INVx2_ASAP7_75t_L g1253 ( 
.A(n_1169),
.Y(n_1253)
);

INVx2_ASAP7_75t_L g1254 ( 
.A(n_1192),
.Y(n_1254)
);

AND2x2_ASAP7_75t_L g1255 ( 
.A(n_1158),
.B(n_867),
.Y(n_1255)
);

INVx1_ASAP7_75t_L g1256 ( 
.A(n_1196),
.Y(n_1256)
);

INVx1_ASAP7_75t_L g1257 ( 
.A(n_1139),
.Y(n_1257)
);

OR2x2_ASAP7_75t_SL g1258 ( 
.A(n_1176),
.B(n_724),
.Y(n_1258)
);

CKINVDCx6p67_ASAP7_75t_R g1259 ( 
.A(n_1183),
.Y(n_1259)
);

INVx1_ASAP7_75t_L g1260 ( 
.A(n_1147),
.Y(n_1260)
);

NAND2xp5_ASAP7_75t_L g1261 ( 
.A(n_1120),
.B(n_1135),
.Y(n_1261)
);

HB1xp67_ASAP7_75t_L g1262 ( 
.A(n_1158),
.Y(n_1262)
);

INVx3_ASAP7_75t_L g1263 ( 
.A(n_1147),
.Y(n_1263)
);

AND2x2_ASAP7_75t_L g1264 ( 
.A(n_1176),
.B(n_938),
.Y(n_1264)
);

BUFx6f_ASAP7_75t_L g1265 ( 
.A(n_1110),
.Y(n_1265)
);

BUFx3_ASAP7_75t_L g1266 ( 
.A(n_1140),
.Y(n_1266)
);

INVx1_ASAP7_75t_L g1267 ( 
.A(n_1166),
.Y(n_1267)
);

NAND2xp5_ASAP7_75t_L g1268 ( 
.A(n_1120),
.B(n_882),
.Y(n_1268)
);

BUFx6f_ASAP7_75t_L g1269 ( 
.A(n_1110),
.Y(n_1269)
);

NAND2xp5_ASAP7_75t_SL g1270 ( 
.A(n_1120),
.B(n_781),
.Y(n_1270)
);

INVx1_ASAP7_75t_L g1271 ( 
.A(n_1168),
.Y(n_1271)
);

HB1xp67_ASAP7_75t_L g1272 ( 
.A(n_1145),
.Y(n_1272)
);

AND2x4_ASAP7_75t_L g1273 ( 
.A(n_1182),
.B(n_976),
.Y(n_1273)
);

NOR2xp33_ASAP7_75t_L g1274 ( 
.A(n_1141),
.B(n_792),
.Y(n_1274)
);

NAND2xp5_ASAP7_75t_SL g1275 ( 
.A(n_1120),
.B(n_807),
.Y(n_1275)
);

HB1xp67_ASAP7_75t_L g1276 ( 
.A(n_1152),
.Y(n_1276)
);

INVx2_ASAP7_75t_L g1277 ( 
.A(n_1144),
.Y(n_1277)
);

NOR2xp33_ASAP7_75t_L g1278 ( 
.A(n_1135),
.B(n_821),
.Y(n_1278)
);

NAND2xp5_ASAP7_75t_SL g1279 ( 
.A(n_1135),
.B(n_837),
.Y(n_1279)
);

BUFx10_ASAP7_75t_L g1280 ( 
.A(n_1100),
.Y(n_1280)
);

NAND2xp5_ASAP7_75t_SL g1281 ( 
.A(n_1135),
.B(n_845),
.Y(n_1281)
);

INVx2_ASAP7_75t_L g1282 ( 
.A(n_1130),
.Y(n_1282)
);

INVx3_ASAP7_75t_L g1283 ( 
.A(n_1182),
.Y(n_1283)
);

OAI22xp5_ASAP7_75t_L g1284 ( 
.A1(n_1190),
.A2(n_750),
.B1(n_798),
.B2(n_786),
.Y(n_1284)
);

BUFx4f_ASAP7_75t_L g1285 ( 
.A(n_1140),
.Y(n_1285)
);

INVx1_ASAP7_75t_L g1286 ( 
.A(n_1163),
.Y(n_1286)
);

INVx2_ASAP7_75t_SL g1287 ( 
.A(n_1164),
.Y(n_1287)
);

INVx1_ASAP7_75t_L g1288 ( 
.A(n_1163),
.Y(n_1288)
);

NAND2xp33_ASAP7_75t_L g1289 ( 
.A(n_1170),
.B(n_1100),
.Y(n_1289)
);

INVx2_ASAP7_75t_L g1290 ( 
.A(n_1130),
.Y(n_1290)
);

NOR2x1p5_ASAP7_75t_L g1291 ( 
.A(n_1151),
.B(n_1099),
.Y(n_1291)
);

OA22x2_ASAP7_75t_L g1292 ( 
.A1(n_1109),
.A2(n_739),
.B1(n_704),
.B2(n_715),
.Y(n_1292)
);

INVx1_ASAP7_75t_L g1293 ( 
.A(n_1171),
.Y(n_1293)
);

AND2x2_ASAP7_75t_L g1294 ( 
.A(n_1167),
.B(n_976),
.Y(n_1294)
);

INVx2_ASAP7_75t_L g1295 ( 
.A(n_1154),
.Y(n_1295)
);

BUFx6f_ASAP7_75t_L g1296 ( 
.A(n_1110),
.Y(n_1296)
);

INVx4_ASAP7_75t_L g1297 ( 
.A(n_1170),
.Y(n_1297)
);

INVx1_ASAP7_75t_L g1298 ( 
.A(n_1171),
.Y(n_1298)
);

NOR2xp33_ASAP7_75t_L g1299 ( 
.A(n_1164),
.B(n_940),
.Y(n_1299)
);

INVx2_ASAP7_75t_SL g1300 ( 
.A(n_1116),
.Y(n_1300)
);

NAND2xp5_ASAP7_75t_L g1301 ( 
.A(n_1180),
.B(n_977),
.Y(n_1301)
);

INVxp67_ASAP7_75t_L g1302 ( 
.A(n_1146),
.Y(n_1302)
);

INVx2_ASAP7_75t_SL g1303 ( 
.A(n_1186),
.Y(n_1303)
);

INVx5_ASAP7_75t_L g1304 ( 
.A(n_1170),
.Y(n_1304)
);

NAND2xp5_ASAP7_75t_SL g1305 ( 
.A(n_1156),
.B(n_1003),
.Y(n_1305)
);

INVx2_ASAP7_75t_L g1306 ( 
.A(n_1157),
.Y(n_1306)
);

INVx4_ASAP7_75t_L g1307 ( 
.A(n_1170),
.Y(n_1307)
);

BUFx10_ASAP7_75t_L g1308 ( 
.A(n_1146),
.Y(n_1308)
);

BUFx10_ASAP7_75t_L g1309 ( 
.A(n_1172),
.Y(n_1309)
);

NAND2xp5_ASAP7_75t_L g1310 ( 
.A(n_1184),
.B(n_1049),
.Y(n_1310)
);

INVx2_ASAP7_75t_L g1311 ( 
.A(n_1157),
.Y(n_1311)
);

INVx1_ASAP7_75t_L g1312 ( 
.A(n_1172),
.Y(n_1312)
);

INVx3_ASAP7_75t_L g1313 ( 
.A(n_1102),
.Y(n_1313)
);

AND2x2_ASAP7_75t_L g1314 ( 
.A(n_1155),
.B(n_1187),
.Y(n_1314)
);

NOR2xp33_ASAP7_75t_L g1315 ( 
.A(n_1165),
.B(n_846),
.Y(n_1315)
);

NAND2xp33_ASAP7_75t_SL g1316 ( 
.A(n_1131),
.B(n_1082),
.Y(n_1316)
);

NOR2xp33_ASAP7_75t_L g1317 ( 
.A(n_1165),
.B(n_947),
.Y(n_1317)
);

BUFx2_ASAP7_75t_L g1318 ( 
.A(n_1123),
.Y(n_1318)
);

INVx2_ASAP7_75t_L g1319 ( 
.A(n_1165),
.Y(n_1319)
);

INVx3_ASAP7_75t_L g1320 ( 
.A(n_1138),
.Y(n_1320)
);

INVx2_ASAP7_75t_L g1321 ( 
.A(n_1184),
.Y(n_1321)
);

OR2x2_ASAP7_75t_L g1322 ( 
.A(n_1160),
.B(n_1090),
.Y(n_1322)
);

AND2x2_ASAP7_75t_L g1323 ( 
.A(n_1155),
.B(n_1187),
.Y(n_1323)
);

NAND2xp5_ASAP7_75t_SL g1324 ( 
.A(n_1118),
.B(n_742),
.Y(n_1324)
);

INVx5_ASAP7_75t_L g1325 ( 
.A(n_1118),
.Y(n_1325)
);

BUFx3_ASAP7_75t_L g1326 ( 
.A(n_1106),
.Y(n_1326)
);

INVx2_ASAP7_75t_L g1327 ( 
.A(n_1184),
.Y(n_1327)
);

NAND2xp5_ASAP7_75t_SL g1328 ( 
.A(n_1122),
.B(n_742),
.Y(n_1328)
);

INVx1_ASAP7_75t_SL g1329 ( 
.A(n_1195),
.Y(n_1329)
);

INVx1_ASAP7_75t_L g1330 ( 
.A(n_1184),
.Y(n_1330)
);

OAI22xp33_ASAP7_75t_L g1331 ( 
.A1(n_1126),
.A2(n_798),
.B1(n_803),
.B2(n_786),
.Y(n_1331)
);

CKINVDCx5p33_ASAP7_75t_R g1332 ( 
.A(n_1107),
.Y(n_1332)
);

NAND2xp5_ASAP7_75t_L g1333 ( 
.A(n_1122),
.B(n_1049),
.Y(n_1333)
);

INVx3_ASAP7_75t_L g1334 ( 
.A(n_1106),
.Y(n_1334)
);

INVx1_ASAP7_75t_L g1335 ( 
.A(n_1127),
.Y(n_1335)
);

INVx1_ASAP7_75t_L g1336 ( 
.A(n_1127),
.Y(n_1336)
);

BUFx10_ASAP7_75t_L g1337 ( 
.A(n_1195),
.Y(n_1337)
);

NAND2xp5_ASAP7_75t_L g1338 ( 
.A(n_1122),
.B(n_1049),
.Y(n_1338)
);

INVx1_ASAP7_75t_L g1339 ( 
.A(n_1137),
.Y(n_1339)
);

INVx2_ASAP7_75t_L g1340 ( 
.A(n_1137),
.Y(n_1340)
);

INVx1_ASAP7_75t_L g1341 ( 
.A(n_1131),
.Y(n_1341)
);

INVx2_ASAP7_75t_SL g1342 ( 
.A(n_1114),
.Y(n_1342)
);

NAND2xp5_ASAP7_75t_L g1343 ( 
.A(n_1174),
.B(n_1049),
.Y(n_1343)
);

BUFx6f_ASAP7_75t_L g1344 ( 
.A(n_1177),
.Y(n_1344)
);

INVx1_ASAP7_75t_L g1345 ( 
.A(n_1179),
.Y(n_1345)
);

OR2x6_ASAP7_75t_L g1346 ( 
.A(n_1107),
.B(n_966),
.Y(n_1346)
);

INVx2_ASAP7_75t_L g1347 ( 
.A(n_1108),
.Y(n_1347)
);

AND2x2_ASAP7_75t_L g1348 ( 
.A(n_1117),
.B(n_1007),
.Y(n_1348)
);

INVx2_ASAP7_75t_L g1349 ( 
.A(n_1108),
.Y(n_1349)
);

INVx1_ASAP7_75t_L g1350 ( 
.A(n_1113),
.Y(n_1350)
);

INVx2_ASAP7_75t_L g1351 ( 
.A(n_1108),
.Y(n_1351)
);

INVx3_ASAP7_75t_L g1352 ( 
.A(n_1113),
.Y(n_1352)
);

INVx2_ASAP7_75t_L g1353 ( 
.A(n_1108),
.Y(n_1353)
);

CKINVDCx5p33_ASAP7_75t_R g1354 ( 
.A(n_1151),
.Y(n_1354)
);

NAND2xp33_ASAP7_75t_SL g1355 ( 
.A(n_1145),
.B(n_747),
.Y(n_1355)
);

CKINVDCx5p33_ASAP7_75t_R g1356 ( 
.A(n_1151),
.Y(n_1356)
);

INVx1_ASAP7_75t_L g1357 ( 
.A(n_1113),
.Y(n_1357)
);

INVxp67_ASAP7_75t_L g1358 ( 
.A(n_1262),
.Y(n_1358)
);

INVx2_ASAP7_75t_L g1359 ( 
.A(n_1236),
.Y(n_1359)
);

AOI221xp5_ASAP7_75t_L g1360 ( 
.A1(n_1341),
.A2(n_1099),
.B1(n_1096),
.B2(n_715),
.C(n_716),
.Y(n_1360)
);

INVx1_ASAP7_75t_L g1361 ( 
.A(n_1205),
.Y(n_1361)
);

INVx2_ASAP7_75t_L g1362 ( 
.A(n_1238),
.Y(n_1362)
);

BUFx2_ASAP7_75t_L g1363 ( 
.A(n_1245),
.Y(n_1363)
);

NAND2xp33_ASAP7_75t_L g1364 ( 
.A(n_1217),
.B(n_1072),
.Y(n_1364)
);

AND2x4_ASAP7_75t_L g1365 ( 
.A(n_1244),
.B(n_782),
.Y(n_1365)
);

HB1xp67_ASAP7_75t_L g1366 ( 
.A(n_1245),
.Y(n_1366)
);

INVx1_ASAP7_75t_L g1367 ( 
.A(n_1205),
.Y(n_1367)
);

NOR2xp67_ASAP7_75t_L g1368 ( 
.A(n_1342),
.B(n_1089),
.Y(n_1368)
);

BUFx6f_ASAP7_75t_L g1369 ( 
.A(n_1266),
.Y(n_1369)
);

INVx1_ASAP7_75t_L g1370 ( 
.A(n_1206),
.Y(n_1370)
);

CKINVDCx5p33_ASAP7_75t_R g1371 ( 
.A(n_1198),
.Y(n_1371)
);

NAND2xp5_ASAP7_75t_SL g1372 ( 
.A(n_1285),
.B(n_1286),
.Y(n_1372)
);

INVx2_ASAP7_75t_L g1373 ( 
.A(n_1197),
.Y(n_1373)
);

INVx2_ASAP7_75t_L g1374 ( 
.A(n_1200),
.Y(n_1374)
);

NOR2xp33_ASAP7_75t_L g1375 ( 
.A(n_1239),
.B(n_1089),
.Y(n_1375)
);

NOR2xp33_ASAP7_75t_L g1376 ( 
.A(n_1248),
.B(n_1092),
.Y(n_1376)
);

NAND2xp5_ASAP7_75t_L g1377 ( 
.A(n_1251),
.B(n_1092),
.Y(n_1377)
);

INVx2_ASAP7_75t_L g1378 ( 
.A(n_1347),
.Y(n_1378)
);

NOR2xp67_ASAP7_75t_L g1379 ( 
.A(n_1234),
.B(n_1097),
.Y(n_1379)
);

A2O1A1Ixp33_ASAP7_75t_L g1380 ( 
.A1(n_1288),
.A2(n_1034),
.B(n_1037),
.C(n_1007),
.Y(n_1380)
);

BUFx8_ASAP7_75t_L g1381 ( 
.A(n_1221),
.Y(n_1381)
);

NAND2xp5_ASAP7_75t_L g1382 ( 
.A(n_1293),
.B(n_1097),
.Y(n_1382)
);

INVx2_ASAP7_75t_L g1383 ( 
.A(n_1349),
.Y(n_1383)
);

INVx2_ASAP7_75t_L g1384 ( 
.A(n_1351),
.Y(n_1384)
);

NAND2xp5_ASAP7_75t_L g1385 ( 
.A(n_1298),
.B(n_815),
.Y(n_1385)
);

NAND2xp5_ASAP7_75t_SL g1386 ( 
.A(n_1266),
.B(n_831),
.Y(n_1386)
);

AOI22xp33_ASAP7_75t_L g1387 ( 
.A1(n_1312),
.A2(n_1037),
.B1(n_1039),
.B2(n_1034),
.Y(n_1387)
);

INVx1_ASAP7_75t_L g1388 ( 
.A(n_1206),
.Y(n_1388)
);

NAND2xp5_ASAP7_75t_L g1389 ( 
.A(n_1264),
.B(n_888),
.Y(n_1389)
);

AND2x2_ASAP7_75t_L g1390 ( 
.A(n_1249),
.B(n_732),
.Y(n_1390)
);

INVxp67_ASAP7_75t_SL g1391 ( 
.A(n_1249),
.Y(n_1391)
);

NAND2x1_ASAP7_75t_L g1392 ( 
.A(n_1217),
.B(n_756),
.Y(n_1392)
);

INVx2_ASAP7_75t_L g1393 ( 
.A(n_1353),
.Y(n_1393)
);

INVxp67_ASAP7_75t_L g1394 ( 
.A(n_1262),
.Y(n_1394)
);

NAND2xp33_ASAP7_75t_R g1395 ( 
.A(n_1247),
.B(n_703),
.Y(n_1395)
);

OAI22xp33_ASAP7_75t_L g1396 ( 
.A1(n_1244),
.A2(n_816),
.B1(n_830),
.B2(n_803),
.Y(n_1396)
);

INVx2_ASAP7_75t_L g1397 ( 
.A(n_1277),
.Y(n_1397)
);

NAND2xp5_ASAP7_75t_SL g1398 ( 
.A(n_1308),
.B(n_1088),
.Y(n_1398)
);

INVx2_ASAP7_75t_SL g1399 ( 
.A(n_1242),
.Y(n_1399)
);

NAND2xp5_ASAP7_75t_L g1400 ( 
.A(n_1274),
.B(n_1049),
.Y(n_1400)
);

NAND2xp5_ASAP7_75t_L g1401 ( 
.A(n_1274),
.B(n_703),
.Y(n_1401)
);

BUFx3_ASAP7_75t_L g1402 ( 
.A(n_1318),
.Y(n_1402)
);

NOR2xp33_ASAP7_75t_L g1403 ( 
.A(n_1302),
.B(n_946),
.Y(n_1403)
);

AOI22xp33_ASAP7_75t_L g1404 ( 
.A1(n_1335),
.A2(n_1067),
.B1(n_1039),
.B2(n_707),
.Y(n_1404)
);

NAND2xp5_ASAP7_75t_L g1405 ( 
.A(n_1294),
.B(n_704),
.Y(n_1405)
);

NAND2xp5_ASAP7_75t_L g1406 ( 
.A(n_1216),
.B(n_716),
.Y(n_1406)
);

BUFx6f_ASAP7_75t_SL g1407 ( 
.A(n_1244),
.Y(n_1407)
);

BUFx3_ASAP7_75t_L g1408 ( 
.A(n_1280),
.Y(n_1408)
);

NAND2xp5_ASAP7_75t_L g1409 ( 
.A(n_1216),
.B(n_728),
.Y(n_1409)
);

NAND2xp5_ASAP7_75t_SL g1410 ( 
.A(n_1302),
.B(n_1287),
.Y(n_1410)
);

OR2x2_ASAP7_75t_L g1411 ( 
.A(n_1207),
.B(n_728),
.Y(n_1411)
);

INVx1_ASAP7_75t_L g1412 ( 
.A(n_1230),
.Y(n_1412)
);

NOR2xp33_ASAP7_75t_L g1413 ( 
.A(n_1300),
.B(n_1021),
.Y(n_1413)
);

AND2x2_ASAP7_75t_L g1414 ( 
.A(n_1210),
.B(n_741),
.Y(n_1414)
);

BUFx6f_ASAP7_75t_SL g1415 ( 
.A(n_1344),
.Y(n_1415)
);

AOI22xp5_ASAP7_75t_L g1416 ( 
.A1(n_1255),
.A2(n_735),
.B1(n_738),
.B2(n_732),
.Y(n_1416)
);

NAND2xp5_ASAP7_75t_L g1417 ( 
.A(n_1352),
.B(n_1067),
.Y(n_1417)
);

AND2x2_ASAP7_75t_L g1418 ( 
.A(n_1246),
.B(n_757),
.Y(n_1418)
);

AND2x2_ASAP7_75t_L g1419 ( 
.A(n_1272),
.B(n_757),
.Y(n_1419)
);

NOR2xp33_ASAP7_75t_L g1420 ( 
.A(n_1303),
.B(n_709),
.Y(n_1420)
);

NAND2xp5_ASAP7_75t_L g1421 ( 
.A(n_1352),
.B(n_735),
.Y(n_1421)
);

NAND2xp5_ASAP7_75t_L g1422 ( 
.A(n_1199),
.B(n_738),
.Y(n_1422)
);

AOI22xp33_ASAP7_75t_L g1423 ( 
.A1(n_1336),
.A2(n_718),
.B1(n_720),
.B2(n_710),
.Y(n_1423)
);

AOI22xp5_ASAP7_75t_L g1424 ( 
.A1(n_1221),
.A2(n_741),
.B1(n_744),
.B2(n_740),
.Y(n_1424)
);

AND2x6_ASAP7_75t_L g1425 ( 
.A(n_1326),
.B(n_743),
.Y(n_1425)
);

INVx2_ASAP7_75t_L g1426 ( 
.A(n_1250),
.Y(n_1426)
);

NAND2xp5_ASAP7_75t_SL g1427 ( 
.A(n_1202),
.B(n_1214),
.Y(n_1427)
);

INVx2_ASAP7_75t_L g1428 ( 
.A(n_1253),
.Y(n_1428)
);

AO221x1_ASAP7_75t_L g1429 ( 
.A1(n_1284),
.A2(n_830),
.B1(n_890),
.B2(n_871),
.C(n_816),
.Y(n_1429)
);

NOR2xp33_ASAP7_75t_L g1430 ( 
.A(n_1232),
.B(n_1237),
.Y(n_1430)
);

NAND2xp5_ASAP7_75t_L g1431 ( 
.A(n_1272),
.B(n_740),
.Y(n_1431)
);

INVx2_ASAP7_75t_L g1432 ( 
.A(n_1254),
.Y(n_1432)
);

NAND2xp5_ASAP7_75t_L g1433 ( 
.A(n_1350),
.B(n_744),
.Y(n_1433)
);

BUFx6f_ASAP7_75t_L g1434 ( 
.A(n_1326),
.Y(n_1434)
);

NOR2xp33_ASAP7_75t_L g1435 ( 
.A(n_1232),
.B(n_711),
.Y(n_1435)
);

NAND2xp5_ASAP7_75t_L g1436 ( 
.A(n_1276),
.B(n_745),
.Y(n_1436)
);

NAND2xp5_ASAP7_75t_L g1437 ( 
.A(n_1276),
.B(n_745),
.Y(n_1437)
);

NAND2xp5_ASAP7_75t_L g1438 ( 
.A(n_1299),
.B(n_752),
.Y(n_1438)
);

NAND2xp5_ASAP7_75t_L g1439 ( 
.A(n_1299),
.B(n_752),
.Y(n_1439)
);

INVx1_ASAP7_75t_L g1440 ( 
.A(n_1201),
.Y(n_1440)
);

AOI22xp5_ASAP7_75t_L g1441 ( 
.A1(n_1355),
.A2(n_758),
.B1(n_761),
.B2(n_753),
.Y(n_1441)
);

INVx1_ASAP7_75t_L g1442 ( 
.A(n_1203),
.Y(n_1442)
);

INVx1_ASAP7_75t_L g1443 ( 
.A(n_1273),
.Y(n_1443)
);

INVx3_ASAP7_75t_R g1444 ( 
.A(n_1322),
.Y(n_1444)
);

AND2x2_ASAP7_75t_L g1445 ( 
.A(n_1348),
.B(n_1086),
.Y(n_1445)
);

OR2x2_ASAP7_75t_L g1446 ( 
.A(n_1284),
.B(n_1258),
.Y(n_1446)
);

INVx1_ASAP7_75t_L g1447 ( 
.A(n_1273),
.Y(n_1447)
);

NAND2xp5_ASAP7_75t_L g1448 ( 
.A(n_1357),
.B(n_753),
.Y(n_1448)
);

NOR2xp33_ASAP7_75t_L g1449 ( 
.A(n_1237),
.B(n_714),
.Y(n_1449)
);

AOI221xp5_ASAP7_75t_L g1450 ( 
.A1(n_1204),
.A2(n_1218),
.B1(n_1331),
.B2(n_1316),
.C(n_1220),
.Y(n_1450)
);

INVxp67_ASAP7_75t_L g1451 ( 
.A(n_1329),
.Y(n_1451)
);

NOR2xp33_ASAP7_75t_L g1452 ( 
.A(n_1243),
.B(n_719),
.Y(n_1452)
);

NAND2xp5_ASAP7_75t_L g1453 ( 
.A(n_1257),
.B(n_761),
.Y(n_1453)
);

BUFx2_ASAP7_75t_L g1454 ( 
.A(n_1235),
.Y(n_1454)
);

NAND2xp5_ASAP7_75t_L g1455 ( 
.A(n_1227),
.B(n_763),
.Y(n_1455)
);

NAND2xp5_ASAP7_75t_L g1456 ( 
.A(n_1260),
.B(n_763),
.Y(n_1456)
);

INVxp67_ASAP7_75t_L g1457 ( 
.A(n_1329),
.Y(n_1457)
);

NAND2xp5_ASAP7_75t_L g1458 ( 
.A(n_1267),
.B(n_764),
.Y(n_1458)
);

AND2x2_ASAP7_75t_L g1459 ( 
.A(n_1222),
.B(n_1259),
.Y(n_1459)
);

INVx1_ASAP7_75t_L g1460 ( 
.A(n_1252),
.Y(n_1460)
);

NAND2xp5_ASAP7_75t_L g1461 ( 
.A(n_1256),
.B(n_1271),
.Y(n_1461)
);

NAND2xp5_ASAP7_75t_L g1462 ( 
.A(n_1263),
.B(n_901),
.Y(n_1462)
);

NAND2xp5_ASAP7_75t_L g1463 ( 
.A(n_1283),
.B(n_1301),
.Y(n_1463)
);

OAI22xp5_ASAP7_75t_L g1464 ( 
.A1(n_1204),
.A2(n_890),
.B1(n_900),
.B2(n_871),
.Y(n_1464)
);

NOR2xp33_ASAP7_75t_L g1465 ( 
.A(n_1219),
.B(n_723),
.Y(n_1465)
);

NAND2xp5_ASAP7_75t_SL g1466 ( 
.A(n_1219),
.B(n_969),
.Y(n_1466)
);

NAND2xp5_ASAP7_75t_SL g1467 ( 
.A(n_1297),
.B(n_969),
.Y(n_1467)
);

OR2x2_ASAP7_75t_L g1468 ( 
.A(n_1218),
.B(n_908),
.Y(n_1468)
);

CKINVDCx20_ASAP7_75t_R g1469 ( 
.A(n_1354),
.Y(n_1469)
);

NOR2xp67_ASAP7_75t_L g1470 ( 
.A(n_1345),
.B(n_908),
.Y(n_1470)
);

INVx1_ASAP7_75t_L g1471 ( 
.A(n_1315),
.Y(n_1471)
);

NOR3xp33_ASAP7_75t_L g1472 ( 
.A(n_1331),
.B(n_1002),
.C(n_861),
.Y(n_1472)
);

INVx2_ASAP7_75t_SL g1473 ( 
.A(n_1280),
.Y(n_1473)
);

NAND2xp5_ASAP7_75t_L g1474 ( 
.A(n_1261),
.B(n_913),
.Y(n_1474)
);

NOR2xp33_ASAP7_75t_L g1475 ( 
.A(n_1309),
.B(n_1247),
.Y(n_1475)
);

AO221x1_ASAP7_75t_L g1476 ( 
.A1(n_1344),
.A2(n_926),
.B1(n_983),
.B2(n_920),
.C(n_900),
.Y(n_1476)
);

AOI22xp33_ASAP7_75t_L g1477 ( 
.A1(n_1355),
.A2(n_727),
.B1(n_731),
.B2(n_730),
.Y(n_1477)
);

BUFx8_ASAP7_75t_L g1478 ( 
.A(n_1344),
.Y(n_1478)
);

INVxp67_ASAP7_75t_SL g1479 ( 
.A(n_1261),
.Y(n_1479)
);

INVx1_ASAP7_75t_L g1480 ( 
.A(n_1315),
.Y(n_1480)
);

INVx1_ASAP7_75t_L g1481 ( 
.A(n_1317),
.Y(n_1481)
);

NAND2xp5_ASAP7_75t_L g1482 ( 
.A(n_1224),
.B(n_913),
.Y(n_1482)
);

NOR2xp33_ASAP7_75t_L g1483 ( 
.A(n_1309),
.B(n_769),
.Y(n_1483)
);

OR2x6_ASAP7_75t_L g1484 ( 
.A(n_1346),
.B(n_1344),
.Y(n_1484)
);

BUFx5_ASAP7_75t_L g1485 ( 
.A(n_1339),
.Y(n_1485)
);

NAND2xp5_ASAP7_75t_L g1486 ( 
.A(n_1268),
.B(n_916),
.Y(n_1486)
);

AOI22xp33_ASAP7_75t_L g1487 ( 
.A1(n_1209),
.A2(n_733),
.B1(n_746),
.B2(n_737),
.Y(n_1487)
);

NAND2xp5_ASAP7_75t_L g1488 ( 
.A(n_1224),
.B(n_916),
.Y(n_1488)
);

INVxp67_ASAP7_75t_L g1489 ( 
.A(n_1314),
.Y(n_1489)
);

INVx1_ASAP7_75t_L g1490 ( 
.A(n_1228),
.Y(n_1490)
);

NOR2xp67_ASAP7_75t_L g1491 ( 
.A(n_1354),
.B(n_1069),
.Y(n_1491)
);

INVxp67_ASAP7_75t_L g1492 ( 
.A(n_1323),
.Y(n_1492)
);

BUFx3_ASAP7_75t_L g1493 ( 
.A(n_1356),
.Y(n_1493)
);

BUFx6f_ASAP7_75t_L g1494 ( 
.A(n_1307),
.Y(n_1494)
);

NAND2xp5_ASAP7_75t_L g1495 ( 
.A(n_1268),
.B(n_1069),
.Y(n_1495)
);

NOR2xp33_ASAP7_75t_L g1496 ( 
.A(n_1356),
.B(n_772),
.Y(n_1496)
);

NOR2xp67_ASAP7_75t_L g1497 ( 
.A(n_1343),
.B(n_1070),
.Y(n_1497)
);

NAND2xp5_ASAP7_75t_L g1498 ( 
.A(n_1278),
.B(n_1070),
.Y(n_1498)
);

INVx2_ASAP7_75t_SL g1499 ( 
.A(n_1235),
.Y(n_1499)
);

INVx2_ASAP7_75t_L g1500 ( 
.A(n_1333),
.Y(n_1500)
);

NAND2xp5_ASAP7_75t_L g1501 ( 
.A(n_1278),
.B(n_1071),
.Y(n_1501)
);

NAND2xp5_ASAP7_75t_SL g1502 ( 
.A(n_1305),
.B(n_770),
.Y(n_1502)
);

NAND2xp5_ASAP7_75t_L g1503 ( 
.A(n_1270),
.B(n_1071),
.Y(n_1503)
);

INVxp33_ASAP7_75t_L g1504 ( 
.A(n_1343),
.Y(n_1504)
);

AND2x2_ASAP7_75t_L g1505 ( 
.A(n_1337),
.B(n_1079),
.Y(n_1505)
);

NOR2xp33_ASAP7_75t_L g1506 ( 
.A(n_1270),
.B(n_777),
.Y(n_1506)
);

NAND2xp5_ASAP7_75t_L g1507 ( 
.A(n_1209),
.B(n_1073),
.Y(n_1507)
);

INVx2_ASAP7_75t_L g1508 ( 
.A(n_1333),
.Y(n_1508)
);

NAND2xp5_ASAP7_75t_SL g1509 ( 
.A(n_1305),
.B(n_785),
.Y(n_1509)
);

OR2x2_ASAP7_75t_L g1510 ( 
.A(n_1316),
.B(n_1073),
.Y(n_1510)
);

INVx2_ASAP7_75t_L g1511 ( 
.A(n_1338),
.Y(n_1511)
);

NAND2xp5_ASAP7_75t_L g1512 ( 
.A(n_1275),
.B(n_1074),
.Y(n_1512)
);

INVx1_ASAP7_75t_L g1513 ( 
.A(n_1310),
.Y(n_1513)
);

NAND2xp5_ASAP7_75t_L g1514 ( 
.A(n_1279),
.B(n_1074),
.Y(n_1514)
);

NAND2xp5_ASAP7_75t_L g1515 ( 
.A(n_1281),
.B(n_1078),
.Y(n_1515)
);

NOR2xp33_ASAP7_75t_L g1516 ( 
.A(n_1281),
.B(n_778),
.Y(n_1516)
);

NOR3xp33_ASAP7_75t_L g1517 ( 
.A(n_1332),
.B(n_929),
.C(n_713),
.Y(n_1517)
);

NAND2xp5_ASAP7_75t_L g1518 ( 
.A(n_1233),
.B(n_1289),
.Y(n_1518)
);

NAND2xp5_ASAP7_75t_L g1519 ( 
.A(n_1233),
.B(n_1078),
.Y(n_1519)
);

NAND2xp5_ASAP7_75t_L g1520 ( 
.A(n_1313),
.B(n_1079),
.Y(n_1520)
);

NOR2xp33_ASAP7_75t_L g1521 ( 
.A(n_1226),
.B(n_779),
.Y(n_1521)
);

HB1xp67_ASAP7_75t_L g1522 ( 
.A(n_1332),
.Y(n_1522)
);

NAND2xp5_ASAP7_75t_L g1523 ( 
.A(n_1313),
.B(n_1081),
.Y(n_1523)
);

NAND2xp5_ASAP7_75t_L g1524 ( 
.A(n_1320),
.B(n_1081),
.Y(n_1524)
);

BUFx6f_ASAP7_75t_SL g1525 ( 
.A(n_1337),
.Y(n_1525)
);

AND2x4_ASAP7_75t_L g1526 ( 
.A(n_1291),
.B(n_751),
.Y(n_1526)
);

NOR2xp33_ASAP7_75t_L g1527 ( 
.A(n_1226),
.B(n_783),
.Y(n_1527)
);

AOI22xp5_ASAP7_75t_L g1528 ( 
.A1(n_1292),
.A2(n_1090),
.B1(n_1094),
.B2(n_1086),
.Y(n_1528)
);

OAI22xp5_ASAP7_75t_L g1529 ( 
.A1(n_1292),
.A2(n_926),
.B1(n_983),
.B2(n_920),
.Y(n_1529)
);

NAND2xp5_ASAP7_75t_L g1530 ( 
.A(n_1289),
.B(n_1324),
.Y(n_1530)
);

INVx2_ASAP7_75t_L g1531 ( 
.A(n_1225),
.Y(n_1531)
);

NOR2xp67_ASAP7_75t_L g1532 ( 
.A(n_1324),
.B(n_1094),
.Y(n_1532)
);

AOI221xp5_ASAP7_75t_L g1533 ( 
.A1(n_1328),
.A2(n_1096),
.B1(n_774),
.B2(n_787),
.C(n_771),
.Y(n_1533)
);

INVx1_ASAP7_75t_L g1534 ( 
.A(n_1320),
.Y(n_1534)
);

INVx1_ASAP7_75t_L g1535 ( 
.A(n_1328),
.Y(n_1535)
);

AND2x2_ASAP7_75t_L g1536 ( 
.A(n_1226),
.B(n_784),
.Y(n_1536)
);

NAND2xp5_ASAP7_75t_L g1537 ( 
.A(n_1208),
.B(n_788),
.Y(n_1537)
);

INVx1_ASAP7_75t_L g1538 ( 
.A(n_1215),
.Y(n_1538)
);

NAND2xp5_ASAP7_75t_L g1539 ( 
.A(n_1212),
.B(n_791),
.Y(n_1539)
);

NAND2xp5_ASAP7_75t_L g1540 ( 
.A(n_1213),
.B(n_793),
.Y(n_1540)
);

INVx2_ASAP7_75t_L g1541 ( 
.A(n_1223),
.Y(n_1541)
);

INVx1_ASAP7_75t_L g1542 ( 
.A(n_1334),
.Y(n_1542)
);

NAND2xp5_ASAP7_75t_L g1543 ( 
.A(n_1229),
.B(n_795),
.Y(n_1543)
);

AOI22xp5_ASAP7_75t_L g1544 ( 
.A1(n_1231),
.A2(n_802),
.B1(n_804),
.B2(n_796),
.Y(n_1544)
);

NAND2xp5_ASAP7_75t_L g1545 ( 
.A(n_1334),
.B(n_805),
.Y(n_1545)
);

INVx1_ASAP7_75t_L g1546 ( 
.A(n_1340),
.Y(n_1546)
);

INVx2_ASAP7_75t_L g1547 ( 
.A(n_1330),
.Y(n_1547)
);

INVx1_ASAP7_75t_L g1548 ( 
.A(n_1231),
.Y(n_1548)
);

BUFx5_ASAP7_75t_L g1549 ( 
.A(n_1304),
.Y(n_1549)
);

NOR2xp33_ASAP7_75t_L g1550 ( 
.A(n_1231),
.B(n_808),
.Y(n_1550)
);

NOR2xp33_ASAP7_75t_L g1551 ( 
.A(n_1304),
.B(n_813),
.Y(n_1551)
);

NAND2xp33_ASAP7_75t_SL g1552 ( 
.A(n_1346),
.B(n_1093),
.Y(n_1552)
);

INVx2_ASAP7_75t_L g1553 ( 
.A(n_1282),
.Y(n_1553)
);

NAND2xp5_ASAP7_75t_L g1554 ( 
.A(n_1325),
.B(n_814),
.Y(n_1554)
);

INVx1_ASAP7_75t_L g1555 ( 
.A(n_1290),
.Y(n_1555)
);

NOR2xp33_ASAP7_75t_SL g1556 ( 
.A(n_1346),
.B(n_847),
.Y(n_1556)
);

NAND2xp5_ASAP7_75t_L g1557 ( 
.A(n_1325),
.B(n_819),
.Y(n_1557)
);

NOR2xp33_ASAP7_75t_L g1558 ( 
.A(n_1295),
.B(n_822),
.Y(n_1558)
);

NAND2xp5_ASAP7_75t_SL g1559 ( 
.A(n_1211),
.B(n_790),
.Y(n_1559)
);

AOI22xp5_ASAP7_75t_L g1560 ( 
.A1(n_1306),
.A2(n_827),
.B1(n_829),
.B2(n_823),
.Y(n_1560)
);

NAND3xp33_ASAP7_75t_L g1561 ( 
.A(n_1211),
.B(n_789),
.C(n_754),
.Y(n_1561)
);

NOR2xp33_ASAP7_75t_L g1562 ( 
.A(n_1311),
.B(n_833),
.Y(n_1562)
);

INVx2_ASAP7_75t_L g1563 ( 
.A(n_1319),
.Y(n_1563)
);

INVx1_ASAP7_75t_L g1564 ( 
.A(n_1321),
.Y(n_1564)
);

NOR2xp33_ASAP7_75t_L g1565 ( 
.A(n_1240),
.B(n_838),
.Y(n_1565)
);

OAI22xp5_ASAP7_75t_L g1566 ( 
.A1(n_1327),
.A2(n_1050),
.B1(n_1093),
.B2(n_1005),
.Y(n_1566)
);

NOR2xp33_ASAP7_75t_L g1567 ( 
.A(n_1240),
.B(n_840),
.Y(n_1567)
);

NOR2xp33_ASAP7_75t_L g1568 ( 
.A(n_1241),
.B(n_842),
.Y(n_1568)
);

OR2x6_ASAP7_75t_L g1569 ( 
.A(n_1241),
.B(n_849),
.Y(n_1569)
);

NOR2xp33_ASAP7_75t_L g1570 ( 
.A(n_1241),
.B(n_843),
.Y(n_1570)
);

BUFx3_ASAP7_75t_L g1571 ( 
.A(n_1241),
.Y(n_1571)
);

BUFx6f_ASAP7_75t_SL g1572 ( 
.A(n_1265),
.Y(n_1572)
);

NAND2xp5_ASAP7_75t_L g1573 ( 
.A(n_1482),
.B(n_853),
.Y(n_1573)
);

NAND2xp5_ASAP7_75t_SL g1574 ( 
.A(n_1363),
.B(n_854),
.Y(n_1574)
);

O2A1O1Ixp33_ASAP7_75t_L g1575 ( 
.A1(n_1446),
.A2(n_801),
.B(n_806),
.C(n_794),
.Y(n_1575)
);

AO21x1_ASAP7_75t_L g1576 ( 
.A1(n_1530),
.A2(n_811),
.B(n_809),
.Y(n_1576)
);

AND2x2_ASAP7_75t_L g1577 ( 
.A(n_1451),
.B(n_1005),
.Y(n_1577)
);

HB1xp67_ASAP7_75t_L g1578 ( 
.A(n_1457),
.Y(n_1578)
);

NAND2xp5_ASAP7_75t_L g1579 ( 
.A(n_1482),
.B(n_855),
.Y(n_1579)
);

BUFx2_ASAP7_75t_L g1580 ( 
.A(n_1391),
.Y(n_1580)
);

NAND2xp5_ASAP7_75t_L g1581 ( 
.A(n_1488),
.B(n_857),
.Y(n_1581)
);

NAND2xp5_ASAP7_75t_L g1582 ( 
.A(n_1488),
.B(n_858),
.Y(n_1582)
);

O2A1O1Ixp33_ASAP7_75t_L g1583 ( 
.A1(n_1411),
.A2(n_825),
.B(n_826),
.C(n_818),
.Y(n_1583)
);

NOR2x1_ASAP7_75t_L g1584 ( 
.A(n_1408),
.B(n_1050),
.Y(n_1584)
);

AOI22xp5_ASAP7_75t_L g1585 ( 
.A1(n_1366),
.A2(n_860),
.B1(n_864),
.B2(n_859),
.Y(n_1585)
);

AOI21xp5_ASAP7_75t_L g1586 ( 
.A1(n_1534),
.A2(n_834),
.B(n_828),
.Y(n_1586)
);

INVx1_ASAP7_75t_L g1587 ( 
.A(n_1443),
.Y(n_1587)
);

AOI21xp5_ASAP7_75t_L g1588 ( 
.A1(n_1542),
.A2(n_836),
.B(n_835),
.Y(n_1588)
);

OAI22xp5_ASAP7_75t_L g1589 ( 
.A1(n_1358),
.A2(n_1394),
.B1(n_1487),
.B2(n_1409),
.Y(n_1589)
);

NAND2xp5_ASAP7_75t_L g1590 ( 
.A(n_1463),
.B(n_868),
.Y(n_1590)
);

AOI21xp5_ASAP7_75t_L g1591 ( 
.A1(n_1520),
.A2(n_844),
.B(n_841),
.Y(n_1591)
);

AOI21xp5_ASAP7_75t_L g1592 ( 
.A1(n_1520),
.A2(n_850),
.B(n_848),
.Y(n_1592)
);

AND2x2_ASAP7_75t_SL g1593 ( 
.A(n_1454),
.B(n_862),
.Y(n_1593)
);

HB1xp67_ASAP7_75t_L g1594 ( 
.A(n_1402),
.Y(n_1594)
);

NAND2xp5_ASAP7_75t_L g1595 ( 
.A(n_1406),
.B(n_869),
.Y(n_1595)
);

NAND2xp5_ASAP7_75t_L g1596 ( 
.A(n_1375),
.B(n_885),
.Y(n_1596)
);

AOI22xp5_ASAP7_75t_L g1597 ( 
.A1(n_1418),
.A2(n_893),
.B1(n_894),
.B2(n_892),
.Y(n_1597)
);

AOI21xp5_ASAP7_75t_L g1598 ( 
.A1(n_1523),
.A2(n_852),
.B(n_851),
.Y(n_1598)
);

NAND2xp5_ASAP7_75t_L g1599 ( 
.A(n_1376),
.B(n_898),
.Y(n_1599)
);

BUFx4f_ASAP7_75t_L g1600 ( 
.A(n_1484),
.Y(n_1600)
);

OR2x6_ASAP7_75t_L g1601 ( 
.A(n_1484),
.B(n_862),
.Y(n_1601)
);

INVx2_ASAP7_75t_L g1602 ( 
.A(n_1546),
.Y(n_1602)
);

OAI21xp5_ASAP7_75t_L g1603 ( 
.A1(n_1531),
.A2(n_863),
.B(n_856),
.Y(n_1603)
);

NAND2xp5_ASAP7_75t_L g1604 ( 
.A(n_1390),
.B(n_899),
.Y(n_1604)
);

INVx1_ASAP7_75t_L g1605 ( 
.A(n_1447),
.Y(n_1605)
);

NAND2xp5_ASAP7_75t_L g1606 ( 
.A(n_1377),
.B(n_919),
.Y(n_1606)
);

AOI21xp5_ASAP7_75t_L g1607 ( 
.A1(n_1523),
.A2(n_866),
.B(n_865),
.Y(n_1607)
);

AOI21x1_ASAP7_75t_L g1608 ( 
.A1(n_1502),
.A2(n_1509),
.B(n_1372),
.Y(n_1608)
);

OAI22xp5_ASAP7_75t_L g1609 ( 
.A1(n_1422),
.A2(n_872),
.B1(n_878),
.B2(n_876),
.Y(n_1609)
);

NAND2xp5_ASAP7_75t_L g1610 ( 
.A(n_1382),
.B(n_921),
.Y(n_1610)
);

INVx1_ASAP7_75t_L g1611 ( 
.A(n_1417),
.Y(n_1611)
);

AOI21xp5_ASAP7_75t_L g1612 ( 
.A1(n_1524),
.A2(n_880),
.B(n_879),
.Y(n_1612)
);

OR2x2_ASAP7_75t_L g1613 ( 
.A(n_1566),
.B(n_991),
.Y(n_1613)
);

O2A1O1Ixp33_ASAP7_75t_L g1614 ( 
.A1(n_1431),
.A2(n_1437),
.B(n_1436),
.C(n_1529),
.Y(n_1614)
);

INVx2_ASAP7_75t_SL g1615 ( 
.A(n_1493),
.Y(n_1615)
);

NAND2xp5_ASAP7_75t_L g1616 ( 
.A(n_1419),
.B(n_930),
.Y(n_1616)
);

OAI21x1_ASAP7_75t_L g1617 ( 
.A1(n_1392),
.A2(n_889),
.B(n_870),
.Y(n_1617)
);

A2O1A1Ixp33_ASAP7_75t_L g1618 ( 
.A1(n_1460),
.A2(n_891),
.B(n_895),
.C(n_884),
.Y(n_1618)
);

INVx1_ASAP7_75t_SL g1619 ( 
.A(n_1425),
.Y(n_1619)
);

INVx1_ASAP7_75t_SL g1620 ( 
.A(n_1425),
.Y(n_1620)
);

AOI21xp5_ASAP7_75t_L g1621 ( 
.A1(n_1524),
.A2(n_905),
.B(n_904),
.Y(n_1621)
);

NAND2xp5_ASAP7_75t_L g1622 ( 
.A(n_1422),
.B(n_931),
.Y(n_1622)
);

INVx2_ASAP7_75t_L g1623 ( 
.A(n_1485),
.Y(n_1623)
);

INVx1_ASAP7_75t_L g1624 ( 
.A(n_1417),
.Y(n_1624)
);

AOI21xp5_ASAP7_75t_L g1625 ( 
.A1(n_1545),
.A2(n_909),
.B(n_906),
.Y(n_1625)
);

NAND2xp5_ASAP7_75t_L g1626 ( 
.A(n_1433),
.B(n_934),
.Y(n_1626)
);

AOI21xp5_ASAP7_75t_L g1627 ( 
.A1(n_1427),
.A2(n_917),
.B(n_914),
.Y(n_1627)
);

AND2x6_ASAP7_75t_SL g1628 ( 
.A(n_1484),
.B(n_923),
.Y(n_1628)
);

AOI21xp5_ASAP7_75t_L g1629 ( 
.A1(n_1479),
.A2(n_925),
.B(n_924),
.Y(n_1629)
);

AOI21xp5_ASAP7_75t_L g1630 ( 
.A1(n_1385),
.A2(n_932),
.B(n_927),
.Y(n_1630)
);

AOI21xp5_ASAP7_75t_L g1631 ( 
.A1(n_1519),
.A2(n_1461),
.B(n_1507),
.Y(n_1631)
);

AOI21xp5_ASAP7_75t_L g1632 ( 
.A1(n_1461),
.A2(n_936),
.B(n_933),
.Y(n_1632)
);

NAND2xp5_ASAP7_75t_L g1633 ( 
.A(n_1433),
.B(n_937),
.Y(n_1633)
);

BUFx2_ASAP7_75t_L g1634 ( 
.A(n_1469),
.Y(n_1634)
);

AND2x2_ASAP7_75t_L g1635 ( 
.A(n_1414),
.B(n_1044),
.Y(n_1635)
);

NAND2xp5_ASAP7_75t_L g1636 ( 
.A(n_1448),
.B(n_939),
.Y(n_1636)
);

NAND2xp33_ASAP7_75t_L g1637 ( 
.A(n_1425),
.B(n_942),
.Y(n_1637)
);

OAI21xp5_ASAP7_75t_L g1638 ( 
.A1(n_1380),
.A2(n_943),
.B(n_941),
.Y(n_1638)
);

AOI21xp5_ASAP7_75t_L g1639 ( 
.A1(n_1507),
.A2(n_948),
.B(n_944),
.Y(n_1639)
);

NOR3xp33_ASAP7_75t_L g1640 ( 
.A(n_1396),
.B(n_1057),
.C(n_949),
.Y(n_1640)
);

NAND2xp5_ASAP7_75t_L g1641 ( 
.A(n_1448),
.B(n_945),
.Y(n_1641)
);

AOI21xp33_ASAP7_75t_L g1642 ( 
.A1(n_1504),
.A2(n_951),
.B(n_950),
.Y(n_1642)
);

BUFx6f_ASAP7_75t_L g1643 ( 
.A(n_1434),
.Y(n_1643)
);

INVx1_ASAP7_75t_L g1644 ( 
.A(n_1440),
.Y(n_1644)
);

AND2x2_ASAP7_75t_L g1645 ( 
.A(n_1445),
.B(n_952),
.Y(n_1645)
);

BUFx8_ASAP7_75t_L g1646 ( 
.A(n_1407),
.Y(n_1646)
);

INVx6_ASAP7_75t_L g1647 ( 
.A(n_1381),
.Y(n_1647)
);

BUFx12f_ASAP7_75t_L g1648 ( 
.A(n_1381),
.Y(n_1648)
);

NAND2xp5_ASAP7_75t_SL g1649 ( 
.A(n_1494),
.B(n_953),
.Y(n_1649)
);

BUFx6f_ASAP7_75t_L g1650 ( 
.A(n_1434),
.Y(n_1650)
);

NAND2x1p5_ASAP7_75t_L g1651 ( 
.A(n_1473),
.B(n_896),
.Y(n_1651)
);

INVx2_ASAP7_75t_SL g1652 ( 
.A(n_1505),
.Y(n_1652)
);

AO21x1_ASAP7_75t_L g1653 ( 
.A1(n_1400),
.A2(n_955),
.B(n_954),
.Y(n_1653)
);

AOI21xp5_ASAP7_75t_L g1654 ( 
.A1(n_1513),
.A2(n_960),
.B(n_959),
.Y(n_1654)
);

INVx1_ASAP7_75t_L g1655 ( 
.A(n_1442),
.Y(n_1655)
);

A2O1A1Ixp33_ASAP7_75t_L g1656 ( 
.A1(n_1471),
.A2(n_965),
.B(n_968),
.C(n_963),
.Y(n_1656)
);

HB1xp67_ASAP7_75t_L g1657 ( 
.A(n_1566),
.Y(n_1657)
);

NAND2xp5_ASAP7_75t_L g1658 ( 
.A(n_1438),
.B(n_956),
.Y(n_1658)
);

A2O1A1Ixp33_ASAP7_75t_L g1659 ( 
.A1(n_1480),
.A2(n_975),
.B(n_985),
.C(n_973),
.Y(n_1659)
);

OAI21xp5_ASAP7_75t_L g1660 ( 
.A1(n_1500),
.A2(n_989),
.B(n_986),
.Y(n_1660)
);

INVx2_ASAP7_75t_SL g1661 ( 
.A(n_1459),
.Y(n_1661)
);

OAI22xp5_ASAP7_75t_L g1662 ( 
.A1(n_1489),
.A2(n_997),
.B1(n_998),
.B2(n_995),
.Y(n_1662)
);

BUFx4f_ASAP7_75t_L g1663 ( 
.A(n_1365),
.Y(n_1663)
);

OAI21xp5_ASAP7_75t_L g1664 ( 
.A1(n_1508),
.A2(n_1011),
.B(n_1004),
.Y(n_1664)
);

AOI21xp5_ASAP7_75t_L g1665 ( 
.A1(n_1421),
.A2(n_1015),
.B(n_1012),
.Y(n_1665)
);

A2O1A1Ixp33_ASAP7_75t_L g1666 ( 
.A1(n_1481),
.A2(n_1020),
.B(n_1035),
.C(n_1017),
.Y(n_1666)
);

OAI21xp5_ASAP7_75t_L g1667 ( 
.A1(n_1511),
.A2(n_1038),
.B(n_1036),
.Y(n_1667)
);

OR2x2_ASAP7_75t_L g1668 ( 
.A(n_1468),
.B(n_958),
.Y(n_1668)
);

BUFx6f_ASAP7_75t_L g1669 ( 
.A(n_1434),
.Y(n_1669)
);

AOI21xp5_ASAP7_75t_L g1670 ( 
.A1(n_1538),
.A2(n_1047),
.B(n_1041),
.Y(n_1670)
);

O2A1O1Ixp33_ASAP7_75t_L g1671 ( 
.A1(n_1529),
.A2(n_1051),
.B(n_1052),
.C(n_1048),
.Y(n_1671)
);

NAND2xp5_ASAP7_75t_L g1672 ( 
.A(n_1439),
.B(n_961),
.Y(n_1672)
);

NOR2xp67_ASAP7_75t_L g1673 ( 
.A(n_1499),
.B(n_30),
.Y(n_1673)
);

INVxp67_ASAP7_75t_L g1674 ( 
.A(n_1395),
.Y(n_1674)
);

AOI22xp33_ASAP7_75t_L g1675 ( 
.A1(n_1450),
.A2(n_1059),
.B1(n_1075),
.B2(n_1058),
.Y(n_1675)
);

NAND2xp5_ASAP7_75t_L g1676 ( 
.A(n_1401),
.B(n_964),
.Y(n_1676)
);

NOR2xp33_ASAP7_75t_L g1677 ( 
.A(n_1399),
.B(n_971),
.Y(n_1677)
);

NOR2xp67_ASAP7_75t_L g1678 ( 
.A(n_1371),
.B(n_1528),
.Y(n_1678)
);

AOI21xp5_ASAP7_75t_L g1679 ( 
.A1(n_1410),
.A2(n_1076),
.B(n_1077),
.Y(n_1679)
);

NAND2xp5_ASAP7_75t_L g1680 ( 
.A(n_1486),
.B(n_970),
.Y(n_1680)
);

INVx1_ASAP7_75t_L g1681 ( 
.A(n_1412),
.Y(n_1681)
);

O2A1O1Ixp33_ASAP7_75t_L g1682 ( 
.A1(n_1405),
.A2(n_1085),
.B(n_1087),
.C(n_1080),
.Y(n_1682)
);

NAND2xp5_ASAP7_75t_L g1683 ( 
.A(n_1495),
.B(n_972),
.Y(n_1683)
);

AOI21xp5_ASAP7_75t_L g1684 ( 
.A1(n_1455),
.A2(n_910),
.B(n_903),
.Y(n_1684)
);

AOI21xp5_ASAP7_75t_L g1685 ( 
.A1(n_1455),
.A2(n_910),
.B(n_903),
.Y(n_1685)
);

BUFx6f_ASAP7_75t_L g1686 ( 
.A(n_1369),
.Y(n_1686)
);

CKINVDCx5p33_ASAP7_75t_R g1687 ( 
.A(n_1525),
.Y(n_1687)
);

OAI21xp33_ASAP7_75t_L g1688 ( 
.A1(n_1465),
.A2(n_1060),
.B(n_1056),
.Y(n_1688)
);

BUFx2_ASAP7_75t_SL g1689 ( 
.A(n_1407),
.Y(n_1689)
);

BUFx2_ASAP7_75t_L g1690 ( 
.A(n_1478),
.Y(n_1690)
);

BUFx6f_ASAP7_75t_L g1691 ( 
.A(n_1369),
.Y(n_1691)
);

NAND2xp5_ASAP7_75t_SL g1692 ( 
.A(n_1491),
.B(n_974),
.Y(n_1692)
);

OAI21x1_ASAP7_75t_L g1693 ( 
.A1(n_1467),
.A2(n_980),
.B(n_967),
.Y(n_1693)
);

INVxp67_ASAP7_75t_L g1694 ( 
.A(n_1474),
.Y(n_1694)
);

AOI22xp5_ASAP7_75t_L g1695 ( 
.A1(n_1492),
.A2(n_979),
.B1(n_981),
.B2(n_978),
.Y(n_1695)
);

AND2x4_ASAP7_75t_L g1696 ( 
.A(n_1497),
.B(n_1018),
.Y(n_1696)
);

INVx4_ASAP7_75t_L g1697 ( 
.A(n_1525),
.Y(n_1697)
);

AOI22xp5_ASAP7_75t_L g1698 ( 
.A1(n_1475),
.A2(n_988),
.B1(n_990),
.B2(n_984),
.Y(n_1698)
);

OAI21xp33_ASAP7_75t_L g1699 ( 
.A1(n_1416),
.A2(n_996),
.B(n_992),
.Y(n_1699)
);

NAND2xp5_ASAP7_75t_L g1700 ( 
.A(n_1403),
.B(n_999),
.Y(n_1700)
);

NOR2xp33_ASAP7_75t_L g1701 ( 
.A(n_1483),
.B(n_1000),
.Y(n_1701)
);

AOI21xp5_ASAP7_75t_L g1702 ( 
.A1(n_1364),
.A2(n_1095),
.B(n_1055),
.Y(n_1702)
);

AOI21xp5_ASAP7_75t_L g1703 ( 
.A1(n_1535),
.A2(n_1456),
.B(n_1453),
.Y(n_1703)
);

AND2x4_ASAP7_75t_L g1704 ( 
.A(n_1526),
.B(n_1095),
.Y(n_1704)
);

AND2x2_ASAP7_75t_L g1705 ( 
.A(n_1510),
.B(n_1001),
.Y(n_1705)
);

AOI21xp5_ASAP7_75t_L g1706 ( 
.A1(n_1458),
.A2(n_1269),
.B(n_1265),
.Y(n_1706)
);

BUFx6f_ASAP7_75t_L g1707 ( 
.A(n_1425),
.Y(n_1707)
);

AND2x2_ASAP7_75t_L g1708 ( 
.A(n_1496),
.B(n_1360),
.Y(n_1708)
);

AOI22xp5_ASAP7_75t_L g1709 ( 
.A1(n_1526),
.A2(n_1008),
.B1(n_1009),
.B2(n_1006),
.Y(n_1709)
);

NAND2xp5_ASAP7_75t_L g1710 ( 
.A(n_1389),
.B(n_1010),
.Y(n_1710)
);

INVx2_ASAP7_75t_SL g1711 ( 
.A(n_1365),
.Y(n_1711)
);

AND2x2_ASAP7_75t_SL g1712 ( 
.A(n_1472),
.B(n_31),
.Y(n_1712)
);

AND2x2_ASAP7_75t_L g1713 ( 
.A(n_1441),
.B(n_1013),
.Y(n_1713)
);

NAND2xp5_ASAP7_75t_L g1714 ( 
.A(n_1477),
.B(n_1016),
.Y(n_1714)
);

BUFx2_ASAP7_75t_L g1715 ( 
.A(n_1478),
.Y(n_1715)
);

NAND2x1_ASAP7_75t_L g1716 ( 
.A(n_1569),
.B(n_1269),
.Y(n_1716)
);

INVx2_ASAP7_75t_L g1717 ( 
.A(n_1426),
.Y(n_1717)
);

AO21x1_ASAP7_75t_L g1718 ( 
.A1(n_1430),
.A2(n_31),
.B(n_32),
.Y(n_1718)
);

AOI22xp5_ASAP7_75t_L g1719 ( 
.A1(n_1466),
.A2(n_1022),
.B1(n_1023),
.B2(n_1019),
.Y(n_1719)
);

NAND2xp5_ASAP7_75t_L g1720 ( 
.A(n_1423),
.B(n_1025),
.Y(n_1720)
);

NOR2xp33_ASAP7_75t_L g1721 ( 
.A(n_1398),
.B(n_1027),
.Y(n_1721)
);

AO21x1_ASAP7_75t_L g1722 ( 
.A1(n_1559),
.A2(n_32),
.B(n_33),
.Y(n_1722)
);

NAND2xp5_ASAP7_75t_L g1723 ( 
.A(n_1361),
.B(n_1028),
.Y(n_1723)
);

BUFx12f_ASAP7_75t_L g1724 ( 
.A(n_1536),
.Y(n_1724)
);

NAND2xp5_ASAP7_75t_L g1725 ( 
.A(n_1367),
.B(n_1030),
.Y(n_1725)
);

NAND2xp5_ASAP7_75t_L g1726 ( 
.A(n_1370),
.B(n_1033),
.Y(n_1726)
);

BUFx2_ASAP7_75t_L g1727 ( 
.A(n_1552),
.Y(n_1727)
);

O2A1O1Ixp33_ASAP7_75t_L g1728 ( 
.A1(n_1462),
.A2(n_1045),
.B(n_1046),
.C(n_1043),
.Y(n_1728)
);

NAND2xp5_ASAP7_75t_L g1729 ( 
.A(n_1388),
.B(n_1054),
.Y(n_1729)
);

AOI21xp5_ASAP7_75t_L g1730 ( 
.A1(n_1386),
.A2(n_1296),
.B(n_1062),
.Y(n_1730)
);

NOR2xp33_ASAP7_75t_L g1731 ( 
.A(n_1548),
.B(n_1061),
.Y(n_1731)
);

AOI22xp5_ASAP7_75t_L g1732 ( 
.A1(n_1413),
.A2(n_1065),
.B1(n_1066),
.B2(n_1064),
.Y(n_1732)
);

AND2x2_ASAP7_75t_L g1733 ( 
.A(n_1424),
.B(n_33),
.Y(n_1733)
);

BUFx6f_ASAP7_75t_L g1734 ( 
.A(n_1569),
.Y(n_1734)
);

NAND2xp5_ASAP7_75t_SL g1735 ( 
.A(n_1532),
.B(n_34),
.Y(n_1735)
);

AOI22xp33_ASAP7_75t_L g1736 ( 
.A1(n_1533),
.A2(n_37),
.B1(n_34),
.B2(n_36),
.Y(n_1736)
);

INVx1_ASAP7_75t_L g1737 ( 
.A(n_1428),
.Y(n_1737)
);

OAI22xp5_ASAP7_75t_L g1738 ( 
.A1(n_1404),
.A2(n_38),
.B1(n_36),
.B2(n_37),
.Y(n_1738)
);

NAND2xp5_ASAP7_75t_L g1739 ( 
.A(n_1435),
.B(n_1449),
.Y(n_1739)
);

NOR2xp33_ASAP7_75t_L g1740 ( 
.A(n_1521),
.B(n_1527),
.Y(n_1740)
);

AOI22xp5_ASAP7_75t_L g1741 ( 
.A1(n_1379),
.A2(n_40),
.B1(n_38),
.B2(n_39),
.Y(n_1741)
);

NAND2xp5_ASAP7_75t_L g1742 ( 
.A(n_1452),
.B(n_39),
.Y(n_1742)
);

A2O1A1Ixp33_ASAP7_75t_L g1743 ( 
.A1(n_1432),
.A2(n_43),
.B(n_41),
.C(n_42),
.Y(n_1743)
);

NAND2xp5_ASAP7_75t_L g1744 ( 
.A(n_1498),
.B(n_42),
.Y(n_1744)
);

A2O1A1Ixp33_ASAP7_75t_L g1745 ( 
.A1(n_1506),
.A2(n_47),
.B(n_44),
.C(n_45),
.Y(n_1745)
);

AND2x2_ASAP7_75t_L g1746 ( 
.A(n_1464),
.B(n_1429),
.Y(n_1746)
);

NAND2xp5_ASAP7_75t_L g1747 ( 
.A(n_1501),
.B(n_44),
.Y(n_1747)
);

INVx3_ASAP7_75t_L g1748 ( 
.A(n_1569),
.Y(n_1748)
);

INVx2_ASAP7_75t_L g1749 ( 
.A(n_1373),
.Y(n_1749)
);

NOR2xp33_ASAP7_75t_L g1750 ( 
.A(n_1550),
.B(n_48),
.Y(n_1750)
);

NAND2xp5_ASAP7_75t_SL g1751 ( 
.A(n_1516),
.B(n_49),
.Y(n_1751)
);

INVx2_ASAP7_75t_L g1752 ( 
.A(n_1374),
.Y(n_1752)
);

AOI22xp5_ASAP7_75t_L g1753 ( 
.A1(n_1420),
.A2(n_52),
.B1(n_49),
.B2(n_50),
.Y(n_1753)
);

NOR2x2_ASAP7_75t_L g1754 ( 
.A(n_1476),
.B(n_52),
.Y(n_1754)
);

INVx3_ASAP7_75t_L g1755 ( 
.A(n_1572),
.Y(n_1755)
);

INVx1_ASAP7_75t_L g1756 ( 
.A(n_1378),
.Y(n_1756)
);

OAI21xp5_ASAP7_75t_L g1757 ( 
.A1(n_1387),
.A2(n_665),
.B(n_663),
.Y(n_1757)
);

AOI21xp5_ASAP7_75t_L g1758 ( 
.A1(n_1537),
.A2(n_700),
.B(n_698),
.Y(n_1758)
);

NAND2xp5_ASAP7_75t_L g1759 ( 
.A(n_1539),
.B(n_53),
.Y(n_1759)
);

INVxp67_ASAP7_75t_L g1760 ( 
.A(n_1415),
.Y(n_1760)
);

INVx2_ASAP7_75t_L g1761 ( 
.A(n_1383),
.Y(n_1761)
);

AOI21xp5_ASAP7_75t_L g1762 ( 
.A1(n_1540),
.A2(n_668),
.B(n_666),
.Y(n_1762)
);

INVx4_ASAP7_75t_L g1763 ( 
.A(n_1415),
.Y(n_1763)
);

NOR2xp33_ASAP7_75t_L g1764 ( 
.A(n_1544),
.B(n_54),
.Y(n_1764)
);

INVx1_ASAP7_75t_L g1765 ( 
.A(n_1384),
.Y(n_1765)
);

AOI21xp5_ASAP7_75t_L g1766 ( 
.A1(n_1543),
.A2(n_696),
.B(n_695),
.Y(n_1766)
);

INVx1_ASAP7_75t_L g1767 ( 
.A(n_1393),
.Y(n_1767)
);

INVx11_ASAP7_75t_L g1768 ( 
.A(n_1444),
.Y(n_1768)
);

A2O1A1Ixp33_ASAP7_75t_L g1769 ( 
.A1(n_1551),
.A2(n_57),
.B(n_55),
.C(n_56),
.Y(n_1769)
);

AOI21xp5_ASAP7_75t_L g1770 ( 
.A1(n_1503),
.A2(n_1514),
.B(n_1512),
.Y(n_1770)
);

NAND2xp5_ASAP7_75t_L g1771 ( 
.A(n_1515),
.B(n_55),
.Y(n_1771)
);

OAI21xp5_ASAP7_75t_L g1772 ( 
.A1(n_1541),
.A2(n_1362),
.B(n_1359),
.Y(n_1772)
);

AOI22xp5_ASAP7_75t_L g1773 ( 
.A1(n_1470),
.A2(n_1368),
.B1(n_1556),
.B2(n_1560),
.Y(n_1773)
);

NOR2xp33_ASAP7_75t_L g1774 ( 
.A(n_1556),
.B(n_57),
.Y(n_1774)
);

NOR2xp33_ASAP7_75t_L g1775 ( 
.A(n_1522),
.B(n_58),
.Y(n_1775)
);

BUFx4f_ASAP7_75t_L g1776 ( 
.A(n_1397),
.Y(n_1776)
);

AOI22xp5_ASAP7_75t_L g1777 ( 
.A1(n_1517),
.A2(n_1464),
.B1(n_1562),
.B2(n_1558),
.Y(n_1777)
);

BUFx4f_ASAP7_75t_L g1778 ( 
.A(n_1555),
.Y(n_1778)
);

O2A1O1Ixp33_ASAP7_75t_L g1779 ( 
.A1(n_1554),
.A2(n_62),
.B(n_60),
.C(n_61),
.Y(n_1779)
);

AOI22xp5_ASAP7_75t_L g1780 ( 
.A1(n_1565),
.A2(n_65),
.B1(n_63),
.B2(n_64),
.Y(n_1780)
);

INVx1_ASAP7_75t_L g1781 ( 
.A(n_1557),
.Y(n_1781)
);

HB1xp67_ASAP7_75t_L g1782 ( 
.A(n_1567),
.Y(n_1782)
);

A2O1A1Ixp33_ASAP7_75t_L g1783 ( 
.A1(n_1568),
.A2(n_67),
.B(n_64),
.C(n_66),
.Y(n_1783)
);

AOI21xp5_ASAP7_75t_L g1784 ( 
.A1(n_1547),
.A2(n_684),
.B(n_683),
.Y(n_1784)
);

O2A1O1Ixp33_ASAP7_75t_L g1785 ( 
.A1(n_1570),
.A2(n_69),
.B(n_67),
.C(n_68),
.Y(n_1785)
);

OAI321xp33_ASAP7_75t_L g1786 ( 
.A1(n_1561),
.A2(n_72),
.A3(n_74),
.B1(n_69),
.B2(n_70),
.C(n_73),
.Y(n_1786)
);

INVx3_ASAP7_75t_L g1787 ( 
.A(n_1572),
.Y(n_1787)
);

NOR2xp33_ASAP7_75t_L g1788 ( 
.A(n_1549),
.B(n_74),
.Y(n_1788)
);

INVxp67_ASAP7_75t_L g1789 ( 
.A(n_1571),
.Y(n_1789)
);

INVx1_ASAP7_75t_SL g1790 ( 
.A(n_1549),
.Y(n_1790)
);

AND2x4_ASAP7_75t_L g1791 ( 
.A(n_1564),
.B(n_76),
.Y(n_1791)
);

BUFx2_ASAP7_75t_L g1792 ( 
.A(n_1553),
.Y(n_1792)
);

AOI21xp5_ASAP7_75t_L g1793 ( 
.A1(n_1563),
.A2(n_678),
.B(n_677),
.Y(n_1793)
);

AOI21xp5_ASAP7_75t_L g1794 ( 
.A1(n_1518),
.A2(n_691),
.B(n_685),
.Y(n_1794)
);

NAND2xp5_ASAP7_75t_L g1795 ( 
.A(n_1490),
.B(n_76),
.Y(n_1795)
);

OAI21xp5_ASAP7_75t_L g1796 ( 
.A1(n_1542),
.A2(n_693),
.B(n_692),
.Y(n_1796)
);

OAI22xp5_ASAP7_75t_L g1797 ( 
.A1(n_1490),
.A2(n_80),
.B1(n_77),
.B2(n_79),
.Y(n_1797)
);

NAND2xp5_ASAP7_75t_L g1798 ( 
.A(n_1490),
.B(n_79),
.Y(n_1798)
);

NOR2xp33_ASAP7_75t_L g1799 ( 
.A(n_1363),
.B(n_81),
.Y(n_1799)
);

INVxp67_ASAP7_75t_L g1800 ( 
.A(n_1363),
.Y(n_1800)
);

AND2x2_ASAP7_75t_L g1801 ( 
.A(n_1363),
.B(n_631),
.Y(n_1801)
);

NAND2xp5_ASAP7_75t_SL g1802 ( 
.A(n_1363),
.B(n_81),
.Y(n_1802)
);

OAI21xp5_ASAP7_75t_L g1803 ( 
.A1(n_1542),
.A2(n_82),
.B(n_83),
.Y(n_1803)
);

OAI21xp5_ASAP7_75t_L g1804 ( 
.A1(n_1542),
.A2(n_82),
.B(n_85),
.Y(n_1804)
);

AOI21xp5_ASAP7_75t_L g1805 ( 
.A1(n_1518),
.A2(n_86),
.B(n_87),
.Y(n_1805)
);

NOR2x1_ASAP7_75t_L g1806 ( 
.A(n_1408),
.B(n_86),
.Y(n_1806)
);

AOI21xp5_ASAP7_75t_L g1807 ( 
.A1(n_1518),
.A2(n_90),
.B(n_91),
.Y(n_1807)
);

OAI21xp5_ASAP7_75t_L g1808 ( 
.A1(n_1542),
.A2(n_90),
.B(n_91),
.Y(n_1808)
);

NAND2xp5_ASAP7_75t_L g1809 ( 
.A(n_1490),
.B(n_92),
.Y(n_1809)
);

INVx1_ASAP7_75t_L g1810 ( 
.A(n_1443),
.Y(n_1810)
);

INVx4_ASAP7_75t_L g1811 ( 
.A(n_1408),
.Y(n_1811)
);

AOI21xp5_ASAP7_75t_L g1812 ( 
.A1(n_1518),
.A2(n_93),
.B(n_94),
.Y(n_1812)
);

NOR2xp33_ASAP7_75t_L g1813 ( 
.A(n_1363),
.B(n_630),
.Y(n_1813)
);

NAND2xp5_ASAP7_75t_L g1814 ( 
.A(n_1490),
.B(n_93),
.Y(n_1814)
);

NAND2xp5_ASAP7_75t_L g1815 ( 
.A(n_1490),
.B(n_95),
.Y(n_1815)
);

NAND2xp5_ASAP7_75t_L g1816 ( 
.A(n_1490),
.B(n_96),
.Y(n_1816)
);

NAND2xp5_ASAP7_75t_L g1817 ( 
.A(n_1490),
.B(n_96),
.Y(n_1817)
);

OAI21xp5_ASAP7_75t_L g1818 ( 
.A1(n_1542),
.A2(n_98),
.B(n_100),
.Y(n_1818)
);

CKINVDCx5p33_ASAP7_75t_R g1819 ( 
.A(n_1525),
.Y(n_1819)
);

O2A1O1Ixp33_ASAP7_75t_L g1820 ( 
.A1(n_1446),
.A2(n_102),
.B(n_100),
.C(n_101),
.Y(n_1820)
);

INVx1_ASAP7_75t_L g1821 ( 
.A(n_1443),
.Y(n_1821)
);

NAND2xp5_ASAP7_75t_SL g1822 ( 
.A(n_1363),
.B(n_102),
.Y(n_1822)
);

AOI21xp5_ASAP7_75t_L g1823 ( 
.A1(n_1518),
.A2(n_103),
.B(n_104),
.Y(n_1823)
);

AND2x4_ASAP7_75t_L g1824 ( 
.A(n_1811),
.B(n_107),
.Y(n_1824)
);

AND2x4_ASAP7_75t_L g1825 ( 
.A(n_1811),
.B(n_107),
.Y(n_1825)
);

AND3x4_ASAP7_75t_L g1826 ( 
.A(n_1640),
.B(n_109),
.C(n_110),
.Y(n_1826)
);

OAI22xp5_ASAP7_75t_L g1827 ( 
.A1(n_1675),
.A2(n_113),
.B1(n_111),
.B2(n_112),
.Y(n_1827)
);

INVx2_ASAP7_75t_SL g1828 ( 
.A(n_1647),
.Y(n_1828)
);

AO22x1_ASAP7_75t_L g1829 ( 
.A1(n_1646),
.A2(n_116),
.B1(n_113),
.B2(n_114),
.Y(n_1829)
);

AOI21x1_ASAP7_75t_SL g1830 ( 
.A1(n_1739),
.A2(n_117),
.B(n_118),
.Y(n_1830)
);

INVx2_ASAP7_75t_SL g1831 ( 
.A(n_1647),
.Y(n_1831)
);

INVx2_ASAP7_75t_SL g1832 ( 
.A(n_1690),
.Y(n_1832)
);

NAND2xp5_ASAP7_75t_L g1833 ( 
.A(n_1708),
.B(n_119),
.Y(n_1833)
);

OAI21x1_ASAP7_75t_L g1834 ( 
.A1(n_1617),
.A2(n_1693),
.B(n_1796),
.Y(n_1834)
);

BUFx4f_ASAP7_75t_L g1835 ( 
.A(n_1648),
.Y(n_1835)
);

OAI21x1_ASAP7_75t_L g1836 ( 
.A1(n_1794),
.A2(n_121),
.B(n_122),
.Y(n_1836)
);

NOR2xp67_ASAP7_75t_SL g1837 ( 
.A(n_1689),
.B(n_123),
.Y(n_1837)
);

OAI21xp5_ASAP7_75t_L g1838 ( 
.A1(n_1770),
.A2(n_125),
.B(n_126),
.Y(n_1838)
);

NOR2x1_ASAP7_75t_SL g1839 ( 
.A(n_1707),
.B(n_127),
.Y(n_1839)
);

AOI22xp5_ASAP7_75t_L g1840 ( 
.A1(n_1800),
.A2(n_129),
.B1(n_127),
.B2(n_128),
.Y(n_1840)
);

NAND3xp33_ASAP7_75t_SL g1841 ( 
.A(n_1773),
.B(n_128),
.C(n_129),
.Y(n_1841)
);

NAND2xp5_ASAP7_75t_L g1842 ( 
.A(n_1575),
.B(n_1705),
.Y(n_1842)
);

AOI211x1_ASAP7_75t_L g1843 ( 
.A1(n_1718),
.A2(n_134),
.B(n_130),
.C(n_133),
.Y(n_1843)
);

INVx1_ASAP7_75t_L g1844 ( 
.A(n_1795),
.Y(n_1844)
);

INVx1_ASAP7_75t_L g1845 ( 
.A(n_1798),
.Y(n_1845)
);

NAND2xp5_ASAP7_75t_L g1846 ( 
.A(n_1611),
.B(n_133),
.Y(n_1846)
);

INVx1_ASAP7_75t_L g1847 ( 
.A(n_1809),
.Y(n_1847)
);

NAND2xp5_ASAP7_75t_L g1848 ( 
.A(n_1624),
.B(n_134),
.Y(n_1848)
);

AOI21x1_ASAP7_75t_SL g1849 ( 
.A1(n_1742),
.A2(n_137),
.B(n_139),
.Y(n_1849)
);

OAI21x1_ASAP7_75t_SL g1850 ( 
.A1(n_1757),
.A2(n_142),
.B(n_143),
.Y(n_1850)
);

OAI21xp5_ASAP7_75t_L g1851 ( 
.A1(n_1591),
.A2(n_142),
.B(n_143),
.Y(n_1851)
);

NAND2xp5_ASAP7_75t_L g1852 ( 
.A(n_1657),
.B(n_144),
.Y(n_1852)
);

NOR2xp33_ASAP7_75t_L g1853 ( 
.A(n_1661),
.B(n_1668),
.Y(n_1853)
);

INVx8_ASAP7_75t_L g1854 ( 
.A(n_1601),
.Y(n_1854)
);

OAI22x1_ASAP7_75t_L g1855 ( 
.A1(n_1791),
.A2(n_147),
.B1(n_145),
.B2(n_146),
.Y(n_1855)
);

A2O1A1Ixp33_ASAP7_75t_L g1856 ( 
.A1(n_1592),
.A2(n_147),
.B(n_145),
.C(n_146),
.Y(n_1856)
);

OAI21xp5_ASAP7_75t_L g1857 ( 
.A1(n_1598),
.A2(n_148),
.B(n_149),
.Y(n_1857)
);

BUFx3_ASAP7_75t_L g1858 ( 
.A(n_1715),
.Y(n_1858)
);

AND2x2_ASAP7_75t_SL g1859 ( 
.A(n_1600),
.B(n_150),
.Y(n_1859)
);

OAI21xp5_ASAP7_75t_L g1860 ( 
.A1(n_1607),
.A2(n_151),
.B(n_153),
.Y(n_1860)
);

NAND2x1p5_ASAP7_75t_L g1861 ( 
.A(n_1734),
.B(n_155),
.Y(n_1861)
);

AOI21xp5_ASAP7_75t_SL g1862 ( 
.A1(n_1707),
.A2(n_156),
.B(n_157),
.Y(n_1862)
);

A2O1A1Ixp33_ASAP7_75t_L g1863 ( 
.A1(n_1612),
.A2(n_161),
.B(n_159),
.C(n_160),
.Y(n_1863)
);

A2O1A1Ixp33_ASAP7_75t_L g1864 ( 
.A1(n_1621),
.A2(n_163),
.B(n_161),
.C(n_162),
.Y(n_1864)
);

OAI21x1_ASAP7_75t_L g1865 ( 
.A1(n_1758),
.A2(n_1766),
.B(n_1762),
.Y(n_1865)
);

OAI21x1_ASAP7_75t_L g1866 ( 
.A1(n_1716),
.A2(n_165),
.B(n_166),
.Y(n_1866)
);

A2O1A1Ixp33_ASAP7_75t_L g1867 ( 
.A1(n_1614),
.A2(n_167),
.B(n_165),
.C(n_166),
.Y(n_1867)
);

AOI22xp5_ASAP7_75t_L g1868 ( 
.A1(n_1577),
.A2(n_172),
.B1(n_170),
.B2(n_171),
.Y(n_1868)
);

INVx1_ASAP7_75t_L g1869 ( 
.A(n_1814),
.Y(n_1869)
);

NAND2xp5_ASAP7_75t_L g1870 ( 
.A(n_1632),
.B(n_173),
.Y(n_1870)
);

NAND2xp5_ASAP7_75t_L g1871 ( 
.A(n_1665),
.B(n_174),
.Y(n_1871)
);

AO31x2_ASAP7_75t_L g1872 ( 
.A1(n_1576),
.A2(n_180),
.A3(n_175),
.B(n_178),
.Y(n_1872)
);

OAI21xp5_ASAP7_75t_L g1873 ( 
.A1(n_1639),
.A2(n_178),
.B(n_180),
.Y(n_1873)
);

NAND2xp5_ASAP7_75t_L g1874 ( 
.A(n_1660),
.B(n_182),
.Y(n_1874)
);

INVx1_ASAP7_75t_L g1875 ( 
.A(n_1815),
.Y(n_1875)
);

OAI21xp5_ASAP7_75t_L g1876 ( 
.A1(n_1603),
.A2(n_185),
.B(n_187),
.Y(n_1876)
);

OAI21x1_ASAP7_75t_L g1877 ( 
.A1(n_1793),
.A2(n_1784),
.B(n_1623),
.Y(n_1877)
);

CKINVDCx5p33_ASAP7_75t_R g1878 ( 
.A(n_1646),
.Y(n_1878)
);

NAND2xp5_ASAP7_75t_L g1879 ( 
.A(n_1660),
.B(n_189),
.Y(n_1879)
);

OAI21xp5_ASAP7_75t_L g1880 ( 
.A1(n_1625),
.A2(n_190),
.B(n_191),
.Y(n_1880)
);

NAND2xp5_ASAP7_75t_L g1881 ( 
.A(n_1664),
.B(n_194),
.Y(n_1881)
);

NAND2xp5_ASAP7_75t_L g1882 ( 
.A(n_1664),
.B(n_194),
.Y(n_1882)
);

NAND2xp5_ASAP7_75t_SL g1883 ( 
.A(n_1578),
.B(n_195),
.Y(n_1883)
);

AOI21x1_ASAP7_75t_SL g1884 ( 
.A1(n_1744),
.A2(n_197),
.B(n_198),
.Y(n_1884)
);

NAND2xp5_ASAP7_75t_L g1885 ( 
.A(n_1667),
.B(n_199),
.Y(n_1885)
);

HB1xp67_ASAP7_75t_L g1886 ( 
.A(n_1594),
.Y(n_1886)
);

AO31x2_ASAP7_75t_L g1887 ( 
.A1(n_1653),
.A2(n_202),
.A3(n_200),
.B(n_201),
.Y(n_1887)
);

NAND2xp5_ASAP7_75t_L g1888 ( 
.A(n_1580),
.B(n_201),
.Y(n_1888)
);

BUFx4f_ASAP7_75t_L g1889 ( 
.A(n_1601),
.Y(n_1889)
);

OAI21x1_ASAP7_75t_SL g1890 ( 
.A1(n_1757),
.A2(n_1804),
.B(n_1803),
.Y(n_1890)
);

INVx1_ASAP7_75t_L g1891 ( 
.A(n_1816),
.Y(n_1891)
);

NAND2xp5_ASAP7_75t_L g1892 ( 
.A(n_1694),
.B(n_1589),
.Y(n_1892)
);

OAI21x1_ASAP7_75t_L g1893 ( 
.A1(n_1608),
.A2(n_203),
.B(n_204),
.Y(n_1893)
);

AOI21xp5_ASAP7_75t_L g1894 ( 
.A1(n_1772),
.A2(n_205),
.B(n_206),
.Y(n_1894)
);

OAI21xp5_ASAP7_75t_L g1895 ( 
.A1(n_1638),
.A2(n_207),
.B(n_208),
.Y(n_1895)
);

NAND2xp5_ASAP7_75t_L g1896 ( 
.A(n_1645),
.B(n_207),
.Y(n_1896)
);

AOI21xp5_ASAP7_75t_L g1897 ( 
.A1(n_1772),
.A2(n_208),
.B(n_210),
.Y(n_1897)
);

NAND2xp5_ASAP7_75t_L g1898 ( 
.A(n_1654),
.B(n_210),
.Y(n_1898)
);

NAND2xp5_ASAP7_75t_L g1899 ( 
.A(n_1667),
.B(n_211),
.Y(n_1899)
);

NAND2xp5_ASAP7_75t_L g1900 ( 
.A(n_1609),
.B(n_211),
.Y(n_1900)
);

INVx1_ASAP7_75t_L g1901 ( 
.A(n_1817),
.Y(n_1901)
);

AND2x2_ASAP7_75t_L g1902 ( 
.A(n_1635),
.B(n_212),
.Y(n_1902)
);

NOR2xp33_ASAP7_75t_L g1903 ( 
.A(n_1711),
.B(n_212),
.Y(n_1903)
);

INVxp67_ASAP7_75t_L g1904 ( 
.A(n_1634),
.Y(n_1904)
);

OAI21xp5_ASAP7_75t_L g1905 ( 
.A1(n_1638),
.A2(n_213),
.B(n_214),
.Y(n_1905)
);

NAND3xp33_ASAP7_75t_SL g1906 ( 
.A(n_1820),
.B(n_217),
.C(n_218),
.Y(n_1906)
);

NAND2x1p5_ASAP7_75t_L g1907 ( 
.A(n_1734),
.B(n_218),
.Y(n_1907)
);

NOR2xp33_ASAP7_75t_L g1908 ( 
.A(n_1663),
.B(n_1652),
.Y(n_1908)
);

AND2x2_ASAP7_75t_L g1909 ( 
.A(n_1593),
.B(n_219),
.Y(n_1909)
);

NAND2xp5_ASAP7_75t_SL g1910 ( 
.A(n_1734),
.B(n_220),
.Y(n_1910)
);

INVx2_ASAP7_75t_L g1911 ( 
.A(n_1602),
.Y(n_1911)
);

BUFx12f_ASAP7_75t_L g1912 ( 
.A(n_1697),
.Y(n_1912)
);

BUFx3_ASAP7_75t_L g1913 ( 
.A(n_1763),
.Y(n_1913)
);

INVx1_ASAP7_75t_L g1914 ( 
.A(n_1681),
.Y(n_1914)
);

A2O1A1Ixp33_ASAP7_75t_L g1915 ( 
.A1(n_1630),
.A2(n_226),
.B(n_222),
.C(n_225),
.Y(n_1915)
);

NAND2xp5_ASAP7_75t_L g1916 ( 
.A(n_1629),
.B(n_225),
.Y(n_1916)
);

AOI21xp5_ASAP7_75t_L g1917 ( 
.A1(n_1573),
.A2(n_226),
.B(n_227),
.Y(n_1917)
);

HB1xp67_ASAP7_75t_L g1918 ( 
.A(n_1663),
.Y(n_1918)
);

NAND2xp5_ASAP7_75t_L g1919 ( 
.A(n_1644),
.B(n_230),
.Y(n_1919)
);

NAND2xp5_ASAP7_75t_L g1920 ( 
.A(n_1655),
.B(n_230),
.Y(n_1920)
);

NAND2xp5_ASAP7_75t_L g1921 ( 
.A(n_1781),
.B(n_231),
.Y(n_1921)
);

OAI22x1_ASAP7_75t_L g1922 ( 
.A1(n_1791),
.A2(n_236),
.B1(n_231),
.B2(n_235),
.Y(n_1922)
);

AND2x2_ASAP7_75t_L g1923 ( 
.A(n_1746),
.B(n_236),
.Y(n_1923)
);

OAI21xp5_ASAP7_75t_L g1924 ( 
.A1(n_1588),
.A2(n_237),
.B(n_238),
.Y(n_1924)
);

OAI21xp33_ASAP7_75t_L g1925 ( 
.A1(n_1579),
.A2(n_237),
.B(n_238),
.Y(n_1925)
);

AOI21xp5_ASAP7_75t_L g1926 ( 
.A1(n_1581),
.A2(n_239),
.B(n_240),
.Y(n_1926)
);

AOI21xp5_ASAP7_75t_L g1927 ( 
.A1(n_1582),
.A2(n_241),
.B(n_242),
.Y(n_1927)
);

AND2x4_ASAP7_75t_L g1928 ( 
.A(n_1601),
.B(n_241),
.Y(n_1928)
);

AOI21xp5_ASAP7_75t_L g1929 ( 
.A1(n_1606),
.A2(n_243),
.B(n_244),
.Y(n_1929)
);

NAND2xp5_ASAP7_75t_SL g1930 ( 
.A(n_1600),
.B(n_243),
.Y(n_1930)
);

AOI21xp5_ASAP7_75t_L g1931 ( 
.A1(n_1610),
.A2(n_245),
.B(n_246),
.Y(n_1931)
);

AOI21xp5_ASAP7_75t_L g1932 ( 
.A1(n_1680),
.A2(n_245),
.B(n_246),
.Y(n_1932)
);

AO31x2_ASAP7_75t_L g1933 ( 
.A1(n_1722),
.A2(n_249),
.A3(n_247),
.B(n_248),
.Y(n_1933)
);

NAND2xp5_ASAP7_75t_L g1934 ( 
.A(n_1670),
.B(n_247),
.Y(n_1934)
);

A2O1A1Ixp33_ASAP7_75t_L g1935 ( 
.A1(n_1682),
.A2(n_251),
.B(n_248),
.C(n_250),
.Y(n_1935)
);

INVx2_ASAP7_75t_SL g1936 ( 
.A(n_1768),
.Y(n_1936)
);

NAND2xp5_ASAP7_75t_L g1937 ( 
.A(n_1684),
.B(n_253),
.Y(n_1937)
);

A2O1A1Ixp33_ASAP7_75t_L g1938 ( 
.A1(n_1785),
.A2(n_255),
.B(n_253),
.C(n_254),
.Y(n_1938)
);

AOI21xp5_ASAP7_75t_L g1939 ( 
.A1(n_1683),
.A2(n_256),
.B(n_257),
.Y(n_1939)
);

NAND2xp5_ASAP7_75t_L g1940 ( 
.A(n_1685),
.B(n_1777),
.Y(n_1940)
);

AOI21xp5_ASAP7_75t_L g1941 ( 
.A1(n_1622),
.A2(n_256),
.B(n_257),
.Y(n_1941)
);

INVx3_ASAP7_75t_L g1942 ( 
.A(n_1755),
.Y(n_1942)
);

NAND2xp5_ASAP7_75t_L g1943 ( 
.A(n_1656),
.B(n_258),
.Y(n_1943)
);

NAND2xp5_ASAP7_75t_SL g1944 ( 
.A(n_1778),
.B(n_261),
.Y(n_1944)
);

AND2x2_ASAP7_75t_L g1945 ( 
.A(n_1613),
.B(n_262),
.Y(n_1945)
);

AO21x1_ASAP7_75t_L g1946 ( 
.A1(n_1803),
.A2(n_1808),
.B(n_1804),
.Y(n_1946)
);

INVx1_ASAP7_75t_L g1947 ( 
.A(n_1737),
.Y(n_1947)
);

BUFx12f_ASAP7_75t_L g1948 ( 
.A(n_1697),
.Y(n_1948)
);

OAI21x1_ASAP7_75t_SL g1949 ( 
.A1(n_1808),
.A2(n_267),
.B(n_268),
.Y(n_1949)
);

AO21x1_ASAP7_75t_L g1950 ( 
.A1(n_1818),
.A2(n_267),
.B(n_268),
.Y(n_1950)
);

AND2x2_ASAP7_75t_L g1951 ( 
.A(n_1713),
.B(n_269),
.Y(n_1951)
);

OAI21xp5_ASAP7_75t_L g1952 ( 
.A1(n_1586),
.A2(n_269),
.B(n_270),
.Y(n_1952)
);

INVx1_ASAP7_75t_L g1953 ( 
.A(n_1587),
.Y(n_1953)
);

AOI21xp5_ASAP7_75t_L g1954 ( 
.A1(n_1626),
.A2(n_271),
.B(n_272),
.Y(n_1954)
);

INVx1_ASAP7_75t_L g1955 ( 
.A(n_1605),
.Y(n_1955)
);

BUFx6f_ASAP7_75t_L g1956 ( 
.A(n_1643),
.Y(n_1956)
);

AND2x4_ASAP7_75t_L g1957 ( 
.A(n_1615),
.B(n_1810),
.Y(n_1957)
);

BUFx12f_ASAP7_75t_L g1958 ( 
.A(n_1687),
.Y(n_1958)
);

NAND2xp5_ASAP7_75t_L g1959 ( 
.A(n_1659),
.B(n_1666),
.Y(n_1959)
);

NAND2xp5_ASAP7_75t_L g1960 ( 
.A(n_1821),
.B(n_1583),
.Y(n_1960)
);

INVx3_ASAP7_75t_L g1961 ( 
.A(n_1755),
.Y(n_1961)
);

OAI21xp5_ASAP7_75t_L g1962 ( 
.A1(n_1618),
.A2(n_279),
.B(n_280),
.Y(n_1962)
);

AND2x4_ASAP7_75t_L g1963 ( 
.A(n_1801),
.B(n_1763),
.Y(n_1963)
);

NAND2x1_ASAP7_75t_SL g1964 ( 
.A(n_1584),
.B(n_1787),
.Y(n_1964)
);

AO31x2_ASAP7_75t_L g1965 ( 
.A1(n_1788),
.A2(n_284),
.A3(n_281),
.B(n_282),
.Y(n_1965)
);

INVx4_ASAP7_75t_L g1966 ( 
.A(n_1787),
.Y(n_1966)
);

INVx1_ASAP7_75t_L g1967 ( 
.A(n_1756),
.Y(n_1967)
);

NAND2xp5_ASAP7_75t_L g1968 ( 
.A(n_1633),
.B(n_281),
.Y(n_1968)
);

NAND2xp5_ASAP7_75t_SL g1969 ( 
.A(n_1778),
.B(n_1707),
.Y(n_1969)
);

AOI21xp5_ASAP7_75t_L g1970 ( 
.A1(n_1636),
.A2(n_1641),
.B(n_1595),
.Y(n_1970)
);

INVx2_ASAP7_75t_SL g1971 ( 
.A(n_1651),
.Y(n_1971)
);

INVx3_ASAP7_75t_L g1972 ( 
.A(n_1748),
.Y(n_1972)
);

AND2x2_ASAP7_75t_L g1973 ( 
.A(n_1704),
.B(n_286),
.Y(n_1973)
);

AOI21xp5_ASAP7_75t_L g1974 ( 
.A1(n_1710),
.A2(n_286),
.B(n_287),
.Y(n_1974)
);

NOR3xp33_ASAP7_75t_L g1975 ( 
.A(n_1740),
.B(n_287),
.C(n_289),
.Y(n_1975)
);

INVx3_ASAP7_75t_L g1976 ( 
.A(n_1748),
.Y(n_1976)
);

AOI21xp5_ASAP7_75t_L g1977 ( 
.A1(n_1658),
.A2(n_289),
.B(n_290),
.Y(n_1977)
);

INVx1_ASAP7_75t_L g1978 ( 
.A(n_1765),
.Y(n_1978)
);

AOI21xp5_ASAP7_75t_L g1979 ( 
.A1(n_1672),
.A2(n_290),
.B(n_291),
.Y(n_1979)
);

AND2x2_ASAP7_75t_L g1980 ( 
.A(n_1704),
.B(n_292),
.Y(n_1980)
);

INVx4_ASAP7_75t_L g1981 ( 
.A(n_1628),
.Y(n_1981)
);

OAI22xp5_ASAP7_75t_L g1982 ( 
.A1(n_1619),
.A2(n_295),
.B1(n_293),
.B2(n_294),
.Y(n_1982)
);

CKINVDCx8_ASAP7_75t_R g1983 ( 
.A(n_1819),
.Y(n_1983)
);

AOI221xp5_ASAP7_75t_L g1984 ( 
.A1(n_1671),
.A2(n_1662),
.B1(n_1764),
.B2(n_1604),
.C(n_1616),
.Y(n_1984)
);

AND2x2_ASAP7_75t_L g1985 ( 
.A(n_1597),
.B(n_298),
.Y(n_1985)
);

NAND2xp5_ASAP7_75t_L g1986 ( 
.A(n_1676),
.B(n_299),
.Y(n_1986)
);

AOI21xp5_ASAP7_75t_SL g1987 ( 
.A1(n_1643),
.A2(n_300),
.B(n_301),
.Y(n_1987)
);

NAND2xp5_ASAP7_75t_L g1988 ( 
.A(n_1590),
.B(n_308),
.Y(n_1988)
);

AOI21x1_ASAP7_75t_SL g1989 ( 
.A1(n_1747),
.A2(n_309),
.B(n_310),
.Y(n_1989)
);

INVx1_ASAP7_75t_L g1990 ( 
.A(n_1767),
.Y(n_1990)
);

AND2x2_ASAP7_75t_L g1991 ( 
.A(n_1733),
.B(n_1585),
.Y(n_1991)
);

INVx3_ASAP7_75t_SL g1992 ( 
.A(n_1754),
.Y(n_1992)
);

BUFx6f_ASAP7_75t_L g1993 ( 
.A(n_1650),
.Y(n_1993)
);

NAND2xp5_ASAP7_75t_L g1994 ( 
.A(n_1627),
.B(n_309),
.Y(n_1994)
);

NAND2xp5_ASAP7_75t_L g1995 ( 
.A(n_1717),
.B(n_310),
.Y(n_1995)
);

NAND2xp5_ASAP7_75t_L g1996 ( 
.A(n_1679),
.B(n_311),
.Y(n_1996)
);

NOR2xp33_ASAP7_75t_L g1997 ( 
.A(n_1674),
.B(n_313),
.Y(n_1997)
);

INVx1_ASAP7_75t_L g1998 ( 
.A(n_1749),
.Y(n_1998)
);

OAI21xp5_ASAP7_75t_L g1999 ( 
.A1(n_1702),
.A2(n_313),
.B(n_314),
.Y(n_1999)
);

NAND2xp5_ASAP7_75t_L g2000 ( 
.A(n_1712),
.B(n_314),
.Y(n_2000)
);

NAND2xp5_ASAP7_75t_L g2001 ( 
.A(n_1771),
.B(n_1750),
.Y(n_2001)
);

OAI21xp5_ASAP7_75t_L g2002 ( 
.A1(n_1805),
.A2(n_1812),
.B(n_1807),
.Y(n_2002)
);

AO31x2_ASAP7_75t_L g2003 ( 
.A1(n_1769),
.A2(n_317),
.A3(n_315),
.B(n_316),
.Y(n_2003)
);

AND2x2_ASAP7_75t_L g2004 ( 
.A(n_1651),
.B(n_1695),
.Y(n_2004)
);

INVx4_ASAP7_75t_L g2005 ( 
.A(n_1650),
.Y(n_2005)
);

AND2x4_ASAP7_75t_L g2006 ( 
.A(n_1692),
.B(n_315),
.Y(n_2006)
);

AO31x2_ASAP7_75t_L g2007 ( 
.A1(n_1783),
.A2(n_319),
.A3(n_316),
.B(n_318),
.Y(n_2007)
);

HB1xp67_ASAP7_75t_L g2008 ( 
.A(n_1760),
.Y(n_2008)
);

NOR2xp67_ASAP7_75t_SL g2009 ( 
.A(n_1786),
.B(n_318),
.Y(n_2009)
);

NOR2xp33_ASAP7_75t_L g2010 ( 
.A(n_1727),
.B(n_320),
.Y(n_2010)
);

OAI21x1_ASAP7_75t_L g2011 ( 
.A1(n_1730),
.A2(n_321),
.B(n_322),
.Y(n_2011)
);

OAI21xp33_ASAP7_75t_L g2012 ( 
.A1(n_1701),
.A2(n_322),
.B(n_323),
.Y(n_2012)
);

INVx1_ASAP7_75t_L g2013 ( 
.A(n_1752),
.Y(n_2013)
);

NAND2xp5_ASAP7_75t_L g2014 ( 
.A(n_1759),
.B(n_323),
.Y(n_2014)
);

OAI21xp5_ASAP7_75t_SL g2015 ( 
.A1(n_1774),
.A2(n_324),
.B(n_325),
.Y(n_2015)
);

NAND2xp5_ASAP7_75t_L g2016 ( 
.A(n_1761),
.B(n_324),
.Y(n_2016)
);

AO31x2_ASAP7_75t_L g2017 ( 
.A1(n_1743),
.A2(n_328),
.A3(n_326),
.B(n_327),
.Y(n_2017)
);

CKINVDCx6p67_ASAP7_75t_R g2018 ( 
.A(n_1724),
.Y(n_2018)
);

AOI21xp5_ASAP7_75t_L g2019 ( 
.A1(n_1596),
.A2(n_330),
.B(n_331),
.Y(n_2019)
);

NOR2xp67_ASAP7_75t_L g2020 ( 
.A(n_1678),
.B(n_332),
.Y(n_2020)
);

OAI22xp5_ASAP7_75t_L g2021 ( 
.A1(n_1619),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2021)
);

OAI22x1_ASAP7_75t_L g2022 ( 
.A1(n_1806),
.A2(n_335),
.B1(n_333),
.B2(n_334),
.Y(n_2022)
);

OAI21xp5_ASAP7_75t_L g2023 ( 
.A1(n_1823),
.A2(n_336),
.B(n_338),
.Y(n_2023)
);

NAND3xp33_ASAP7_75t_L g2024 ( 
.A(n_1677),
.B(n_338),
.C(n_339),
.Y(n_2024)
);

NAND2x1p5_ASAP7_75t_L g2025 ( 
.A(n_1776),
.B(n_339),
.Y(n_2025)
);

NAND2xp5_ASAP7_75t_L g2026 ( 
.A(n_1799),
.B(n_1813),
.Y(n_2026)
);

INVx1_ASAP7_75t_L g2027 ( 
.A(n_1797),
.Y(n_2027)
);

OAI21x1_ASAP7_75t_SL g2028 ( 
.A1(n_1818),
.A2(n_340),
.B(n_341),
.Y(n_2028)
);

NAND2xp5_ASAP7_75t_SL g2029 ( 
.A(n_1776),
.B(n_341),
.Y(n_2029)
);

OAI21xp33_ASAP7_75t_L g2030 ( 
.A1(n_1599),
.A2(n_344),
.B(n_345),
.Y(n_2030)
);

BUFx3_ASAP7_75t_L g2031 ( 
.A(n_1792),
.Y(n_2031)
);

A2O1A1Ixp33_ASAP7_75t_L g2032 ( 
.A1(n_1779),
.A2(n_348),
.B(n_346),
.C(n_347),
.Y(n_2032)
);

AOI21xp5_ASAP7_75t_L g2033 ( 
.A1(n_1723),
.A2(n_348),
.B(n_349),
.Y(n_2033)
);

INVx2_ASAP7_75t_SL g2034 ( 
.A(n_1649),
.Y(n_2034)
);

NAND2xp5_ASAP7_75t_SL g2035 ( 
.A(n_1642),
.B(n_350),
.Y(n_2035)
);

OAI22xp5_ASAP7_75t_L g2036 ( 
.A1(n_1620),
.A2(n_352),
.B1(n_350),
.B2(n_351),
.Y(n_2036)
);

OAI22xp5_ASAP7_75t_L g2037 ( 
.A1(n_1620),
.A2(n_1736),
.B1(n_1753),
.B2(n_1780),
.Y(n_2037)
);

AO31x2_ASAP7_75t_L g2038 ( 
.A1(n_1745),
.A2(n_357),
.A3(n_354),
.B(n_356),
.Y(n_2038)
);

BUFx2_ASAP7_75t_SL g2039 ( 
.A(n_1673),
.Y(n_2039)
);

INVx8_ASAP7_75t_L g2040 ( 
.A(n_1650),
.Y(n_2040)
);

OAI21xp5_ASAP7_75t_L g2041 ( 
.A1(n_1751),
.A2(n_354),
.B(n_356),
.Y(n_2041)
);

INVx1_ASAP7_75t_L g2042 ( 
.A(n_1696),
.Y(n_2042)
);

OAI22xp5_ASAP7_75t_L g2043 ( 
.A1(n_1741),
.A2(n_360),
.B1(n_358),
.B2(n_359),
.Y(n_2043)
);

NAND2xp5_ASAP7_75t_L g2044 ( 
.A(n_1696),
.B(n_361),
.Y(n_2044)
);

OAI21x1_ASAP7_75t_L g2045 ( 
.A1(n_1735),
.A2(n_364),
.B(n_365),
.Y(n_2045)
);

INVx1_ASAP7_75t_L g2046 ( 
.A(n_1725),
.Y(n_2046)
);

BUFx4_ASAP7_75t_R g2047 ( 
.A(n_1637),
.Y(n_2047)
);

NAND2xp5_ASAP7_75t_L g2048 ( 
.A(n_1782),
.B(n_365),
.Y(n_2048)
);

AOI21xp5_ASAP7_75t_L g2049 ( 
.A1(n_1726),
.A2(n_366),
.B(n_367),
.Y(n_2049)
);

NAND2xp5_ASAP7_75t_L g2050 ( 
.A(n_1720),
.B(n_367),
.Y(n_2050)
);

HB1xp67_ASAP7_75t_L g2051 ( 
.A(n_1738),
.Y(n_2051)
);

AND2x2_ASAP7_75t_L g2052 ( 
.A(n_1709),
.B(n_368),
.Y(n_2052)
);

NAND2xp5_ASAP7_75t_L g2053 ( 
.A(n_1714),
.B(n_368),
.Y(n_2053)
);

HB1xp67_ASAP7_75t_L g2054 ( 
.A(n_1802),
.Y(n_2054)
);

OAI21xp5_ASAP7_75t_L g2055 ( 
.A1(n_1728),
.A2(n_370),
.B(n_371),
.Y(n_2055)
);

CKINVDCx5p33_ASAP7_75t_R g2056 ( 
.A(n_1775),
.Y(n_2056)
);

AND2x2_ASAP7_75t_L g2057 ( 
.A(n_1698),
.B(n_370),
.Y(n_2057)
);

AOI21xp5_ASAP7_75t_L g2058 ( 
.A1(n_1729),
.A2(n_372),
.B(n_374),
.Y(n_2058)
);

AOI21xp5_ASAP7_75t_L g2059 ( 
.A1(n_1700),
.A2(n_375),
.B(n_377),
.Y(n_2059)
);

INVx1_ASAP7_75t_SL g2060 ( 
.A(n_1790),
.Y(n_2060)
);

OAI22x1_ASAP7_75t_L g2061 ( 
.A1(n_1822),
.A2(n_378),
.B1(n_375),
.B2(n_377),
.Y(n_2061)
);

NOR2xp33_ASAP7_75t_SL g2062 ( 
.A(n_1669),
.B(n_1790),
.Y(n_2062)
);

NAND2xp5_ASAP7_75t_L g2063 ( 
.A(n_1721),
.B(n_379),
.Y(n_2063)
);

AOI21xp33_ASAP7_75t_L g2064 ( 
.A1(n_1786),
.A2(n_381),
.B(n_382),
.Y(n_2064)
);

OAI21xp5_ASAP7_75t_L g2065 ( 
.A1(n_1719),
.A2(n_383),
.B(n_384),
.Y(n_2065)
);

OAI21xp5_ASAP7_75t_L g2066 ( 
.A1(n_1574),
.A2(n_384),
.B(n_385),
.Y(n_2066)
);

OAI22xp5_ASAP7_75t_L g2067 ( 
.A1(n_1686),
.A2(n_387),
.B1(n_385),
.B2(n_386),
.Y(n_2067)
);

NAND2xp5_ASAP7_75t_L g2068 ( 
.A(n_1688),
.B(n_388),
.Y(n_2068)
);

BUFx6f_ASAP7_75t_L g2069 ( 
.A(n_1686),
.Y(n_2069)
);

AND2x2_ASAP7_75t_L g2070 ( 
.A(n_1732),
.B(n_389),
.Y(n_2070)
);

OAI21xp5_ASAP7_75t_L g2071 ( 
.A1(n_1699),
.A2(n_390),
.B(n_391),
.Y(n_2071)
);

INVx1_ASAP7_75t_L g2072 ( 
.A(n_1731),
.Y(n_2072)
);

AND3x4_ASAP7_75t_L g2073 ( 
.A(n_1789),
.B(n_390),
.C(n_392),
.Y(n_2073)
);

AND2x4_ASAP7_75t_L g2074 ( 
.A(n_1691),
.B(n_394),
.Y(n_2074)
);

OAI21x1_ASAP7_75t_SL g2075 ( 
.A1(n_1757),
.A2(n_395),
.B(n_396),
.Y(n_2075)
);

NAND2xp5_ASAP7_75t_L g2076 ( 
.A(n_1675),
.B(n_397),
.Y(n_2076)
);

AO31x2_ASAP7_75t_L g2077 ( 
.A1(n_1718),
.A2(n_401),
.A3(n_399),
.B(n_400),
.Y(n_2077)
);

OAI21x1_ASAP7_75t_L g2078 ( 
.A1(n_1706),
.A2(n_399),
.B(n_401),
.Y(n_2078)
);

NAND2xp5_ASAP7_75t_L g2079 ( 
.A(n_1675),
.B(n_402),
.Y(n_2079)
);

INVx1_ASAP7_75t_L g2080 ( 
.A(n_1795),
.Y(n_2080)
);

INVx2_ASAP7_75t_SL g2081 ( 
.A(n_1647),
.Y(n_2081)
);

NOR2xp67_ASAP7_75t_L g2082 ( 
.A(n_1648),
.B(n_404),
.Y(n_2082)
);

INVxp67_ASAP7_75t_SL g2083 ( 
.A(n_1734),
.Y(n_2083)
);

INVx1_ASAP7_75t_L g2084 ( 
.A(n_1795),
.Y(n_2084)
);

NAND2x1p5_ASAP7_75t_L g2085 ( 
.A(n_1734),
.B(n_405),
.Y(n_2085)
);

NAND2xp5_ASAP7_75t_L g2086 ( 
.A(n_1675),
.B(n_406),
.Y(n_2086)
);

INVx2_ASAP7_75t_L g2087 ( 
.A(n_1602),
.Y(n_2087)
);

HB1xp67_ASAP7_75t_L g2088 ( 
.A(n_1800),
.Y(n_2088)
);

A2O1A1Ixp33_ASAP7_75t_L g2089 ( 
.A1(n_1703),
.A2(n_408),
.B(n_406),
.C(n_407),
.Y(n_2089)
);

OAI21x1_ASAP7_75t_L g2090 ( 
.A1(n_1706),
.A2(n_408),
.B(n_409),
.Y(n_2090)
);

NAND2xp5_ASAP7_75t_L g2091 ( 
.A(n_1675),
.B(n_409),
.Y(n_2091)
);

AOI21xp33_ASAP7_75t_L g2092 ( 
.A1(n_1742),
.A2(n_410),
.B(n_411),
.Y(n_2092)
);

BUFx6f_ASAP7_75t_L g2093 ( 
.A(n_1643),
.Y(n_2093)
);

NAND2xp5_ASAP7_75t_SL g2094 ( 
.A(n_1800),
.B(n_410),
.Y(n_2094)
);

INVx2_ASAP7_75t_L g2095 ( 
.A(n_1602),
.Y(n_2095)
);

NAND3xp33_ASAP7_75t_L g2096 ( 
.A(n_1701),
.B(n_411),
.C(n_412),
.Y(n_2096)
);

NOR2xp33_ASAP7_75t_L g2097 ( 
.A(n_1800),
.B(n_413),
.Y(n_2097)
);

INVx1_ASAP7_75t_L g2098 ( 
.A(n_1795),
.Y(n_2098)
);

NAND2xp5_ASAP7_75t_SL g2099 ( 
.A(n_1800),
.B(n_414),
.Y(n_2099)
);

A2O1A1Ixp33_ASAP7_75t_L g2100 ( 
.A1(n_1703),
.A2(n_416),
.B(n_414),
.C(n_415),
.Y(n_2100)
);

OAI21x1_ASAP7_75t_SL g2101 ( 
.A1(n_1757),
.A2(n_415),
.B(n_416),
.Y(n_2101)
);

AND2x2_ASAP7_75t_L g2102 ( 
.A(n_1578),
.B(n_417),
.Y(n_2102)
);

NAND2xp5_ASAP7_75t_L g2103 ( 
.A(n_1675),
.B(n_420),
.Y(n_2103)
);

OAI21x1_ASAP7_75t_L g2104 ( 
.A1(n_1706),
.A2(n_421),
.B(n_423),
.Y(n_2104)
);

NAND2xp5_ASAP7_75t_L g2105 ( 
.A(n_1675),
.B(n_424),
.Y(n_2105)
);

NAND2xp5_ASAP7_75t_L g2106 ( 
.A(n_1675),
.B(n_424),
.Y(n_2106)
);

INVx1_ASAP7_75t_L g2107 ( 
.A(n_1795),
.Y(n_2107)
);

NOR3xp33_ASAP7_75t_L g2108 ( 
.A(n_1740),
.B(n_427),
.C(n_428),
.Y(n_2108)
);

NAND2xp5_ASAP7_75t_L g2109 ( 
.A(n_1675),
.B(n_427),
.Y(n_2109)
);

AO22x2_ASAP7_75t_L g2110 ( 
.A1(n_1791),
.A2(n_428),
.B1(n_429),
.B2(n_430),
.Y(n_2110)
);

OAI21xp5_ASAP7_75t_SL g2111 ( 
.A1(n_1800),
.A2(n_429),
.B(n_431),
.Y(n_2111)
);

A2O1A1Ixp33_ASAP7_75t_L g2112 ( 
.A1(n_1703),
.A2(n_432),
.B(n_433),
.C(n_434),
.Y(n_2112)
);

CKINVDCx5p33_ASAP7_75t_R g2113 ( 
.A(n_1648),
.Y(n_2113)
);

OAI21x1_ASAP7_75t_L g2114 ( 
.A1(n_1706),
.A2(n_432),
.B(n_433),
.Y(n_2114)
);

AND2x2_ASAP7_75t_L g2115 ( 
.A(n_1578),
.B(n_436),
.Y(n_2115)
);

OR2x2_ASAP7_75t_L g2116 ( 
.A(n_1800),
.B(n_436),
.Y(n_2116)
);

A2O1A1Ixp33_ASAP7_75t_L g2117 ( 
.A1(n_1703),
.A2(n_437),
.B(n_438),
.C(n_439),
.Y(n_2117)
);

OAI21x1_ASAP7_75t_L g2118 ( 
.A1(n_1706),
.A2(n_440),
.B(n_441),
.Y(n_2118)
);

INVx1_ASAP7_75t_L g2119 ( 
.A(n_1795),
.Y(n_2119)
);

NAND3xp33_ASAP7_75t_L g2120 ( 
.A(n_1701),
.B(n_440),
.C(n_442),
.Y(n_2120)
);

INVx2_ASAP7_75t_L g2121 ( 
.A(n_1602),
.Y(n_2121)
);

INVx1_ASAP7_75t_L g2122 ( 
.A(n_1795),
.Y(n_2122)
);

INVx2_ASAP7_75t_L g2123 ( 
.A(n_1602),
.Y(n_2123)
);

BUFx3_ASAP7_75t_L g2124 ( 
.A(n_1648),
.Y(n_2124)
);

INVx1_ASAP7_75t_L g2125 ( 
.A(n_1795),
.Y(n_2125)
);

INVx1_ASAP7_75t_L g2126 ( 
.A(n_1795),
.Y(n_2126)
);

AND2x2_ASAP7_75t_L g2127 ( 
.A(n_1578),
.B(n_445),
.Y(n_2127)
);

AO21x1_ASAP7_75t_L g2128 ( 
.A1(n_1757),
.A2(n_446),
.B(n_447),
.Y(n_2128)
);

A2O1A1Ixp33_ASAP7_75t_L g2129 ( 
.A1(n_1703),
.A2(n_446),
.B(n_447),
.C(n_448),
.Y(n_2129)
);

HB1xp67_ASAP7_75t_L g2130 ( 
.A(n_1800),
.Y(n_2130)
);

NAND2xp5_ASAP7_75t_L g2131 ( 
.A(n_1675),
.B(n_448),
.Y(n_2131)
);

NAND3xp33_ASAP7_75t_L g2132 ( 
.A(n_1701),
.B(n_449),
.C(n_450),
.Y(n_2132)
);

AND2x2_ASAP7_75t_L g2133 ( 
.A(n_1578),
.B(n_449),
.Y(n_2133)
);

OAI21xp5_ASAP7_75t_L g2134 ( 
.A1(n_1631),
.A2(n_450),
.B(n_451),
.Y(n_2134)
);

NAND2xp5_ASAP7_75t_L g2135 ( 
.A(n_1675),
.B(n_451),
.Y(n_2135)
);

OAI21x1_ASAP7_75t_L g2136 ( 
.A1(n_1706),
.A2(n_452),
.B(n_453),
.Y(n_2136)
);

NAND2xp5_ASAP7_75t_L g2137 ( 
.A(n_1675),
.B(n_454),
.Y(n_2137)
);

INVx2_ASAP7_75t_L g2138 ( 
.A(n_1602),
.Y(n_2138)
);

NAND2xp5_ASAP7_75t_L g2139 ( 
.A(n_1675),
.B(n_456),
.Y(n_2139)
);

OA21x2_ASAP7_75t_L g2140 ( 
.A1(n_1796),
.A2(n_456),
.B(n_457),
.Y(n_2140)
);

A2O1A1Ixp33_ASAP7_75t_L g2141 ( 
.A1(n_1703),
.A2(n_457),
.B(n_458),
.C(n_459),
.Y(n_2141)
);

OAI21xp5_ASAP7_75t_L g2142 ( 
.A1(n_1631),
.A2(n_460),
.B(n_461),
.Y(n_2142)
);

A2O1A1Ixp33_ASAP7_75t_L g2143 ( 
.A1(n_1703),
.A2(n_462),
.B(n_463),
.C(n_464),
.Y(n_2143)
);

NAND2xp5_ASAP7_75t_L g2144 ( 
.A(n_1675),
.B(n_462),
.Y(n_2144)
);

NAND2xp5_ASAP7_75t_L g2145 ( 
.A(n_1675),
.B(n_465),
.Y(n_2145)
);

O2A1O1Ixp33_ASAP7_75t_L g2146 ( 
.A1(n_1614),
.A2(n_465),
.B(n_466),
.C(n_467),
.Y(n_2146)
);

NAND2xp5_ASAP7_75t_SL g2147 ( 
.A(n_1800),
.B(n_466),
.Y(n_2147)
);

BUFx6f_ASAP7_75t_L g2148 ( 
.A(n_1643),
.Y(n_2148)
);

BUFx4f_ASAP7_75t_L g2149 ( 
.A(n_1648),
.Y(n_2149)
);

NAND2xp5_ASAP7_75t_L g2150 ( 
.A(n_1675),
.B(n_470),
.Y(n_2150)
);

NAND2xp5_ASAP7_75t_L g2151 ( 
.A(n_1675),
.B(n_472),
.Y(n_2151)
);

OAI21xp5_ASAP7_75t_SL g2152 ( 
.A1(n_1800),
.A2(n_473),
.B(n_474),
.Y(n_2152)
);

NAND2xp5_ASAP7_75t_L g2153 ( 
.A(n_1675),
.B(n_475),
.Y(n_2153)
);

NAND2xp5_ASAP7_75t_L g2154 ( 
.A(n_1675),
.B(n_475),
.Y(n_2154)
);

INVx2_ASAP7_75t_SL g2155 ( 
.A(n_1647),
.Y(n_2155)
);

NAND2xp5_ASAP7_75t_L g2156 ( 
.A(n_1675),
.B(n_478),
.Y(n_2156)
);

OAI22x1_ASAP7_75t_L g2157 ( 
.A1(n_1657),
.A2(n_480),
.B1(n_481),
.B2(n_483),
.Y(n_2157)
);

INVx2_ASAP7_75t_L g2158 ( 
.A(n_1602),
.Y(n_2158)
);

INVx2_ASAP7_75t_L g2159 ( 
.A(n_1602),
.Y(n_2159)
);

INVx3_ASAP7_75t_L g2160 ( 
.A(n_1734),
.Y(n_2160)
);

CKINVDCx20_ASAP7_75t_R g2161 ( 
.A(n_1646),
.Y(n_2161)
);

NOR2xp33_ASAP7_75t_L g2162 ( 
.A(n_1800),
.B(n_484),
.Y(n_2162)
);

OA21x2_ASAP7_75t_L g2163 ( 
.A1(n_1796),
.A2(n_485),
.B(n_486),
.Y(n_2163)
);

A2O1A1Ixp33_ASAP7_75t_L g2164 ( 
.A1(n_1703),
.A2(n_486),
.B(n_487),
.C(n_488),
.Y(n_2164)
);

NAND2xp5_ASAP7_75t_L g2165 ( 
.A(n_1675),
.B(n_489),
.Y(n_2165)
);

INVx5_ASAP7_75t_L g2166 ( 
.A(n_1734),
.Y(n_2166)
);

NAND2xp5_ASAP7_75t_L g2167 ( 
.A(n_1675),
.B(n_491),
.Y(n_2167)
);

NOR2xp33_ASAP7_75t_L g2168 ( 
.A(n_1800),
.B(n_493),
.Y(n_2168)
);

AND2x2_ASAP7_75t_L g2169 ( 
.A(n_1578),
.B(n_494),
.Y(n_2169)
);

AND2x6_ASAP7_75t_L g2170 ( 
.A(n_1707),
.B(n_495),
.Y(n_2170)
);

OAI21xp5_ASAP7_75t_L g2171 ( 
.A1(n_1631),
.A2(n_495),
.B(n_496),
.Y(n_2171)
);

AO31x2_ASAP7_75t_L g2172 ( 
.A1(n_1718),
.A2(n_496),
.A3(n_497),
.B(n_498),
.Y(n_2172)
);

NAND2x1p5_ASAP7_75t_L g2173 ( 
.A(n_1734),
.B(n_499),
.Y(n_2173)
);

NAND2xp5_ASAP7_75t_L g2174 ( 
.A(n_1675),
.B(n_500),
.Y(n_2174)
);

OAI21xp5_ASAP7_75t_L g2175 ( 
.A1(n_1631),
.A2(n_501),
.B(n_502),
.Y(n_2175)
);

OAI21x1_ASAP7_75t_SL g2176 ( 
.A1(n_1757),
.A2(n_501),
.B(n_502),
.Y(n_2176)
);

INVx3_ASAP7_75t_L g2177 ( 
.A(n_1734),
.Y(n_2177)
);

NAND2xp5_ASAP7_75t_SL g2178 ( 
.A(n_1800),
.B(n_503),
.Y(n_2178)
);

AO31x2_ASAP7_75t_L g2179 ( 
.A1(n_1718),
.A2(n_504),
.A3(n_506),
.B(n_507),
.Y(n_2179)
);

OAI21x1_ASAP7_75t_L g2180 ( 
.A1(n_1706),
.A2(n_504),
.B(n_508),
.Y(n_2180)
);

OAI21xp5_ASAP7_75t_L g2181 ( 
.A1(n_1631),
.A2(n_509),
.B(n_510),
.Y(n_2181)
);

INVx1_ASAP7_75t_L g2182 ( 
.A(n_1795),
.Y(n_2182)
);

OAI21x1_ASAP7_75t_L g2183 ( 
.A1(n_1706),
.A2(n_510),
.B(n_511),
.Y(n_2183)
);

AOI21xp5_ASAP7_75t_L g2184 ( 
.A1(n_1631),
.A2(n_512),
.B(n_513),
.Y(n_2184)
);

NAND2xp5_ASAP7_75t_L g2185 ( 
.A(n_1675),
.B(n_512),
.Y(n_2185)
);

OAI21x1_ASAP7_75t_L g2186 ( 
.A1(n_1706),
.A2(n_513),
.B(n_514),
.Y(n_2186)
);

NAND2xp5_ASAP7_75t_SL g2187 ( 
.A(n_1800),
.B(n_515),
.Y(n_2187)
);

INVx1_ASAP7_75t_L g2188 ( 
.A(n_1795),
.Y(n_2188)
);

AOI21xp5_ASAP7_75t_SL g2189 ( 
.A1(n_1707),
.A2(n_516),
.B(n_518),
.Y(n_2189)
);

AND2x4_ASAP7_75t_L g2190 ( 
.A(n_1811),
.B(n_518),
.Y(n_2190)
);

NAND2xp5_ASAP7_75t_L g2191 ( 
.A(n_1675),
.B(n_519),
.Y(n_2191)
);

NOR2xp33_ASAP7_75t_L g2192 ( 
.A(n_1800),
.B(n_520),
.Y(n_2192)
);

NAND2xp5_ASAP7_75t_L g2193 ( 
.A(n_1675),
.B(n_520),
.Y(n_2193)
);

HB1xp67_ASAP7_75t_L g2194 ( 
.A(n_1800),
.Y(n_2194)
);

NAND2xp5_ASAP7_75t_L g2195 ( 
.A(n_1675),
.B(n_521),
.Y(n_2195)
);

INVx2_ASAP7_75t_L g2196 ( 
.A(n_1602),
.Y(n_2196)
);

OA21x2_ASAP7_75t_L g2197 ( 
.A1(n_1890),
.A2(n_523),
.B(n_524),
.Y(n_2197)
);

BUFx2_ASAP7_75t_L g2198 ( 
.A(n_1889),
.Y(n_2198)
);

OA21x2_ASAP7_75t_L g2199 ( 
.A1(n_2002),
.A2(n_525),
.B(n_527),
.Y(n_2199)
);

AO21x2_ASAP7_75t_L g2200 ( 
.A1(n_1850),
.A2(n_2101),
.B(n_2075),
.Y(n_2200)
);

BUFx2_ASAP7_75t_R g2201 ( 
.A(n_1878),
.Y(n_2201)
);

BUFx5_ASAP7_75t_L g2202 ( 
.A(n_2170),
.Y(n_2202)
);

AOI22x1_ASAP7_75t_L g2203 ( 
.A1(n_1970),
.A2(n_529),
.B1(n_530),
.B2(n_531),
.Y(n_2203)
);

BUFx3_ASAP7_75t_L g2204 ( 
.A(n_2040),
.Y(n_2204)
);

CKINVDCx5p33_ASAP7_75t_R g2205 ( 
.A(n_1835),
.Y(n_2205)
);

CKINVDCx11_ASAP7_75t_R g2206 ( 
.A(n_2161),
.Y(n_2206)
);

NAND2xp5_ASAP7_75t_L g2207 ( 
.A(n_1984),
.B(n_532),
.Y(n_2207)
);

INVx6_ASAP7_75t_L g2208 ( 
.A(n_2166),
.Y(n_2208)
);

AO21x2_ASAP7_75t_L g2209 ( 
.A1(n_2176),
.A2(n_534),
.B(n_536),
.Y(n_2209)
);

INVx1_ASAP7_75t_L g2210 ( 
.A(n_1914),
.Y(n_2210)
);

AO21x2_ASAP7_75t_L g2211 ( 
.A1(n_1946),
.A2(n_537),
.B(n_538),
.Y(n_2211)
);

BUFx3_ASAP7_75t_L g2212 ( 
.A(n_2040),
.Y(n_2212)
);

INVx1_ASAP7_75t_L g2213 ( 
.A(n_1919),
.Y(n_2213)
);

NAND3xp33_ASAP7_75t_L g2214 ( 
.A(n_1843),
.B(n_538),
.C(n_539),
.Y(n_2214)
);

OAI21x1_ASAP7_75t_L g2215 ( 
.A1(n_1830),
.A2(n_539),
.B(n_540),
.Y(n_2215)
);

INVx1_ASAP7_75t_L g2216 ( 
.A(n_1919),
.Y(n_2216)
);

AO21x2_ASAP7_75t_L g2217 ( 
.A1(n_2002),
.A2(n_542),
.B(n_543),
.Y(n_2217)
);

AND2x4_ASAP7_75t_L g2218 ( 
.A(n_1971),
.B(n_630),
.Y(n_2218)
);

OAI21x1_ASAP7_75t_L g2219 ( 
.A1(n_1884),
.A2(n_543),
.B(n_545),
.Y(n_2219)
);

AO21x2_ASAP7_75t_L g2220 ( 
.A1(n_1838),
.A2(n_547),
.B(n_549),
.Y(n_2220)
);

AO21x1_ASAP7_75t_L g2221 ( 
.A1(n_2064),
.A2(n_2071),
.B(n_2134),
.Y(n_2221)
);

INVx1_ASAP7_75t_L g2222 ( 
.A(n_1920),
.Y(n_2222)
);

NAND2x1p5_ASAP7_75t_L g2223 ( 
.A(n_1889),
.B(n_547),
.Y(n_2223)
);

INVx1_ASAP7_75t_L g2224 ( 
.A(n_1920),
.Y(n_2224)
);

BUFx3_ASAP7_75t_L g2225 ( 
.A(n_2040),
.Y(n_2225)
);

AOI21x1_ASAP7_75t_L g2226 ( 
.A1(n_1940),
.A2(n_550),
.B(n_552),
.Y(n_2226)
);

AND2x2_ASAP7_75t_L g2227 ( 
.A(n_1911),
.B(n_628),
.Y(n_2227)
);

NOR2x1_ASAP7_75t_R g2228 ( 
.A(n_2113),
.B(n_550),
.Y(n_2228)
);

OAI21x1_ASAP7_75t_L g2229 ( 
.A1(n_1989),
.A2(n_552),
.B(n_553),
.Y(n_2229)
);

INVx6_ASAP7_75t_L g2230 ( 
.A(n_2166),
.Y(n_2230)
);

INVx1_ASAP7_75t_L g2231 ( 
.A(n_1947),
.Y(n_2231)
);

CKINVDCx5p33_ASAP7_75t_R g2232 ( 
.A(n_1835),
.Y(n_2232)
);

BUFx3_ASAP7_75t_L g2233 ( 
.A(n_2166),
.Y(n_2233)
);

INVx1_ASAP7_75t_L g2234 ( 
.A(n_1967),
.Y(n_2234)
);

OAI21x1_ASAP7_75t_L g2235 ( 
.A1(n_1849),
.A2(n_553),
.B(n_554),
.Y(n_2235)
);

INVx1_ASAP7_75t_L g2236 ( 
.A(n_1978),
.Y(n_2236)
);

CKINVDCx6p67_ASAP7_75t_R g2237 ( 
.A(n_2124),
.Y(n_2237)
);

INVx3_ASAP7_75t_L g2238 ( 
.A(n_2005),
.Y(n_2238)
);

INVx3_ASAP7_75t_L g2239 ( 
.A(n_2005),
.Y(n_2239)
);

OA21x2_ASAP7_75t_L g2240 ( 
.A1(n_1893),
.A2(n_554),
.B(n_556),
.Y(n_2240)
);

AND2x4_ASAP7_75t_L g2241 ( 
.A(n_2046),
.B(n_556),
.Y(n_2241)
);

BUFx2_ASAP7_75t_L g2242 ( 
.A(n_1858),
.Y(n_2242)
);

OAI21x1_ASAP7_75t_SL g2243 ( 
.A1(n_1949),
.A2(n_2028),
.B(n_1905),
.Y(n_2243)
);

AND2x2_ASAP7_75t_L g2244 ( 
.A(n_2087),
.B(n_627),
.Y(n_2244)
);

NAND2xp5_ASAP7_75t_L g2245 ( 
.A(n_1991),
.B(n_557),
.Y(n_2245)
);

AOI22xp33_ASAP7_75t_L g2246 ( 
.A1(n_1842),
.A2(n_559),
.B1(n_561),
.B2(n_562),
.Y(n_2246)
);

OAI21xp5_ASAP7_75t_L g2247 ( 
.A1(n_1892),
.A2(n_564),
.B(n_565),
.Y(n_2247)
);

AO21x2_ASAP7_75t_L g2248 ( 
.A1(n_1838),
.A2(n_564),
.B(n_565),
.Y(n_2248)
);

AO21x2_ASAP7_75t_L g2249 ( 
.A1(n_2128),
.A2(n_566),
.B(n_567),
.Y(n_2249)
);

AOI21xp33_ASAP7_75t_SL g2250 ( 
.A1(n_1992),
.A2(n_566),
.B(n_567),
.Y(n_2250)
);

HB1xp67_ASAP7_75t_L g2251 ( 
.A(n_2031),
.Y(n_2251)
);

AO21x2_ASAP7_75t_L g2252 ( 
.A1(n_2134),
.A2(n_568),
.B(n_569),
.Y(n_2252)
);

OAI21xp5_ASAP7_75t_L g2253 ( 
.A1(n_2001),
.A2(n_568),
.B(n_569),
.Y(n_2253)
);

AND2x2_ASAP7_75t_L g2254 ( 
.A(n_2095),
.B(n_570),
.Y(n_2254)
);

OAI21xp5_ASAP7_75t_L g2255 ( 
.A1(n_2001),
.A2(n_570),
.B(n_571),
.Y(n_2255)
);

AO21x2_ASAP7_75t_L g2256 ( 
.A1(n_2142),
.A2(n_2175),
.B(n_2171),
.Y(n_2256)
);

NAND2xp5_ASAP7_75t_L g2257 ( 
.A(n_1960),
.B(n_571),
.Y(n_2257)
);

AOI22xp5_ASAP7_75t_L g2258 ( 
.A1(n_1853),
.A2(n_572),
.B1(n_573),
.B2(n_574),
.Y(n_2258)
);

INVx4_ASAP7_75t_L g2259 ( 
.A(n_2166),
.Y(n_2259)
);

BUFx3_ASAP7_75t_L g2260 ( 
.A(n_1854),
.Y(n_2260)
);

HB1xp67_ASAP7_75t_L g2261 ( 
.A(n_2088),
.Y(n_2261)
);

HB1xp67_ASAP7_75t_L g2262 ( 
.A(n_2130),
.Y(n_2262)
);

INVx1_ASAP7_75t_SL g2263 ( 
.A(n_2194),
.Y(n_2263)
);

INVx1_ASAP7_75t_L g2264 ( 
.A(n_1990),
.Y(n_2264)
);

CKINVDCx14_ASAP7_75t_R g2265 ( 
.A(n_2149),
.Y(n_2265)
);

OAI21xp5_ASAP7_75t_L g2266 ( 
.A1(n_1833),
.A2(n_575),
.B(n_576),
.Y(n_2266)
);

OR2x2_ASAP7_75t_L g2267 ( 
.A(n_1886),
.B(n_578),
.Y(n_2267)
);

INVx1_ASAP7_75t_L g2268 ( 
.A(n_1953),
.Y(n_2268)
);

BUFx12f_ASAP7_75t_L g2269 ( 
.A(n_1912),
.Y(n_2269)
);

OA21x2_ASAP7_75t_L g2270 ( 
.A1(n_2142),
.A2(n_578),
.B(n_579),
.Y(n_2270)
);

INVx2_ASAP7_75t_L g2271 ( 
.A(n_2121),
.Y(n_2271)
);

OAI21x1_ASAP7_75t_L g2272 ( 
.A1(n_1836),
.A2(n_579),
.B(n_580),
.Y(n_2272)
);

INVx2_ASAP7_75t_L g2273 ( 
.A(n_2123),
.Y(n_2273)
);

INVx1_ASAP7_75t_L g2274 ( 
.A(n_1955),
.Y(n_2274)
);

INVx2_ASAP7_75t_L g2275 ( 
.A(n_2138),
.Y(n_2275)
);

INVx2_ASAP7_75t_L g2276 ( 
.A(n_2158),
.Y(n_2276)
);

BUFx2_ASAP7_75t_L g2277 ( 
.A(n_1854),
.Y(n_2277)
);

AO31x2_ASAP7_75t_L g2278 ( 
.A1(n_1950),
.A2(n_581),
.A3(n_582),
.B(n_583),
.Y(n_2278)
);

CKINVDCx5p33_ASAP7_75t_R g2279 ( 
.A(n_2149),
.Y(n_2279)
);

BUFx2_ASAP7_75t_L g2280 ( 
.A(n_1854),
.Y(n_2280)
);

INVx6_ASAP7_75t_L g2281 ( 
.A(n_1948),
.Y(n_2281)
);

NAND2x1p5_ASAP7_75t_L g2282 ( 
.A(n_1928),
.B(n_582),
.Y(n_2282)
);

INVx1_ASAP7_75t_L g2283 ( 
.A(n_2159),
.Y(n_2283)
);

NAND2xp5_ASAP7_75t_L g2284 ( 
.A(n_1960),
.B(n_584),
.Y(n_2284)
);

INVx2_ASAP7_75t_L g2285 ( 
.A(n_2196),
.Y(n_2285)
);

NAND3xp33_ASAP7_75t_L g2286 ( 
.A(n_1867),
.B(n_2108),
.C(n_1975),
.Y(n_2286)
);

CKINVDCx8_ASAP7_75t_R g2287 ( 
.A(n_2170),
.Y(n_2287)
);

OAI22xp5_ASAP7_75t_L g2288 ( 
.A1(n_1928),
.A2(n_585),
.B1(n_587),
.B2(n_588),
.Y(n_2288)
);

AO21x2_ASAP7_75t_L g2289 ( 
.A1(n_2171),
.A2(n_587),
.B(n_588),
.Y(n_2289)
);

AND2x4_ASAP7_75t_L g2290 ( 
.A(n_1844),
.B(n_591),
.Y(n_2290)
);

HB1xp67_ASAP7_75t_L g2291 ( 
.A(n_1832),
.Y(n_2291)
);

AOI22xp33_ASAP7_75t_L g2292 ( 
.A1(n_1859),
.A2(n_594),
.B1(n_595),
.B2(n_597),
.Y(n_2292)
);

INVx1_ASAP7_75t_SL g2293 ( 
.A(n_2018),
.Y(n_2293)
);

AO21x2_ASAP7_75t_L g2294 ( 
.A1(n_2175),
.A2(n_594),
.B(n_599),
.Y(n_2294)
);

INVx6_ASAP7_75t_L g2295 ( 
.A(n_1966),
.Y(n_2295)
);

OA21x2_ASAP7_75t_L g2296 ( 
.A1(n_2181),
.A2(n_1940),
.B(n_2078),
.Y(n_2296)
);

INVx1_ASAP7_75t_L g2297 ( 
.A(n_2110),
.Y(n_2297)
);

BUFx6f_ASAP7_75t_SL g2298 ( 
.A(n_2170),
.Y(n_2298)
);

A2O1A1Ixp33_ASAP7_75t_L g2299 ( 
.A1(n_2146),
.A2(n_600),
.B(n_601),
.C(n_602),
.Y(n_2299)
);

BUFx2_ASAP7_75t_SL g2300 ( 
.A(n_1983),
.Y(n_2300)
);

OAI21x1_ASAP7_75t_L g2301 ( 
.A1(n_2090),
.A2(n_600),
.B(n_601),
.Y(n_2301)
);

OR2x6_ASAP7_75t_L g2302 ( 
.A(n_2025),
.B(n_602),
.Y(n_2302)
);

OA21x2_ASAP7_75t_L g2303 ( 
.A1(n_2181),
.A2(n_603),
.B(n_604),
.Y(n_2303)
);

NOR2x1_ASAP7_75t_SL g2304 ( 
.A(n_1969),
.B(n_603),
.Y(n_2304)
);

AOI21x1_ASAP7_75t_L g2305 ( 
.A1(n_2009),
.A2(n_604),
.B(n_605),
.Y(n_2305)
);

INVxp67_ASAP7_75t_SL g2306 ( 
.A(n_1861),
.Y(n_2306)
);

BUFx3_ASAP7_75t_L g2307 ( 
.A(n_1913),
.Y(n_2307)
);

INVx1_ASAP7_75t_SL g2308 ( 
.A(n_1824),
.Y(n_2308)
);

AO21x2_ASAP7_75t_L g2309 ( 
.A1(n_2064),
.A2(n_605),
.B(n_606),
.Y(n_2309)
);

BUFx3_ASAP7_75t_L g2310 ( 
.A(n_1956),
.Y(n_2310)
);

INVx1_ASAP7_75t_L g2311 ( 
.A(n_2110),
.Y(n_2311)
);

OAI21x1_ASAP7_75t_L g2312 ( 
.A1(n_2104),
.A2(n_606),
.B(n_607),
.Y(n_2312)
);

INVx1_ASAP7_75t_L g2313 ( 
.A(n_1846),
.Y(n_2313)
);

INVx1_ASAP7_75t_L g2314 ( 
.A(n_1846),
.Y(n_2314)
);

OAI21x1_ASAP7_75t_L g2315 ( 
.A1(n_2114),
.A2(n_607),
.B(n_608),
.Y(n_2315)
);

INVx2_ASAP7_75t_L g2316 ( 
.A(n_1998),
.Y(n_2316)
);

OR2x2_ASAP7_75t_L g2317 ( 
.A(n_2116),
.B(n_609),
.Y(n_2317)
);

AO31x2_ASAP7_75t_L g2318 ( 
.A1(n_2089),
.A2(n_610),
.A3(n_611),
.B(n_612),
.Y(n_2318)
);

BUFx6f_ASAP7_75t_SL g2319 ( 
.A(n_2170),
.Y(n_2319)
);

CKINVDCx5p33_ASAP7_75t_R g2320 ( 
.A(n_1958),
.Y(n_2320)
);

CKINVDCx20_ASAP7_75t_R g2321 ( 
.A(n_1981),
.Y(n_2321)
);

OAI21xp5_ASAP7_75t_L g2322 ( 
.A1(n_2037),
.A2(n_610),
.B(n_612),
.Y(n_2322)
);

INVx1_ASAP7_75t_SL g2323 ( 
.A(n_1824),
.Y(n_2323)
);

BUFx8_ASAP7_75t_L g2324 ( 
.A(n_1828),
.Y(n_2324)
);

OAI21x1_ASAP7_75t_L g2325 ( 
.A1(n_2118),
.A2(n_613),
.B(n_614),
.Y(n_2325)
);

BUFx3_ASAP7_75t_L g2326 ( 
.A(n_1993),
.Y(n_2326)
);

BUFx3_ASAP7_75t_L g2327 ( 
.A(n_1993),
.Y(n_2327)
);

INVx1_ASAP7_75t_L g2328 ( 
.A(n_1848),
.Y(n_2328)
);

OAI21x1_ASAP7_75t_L g2329 ( 
.A1(n_2136),
.A2(n_615),
.B(n_616),
.Y(n_2329)
);

NAND2xp5_ASAP7_75t_L g2330 ( 
.A(n_2027),
.B(n_617),
.Y(n_2330)
);

AOI22xp5_ASAP7_75t_L g2331 ( 
.A1(n_2056),
.A2(n_617),
.B1(n_618),
.B2(n_619),
.Y(n_2331)
);

OA21x2_ASAP7_75t_L g2332 ( 
.A1(n_2180),
.A2(n_618),
.B(n_620),
.Y(n_2332)
);

OAI21x1_ASAP7_75t_L g2333 ( 
.A1(n_2183),
.A2(n_622),
.B(n_623),
.Y(n_2333)
);

CKINVDCx6p67_ASAP7_75t_R g2334 ( 
.A(n_1981),
.Y(n_2334)
);

AO21x2_ASAP7_75t_L g2335 ( 
.A1(n_2023),
.A2(n_622),
.B(n_623),
.Y(n_2335)
);

INVx1_ASAP7_75t_L g2336 ( 
.A(n_1848),
.Y(n_2336)
);

NAND2x1p5_ASAP7_75t_L g2337 ( 
.A(n_2160),
.B(n_624),
.Y(n_2337)
);

INVx2_ASAP7_75t_L g2338 ( 
.A(n_2013),
.Y(n_2338)
);

NAND2xp5_ASAP7_75t_L g2339 ( 
.A(n_1959),
.B(n_626),
.Y(n_2339)
);

AO21x2_ASAP7_75t_L g2340 ( 
.A1(n_2023),
.A2(n_624),
.B(n_625),
.Y(n_2340)
);

OAI21x1_ASAP7_75t_L g2341 ( 
.A1(n_2186),
.A2(n_625),
.B(n_626),
.Y(n_2341)
);

INVx2_ASAP7_75t_L g2342 ( 
.A(n_2069),
.Y(n_2342)
);

BUFx3_ASAP7_75t_L g2343 ( 
.A(n_2069),
.Y(n_2343)
);

INVx1_ASAP7_75t_L g2344 ( 
.A(n_1921),
.Y(n_2344)
);

BUFx2_ASAP7_75t_SL g2345 ( 
.A(n_1825),
.Y(n_2345)
);

HB1xp67_ASAP7_75t_SL g2346 ( 
.A(n_1936),
.Y(n_2346)
);

INVx2_ASAP7_75t_L g2347 ( 
.A(n_2093),
.Y(n_2347)
);

BUFx2_ASAP7_75t_R g2348 ( 
.A(n_2000),
.Y(n_2348)
);

AO21x2_ASAP7_75t_L g2349 ( 
.A1(n_2071),
.A2(n_1999),
.B(n_1852),
.Y(n_2349)
);

OR2x6_ASAP7_75t_L g2350 ( 
.A(n_2025),
.B(n_1861),
.Y(n_2350)
);

INVx1_ASAP7_75t_L g2351 ( 
.A(n_1921),
.Y(n_2351)
);

BUFx3_ASAP7_75t_L g2352 ( 
.A(n_2093),
.Y(n_2352)
);

OR2x2_ASAP7_75t_L g2353 ( 
.A(n_1902),
.B(n_1904),
.Y(n_2353)
);

INVx1_ASAP7_75t_L g2354 ( 
.A(n_1995),
.Y(n_2354)
);

BUFx8_ASAP7_75t_SL g2355 ( 
.A(n_1963),
.Y(n_2355)
);

AND2x2_ASAP7_75t_L g2356 ( 
.A(n_1909),
.B(n_2004),
.Y(n_2356)
);

BUFx3_ASAP7_75t_L g2357 ( 
.A(n_2148),
.Y(n_2357)
);

BUFx2_ASAP7_75t_SL g2358 ( 
.A(n_1825),
.Y(n_2358)
);

INVx1_ASAP7_75t_L g2359 ( 
.A(n_1995),
.Y(n_2359)
);

HB1xp67_ASAP7_75t_L g2360 ( 
.A(n_2190),
.Y(n_2360)
);

INVx1_ASAP7_75t_L g2361 ( 
.A(n_2016),
.Y(n_2361)
);

INVx1_ASAP7_75t_L g2362 ( 
.A(n_2016),
.Y(n_2362)
);

BUFx3_ASAP7_75t_L g2363 ( 
.A(n_2148),
.Y(n_2363)
);

BUFx2_ASAP7_75t_SL g2364 ( 
.A(n_2190),
.Y(n_2364)
);

INVx3_ASAP7_75t_L g2365 ( 
.A(n_2074),
.Y(n_2365)
);

NAND2xp5_ASAP7_75t_L g2366 ( 
.A(n_1959),
.B(n_2072),
.Y(n_2366)
);

BUFx3_ASAP7_75t_L g2367 ( 
.A(n_2160),
.Y(n_2367)
);

INVx1_ASAP7_75t_L g2368 ( 
.A(n_1870),
.Y(n_2368)
);

BUFx3_ASAP7_75t_L g2369 ( 
.A(n_2177),
.Y(n_2369)
);

NAND2xp5_ASAP7_75t_L g2370 ( 
.A(n_1951),
.B(n_1945),
.Y(n_2370)
);

BUFx6f_ASAP7_75t_L g2371 ( 
.A(n_2177),
.Y(n_2371)
);

CKINVDCx20_ASAP7_75t_R g2372 ( 
.A(n_1831),
.Y(n_2372)
);

AND2x4_ASAP7_75t_L g2373 ( 
.A(n_1845),
.B(n_1847),
.Y(n_2373)
);

INVxp67_ASAP7_75t_L g2374 ( 
.A(n_2102),
.Y(n_2374)
);

AO21x2_ASAP7_75t_L g2375 ( 
.A1(n_1999),
.A2(n_1852),
.B(n_2055),
.Y(n_2375)
);

OAI21x1_ASAP7_75t_SL g2376 ( 
.A1(n_1895),
.A2(n_1905),
.B(n_1876),
.Y(n_2376)
);

NOR2xp67_ASAP7_75t_L g2377 ( 
.A(n_2081),
.B(n_2155),
.Y(n_2377)
);

BUFx6f_ASAP7_75t_L g2378 ( 
.A(n_2074),
.Y(n_2378)
);

AND2x2_ASAP7_75t_L g2379 ( 
.A(n_1869),
.B(n_1875),
.Y(n_2379)
);

AO21x2_ASAP7_75t_L g2380 ( 
.A1(n_2055),
.A2(n_1895),
.B(n_1937),
.Y(n_2380)
);

BUFx10_ASAP7_75t_L g2381 ( 
.A(n_1963),
.Y(n_2381)
);

INVx1_ASAP7_75t_L g2382 ( 
.A(n_1870),
.Y(n_2382)
);

OAI21x1_ASAP7_75t_L g2383 ( 
.A1(n_2011),
.A2(n_2163),
.B(n_2140),
.Y(n_2383)
);

BUFx2_ASAP7_75t_L g2384 ( 
.A(n_1964),
.Y(n_2384)
);

BUFx2_ASAP7_75t_L g2385 ( 
.A(n_2008),
.Y(n_2385)
);

NOR2xp67_ASAP7_75t_L g2386 ( 
.A(n_1966),
.B(n_1942),
.Y(n_2386)
);

OAI21xp5_ASAP7_75t_L g2387 ( 
.A1(n_2037),
.A2(n_1968),
.B(n_2050),
.Y(n_2387)
);

OAI21xp5_ASAP7_75t_L g2388 ( 
.A1(n_1968),
.A2(n_2050),
.B(n_1901),
.Y(n_2388)
);

OAI21x1_ASAP7_75t_L g2389 ( 
.A1(n_2140),
.A2(n_2163),
.B(n_1866),
.Y(n_2389)
);

HB1xp67_ASAP7_75t_L g2390 ( 
.A(n_1973),
.Y(n_2390)
);

INVx1_ASAP7_75t_L g2391 ( 
.A(n_1871),
.Y(n_2391)
);

BUFx2_ASAP7_75t_L g2392 ( 
.A(n_1918),
.Y(n_2392)
);

OAI21x1_ASAP7_75t_SL g2393 ( 
.A1(n_1876),
.A2(n_1839),
.B(n_1962),
.Y(n_2393)
);

INVx1_ASAP7_75t_L g2394 ( 
.A(n_1871),
.Y(n_2394)
);

AO21x1_ASAP7_75t_L g2395 ( 
.A1(n_1907),
.A2(n_2173),
.B(n_2085),
.Y(n_2395)
);

INVx1_ASAP7_75t_L g2396 ( 
.A(n_1827),
.Y(n_2396)
);

AND2x2_ASAP7_75t_L g2397 ( 
.A(n_2115),
.B(n_2127),
.Y(n_2397)
);

NAND2xp5_ASAP7_75t_L g2398 ( 
.A(n_1985),
.B(n_2070),
.Y(n_2398)
);

BUFx3_ASAP7_75t_L g2399 ( 
.A(n_2060),
.Y(n_2399)
);

HB1xp67_ASAP7_75t_L g2400 ( 
.A(n_1980),
.Y(n_2400)
);

BUFx5_ASAP7_75t_L g2401 ( 
.A(n_1891),
.Y(n_2401)
);

INVx2_ASAP7_75t_SL g2402 ( 
.A(n_2060),
.Y(n_2402)
);

INVx1_ASAP7_75t_L g2403 ( 
.A(n_1827),
.Y(n_2403)
);

INVx1_ASAP7_75t_L g2404 ( 
.A(n_1916),
.Y(n_2404)
);

INVx1_ASAP7_75t_SL g2405 ( 
.A(n_2133),
.Y(n_2405)
);

AOI21x1_ASAP7_75t_L g2406 ( 
.A1(n_2014),
.A2(n_2051),
.B(n_1937),
.Y(n_2406)
);

NOR2xp33_ASAP7_75t_L g2407 ( 
.A(n_2026),
.B(n_2042),
.Y(n_2407)
);

INVx1_ASAP7_75t_L g2408 ( 
.A(n_1916),
.Y(n_2408)
);

NAND2x1p5_ASAP7_75t_L g2409 ( 
.A(n_1837),
.B(n_1972),
.Y(n_2409)
);

INVx1_ASAP7_75t_L g2410 ( 
.A(n_1855),
.Y(n_2410)
);

INVx3_ASAP7_75t_SL g2411 ( 
.A(n_1957),
.Y(n_2411)
);

NOR2xp67_ASAP7_75t_L g2412 ( 
.A(n_1942),
.B(n_1961),
.Y(n_2412)
);

OA21x2_ASAP7_75t_L g2413 ( 
.A1(n_1894),
.A2(n_1897),
.B(n_2184),
.Y(n_2413)
);

BUFx3_ASAP7_75t_L g2414 ( 
.A(n_1972),
.Y(n_2414)
);

NAND2xp5_ASAP7_75t_L g2415 ( 
.A(n_2052),
.B(n_2057),
.Y(n_2415)
);

OAI21x1_ASAP7_75t_L g2416 ( 
.A1(n_2085),
.A2(n_2173),
.B(n_2045),
.Y(n_2416)
);

BUFx12f_ASAP7_75t_L g2417 ( 
.A(n_2034),
.Y(n_2417)
);

NAND2xp5_ASAP7_75t_L g2418 ( 
.A(n_2195),
.B(n_2076),
.Y(n_2418)
);

BUFx2_ASAP7_75t_R g2419 ( 
.A(n_2000),
.Y(n_2419)
);

OAI21x1_ASAP7_75t_SL g2420 ( 
.A1(n_1962),
.A2(n_2065),
.B(n_1879),
.Y(n_2420)
);

BUFx3_ASAP7_75t_L g2421 ( 
.A(n_1976),
.Y(n_2421)
);

OR2x2_ASAP7_75t_L g2422 ( 
.A(n_2048),
.B(n_2169),
.Y(n_2422)
);

BUFx2_ASAP7_75t_L g2423 ( 
.A(n_2083),
.Y(n_2423)
);

NOR2xp33_ASAP7_75t_L g2424 ( 
.A(n_2026),
.B(n_2054),
.Y(n_2424)
);

BUFx2_ASAP7_75t_R g2425 ( 
.A(n_1930),
.Y(n_2425)
);

AO221x1_ASAP7_75t_L g2426 ( 
.A1(n_1922),
.A2(n_2022),
.B1(n_1982),
.B2(n_2021),
.C(n_2036),
.Y(n_2426)
);

OR2x6_ASAP7_75t_L g2427 ( 
.A(n_2039),
.B(n_2047),
.Y(n_2427)
);

NOR2xp67_ASAP7_75t_L g2428 ( 
.A(n_1961),
.B(n_2020),
.Y(n_2428)
);

BUFx3_ASAP7_75t_L g2429 ( 
.A(n_1976),
.Y(n_2429)
);

AOI22x1_ASAP7_75t_L g2430 ( 
.A1(n_2061),
.A2(n_1929),
.B1(n_1931),
.B2(n_1932),
.Y(n_2430)
);

OA21x2_ASAP7_75t_L g2431 ( 
.A1(n_2032),
.A2(n_2030),
.B(n_1925),
.Y(n_2431)
);

BUFx3_ASAP7_75t_L g2432 ( 
.A(n_1957),
.Y(n_2432)
);

NAND2xp5_ASAP7_75t_L g2433 ( 
.A(n_2195),
.B(n_2076),
.Y(n_2433)
);

INVx4_ASAP7_75t_SL g2434 ( 
.A(n_2003),
.Y(n_2434)
);

AOI22x1_ASAP7_75t_L g2435 ( 
.A1(n_1939),
.A2(n_1979),
.B1(n_1977),
.B2(n_1941),
.Y(n_2435)
);

BUFx3_ASAP7_75t_L g2436 ( 
.A(n_1908),
.Y(n_2436)
);

NAND2x1p5_ASAP7_75t_L g2437 ( 
.A(n_1944),
.B(n_2006),
.Y(n_2437)
);

AO21x2_ASAP7_75t_L g2438 ( 
.A1(n_1841),
.A2(n_1879),
.B(n_1874),
.Y(n_2438)
);

AND2x4_ASAP7_75t_L g2439 ( 
.A(n_2080),
.B(n_2084),
.Y(n_2439)
);

NAND2xp5_ASAP7_75t_L g2440 ( 
.A(n_2193),
.B(n_2079),
.Y(n_2440)
);

OAI22xp5_ASAP7_75t_L g2441 ( 
.A1(n_1881),
.A2(n_1882),
.B1(n_1885),
.B2(n_1899),
.Y(n_2441)
);

INVx5_ASAP7_75t_SL g2442 ( 
.A(n_2006),
.Y(n_2442)
);

BUFx8_ASAP7_75t_L g2443 ( 
.A(n_1923),
.Y(n_2443)
);

INVx1_ASAP7_75t_L g2444 ( 
.A(n_1996),
.Y(n_2444)
);

AND2x4_ASAP7_75t_L g2445 ( 
.A(n_2098),
.B(n_2107),
.Y(n_2445)
);

NAND2x1p5_ASAP7_75t_L g2446 ( 
.A(n_2029),
.B(n_1910),
.Y(n_2446)
);

AOI22x1_ASAP7_75t_L g2447 ( 
.A1(n_1954),
.A2(n_1917),
.B1(n_1926),
.B2(n_1927),
.Y(n_2447)
);

AOI21xp5_ASAP7_75t_L g2448 ( 
.A1(n_2119),
.A2(n_2125),
.B(n_2122),
.Y(n_2448)
);

OAI21xp5_ASAP7_75t_L g2449 ( 
.A1(n_2126),
.A2(n_2188),
.B(n_2182),
.Y(n_2449)
);

BUFx3_ASAP7_75t_L g2450 ( 
.A(n_2073),
.Y(n_2450)
);

NAND2xp5_ASAP7_75t_L g2451 ( 
.A(n_2193),
.B(n_2079),
.Y(n_2451)
);

OA21x2_ASAP7_75t_L g2452 ( 
.A1(n_2100),
.A2(n_2129),
.B(n_2117),
.Y(n_2452)
);

AND2x4_ASAP7_75t_L g2453 ( 
.A(n_1988),
.B(n_1896),
.Y(n_2453)
);

BUFx2_ASAP7_75t_L g2454 ( 
.A(n_2066),
.Y(n_2454)
);

OAI21x1_ASAP7_75t_L g2455 ( 
.A1(n_1873),
.A2(n_1857),
.B(n_1860),
.Y(n_2455)
);

INVx5_ASAP7_75t_L g2456 ( 
.A(n_2062),
.Y(n_2456)
);

OAI21x1_ASAP7_75t_L g2457 ( 
.A1(n_1851),
.A2(n_1857),
.B(n_1860),
.Y(n_2457)
);

BUFx3_ASAP7_75t_L g2458 ( 
.A(n_2131),
.Y(n_2458)
);

BUFx3_ASAP7_75t_L g2459 ( 
.A(n_2135),
.Y(n_2459)
);

NAND2xp5_ASAP7_75t_L g2460 ( 
.A(n_2086),
.B(n_2091),
.Y(n_2460)
);

BUFx3_ASAP7_75t_L g2461 ( 
.A(n_2137),
.Y(n_2461)
);

AO21x2_ASAP7_75t_L g2462 ( 
.A1(n_1881),
.A2(n_1882),
.B(n_1885),
.Y(n_2462)
);

AND2x2_ASAP7_75t_L g2463 ( 
.A(n_1924),
.B(n_1952),
.Y(n_2463)
);

NAND2xp5_ASAP7_75t_L g2464 ( 
.A(n_2086),
.B(n_2091),
.Y(n_2464)
);

INVx1_ASAP7_75t_L g2465 ( 
.A(n_1996),
.Y(n_2465)
);

OA21x2_ASAP7_75t_L g2466 ( 
.A1(n_2112),
.A2(n_2141),
.B(n_2143),
.Y(n_2466)
);

AO21x2_ASAP7_75t_L g2467 ( 
.A1(n_1906),
.A2(n_2164),
.B(n_2065),
.Y(n_2467)
);

OA21x2_ASAP7_75t_L g2468 ( 
.A1(n_2012),
.A2(n_1938),
.B(n_1880),
.Y(n_2468)
);

OR2x6_ASAP7_75t_L g2469 ( 
.A(n_1862),
.B(n_2189),
.Y(n_2469)
);

AOI21xp5_ASAP7_75t_L g2470 ( 
.A1(n_1986),
.A2(n_2053),
.B(n_2063),
.Y(n_2470)
);

BUFx3_ASAP7_75t_L g2471 ( 
.A(n_2103),
.Y(n_2471)
);

INVx1_ASAP7_75t_L g2472 ( 
.A(n_1994),
.Y(n_2472)
);

INVx2_ASAP7_75t_SL g2473 ( 
.A(n_1888),
.Y(n_2473)
);

OA21x2_ASAP7_75t_L g2474 ( 
.A1(n_1880),
.A2(n_2041),
.B(n_1924),
.Y(n_2474)
);

NOR2xp33_ASAP7_75t_L g2475 ( 
.A(n_2063),
.B(n_2097),
.Y(n_2475)
);

AO31x2_ASAP7_75t_L g2476 ( 
.A1(n_2157),
.A2(n_2043),
.A3(n_1935),
.B(n_1856),
.Y(n_2476)
);

BUFx3_ASAP7_75t_L g2477 ( 
.A(n_2103),
.Y(n_2477)
);

OAI22xp5_ASAP7_75t_L g2478 ( 
.A1(n_2053),
.A2(n_2150),
.B1(n_2191),
.B2(n_2105),
.Y(n_2478)
);

OAI21x1_ASAP7_75t_L g2479 ( 
.A1(n_2033),
.A2(n_2049),
.B(n_2058),
.Y(n_2479)
);

NAND2xp5_ASAP7_75t_L g2480 ( 
.A(n_2105),
.B(n_2106),
.Y(n_2480)
);

NAND2xp5_ASAP7_75t_L g2481 ( 
.A(n_2106),
.B(n_2109),
.Y(n_2481)
);

INVx1_ASAP7_75t_L g2482 ( 
.A(n_1994),
.Y(n_2482)
);

CKINVDCx5p33_ASAP7_75t_R g2483 ( 
.A(n_1829),
.Y(n_2483)
);

NAND2x1p5_ASAP7_75t_L g2484 ( 
.A(n_2035),
.B(n_2094),
.Y(n_2484)
);

BUFx3_ASAP7_75t_L g2485 ( 
.A(n_2109),
.Y(n_2485)
);

NOR2xp33_ASAP7_75t_L g2486 ( 
.A(n_2162),
.B(n_2168),
.Y(n_2486)
);

OAI21x1_ASAP7_75t_L g2487 ( 
.A1(n_2019),
.A2(n_1974),
.B(n_2059),
.Y(n_2487)
);

OA21x2_ASAP7_75t_L g2488 ( 
.A1(n_1952),
.A2(n_2092),
.B(n_2015),
.Y(n_2488)
);

OAI21x1_ASAP7_75t_L g2489 ( 
.A1(n_2068),
.A2(n_1934),
.B(n_2066),
.Y(n_2489)
);

AO21x2_ASAP7_75t_L g2490 ( 
.A1(n_2068),
.A2(n_2092),
.B(n_1934),
.Y(n_2490)
);

AO21x2_ASAP7_75t_L g2491 ( 
.A1(n_2096),
.A2(n_2120),
.B(n_2132),
.Y(n_2491)
);

OR2x2_ASAP7_75t_SL g2492 ( 
.A(n_1826),
.B(n_2024),
.Y(n_2492)
);

AOI21xp33_ASAP7_75t_L g2493 ( 
.A1(n_1903),
.A2(n_2192),
.B(n_2044),
.Y(n_2493)
);

OAI21x1_ASAP7_75t_L g2494 ( 
.A1(n_2067),
.A2(n_1898),
.B(n_2036),
.Y(n_2494)
);

NAND3xp33_ASAP7_75t_L g2495 ( 
.A(n_1863),
.B(n_1864),
.C(n_1915),
.Y(n_2495)
);

CKINVDCx16_ASAP7_75t_R g2496 ( 
.A(n_2067),
.Y(n_2496)
);

BUFx2_ASAP7_75t_R g2497 ( 
.A(n_2139),
.Y(n_2497)
);

BUFx3_ASAP7_75t_L g2498 ( 
.A(n_2139),
.Y(n_2498)
);

OAI21x1_ASAP7_75t_L g2499 ( 
.A1(n_1982),
.A2(n_2021),
.B(n_1987),
.Y(n_2499)
);

BUFx6f_ASAP7_75t_L g2500 ( 
.A(n_2144),
.Y(n_2500)
);

INVx1_ASAP7_75t_L g2501 ( 
.A(n_1943),
.Y(n_2501)
);

INVx1_ASAP7_75t_L g2502 ( 
.A(n_1943),
.Y(n_2502)
);

NAND2xp5_ASAP7_75t_L g2503 ( 
.A(n_2191),
.B(n_2156),
.Y(n_2503)
);

INVx1_ASAP7_75t_L g2504 ( 
.A(n_1868),
.Y(n_2504)
);

INVx2_ASAP7_75t_R g2505 ( 
.A(n_1933),
.Y(n_2505)
);

INVxp67_ASAP7_75t_SL g2506 ( 
.A(n_2144),
.Y(n_2506)
);

OAI21x1_ASAP7_75t_L g2507 ( 
.A1(n_2043),
.A2(n_2156),
.B(n_2185),
.Y(n_2507)
);

AOI221xp5_ASAP7_75t_L g2508 ( 
.A1(n_2145),
.A2(n_2185),
.B1(n_2174),
.B2(n_2150),
.C(n_2167),
.Y(n_2508)
);

OAI21x1_ASAP7_75t_L g2509 ( 
.A1(n_2145),
.A2(n_2154),
.B(n_2151),
.Y(n_2509)
);

CKINVDCx6p67_ASAP7_75t_R g2510 ( 
.A(n_1883),
.Y(n_2510)
);

OA21x2_ASAP7_75t_L g2511 ( 
.A1(n_2111),
.A2(n_2152),
.B(n_2174),
.Y(n_2511)
);

NOR2xp33_ASAP7_75t_L g2512 ( 
.A(n_2151),
.B(n_2154),
.Y(n_2512)
);

INVx1_ASAP7_75t_L g2513 ( 
.A(n_1900),
.Y(n_2513)
);

OAI21xp5_ASAP7_75t_L g2514 ( 
.A1(n_2153),
.A2(n_2167),
.B(n_2165),
.Y(n_2514)
);

HB1xp67_ASAP7_75t_L g2515 ( 
.A(n_2153),
.Y(n_2515)
);

OAI21x1_ASAP7_75t_L g2516 ( 
.A1(n_2165),
.A2(n_2187),
.B(n_2178),
.Y(n_2516)
);

OR2x2_ASAP7_75t_L g2517 ( 
.A(n_2099),
.B(n_2147),
.Y(n_2517)
);

INVx1_ASAP7_75t_L g2518 ( 
.A(n_1887),
.Y(n_2518)
);

INVx1_ASAP7_75t_SL g2519 ( 
.A(n_1997),
.Y(n_2519)
);

OAI21x1_ASAP7_75t_L g2520 ( 
.A1(n_1840),
.A2(n_2010),
.B(n_2172),
.Y(n_2520)
);

INVx3_ASAP7_75t_L g2521 ( 
.A(n_2017),
.Y(n_2521)
);

OAI21x1_ASAP7_75t_L g2522 ( 
.A1(n_2077),
.A2(n_2179),
.B(n_2172),
.Y(n_2522)
);

OAI21x1_ASAP7_75t_L g2523 ( 
.A1(n_2077),
.A2(n_2179),
.B(n_2017),
.Y(n_2523)
);

BUFx4f_ASAP7_75t_SL g2524 ( 
.A(n_2082),
.Y(n_2524)
);

INVx3_ASAP7_75t_L g2525 ( 
.A(n_2017),
.Y(n_2525)
);

INVx1_ASAP7_75t_SL g2526 ( 
.A(n_1965),
.Y(n_2526)
);

OA21x2_ASAP7_75t_L g2527 ( 
.A1(n_2007),
.A2(n_2038),
.B(n_2003),
.Y(n_2527)
);

AND2x2_ASAP7_75t_L g2528 ( 
.A(n_2007),
.B(n_1887),
.Y(n_2528)
);

AO21x1_ASAP7_75t_L g2529 ( 
.A1(n_1887),
.A2(n_1872),
.B(n_1965),
.Y(n_2529)
);

AO21x2_ASAP7_75t_L g2530 ( 
.A1(n_1965),
.A2(n_1890),
.B(n_1850),
.Y(n_2530)
);

AO21x2_ASAP7_75t_L g2531 ( 
.A1(n_1890),
.A2(n_2075),
.B(n_1850),
.Y(n_2531)
);

BUFx4f_ASAP7_75t_SL g2532 ( 
.A(n_2161),
.Y(n_2532)
);

AOI22xp5_ASAP7_75t_L g2533 ( 
.A1(n_1853),
.A2(n_1284),
.B1(n_1187),
.B2(n_1195),
.Y(n_2533)
);

OAI21x1_ASAP7_75t_L g2534 ( 
.A1(n_1834),
.A2(n_1865),
.B(n_1877),
.Y(n_2534)
);

BUFx3_ASAP7_75t_L g2535 ( 
.A(n_2040),
.Y(n_2535)
);

OR2x2_ASAP7_75t_L g2536 ( 
.A(n_2088),
.B(n_1284),
.Y(n_2536)
);

AO21x2_ASAP7_75t_L g2537 ( 
.A1(n_2534),
.A2(n_2420),
.B(n_2529),
.Y(n_2537)
);

NOR2x1_ASAP7_75t_SL g2538 ( 
.A(n_2302),
.B(n_2345),
.Y(n_2538)
);

OAI22xp33_ASAP7_75t_L g2539 ( 
.A1(n_2496),
.A2(n_2302),
.B1(n_2282),
.B2(n_2287),
.Y(n_2539)
);

OAI21xp5_ASAP7_75t_L g2540 ( 
.A1(n_2507),
.A2(n_2387),
.B(n_2478),
.Y(n_2540)
);

INVx1_ASAP7_75t_L g2541 ( 
.A(n_2379),
.Y(n_2541)
);

AOI21x1_ASAP7_75t_L g2542 ( 
.A1(n_2406),
.A2(n_2518),
.B(n_2389),
.Y(n_2542)
);

NAND2x1p5_ASAP7_75t_L g2543 ( 
.A(n_2259),
.B(n_2204),
.Y(n_2543)
);

AO21x2_ASAP7_75t_L g2544 ( 
.A1(n_2243),
.A2(n_2376),
.B(n_2389),
.Y(n_2544)
);

INVx1_ASAP7_75t_L g2545 ( 
.A(n_2379),
.Y(n_2545)
);

INVx2_ASAP7_75t_L g2546 ( 
.A(n_2271),
.Y(n_2546)
);

AO21x2_ASAP7_75t_L g2547 ( 
.A1(n_2383),
.A2(n_2393),
.B(n_2522),
.Y(n_2547)
);

AO21x2_ASAP7_75t_L g2548 ( 
.A1(n_2383),
.A2(n_2522),
.B(n_2523),
.Y(n_2548)
);

INVx6_ASAP7_75t_L g2549 ( 
.A(n_2324),
.Y(n_2549)
);

OAI22xp33_ASAP7_75t_L g2550 ( 
.A1(n_2302),
.A2(n_2282),
.B1(n_2287),
.B2(n_2450),
.Y(n_2550)
);

OR2x2_ASAP7_75t_L g2551 ( 
.A(n_2263),
.B(n_2415),
.Y(n_2551)
);

INVx1_ASAP7_75t_L g2552 ( 
.A(n_2210),
.Y(n_2552)
);

INVx1_ASAP7_75t_L g2553 ( 
.A(n_2268),
.Y(n_2553)
);

INVx1_ASAP7_75t_L g2554 ( 
.A(n_2274),
.Y(n_2554)
);

INVx2_ASAP7_75t_L g2555 ( 
.A(n_2273),
.Y(n_2555)
);

INVx1_ASAP7_75t_L g2556 ( 
.A(n_2231),
.Y(n_2556)
);

INVx3_ASAP7_75t_L g2557 ( 
.A(n_2259),
.Y(n_2557)
);

OAI22xp5_ASAP7_75t_L g2558 ( 
.A1(n_2302),
.A2(n_2442),
.B1(n_2463),
.B2(n_2290),
.Y(n_2558)
);

INVx1_ASAP7_75t_L g2559 ( 
.A(n_2234),
.Y(n_2559)
);

INVx1_ASAP7_75t_L g2560 ( 
.A(n_2236),
.Y(n_2560)
);

INVx1_ASAP7_75t_SL g2561 ( 
.A(n_2532),
.Y(n_2561)
);

INVx1_ASAP7_75t_L g2562 ( 
.A(n_2264),
.Y(n_2562)
);

INVx1_ASAP7_75t_L g2563 ( 
.A(n_2283),
.Y(n_2563)
);

INVx1_ASAP7_75t_L g2564 ( 
.A(n_2316),
.Y(n_2564)
);

INVx1_ASAP7_75t_L g2565 ( 
.A(n_2316),
.Y(n_2565)
);

INVx2_ASAP7_75t_SL g2566 ( 
.A(n_2281),
.Y(n_2566)
);

INVx1_ASAP7_75t_L g2567 ( 
.A(n_2338),
.Y(n_2567)
);

NAND2x1p5_ASAP7_75t_L g2568 ( 
.A(n_2259),
.B(n_2204),
.Y(n_2568)
);

INVx1_ASAP7_75t_L g2569 ( 
.A(n_2338),
.Y(n_2569)
);

INVx2_ASAP7_75t_L g2570 ( 
.A(n_2273),
.Y(n_2570)
);

INVxp33_ASAP7_75t_L g2571 ( 
.A(n_2251),
.Y(n_2571)
);

INVx2_ASAP7_75t_L g2572 ( 
.A(n_2275),
.Y(n_2572)
);

INVx4_ASAP7_75t_L g2573 ( 
.A(n_2205),
.Y(n_2573)
);

AND2x2_ASAP7_75t_L g2574 ( 
.A(n_2356),
.B(n_2450),
.Y(n_2574)
);

HB1xp67_ASAP7_75t_L g2575 ( 
.A(n_2399),
.Y(n_2575)
);

AND2x4_ASAP7_75t_L g2576 ( 
.A(n_2373),
.B(n_2439),
.Y(n_2576)
);

INVx1_ASAP7_75t_L g2577 ( 
.A(n_2227),
.Y(n_2577)
);

INVx2_ASAP7_75t_L g2578 ( 
.A(n_2276),
.Y(n_2578)
);

OAI22xp33_ASAP7_75t_L g2579 ( 
.A1(n_2483),
.A2(n_2323),
.B1(n_2308),
.B2(n_2350),
.Y(n_2579)
);

BUFx3_ASAP7_75t_L g2580 ( 
.A(n_2212),
.Y(n_2580)
);

INVx2_ASAP7_75t_L g2581 ( 
.A(n_2285),
.Y(n_2581)
);

INVx1_ASAP7_75t_L g2582 ( 
.A(n_2227),
.Y(n_2582)
);

AND2x4_ASAP7_75t_L g2583 ( 
.A(n_2373),
.B(n_2439),
.Y(n_2583)
);

AND2x2_ASAP7_75t_L g2584 ( 
.A(n_2411),
.B(n_2373),
.Y(n_2584)
);

INVx1_ASAP7_75t_L g2585 ( 
.A(n_2244),
.Y(n_2585)
);

INVx2_ASAP7_75t_L g2586 ( 
.A(n_2285),
.Y(n_2586)
);

OAI21xp5_ASAP7_75t_L g2587 ( 
.A1(n_2507),
.A2(n_2457),
.B(n_2455),
.Y(n_2587)
);

INVx1_ASAP7_75t_L g2588 ( 
.A(n_2244),
.Y(n_2588)
);

INVx1_ASAP7_75t_L g2589 ( 
.A(n_2254),
.Y(n_2589)
);

BUFx3_ASAP7_75t_L g2590 ( 
.A(n_2212),
.Y(n_2590)
);

INVx3_ASAP7_75t_L g2591 ( 
.A(n_2233),
.Y(n_2591)
);

BUFx2_ASAP7_75t_R g2592 ( 
.A(n_2205),
.Y(n_2592)
);

INVx11_ASAP7_75t_L g2593 ( 
.A(n_2269),
.Y(n_2593)
);

NAND2x1p5_ASAP7_75t_L g2594 ( 
.A(n_2225),
.B(n_2535),
.Y(n_2594)
);

INVx11_ASAP7_75t_L g2595 ( 
.A(n_2269),
.Y(n_2595)
);

BUFx3_ASAP7_75t_L g2596 ( 
.A(n_2225),
.Y(n_2596)
);

AOI22xp5_ASAP7_75t_L g2597 ( 
.A1(n_2486),
.A2(n_2533),
.B1(n_2475),
.B2(n_2424),
.Y(n_2597)
);

BUFx4f_ASAP7_75t_SL g2598 ( 
.A(n_2237),
.Y(n_2598)
);

INVx3_ASAP7_75t_L g2599 ( 
.A(n_2233),
.Y(n_2599)
);

AOI22xp33_ASAP7_75t_SL g2600 ( 
.A1(n_2358),
.A2(n_2364),
.B1(n_2426),
.B2(n_2442),
.Y(n_2600)
);

OAI22xp33_ASAP7_75t_L g2601 ( 
.A1(n_2483),
.A2(n_2350),
.B1(n_2297),
.B2(n_2311),
.Y(n_2601)
);

OAI22xp33_ASAP7_75t_L g2602 ( 
.A1(n_2350),
.A2(n_2322),
.B1(n_2360),
.B2(n_2223),
.Y(n_2602)
);

BUFx2_ASAP7_75t_L g2603 ( 
.A(n_2355),
.Y(n_2603)
);

INVx4_ASAP7_75t_L g2604 ( 
.A(n_2232),
.Y(n_2604)
);

INVx3_ASAP7_75t_L g2605 ( 
.A(n_2208),
.Y(n_2605)
);

AOI22xp33_ASAP7_75t_L g2606 ( 
.A1(n_2504),
.A2(n_2511),
.B1(n_2475),
.B2(n_2410),
.Y(n_2606)
);

AOI22xp33_ASAP7_75t_L g2607 ( 
.A1(n_2511),
.A2(n_2286),
.B1(n_2463),
.B2(n_2512),
.Y(n_2607)
);

BUFx2_ASAP7_75t_L g2608 ( 
.A(n_2355),
.Y(n_2608)
);

CKINVDCx20_ASAP7_75t_R g2609 ( 
.A(n_2206),
.Y(n_2609)
);

BUFx3_ASAP7_75t_L g2610 ( 
.A(n_2535),
.Y(n_2610)
);

AND2x2_ASAP7_75t_L g2611 ( 
.A(n_2411),
.B(n_2445),
.Y(n_2611)
);

OAI22xp5_ASAP7_75t_L g2612 ( 
.A1(n_2442),
.A2(n_2290),
.B1(n_2319),
.B2(n_2298),
.Y(n_2612)
);

INVx1_ASAP7_75t_L g2613 ( 
.A(n_2218),
.Y(n_2613)
);

INVx2_ASAP7_75t_L g2614 ( 
.A(n_2401),
.Y(n_2614)
);

HB1xp67_ASAP7_75t_L g2615 ( 
.A(n_2399),
.Y(n_2615)
);

INVx2_ASAP7_75t_SL g2616 ( 
.A(n_2281),
.Y(n_2616)
);

INVx2_ASAP7_75t_SL g2617 ( 
.A(n_2281),
.Y(n_2617)
);

NAND2x1p5_ASAP7_75t_L g2618 ( 
.A(n_2260),
.B(n_2456),
.Y(n_2618)
);

INVx2_ASAP7_75t_L g2619 ( 
.A(n_2401),
.Y(n_2619)
);

HB1xp67_ASAP7_75t_L g2620 ( 
.A(n_2402),
.Y(n_2620)
);

OR2x2_ASAP7_75t_L g2621 ( 
.A(n_2398),
.B(n_2536),
.Y(n_2621)
);

INVx1_ASAP7_75t_L g2622 ( 
.A(n_2218),
.Y(n_2622)
);

BUFx2_ASAP7_75t_L g2623 ( 
.A(n_2307),
.Y(n_2623)
);

AOI22xp33_ASAP7_75t_L g2624 ( 
.A1(n_2511),
.A2(n_2512),
.B1(n_2292),
.B2(n_2403),
.Y(n_2624)
);

INVx1_ASAP7_75t_L g2625 ( 
.A(n_2449),
.Y(n_2625)
);

OAI22xp5_ASAP7_75t_L g2626 ( 
.A1(n_2290),
.A2(n_2319),
.B1(n_2298),
.B2(n_2241),
.Y(n_2626)
);

INVx2_ASAP7_75t_L g2627 ( 
.A(n_2401),
.Y(n_2627)
);

INVx1_ASAP7_75t_L g2628 ( 
.A(n_2241),
.Y(n_2628)
);

INVx2_ASAP7_75t_L g2629 ( 
.A(n_2401),
.Y(n_2629)
);

BUFx2_ASAP7_75t_L g2630 ( 
.A(n_2307),
.Y(n_2630)
);

AOI22xp33_ASAP7_75t_L g2631 ( 
.A1(n_2292),
.A2(n_2396),
.B1(n_2424),
.B2(n_2207),
.Y(n_2631)
);

BUFx2_ASAP7_75t_L g2632 ( 
.A(n_2260),
.Y(n_2632)
);

OAI22xp5_ASAP7_75t_L g2633 ( 
.A1(n_2298),
.A2(n_2319),
.B1(n_2241),
.B2(n_2350),
.Y(n_2633)
);

INVx1_ASAP7_75t_L g2634 ( 
.A(n_2330),
.Y(n_2634)
);

AND2x2_ASAP7_75t_L g2635 ( 
.A(n_2397),
.B(n_2390),
.Y(n_2635)
);

INVx2_ASAP7_75t_SL g2636 ( 
.A(n_2532),
.Y(n_2636)
);

INVx2_ASAP7_75t_L g2637 ( 
.A(n_2401),
.Y(n_2637)
);

INVx1_ASAP7_75t_L g2638 ( 
.A(n_2267),
.Y(n_2638)
);

NAND2x1p5_ASAP7_75t_L g2639 ( 
.A(n_2456),
.B(n_2198),
.Y(n_2639)
);

OAI22xp5_ASAP7_75t_L g2640 ( 
.A1(n_2515),
.A2(n_2433),
.B1(n_2440),
.B2(n_2418),
.Y(n_2640)
);

HB1xp67_ASAP7_75t_L g2641 ( 
.A(n_2402),
.Y(n_2641)
);

INVx2_ASAP7_75t_L g2642 ( 
.A(n_2401),
.Y(n_2642)
);

INVx11_ASAP7_75t_L g2643 ( 
.A(n_2324),
.Y(n_2643)
);

INVx1_ASAP7_75t_L g2644 ( 
.A(n_2261),
.Y(n_2644)
);

INVx1_ASAP7_75t_L g2645 ( 
.A(n_2262),
.Y(n_2645)
);

AOI21x1_ASAP7_75t_L g2646 ( 
.A1(n_2395),
.A2(n_2221),
.B(n_2470),
.Y(n_2646)
);

INVx2_ASAP7_75t_L g2647 ( 
.A(n_2401),
.Y(n_2647)
);

INVx3_ASAP7_75t_L g2648 ( 
.A(n_2208),
.Y(n_2648)
);

INVx1_ASAP7_75t_L g2649 ( 
.A(n_2223),
.Y(n_2649)
);

BUFx2_ASAP7_75t_L g2650 ( 
.A(n_2277),
.Y(n_2650)
);

OAI221xp5_ASAP7_75t_L g2651 ( 
.A1(n_2370),
.A2(n_2299),
.B1(n_2388),
.B2(n_2513),
.C(n_2486),
.Y(n_2651)
);

INVx1_ASAP7_75t_L g2652 ( 
.A(n_2337),
.Y(n_2652)
);

AOI22xp33_ASAP7_75t_SL g2653 ( 
.A1(n_2443),
.A2(n_2454),
.B1(n_2488),
.B2(n_2474),
.Y(n_2653)
);

AOI22xp33_ASAP7_75t_L g2654 ( 
.A1(n_2453),
.A2(n_2408),
.B1(n_2404),
.B2(n_2471),
.Y(n_2654)
);

HB1xp67_ASAP7_75t_L g2655 ( 
.A(n_2500),
.Y(n_2655)
);

INVx1_ASAP7_75t_L g2656 ( 
.A(n_2337),
.Y(n_2656)
);

INVx2_ASAP7_75t_SL g2657 ( 
.A(n_2237),
.Y(n_2657)
);

INVx1_ASAP7_75t_L g2658 ( 
.A(n_2317),
.Y(n_2658)
);

HB1xp67_ASAP7_75t_L g2659 ( 
.A(n_2500),
.Y(n_2659)
);

INVx1_ASAP7_75t_L g2660 ( 
.A(n_2448),
.Y(n_2660)
);

INVx3_ASAP7_75t_L g2661 ( 
.A(n_2208),
.Y(n_2661)
);

BUFx3_ASAP7_75t_L g2662 ( 
.A(n_2324),
.Y(n_2662)
);

NAND2xp5_ASAP7_75t_L g2663 ( 
.A(n_2368),
.B(n_2382),
.Y(n_2663)
);

NOR2xp33_ASAP7_75t_L g2664 ( 
.A(n_2400),
.B(n_2245),
.Y(n_2664)
);

OAI22xp33_ASAP7_75t_L g2665 ( 
.A1(n_2427),
.A2(n_2253),
.B1(n_2255),
.B2(n_2258),
.Y(n_2665)
);

HB1xp67_ASAP7_75t_L g2666 ( 
.A(n_2500),
.Y(n_2666)
);

CKINVDCx20_ASAP7_75t_R g2667 ( 
.A(n_2206),
.Y(n_2667)
);

CKINVDCx20_ASAP7_75t_R g2668 ( 
.A(n_2265),
.Y(n_2668)
);

INVx1_ASAP7_75t_L g2669 ( 
.A(n_2366),
.Y(n_2669)
);

INVx1_ASAP7_75t_L g2670 ( 
.A(n_2339),
.Y(n_2670)
);

OAI22xp5_ASAP7_75t_L g2671 ( 
.A1(n_2451),
.A2(n_2460),
.B1(n_2480),
.B2(n_2464),
.Y(n_2671)
);

INVx1_ASAP7_75t_L g2672 ( 
.A(n_2409),
.Y(n_2672)
);

AOI22xp33_ASAP7_75t_SL g2673 ( 
.A1(n_2443),
.A2(n_2488),
.B1(n_2474),
.B2(n_2203),
.Y(n_2673)
);

INVx1_ASAP7_75t_L g2674 ( 
.A(n_2409),
.Y(n_2674)
);

INVx1_ASAP7_75t_L g2675 ( 
.A(n_2385),
.Y(n_2675)
);

INVx1_ASAP7_75t_L g2676 ( 
.A(n_2407),
.Y(n_2676)
);

AND2x2_ASAP7_75t_L g2677 ( 
.A(n_2432),
.B(n_2405),
.Y(n_2677)
);

INVx3_ASAP7_75t_L g2678 ( 
.A(n_2230),
.Y(n_2678)
);

BUFx3_ASAP7_75t_L g2679 ( 
.A(n_2242),
.Y(n_2679)
);

INVx1_ASAP7_75t_L g2680 ( 
.A(n_2407),
.Y(n_2680)
);

INVx1_ASAP7_75t_L g2681 ( 
.A(n_2278),
.Y(n_2681)
);

INVx1_ASAP7_75t_L g2682 ( 
.A(n_2278),
.Y(n_2682)
);

AND2x2_ASAP7_75t_L g2683 ( 
.A(n_2432),
.B(n_2381),
.Y(n_2683)
);

INVx1_ASAP7_75t_L g2684 ( 
.A(n_2278),
.Y(n_2684)
);

INVx1_ASAP7_75t_L g2685 ( 
.A(n_2278),
.Y(n_2685)
);

AND2x2_ASAP7_75t_L g2686 ( 
.A(n_2381),
.B(n_2436),
.Y(n_2686)
);

AND2x2_ASAP7_75t_L g2687 ( 
.A(n_2381),
.B(n_2436),
.Y(n_2687)
);

INVx1_ASAP7_75t_L g2688 ( 
.A(n_2257),
.Y(n_2688)
);

INVx2_ASAP7_75t_SL g2689 ( 
.A(n_2232),
.Y(n_2689)
);

BUFx2_ASAP7_75t_L g2690 ( 
.A(n_2280),
.Y(n_2690)
);

INVx1_ASAP7_75t_L g2691 ( 
.A(n_2284),
.Y(n_2691)
);

AND2x2_ASAP7_75t_L g2692 ( 
.A(n_2374),
.B(n_2291),
.Y(n_2692)
);

INVx1_ASAP7_75t_L g2693 ( 
.A(n_2272),
.Y(n_2693)
);

INVx3_ASAP7_75t_L g2694 ( 
.A(n_2230),
.Y(n_2694)
);

INVx1_ASAP7_75t_L g2695 ( 
.A(n_2272),
.Y(n_2695)
);

INVx3_ASAP7_75t_L g2696 ( 
.A(n_2230),
.Y(n_2696)
);

CKINVDCx5p33_ASAP7_75t_R g2697 ( 
.A(n_2265),
.Y(n_2697)
);

OAI21xp5_ASAP7_75t_L g2698 ( 
.A1(n_2455),
.A2(n_2457),
.B(n_2509),
.Y(n_2698)
);

AND2x4_ASAP7_75t_L g2699 ( 
.A(n_2386),
.B(n_2427),
.Y(n_2699)
);

INVx1_ASAP7_75t_L g2700 ( 
.A(n_2344),
.Y(n_2700)
);

HB1xp67_ASAP7_75t_L g2701 ( 
.A(n_2378),
.Y(n_2701)
);

INVx1_ASAP7_75t_L g2702 ( 
.A(n_2351),
.Y(n_2702)
);

INVx1_ASAP7_75t_L g2703 ( 
.A(n_2226),
.Y(n_2703)
);

INVx1_ASAP7_75t_L g2704 ( 
.A(n_2301),
.Y(n_2704)
);

INVx1_ASAP7_75t_L g2705 ( 
.A(n_2301),
.Y(n_2705)
);

INVx1_ASAP7_75t_SL g2706 ( 
.A(n_2372),
.Y(n_2706)
);

INVx1_ASAP7_75t_L g2707 ( 
.A(n_2312),
.Y(n_2707)
);

INVx1_ASAP7_75t_SL g2708 ( 
.A(n_2372),
.Y(n_2708)
);

OR2x2_ASAP7_75t_L g2709 ( 
.A(n_2353),
.B(n_2422),
.Y(n_2709)
);

INVx1_ASAP7_75t_L g2710 ( 
.A(n_2312),
.Y(n_2710)
);

INVx1_ASAP7_75t_L g2711 ( 
.A(n_2315),
.Y(n_2711)
);

INVx1_ASAP7_75t_L g2712 ( 
.A(n_2325),
.Y(n_2712)
);

INVx1_ASAP7_75t_L g2713 ( 
.A(n_2325),
.Y(n_2713)
);

BUFx2_ASAP7_75t_L g2714 ( 
.A(n_2427),
.Y(n_2714)
);

OR2x2_ASAP7_75t_L g2715 ( 
.A(n_2392),
.B(n_2492),
.Y(n_2715)
);

INVx3_ASAP7_75t_L g2716 ( 
.A(n_2295),
.Y(n_2716)
);

NAND2xp5_ASAP7_75t_L g2717 ( 
.A(n_2391),
.B(n_2394),
.Y(n_2717)
);

INVx1_ASAP7_75t_L g2718 ( 
.A(n_2329),
.Y(n_2718)
);

INVx1_ASAP7_75t_L g2719 ( 
.A(n_2333),
.Y(n_2719)
);

AOI22xp33_ASAP7_75t_L g2720 ( 
.A1(n_2453),
.A2(n_2471),
.B1(n_2485),
.B2(n_2477),
.Y(n_2720)
);

INVx3_ASAP7_75t_L g2721 ( 
.A(n_2295),
.Y(n_2721)
);

HB1xp67_ASAP7_75t_L g2722 ( 
.A(n_2378),
.Y(n_2722)
);

OR2x2_ASAP7_75t_L g2723 ( 
.A(n_2427),
.B(n_2519),
.Y(n_2723)
);

BUFx2_ASAP7_75t_L g2724 ( 
.A(n_2443),
.Y(n_2724)
);

NAND2xp5_ASAP7_75t_L g2725 ( 
.A(n_2444),
.B(n_2465),
.Y(n_2725)
);

BUFx8_ASAP7_75t_SL g2726 ( 
.A(n_2279),
.Y(n_2726)
);

INVx1_ASAP7_75t_L g2727 ( 
.A(n_2341),
.Y(n_2727)
);

INVx1_ASAP7_75t_L g2728 ( 
.A(n_2213),
.Y(n_2728)
);

INVx2_ASAP7_75t_L g2729 ( 
.A(n_2332),
.Y(n_2729)
);

AOI21x1_ASAP7_75t_L g2730 ( 
.A1(n_2528),
.A2(n_2431),
.B(n_2296),
.Y(n_2730)
);

AOI22xp33_ASAP7_75t_L g2731 ( 
.A1(n_2453),
.A2(n_2485),
.B1(n_2498),
.B2(n_2477),
.Y(n_2731)
);

CKINVDCx11_ASAP7_75t_R g2732 ( 
.A(n_2293),
.Y(n_2732)
);

OAI21xp5_ASAP7_75t_L g2733 ( 
.A1(n_2509),
.A2(n_2506),
.B(n_2514),
.Y(n_2733)
);

NAND2xp5_ASAP7_75t_L g2734 ( 
.A(n_2472),
.B(n_2482),
.Y(n_2734)
);

AOI22xp33_ASAP7_75t_L g2735 ( 
.A1(n_2498),
.A2(n_2508),
.B1(n_2214),
.B2(n_2313),
.Y(n_2735)
);

HB1xp67_ASAP7_75t_L g2736 ( 
.A(n_2378),
.Y(n_2736)
);

INVx1_ASAP7_75t_L g2737 ( 
.A(n_2216),
.Y(n_2737)
);

BUFx2_ASAP7_75t_L g2738 ( 
.A(n_2417),
.Y(n_2738)
);

BUFx2_ASAP7_75t_L g2739 ( 
.A(n_2417),
.Y(n_2739)
);

INVxp33_ASAP7_75t_L g2740 ( 
.A(n_2378),
.Y(n_2740)
);

AOI322xp5_ASAP7_75t_L g2741 ( 
.A1(n_2246),
.A2(n_2321),
.A3(n_2331),
.B1(n_2528),
.B2(n_2224),
.C1(n_2222),
.C2(n_2279),
.Y(n_2741)
);

INVx2_ASAP7_75t_SL g2742 ( 
.A(n_2295),
.Y(n_2742)
);

NAND2xp5_ASAP7_75t_L g2743 ( 
.A(n_2501),
.B(n_2502),
.Y(n_2743)
);

INVx1_ASAP7_75t_L g2744 ( 
.A(n_2288),
.Y(n_2744)
);

INVx1_ASAP7_75t_L g2745 ( 
.A(n_2314),
.Y(n_2745)
);

INVx1_ASAP7_75t_L g2746 ( 
.A(n_2328),
.Y(n_2746)
);

INVx2_ASAP7_75t_L g2747 ( 
.A(n_2199),
.Y(n_2747)
);

NOR2xp33_ASAP7_75t_L g2748 ( 
.A(n_2497),
.B(n_2493),
.Y(n_2748)
);

BUFx3_ASAP7_75t_L g2749 ( 
.A(n_2423),
.Y(n_2749)
);

INVx1_ASAP7_75t_L g2750 ( 
.A(n_2336),
.Y(n_2750)
);

INVx1_ASAP7_75t_L g2751 ( 
.A(n_2384),
.Y(n_2751)
);

INVx2_ASAP7_75t_L g2752 ( 
.A(n_2199),
.Y(n_2752)
);

INVx2_ASAP7_75t_L g2753 ( 
.A(n_2199),
.Y(n_2753)
);

INVx1_ASAP7_75t_L g2754 ( 
.A(n_2318),
.Y(n_2754)
);

HB1xp67_ASAP7_75t_L g2755 ( 
.A(n_2365),
.Y(n_2755)
);

AOI22xp5_ASAP7_75t_L g2756 ( 
.A1(n_2473),
.A2(n_2481),
.B1(n_2503),
.B2(n_2510),
.Y(n_2756)
);

BUFx3_ASAP7_75t_L g2757 ( 
.A(n_2238),
.Y(n_2757)
);

INVx2_ASAP7_75t_SL g2758 ( 
.A(n_2320),
.Y(n_2758)
);

OAI22xp33_ASAP7_75t_L g2759 ( 
.A1(n_2247),
.A2(n_2437),
.B1(n_2474),
.B2(n_2266),
.Y(n_2759)
);

INVx1_ASAP7_75t_L g2760 ( 
.A(n_2318),
.Y(n_2760)
);

INVx1_ASAP7_75t_L g2761 ( 
.A(n_2318),
.Y(n_2761)
);

CKINVDCx20_ASAP7_75t_R g2762 ( 
.A(n_2320),
.Y(n_2762)
);

OR2x2_ASAP7_75t_L g2763 ( 
.A(n_2473),
.B(n_2517),
.Y(n_2763)
);

HB1xp67_ASAP7_75t_L g2764 ( 
.A(n_2365),
.Y(n_2764)
);

BUFx2_ASAP7_75t_L g2765 ( 
.A(n_2238),
.Y(n_2765)
);

BUFx3_ASAP7_75t_L g2766 ( 
.A(n_2238),
.Y(n_2766)
);

CKINVDCx5p33_ASAP7_75t_R g2767 ( 
.A(n_2201),
.Y(n_2767)
);

BUFx3_ASAP7_75t_L g2768 ( 
.A(n_2239),
.Y(n_2768)
);

AND2x4_ASAP7_75t_L g2769 ( 
.A(n_2239),
.B(n_2414),
.Y(n_2769)
);

INVx1_ASAP7_75t_L g2770 ( 
.A(n_2318),
.Y(n_2770)
);

INVx1_ASAP7_75t_L g2771 ( 
.A(n_2304),
.Y(n_2771)
);

OR2x2_ASAP7_75t_L g2772 ( 
.A(n_2510),
.B(n_2437),
.Y(n_2772)
);

AOI21xp33_ASAP7_75t_L g2773 ( 
.A1(n_2488),
.A2(n_2467),
.B(n_2438),
.Y(n_2773)
);

AO21x2_ASAP7_75t_L g2774 ( 
.A1(n_2530),
.A2(n_2215),
.B(n_2235),
.Y(n_2774)
);

AOI22xp33_ASAP7_75t_SL g2775 ( 
.A1(n_2270),
.A2(n_2303),
.B1(n_2256),
.B2(n_2202),
.Y(n_2775)
);

BUFx2_ASAP7_75t_L g2776 ( 
.A(n_2239),
.Y(n_2776)
);

OAI22xp5_ASAP7_75t_L g2777 ( 
.A1(n_2246),
.A2(n_2299),
.B1(n_2270),
.B2(n_2303),
.Y(n_2777)
);

INVx1_ASAP7_75t_L g2778 ( 
.A(n_2354),
.Y(n_2778)
);

INVx3_ASAP7_75t_L g2779 ( 
.A(n_2310),
.Y(n_2779)
);

NAND2xp5_ASAP7_75t_L g2780 ( 
.A(n_2671),
.B(n_2625),
.Y(n_2780)
);

AND2x2_ASAP7_75t_L g2781 ( 
.A(n_2635),
.B(n_2414),
.Y(n_2781)
);

INVx1_ASAP7_75t_L g2782 ( 
.A(n_2552),
.Y(n_2782)
);

INVx2_ASAP7_75t_SL g2783 ( 
.A(n_2643),
.Y(n_2783)
);

AOI22xp33_ASAP7_75t_L g2784 ( 
.A1(n_2550),
.A2(n_2458),
.B1(n_2459),
.B2(n_2461),
.Y(n_2784)
);

AND2x2_ASAP7_75t_L g2785 ( 
.A(n_2584),
.B(n_2421),
.Y(n_2785)
);

AND2x2_ASAP7_75t_L g2786 ( 
.A(n_2611),
.B(n_2421),
.Y(n_2786)
);

NAND2xp5_ASAP7_75t_L g2787 ( 
.A(n_2671),
.B(n_2462),
.Y(n_2787)
);

OAI22xp5_ASAP7_75t_L g2788 ( 
.A1(n_2539),
.A2(n_2303),
.B1(n_2270),
.B2(n_2361),
.Y(n_2788)
);

BUFx2_ASAP7_75t_L g2789 ( 
.A(n_2749),
.Y(n_2789)
);

OAI22xp5_ASAP7_75t_L g2790 ( 
.A1(n_2539),
.A2(n_2362),
.B1(n_2359),
.B2(n_2441),
.Y(n_2790)
);

AND2x2_ASAP7_75t_L g2791 ( 
.A(n_2574),
.B(n_2429),
.Y(n_2791)
);

AOI22xp33_ASAP7_75t_L g2792 ( 
.A1(n_2550),
.A2(n_2458),
.B1(n_2459),
.B2(n_2461),
.Y(n_2792)
);

INVx1_ASAP7_75t_L g2793 ( 
.A(n_2553),
.Y(n_2793)
);

INVx3_ASAP7_75t_L g2794 ( 
.A(n_2557),
.Y(n_2794)
);

AOI22xp33_ASAP7_75t_SL g2795 ( 
.A1(n_2558),
.A2(n_2202),
.B1(n_2256),
.B2(n_2220),
.Y(n_2795)
);

INVx2_ASAP7_75t_SL g2796 ( 
.A(n_2598),
.Y(n_2796)
);

INVx1_ASAP7_75t_L g2797 ( 
.A(n_2554),
.Y(n_2797)
);

OAI22xp5_ASAP7_75t_L g2798 ( 
.A1(n_2558),
.A2(n_2306),
.B1(n_2365),
.B2(n_2456),
.Y(n_2798)
);

BUFx2_ASAP7_75t_L g2799 ( 
.A(n_2749),
.Y(n_2799)
);

NAND2xp5_ASAP7_75t_L g2800 ( 
.A(n_2640),
.B(n_2462),
.Y(n_2800)
);

AND2x4_ASAP7_75t_L g2801 ( 
.A(n_2538),
.B(n_2367),
.Y(n_2801)
);

AND2x4_ASAP7_75t_L g2802 ( 
.A(n_2576),
.B(n_2367),
.Y(n_2802)
);

INVx1_ASAP7_75t_L g2803 ( 
.A(n_2556),
.Y(n_2803)
);

OR2x2_ASAP7_75t_L g2804 ( 
.A(n_2551),
.B(n_2709),
.Y(n_2804)
);

INVx2_ASAP7_75t_SL g2805 ( 
.A(n_2598),
.Y(n_2805)
);

INVx2_ASAP7_75t_SL g2806 ( 
.A(n_2593),
.Y(n_2806)
);

AND2x2_ASAP7_75t_L g2807 ( 
.A(n_2576),
.B(n_2429),
.Y(n_2807)
);

NAND2xp5_ASAP7_75t_L g2808 ( 
.A(n_2640),
.B(n_2526),
.Y(n_2808)
);

INVx2_ASAP7_75t_SL g2809 ( 
.A(n_2595),
.Y(n_2809)
);

INVx1_ASAP7_75t_L g2810 ( 
.A(n_2559),
.Y(n_2810)
);

INVx1_ASAP7_75t_L g2811 ( 
.A(n_2560),
.Y(n_2811)
);

HB1xp67_ASAP7_75t_L g2812 ( 
.A(n_2575),
.Y(n_2812)
);

AND2x2_ASAP7_75t_L g2813 ( 
.A(n_2583),
.B(n_2369),
.Y(n_2813)
);

AND2x2_ASAP7_75t_L g2814 ( 
.A(n_2583),
.B(n_2369),
.Y(n_2814)
);

INVx1_ASAP7_75t_L g2815 ( 
.A(n_2562),
.Y(n_2815)
);

HB1xp67_ASAP7_75t_L g2816 ( 
.A(n_2575),
.Y(n_2816)
);

INVx1_ASAP7_75t_L g2817 ( 
.A(n_2563),
.Y(n_2817)
);

INVx1_ASAP7_75t_L g2818 ( 
.A(n_2541),
.Y(n_2818)
);

INVx1_ASAP7_75t_L g2819 ( 
.A(n_2545),
.Y(n_2819)
);

AND2x2_ASAP7_75t_L g2820 ( 
.A(n_2621),
.B(n_2476),
.Y(n_2820)
);

INVx1_ASAP7_75t_L g2821 ( 
.A(n_2700),
.Y(n_2821)
);

INVx1_ASAP7_75t_L g2822 ( 
.A(n_2702),
.Y(n_2822)
);

NAND2xp5_ASAP7_75t_L g2823 ( 
.A(n_2669),
.B(n_2676),
.Y(n_2823)
);

INVx1_ASAP7_75t_L g2824 ( 
.A(n_2728),
.Y(n_2824)
);

AND2x2_ASAP7_75t_L g2825 ( 
.A(n_2623),
.B(n_2476),
.Y(n_2825)
);

INVx1_ASAP7_75t_SL g2826 ( 
.A(n_2765),
.Y(n_2826)
);

INVx1_ASAP7_75t_L g2827 ( 
.A(n_2737),
.Y(n_2827)
);

AND2x4_ASAP7_75t_L g2828 ( 
.A(n_2557),
.B(n_2434),
.Y(n_2828)
);

HB1xp67_ASAP7_75t_L g2829 ( 
.A(n_2615),
.Y(n_2829)
);

INVx1_ASAP7_75t_L g2830 ( 
.A(n_2745),
.Y(n_2830)
);

NAND2xp5_ASAP7_75t_L g2831 ( 
.A(n_2680),
.B(n_2527),
.Y(n_2831)
);

AND2x2_ASAP7_75t_L g2832 ( 
.A(n_2630),
.B(n_2476),
.Y(n_2832)
);

INVx1_ASAP7_75t_L g2833 ( 
.A(n_2746),
.Y(n_2833)
);

INVx3_ASAP7_75t_L g2834 ( 
.A(n_2543),
.Y(n_2834)
);

INVx1_ASAP7_75t_L g2835 ( 
.A(n_2750),
.Y(n_2835)
);

AND2x4_ASAP7_75t_L g2836 ( 
.A(n_2757),
.B(n_2434),
.Y(n_2836)
);

INVx1_ASAP7_75t_L g2837 ( 
.A(n_2778),
.Y(n_2837)
);

HB1xp67_ASAP7_75t_L g2838 ( 
.A(n_2615),
.Y(n_2838)
);

OAI21xp5_ASAP7_75t_SL g2839 ( 
.A1(n_2600),
.A2(n_2250),
.B(n_2446),
.Y(n_2839)
);

INVx1_ASAP7_75t_L g2840 ( 
.A(n_2564),
.Y(n_2840)
);

OR2x2_ASAP7_75t_L g2841 ( 
.A(n_2679),
.B(n_2527),
.Y(n_2841)
);

INVx1_ASAP7_75t_L g2842 ( 
.A(n_2565),
.Y(n_2842)
);

AND2x2_ASAP7_75t_L g2843 ( 
.A(n_2677),
.B(n_2476),
.Y(n_2843)
);

AND2x2_ASAP7_75t_L g2844 ( 
.A(n_2658),
.B(n_2348),
.Y(n_2844)
);

AO31x2_ASAP7_75t_L g2845 ( 
.A1(n_2777),
.A2(n_2347),
.A3(n_2342),
.B(n_2505),
.Y(n_2845)
);

AND2x4_ASAP7_75t_SL g2846 ( 
.A(n_2668),
.B(n_2334),
.Y(n_2846)
);

INVx1_ASAP7_75t_L g2847 ( 
.A(n_2567),
.Y(n_2847)
);

INVx1_ASAP7_75t_L g2848 ( 
.A(n_2569),
.Y(n_2848)
);

INVx1_ASAP7_75t_L g2849 ( 
.A(n_2644),
.Y(n_2849)
);

NOR2xp33_ASAP7_75t_R g2850 ( 
.A(n_2668),
.B(n_2202),
.Y(n_2850)
);

INVx1_ASAP7_75t_L g2851 ( 
.A(n_2645),
.Y(n_2851)
);

AND2x2_ASAP7_75t_L g2852 ( 
.A(n_2679),
.B(n_2419),
.Y(n_2852)
);

BUFx5_ASAP7_75t_L g2853 ( 
.A(n_2757),
.Y(n_2853)
);

OR2x2_ASAP7_75t_L g2854 ( 
.A(n_2675),
.B(n_2527),
.Y(n_2854)
);

INVxp67_ASAP7_75t_L g2855 ( 
.A(n_2620),
.Y(n_2855)
);

OAI21xp33_ASAP7_75t_L g2856 ( 
.A1(n_2606),
.A2(n_2525),
.B(n_2521),
.Y(n_2856)
);

AND2x4_ASAP7_75t_L g2857 ( 
.A(n_2766),
.B(n_2434),
.Y(n_2857)
);

OR2x2_ASAP7_75t_L g2858 ( 
.A(n_2763),
.B(n_2530),
.Y(n_2858)
);

INVx2_ASAP7_75t_SL g2859 ( 
.A(n_2549),
.Y(n_2859)
);

NOR2x1_ASAP7_75t_SL g2860 ( 
.A(n_2626),
.B(n_2300),
.Y(n_2860)
);

AND2x4_ASAP7_75t_SL g2861 ( 
.A(n_2609),
.B(n_2334),
.Y(n_2861)
);

INVx1_ASAP7_75t_L g2862 ( 
.A(n_2663),
.Y(n_2862)
);

AOI22xp33_ASAP7_75t_SL g2863 ( 
.A1(n_2626),
.A2(n_2202),
.B1(n_2220),
.B2(n_2248),
.Y(n_2863)
);

NAND2xp5_ASAP7_75t_L g2864 ( 
.A(n_2663),
.B(n_2490),
.Y(n_2864)
);

INVx1_ASAP7_75t_L g2865 ( 
.A(n_2717),
.Y(n_2865)
);

NOR2xp33_ASAP7_75t_L g2866 ( 
.A(n_2597),
.B(n_2425),
.Y(n_2866)
);

BUFx2_ASAP7_75t_L g2867 ( 
.A(n_2662),
.Y(n_2867)
);

INVx1_ASAP7_75t_SL g2868 ( 
.A(n_2776),
.Y(n_2868)
);

OAI22xp5_ASAP7_75t_L g2869 ( 
.A1(n_2602),
.A2(n_2651),
.B1(n_2612),
.B2(n_2633),
.Y(n_2869)
);

AND2x2_ASAP7_75t_L g2870 ( 
.A(n_2692),
.B(n_2412),
.Y(n_2870)
);

NAND2xp5_ASAP7_75t_L g2871 ( 
.A(n_2717),
.B(n_2490),
.Y(n_2871)
);

INVx1_ASAP7_75t_L g2872 ( 
.A(n_2725),
.Y(n_2872)
);

AND2x2_ASAP7_75t_L g2873 ( 
.A(n_2580),
.B(n_2516),
.Y(n_2873)
);

AND2x2_ASAP7_75t_L g2874 ( 
.A(n_2580),
.B(n_2516),
.Y(n_2874)
);

INVx1_ASAP7_75t_L g2875 ( 
.A(n_2725),
.Y(n_2875)
);

AND2x2_ASAP7_75t_L g2876 ( 
.A(n_2590),
.B(n_2596),
.Y(n_2876)
);

INVx3_ASAP7_75t_L g2877 ( 
.A(n_2543),
.Y(n_2877)
);

NAND2xp5_ASAP7_75t_L g2878 ( 
.A(n_2734),
.B(n_2349),
.Y(n_2878)
);

OR2x2_ASAP7_75t_L g2879 ( 
.A(n_2638),
.B(n_2521),
.Y(n_2879)
);

INVx1_ASAP7_75t_L g2880 ( 
.A(n_2734),
.Y(n_2880)
);

BUFx3_ASAP7_75t_L g2881 ( 
.A(n_2662),
.Y(n_2881)
);

HB1xp67_ASAP7_75t_L g2882 ( 
.A(n_2655),
.Y(n_2882)
);

BUFx2_ASAP7_75t_L g2883 ( 
.A(n_2590),
.Y(n_2883)
);

OR2x2_ASAP7_75t_L g2884 ( 
.A(n_2706),
.B(n_2521),
.Y(n_2884)
);

AND2x4_ASAP7_75t_L g2885 ( 
.A(n_2766),
.B(n_2768),
.Y(n_2885)
);

INVx3_ASAP7_75t_L g2886 ( 
.A(n_2568),
.Y(n_2886)
);

AND2x2_ASAP7_75t_L g2887 ( 
.A(n_2596),
.B(n_2484),
.Y(n_2887)
);

NAND2xp5_ASAP7_75t_L g2888 ( 
.A(n_2606),
.B(n_2349),
.Y(n_2888)
);

INVx1_ASAP7_75t_SL g2889 ( 
.A(n_2768),
.Y(n_2889)
);

OAI221xp5_ASAP7_75t_L g2890 ( 
.A1(n_2631),
.A2(n_2430),
.B1(n_2495),
.B2(n_2435),
.C(n_2447),
.Y(n_2890)
);

INVx1_ASAP7_75t_SL g2891 ( 
.A(n_2769),
.Y(n_2891)
);

AND2x2_ASAP7_75t_L g2892 ( 
.A(n_2610),
.B(n_2484),
.Y(n_2892)
);

HB1xp67_ASAP7_75t_L g2893 ( 
.A(n_2655),
.Y(n_2893)
);

NAND2xp5_ASAP7_75t_L g2894 ( 
.A(n_2607),
.B(n_2743),
.Y(n_2894)
);

AOI22xp33_ASAP7_75t_L g2895 ( 
.A1(n_2665),
.A2(n_2438),
.B1(n_2294),
.B2(n_2252),
.Y(n_2895)
);

AND2x2_ASAP7_75t_L g2896 ( 
.A(n_2610),
.B(n_2209),
.Y(n_2896)
);

INVx2_ASAP7_75t_L g2897 ( 
.A(n_2546),
.Y(n_2897)
);

OR2x2_ASAP7_75t_L g2898 ( 
.A(n_2708),
.B(n_2525),
.Y(n_2898)
);

INVx2_ASAP7_75t_SL g2899 ( 
.A(n_2549),
.Y(n_2899)
);

INVx1_ASAP7_75t_L g2900 ( 
.A(n_2743),
.Y(n_2900)
);

NAND2xp5_ASAP7_75t_L g2901 ( 
.A(n_2607),
.B(n_2525),
.Y(n_2901)
);

INVx1_ASAP7_75t_L g2902 ( 
.A(n_2751),
.Y(n_2902)
);

INVx3_ASAP7_75t_L g2903 ( 
.A(n_2568),
.Y(n_2903)
);

AND2x4_ASAP7_75t_L g2904 ( 
.A(n_2769),
.B(n_2699),
.Y(n_2904)
);

INVx1_ASAP7_75t_L g2905 ( 
.A(n_2555),
.Y(n_2905)
);

CKINVDCx5p33_ASAP7_75t_R g2906 ( 
.A(n_2726),
.Y(n_2906)
);

BUFx3_ASAP7_75t_L g2907 ( 
.A(n_2549),
.Y(n_2907)
);

INVx1_ASAP7_75t_L g2908 ( 
.A(n_2570),
.Y(n_2908)
);

HB1xp67_ASAP7_75t_L g2909 ( 
.A(n_2659),
.Y(n_2909)
);

INVx1_ASAP7_75t_L g2910 ( 
.A(n_2572),
.Y(n_2910)
);

AND2x2_ASAP7_75t_L g2911 ( 
.A(n_2686),
.B(n_2209),
.Y(n_2911)
);

OAI22xp33_ASAP7_75t_L g2912 ( 
.A1(n_2651),
.A2(n_2456),
.B1(n_2468),
.B2(n_2197),
.Y(n_2912)
);

AND2x2_ASAP7_75t_L g2913 ( 
.A(n_2687),
.B(n_2335),
.Y(n_2913)
);

AND2x2_ASAP7_75t_L g2914 ( 
.A(n_2664),
.B(n_2632),
.Y(n_2914)
);

HB1xp67_ASAP7_75t_L g2915 ( 
.A(n_2659),
.Y(n_2915)
);

AND2x2_ASAP7_75t_L g2916 ( 
.A(n_2664),
.B(n_2335),
.Y(n_2916)
);

AND2x2_ASAP7_75t_L g2917 ( 
.A(n_2571),
.B(n_2340),
.Y(n_2917)
);

BUFx2_ASAP7_75t_L g2918 ( 
.A(n_2699),
.Y(n_2918)
);

INVxp67_ASAP7_75t_SL g2919 ( 
.A(n_2729),
.Y(n_2919)
);

NAND2xp5_ASAP7_75t_L g2920 ( 
.A(n_2654),
.B(n_2375),
.Y(n_2920)
);

BUFx6f_ASAP7_75t_L g2921 ( 
.A(n_2594),
.Y(n_2921)
);

AND2x2_ASAP7_75t_L g2922 ( 
.A(n_2571),
.B(n_2340),
.Y(n_2922)
);

AND2x2_ASAP7_75t_L g2923 ( 
.A(n_2724),
.B(n_2594),
.Y(n_2923)
);

INVx1_ASAP7_75t_L g2924 ( 
.A(n_2578),
.Y(n_2924)
);

AND2x2_ASAP7_75t_L g2925 ( 
.A(n_2650),
.B(n_2520),
.Y(n_2925)
);

AOI22xp33_ASAP7_75t_L g2926 ( 
.A1(n_2665),
.A2(n_2289),
.B1(n_2252),
.B2(n_2294),
.Y(n_2926)
);

AOI21xp33_ASAP7_75t_L g2927 ( 
.A1(n_2602),
.A2(n_2467),
.B(n_2491),
.Y(n_2927)
);

AND2x2_ASAP7_75t_L g2928 ( 
.A(n_2690),
.B(n_2520),
.Y(n_2928)
);

AND2x2_ASAP7_75t_L g2929 ( 
.A(n_2683),
.B(n_2217),
.Y(n_2929)
);

INVx2_ASAP7_75t_SL g2930 ( 
.A(n_2657),
.Y(n_2930)
);

AND2x2_ASAP7_75t_L g2931 ( 
.A(n_2748),
.B(n_2249),
.Y(n_2931)
);

INVx1_ASAP7_75t_L g2932 ( 
.A(n_2581),
.Y(n_2932)
);

AND2x2_ASAP7_75t_L g2933 ( 
.A(n_2748),
.B(n_2249),
.Y(n_2933)
);

AND2x2_ASAP7_75t_L g2934 ( 
.A(n_2723),
.B(n_2211),
.Y(n_2934)
);

INVx1_ASAP7_75t_L g2935 ( 
.A(n_2586),
.Y(n_2935)
);

HB1xp67_ASAP7_75t_L g2936 ( 
.A(n_2666),
.Y(n_2936)
);

INVx4_ASAP7_75t_L g2937 ( 
.A(n_2618),
.Y(n_2937)
);

INVx1_ASAP7_75t_L g2938 ( 
.A(n_2649),
.Y(n_2938)
);

INVx3_ASAP7_75t_L g2939 ( 
.A(n_2618),
.Y(n_2939)
);

NAND2xp5_ASAP7_75t_L g2940 ( 
.A(n_2654),
.B(n_2375),
.Y(n_2940)
);

INVx2_ASAP7_75t_SL g2941 ( 
.A(n_2697),
.Y(n_2941)
);

OAI22xp5_ASAP7_75t_SL g2942 ( 
.A1(n_2609),
.A2(n_2321),
.B1(n_2524),
.B2(n_2197),
.Y(n_2942)
);

INVx1_ASAP7_75t_L g2943 ( 
.A(n_2620),
.Y(n_2943)
);

INVx3_ASAP7_75t_L g2944 ( 
.A(n_2591),
.Y(n_2944)
);

INVx1_ASAP7_75t_L g2945 ( 
.A(n_2641),
.Y(n_2945)
);

INVx1_ASAP7_75t_L g2946 ( 
.A(n_2641),
.Y(n_2946)
);

INVx1_ASAP7_75t_L g2947 ( 
.A(n_2577),
.Y(n_2947)
);

OR2x2_ASAP7_75t_L g2948 ( 
.A(n_2582),
.B(n_2289),
.Y(n_2948)
);

AND2x2_ASAP7_75t_L g2949 ( 
.A(n_2591),
.B(n_2211),
.Y(n_2949)
);

INVx1_ASAP7_75t_L g2950 ( 
.A(n_2585),
.Y(n_2950)
);

INVx4_ASAP7_75t_L g2951 ( 
.A(n_2603),
.Y(n_2951)
);

OAI22xp5_ASAP7_75t_L g2952 ( 
.A1(n_2612),
.A2(n_2468),
.B1(n_2197),
.B2(n_2446),
.Y(n_2952)
);

AND2x2_ASAP7_75t_L g2953 ( 
.A(n_2599),
.B(n_2248),
.Y(n_2953)
);

BUFx3_ASAP7_75t_L g2954 ( 
.A(n_2726),
.Y(n_2954)
);

INVx4_ASAP7_75t_R g2955 ( 
.A(n_2561),
.Y(n_2955)
);

NAND2xp5_ASAP7_75t_L g2956 ( 
.A(n_2588),
.B(n_2380),
.Y(n_2956)
);

INVx1_ASAP7_75t_L g2957 ( 
.A(n_2589),
.Y(n_2957)
);

INVx1_ASAP7_75t_L g2958 ( 
.A(n_2715),
.Y(n_2958)
);

INVx3_ASAP7_75t_L g2959 ( 
.A(n_2639),
.Y(n_2959)
);

INVx1_ASAP7_75t_L g2960 ( 
.A(n_2670),
.Y(n_2960)
);

AND2x2_ASAP7_75t_L g2961 ( 
.A(n_2742),
.B(n_2377),
.Y(n_2961)
);

INVx1_ASAP7_75t_L g2962 ( 
.A(n_2613),
.Y(n_2962)
);

INVx2_ASAP7_75t_SL g2963 ( 
.A(n_2608),
.Y(n_2963)
);

NOR2x1_ASAP7_75t_L g2964 ( 
.A(n_2633),
.B(n_2772),
.Y(n_2964)
);

HB1xp67_ASAP7_75t_L g2965 ( 
.A(n_2666),
.Y(n_2965)
);

AND2x4_ASAP7_75t_L g2966 ( 
.A(n_2714),
.B(n_2327),
.Y(n_2966)
);

AND2x4_ASAP7_75t_L g2967 ( 
.A(n_2701),
.B(n_2327),
.Y(n_2967)
);

AND2x2_ASAP7_75t_L g2968 ( 
.A(n_2716),
.B(n_2721),
.Y(n_2968)
);

AND2x2_ASAP7_75t_L g2969 ( 
.A(n_2716),
.B(n_2721),
.Y(n_2969)
);

AND2x2_ASAP7_75t_L g2970 ( 
.A(n_2634),
.B(n_2309),
.Y(n_2970)
);

AOI22xp5_ASAP7_75t_L g2971 ( 
.A1(n_2631),
.A2(n_2452),
.B1(n_2466),
.B2(n_2380),
.Y(n_2971)
);

AND2x4_ASAP7_75t_L g2972 ( 
.A(n_2701),
.B(n_2326),
.Y(n_2972)
);

NAND2xp5_ASAP7_75t_L g2973 ( 
.A(n_2624),
.B(n_2735),
.Y(n_2973)
);

INVx1_ASAP7_75t_L g2974 ( 
.A(n_2622),
.Y(n_2974)
);

NOR2xp33_ASAP7_75t_L g2975 ( 
.A(n_2756),
.B(n_2228),
.Y(n_2975)
);

CKINVDCx14_ASAP7_75t_R g2976 ( 
.A(n_2667),
.Y(n_2976)
);

CKINVDCx6p67_ASAP7_75t_R g2977 ( 
.A(n_2667),
.Y(n_2977)
);

AND2x2_ASAP7_75t_L g2978 ( 
.A(n_2744),
.B(n_2309),
.Y(n_2978)
);

OAI21xp33_ASAP7_75t_L g2979 ( 
.A1(n_2624),
.A2(n_2499),
.B(n_2235),
.Y(n_2979)
);

INVx1_ASAP7_75t_L g2980 ( 
.A(n_2672),
.Y(n_2980)
);

AND2x2_ASAP7_75t_L g2981 ( 
.A(n_2688),
.B(n_2428),
.Y(n_2981)
);

AND2x4_ASAP7_75t_L g2982 ( 
.A(n_2722),
.B(n_2343),
.Y(n_2982)
);

AND2x2_ASAP7_75t_L g2983 ( 
.A(n_2691),
.B(n_2494),
.Y(n_2983)
);

NAND2xp5_ASAP7_75t_L g2984 ( 
.A(n_2735),
.B(n_2489),
.Y(n_2984)
);

INVx1_ASAP7_75t_L g2985 ( 
.A(n_2674),
.Y(n_2985)
);

BUFx3_ASAP7_75t_L g2986 ( 
.A(n_2762),
.Y(n_2986)
);

AND2x2_ASAP7_75t_L g2987 ( 
.A(n_2605),
.B(n_2494),
.Y(n_2987)
);

AND2x2_ASAP7_75t_L g2988 ( 
.A(n_2605),
.B(n_2371),
.Y(n_2988)
);

AND2x4_ASAP7_75t_L g2989 ( 
.A(n_2722),
.B(n_2343),
.Y(n_2989)
);

OAI22xp5_ASAP7_75t_L g2990 ( 
.A1(n_2600),
.A2(n_2468),
.B1(n_2469),
.B2(n_2466),
.Y(n_2990)
);

INVx3_ASAP7_75t_L g2991 ( 
.A(n_2639),
.Y(n_2991)
);

INVx1_ASAP7_75t_L g2992 ( 
.A(n_2755),
.Y(n_2992)
);

AND2x2_ASAP7_75t_L g2993 ( 
.A(n_2648),
.B(n_2371),
.Y(n_2993)
);

INVx2_ASAP7_75t_SL g2994 ( 
.A(n_2573),
.Y(n_2994)
);

BUFx2_ASAP7_75t_L g2995 ( 
.A(n_2779),
.Y(n_2995)
);

INVx1_ASAP7_75t_L g2996 ( 
.A(n_2755),
.Y(n_2996)
);

NOR2xp33_ASAP7_75t_L g2997 ( 
.A(n_2601),
.B(n_2524),
.Y(n_2997)
);

INVx1_ASAP7_75t_L g2998 ( 
.A(n_2764),
.Y(n_2998)
);

AND2x2_ASAP7_75t_L g2999 ( 
.A(n_2648),
.B(n_2661),
.Y(n_2999)
);

INVx4_ASAP7_75t_L g3000 ( 
.A(n_2573),
.Y(n_3000)
);

AND2x2_ASAP7_75t_L g3001 ( 
.A(n_2661),
.B(n_2371),
.Y(n_3001)
);

AND2x2_ASAP7_75t_L g3002 ( 
.A(n_2678),
.B(n_2371),
.Y(n_3002)
);

HB1xp67_ASAP7_75t_L g3003 ( 
.A(n_2764),
.Y(n_3003)
);

INVx1_ASAP7_75t_L g3004 ( 
.A(n_2628),
.Y(n_3004)
);

INVx1_ASAP7_75t_L g3005 ( 
.A(n_2652),
.Y(n_3005)
);

AND2x4_ASAP7_75t_SL g3006 ( 
.A(n_2937),
.B(n_2876),
.Y(n_3006)
);

INVx1_ASAP7_75t_L g3007 ( 
.A(n_2782),
.Y(n_3007)
);

AND2x2_ASAP7_75t_L g3008 ( 
.A(n_2914),
.B(n_2736),
.Y(n_3008)
);

OR2x2_ASAP7_75t_L g3009 ( 
.A(n_2804),
.B(n_2720),
.Y(n_3009)
);

NAND2xp5_ASAP7_75t_L g3010 ( 
.A(n_2780),
.B(n_2681),
.Y(n_3010)
);

AND2x2_ASAP7_75t_L g3011 ( 
.A(n_2781),
.B(n_2720),
.Y(n_3011)
);

NAND2xp5_ASAP7_75t_L g3012 ( 
.A(n_2780),
.B(n_2682),
.Y(n_3012)
);

AND2x4_ASAP7_75t_L g3013 ( 
.A(n_2860),
.B(n_2731),
.Y(n_3013)
);

INVx1_ASAP7_75t_L g3014 ( 
.A(n_2793),
.Y(n_3014)
);

AND2x2_ASAP7_75t_L g3015 ( 
.A(n_2958),
.B(n_2731),
.Y(n_3015)
);

INVx1_ASAP7_75t_L g3016 ( 
.A(n_2797),
.Y(n_3016)
);

NAND2xp5_ASAP7_75t_L g3017 ( 
.A(n_2894),
.B(n_2684),
.Y(n_3017)
);

OR2x2_ASAP7_75t_L g3018 ( 
.A(n_2789),
.B(n_2540),
.Y(n_3018)
);

NAND2xp5_ASAP7_75t_L g3019 ( 
.A(n_2894),
.B(n_2685),
.Y(n_3019)
);

INVx1_ASAP7_75t_L g3020 ( 
.A(n_2803),
.Y(n_3020)
);

AND2x2_ASAP7_75t_L g3021 ( 
.A(n_2799),
.B(n_2653),
.Y(n_3021)
);

INVx2_ASAP7_75t_L g3022 ( 
.A(n_2897),
.Y(n_3022)
);

AND2x2_ASAP7_75t_L g3023 ( 
.A(n_2870),
.B(n_2653),
.Y(n_3023)
);

INVx1_ASAP7_75t_L g3024 ( 
.A(n_2810),
.Y(n_3024)
);

AND2x2_ASAP7_75t_L g3025 ( 
.A(n_2843),
.B(n_2740),
.Y(n_3025)
);

NAND2xp5_ASAP7_75t_L g3026 ( 
.A(n_2983),
.B(n_2754),
.Y(n_3026)
);

INVx1_ASAP7_75t_L g3027 ( 
.A(n_2811),
.Y(n_3027)
);

INVx2_ASAP7_75t_SL g3028 ( 
.A(n_2846),
.Y(n_3028)
);

INVx1_ASAP7_75t_L g3029 ( 
.A(n_2815),
.Y(n_3029)
);

INVxp67_ASAP7_75t_SL g3030 ( 
.A(n_2919),
.Y(n_3030)
);

AND2x2_ASAP7_75t_L g3031 ( 
.A(n_2883),
.B(n_2791),
.Y(n_3031)
);

INVx1_ASAP7_75t_L g3032 ( 
.A(n_2817),
.Y(n_3032)
);

AND2x4_ASAP7_75t_L g3033 ( 
.A(n_2891),
.B(n_2544),
.Y(n_3033)
);

INVx1_ASAP7_75t_L g3034 ( 
.A(n_2849),
.Y(n_3034)
);

NAND2xp5_ASAP7_75t_L g3035 ( 
.A(n_2820),
.B(n_2760),
.Y(n_3035)
);

AND2x4_ASAP7_75t_L g3036 ( 
.A(n_2891),
.B(n_2544),
.Y(n_3036)
);

INVxp67_ASAP7_75t_SL g3037 ( 
.A(n_2919),
.Y(n_3037)
);

NAND2xp5_ASAP7_75t_L g3038 ( 
.A(n_2916),
.B(n_2761),
.Y(n_3038)
);

INVx1_ASAP7_75t_L g3039 ( 
.A(n_2851),
.Y(n_3039)
);

AND2x2_ASAP7_75t_L g3040 ( 
.A(n_2785),
.B(n_2740),
.Y(n_3040)
);

OAI222xp33_ASAP7_75t_L g3041 ( 
.A1(n_2790),
.A2(n_2601),
.B1(n_2673),
.B2(n_2579),
.C1(n_2775),
.C2(n_2759),
.Y(n_3041)
);

AND2x2_ASAP7_75t_L g3042 ( 
.A(n_2786),
.B(n_2779),
.Y(n_3042)
);

HB1xp67_ASAP7_75t_L g3043 ( 
.A(n_3003),
.Y(n_3043)
);

INVx1_ASAP7_75t_L g3044 ( 
.A(n_2821),
.Y(n_3044)
);

INVx1_ASAP7_75t_L g3045 ( 
.A(n_2822),
.Y(n_3045)
);

INVx1_ASAP7_75t_L g3046 ( 
.A(n_2824),
.Y(n_3046)
);

INVx1_ASAP7_75t_L g3047 ( 
.A(n_2827),
.Y(n_3047)
);

INVx1_ASAP7_75t_L g3048 ( 
.A(n_2830),
.Y(n_3048)
);

AND2x2_ASAP7_75t_L g3049 ( 
.A(n_2902),
.B(n_2540),
.Y(n_3049)
);

AOI22xp33_ASAP7_75t_L g3050 ( 
.A1(n_2790),
.A2(n_2759),
.B1(n_2579),
.B2(n_2452),
.Y(n_3050)
);

INVx1_ASAP7_75t_L g3051 ( 
.A(n_2833),
.Y(n_3051)
);

AND2x2_ASAP7_75t_L g3052 ( 
.A(n_2960),
.B(n_2614),
.Y(n_3052)
);

INVx1_ASAP7_75t_L g3053 ( 
.A(n_2835),
.Y(n_3053)
);

OAI22xp33_ASAP7_75t_SL g3054 ( 
.A1(n_2867),
.A2(n_2656),
.B1(n_2771),
.B2(n_2767),
.Y(n_3054)
);

INVx1_ASAP7_75t_L g3055 ( 
.A(n_2837),
.Y(n_3055)
);

INVx1_ASAP7_75t_L g3056 ( 
.A(n_2818),
.Y(n_3056)
);

INVx1_ASAP7_75t_L g3057 ( 
.A(n_2819),
.Y(n_3057)
);

INVx2_ASAP7_75t_SL g3058 ( 
.A(n_2861),
.Y(n_3058)
);

AND2x2_ASAP7_75t_L g3059 ( 
.A(n_2825),
.B(n_2619),
.Y(n_3059)
);

OR2x2_ASAP7_75t_L g3060 ( 
.A(n_2826),
.B(n_2770),
.Y(n_3060)
);

INVx1_ASAP7_75t_L g3061 ( 
.A(n_2947),
.Y(n_3061)
);

NAND2xp33_ASAP7_75t_L g3062 ( 
.A(n_2850),
.B(n_2202),
.Y(n_3062)
);

OR2x2_ASAP7_75t_L g3063 ( 
.A(n_2826),
.B(n_2660),
.Y(n_3063)
);

INVx1_ASAP7_75t_L g3064 ( 
.A(n_2950),
.Y(n_3064)
);

AND2x2_ASAP7_75t_L g3065 ( 
.A(n_2832),
.B(n_2627),
.Y(n_3065)
);

AOI22xp33_ASAP7_75t_L g3066 ( 
.A1(n_2866),
.A2(n_2452),
.B1(n_2466),
.B2(n_2673),
.Y(n_3066)
);

AND2x2_ASAP7_75t_L g3067 ( 
.A(n_2868),
.B(n_2629),
.Y(n_3067)
);

BUFx3_ASAP7_75t_L g3068 ( 
.A(n_2881),
.Y(n_3068)
);

AND2x4_ASAP7_75t_L g3069 ( 
.A(n_2828),
.B(n_2925),
.Y(n_3069)
);

INVx1_ASAP7_75t_L g3070 ( 
.A(n_2957),
.Y(n_3070)
);

AND2x2_ASAP7_75t_L g3071 ( 
.A(n_2868),
.B(n_2637),
.Y(n_3071)
);

HB1xp67_ASAP7_75t_L g3072 ( 
.A(n_3003),
.Y(n_3072)
);

AND2x2_ASAP7_75t_L g3073 ( 
.A(n_2931),
.B(n_2642),
.Y(n_3073)
);

INVx1_ASAP7_75t_L g3074 ( 
.A(n_2823),
.Y(n_3074)
);

HB1xp67_ASAP7_75t_L g3075 ( 
.A(n_2812),
.Y(n_3075)
);

OR2x2_ASAP7_75t_L g3076 ( 
.A(n_2862),
.B(n_2647),
.Y(n_3076)
);

INVx1_ASAP7_75t_L g3077 ( 
.A(n_2823),
.Y(n_3077)
);

BUFx2_ASAP7_75t_L g3078 ( 
.A(n_2850),
.Y(n_3078)
);

AND2x2_ASAP7_75t_L g3079 ( 
.A(n_2933),
.B(n_2678),
.Y(n_3079)
);

NAND2xp5_ASAP7_75t_L g3080 ( 
.A(n_2865),
.B(n_2741),
.Y(n_3080)
);

AOI22xp33_ASAP7_75t_SL g3081 ( 
.A1(n_2869),
.A2(n_2202),
.B1(n_2499),
.B2(n_2200),
.Y(n_3081)
);

INVx1_ASAP7_75t_L g3082 ( 
.A(n_2840),
.Y(n_3082)
);

INVx1_ASAP7_75t_L g3083 ( 
.A(n_2842),
.Y(n_3083)
);

OAI222xp33_ASAP7_75t_L g3084 ( 
.A1(n_2869),
.A2(n_2775),
.B1(n_2646),
.B2(n_2703),
.C1(n_2710),
.C2(n_2711),
.Y(n_3084)
);

AND2x2_ASAP7_75t_L g3085 ( 
.A(n_2938),
.B(n_2981),
.Y(n_3085)
);

HB1xp67_ASAP7_75t_L g3086 ( 
.A(n_2812),
.Y(n_3086)
);

HB1xp67_ASAP7_75t_L g3087 ( 
.A(n_2816),
.Y(n_3087)
);

OR2x2_ASAP7_75t_L g3088 ( 
.A(n_2872),
.B(n_2738),
.Y(n_3088)
);

INVx1_ASAP7_75t_L g3089 ( 
.A(n_2847),
.Y(n_3089)
);

AND2x2_ASAP7_75t_L g3090 ( 
.A(n_2923),
.B(n_2694),
.Y(n_3090)
);

OR2x2_ASAP7_75t_L g3091 ( 
.A(n_2875),
.B(n_2739),
.Y(n_3091)
);

NAND2xp5_ASAP7_75t_L g3092 ( 
.A(n_2880),
.B(n_2733),
.Y(n_3092)
);

BUFx3_ASAP7_75t_L g3093 ( 
.A(n_2885),
.Y(n_3093)
);

INVx1_ASAP7_75t_L g3094 ( 
.A(n_2848),
.Y(n_3094)
);

AND2x2_ASAP7_75t_L g3095 ( 
.A(n_2904),
.B(n_2694),
.Y(n_3095)
);

INVx1_ASAP7_75t_L g3096 ( 
.A(n_2900),
.Y(n_3096)
);

AND2x2_ASAP7_75t_L g3097 ( 
.A(n_2904),
.B(n_2696),
.Y(n_3097)
);

OAI22xp5_ASAP7_75t_L g3098 ( 
.A1(n_2784),
.A2(n_2747),
.B1(n_2752),
.B2(n_2753),
.Y(n_3098)
);

OR2x2_ASAP7_75t_L g3099 ( 
.A(n_2884),
.B(n_2566),
.Y(n_3099)
);

AND2x2_ASAP7_75t_L g3100 ( 
.A(n_3005),
.B(n_2696),
.Y(n_3100)
);

AND2x2_ASAP7_75t_L g3101 ( 
.A(n_2813),
.B(n_2733),
.Y(n_3101)
);

INVx4_ASAP7_75t_L g3102 ( 
.A(n_2937),
.Y(n_3102)
);

NAND2xp5_ASAP7_75t_L g3103 ( 
.A(n_2956),
.B(n_2773),
.Y(n_3103)
);

INVx1_ASAP7_75t_L g3104 ( 
.A(n_2943),
.Y(n_3104)
);

AND2x2_ASAP7_75t_L g3105 ( 
.A(n_2814),
.B(n_2531),
.Y(n_3105)
);

AND2x4_ASAP7_75t_L g3106 ( 
.A(n_2828),
.B(n_2547),
.Y(n_3106)
);

BUFx6f_ASAP7_75t_L g3107 ( 
.A(n_2921),
.Y(n_3107)
);

INVxp67_ASAP7_75t_SL g3108 ( 
.A(n_2882),
.Y(n_3108)
);

INVx3_ASAP7_75t_L g3109 ( 
.A(n_2794),
.Y(n_3109)
);

AOI22xp33_ASAP7_75t_L g3110 ( 
.A1(n_2866),
.A2(n_2997),
.B1(n_2975),
.B2(n_2973),
.Y(n_3110)
);

AND2x2_ASAP7_75t_L g3111 ( 
.A(n_2807),
.B(n_2531),
.Y(n_3111)
);

NAND2xp5_ASAP7_75t_L g3112 ( 
.A(n_2956),
.B(n_2773),
.Y(n_3112)
);

INVx1_ASAP7_75t_L g3113 ( 
.A(n_2945),
.Y(n_3113)
);

OR2x6_ASAP7_75t_SL g3114 ( 
.A(n_2906),
.B(n_2732),
.Y(n_3114)
);

INVxp67_ASAP7_75t_SL g3115 ( 
.A(n_2882),
.Y(n_3115)
);

INVx2_ASAP7_75t_SL g3116 ( 
.A(n_2955),
.Y(n_3116)
);

NAND2xp5_ASAP7_75t_L g3117 ( 
.A(n_2973),
.B(n_2587),
.Y(n_3117)
);

HB1xp67_ASAP7_75t_L g3118 ( 
.A(n_2816),
.Y(n_3118)
);

INVx1_ASAP7_75t_L g3119 ( 
.A(n_2946),
.Y(n_3119)
);

AND2x2_ASAP7_75t_L g3120 ( 
.A(n_2980),
.B(n_2689),
.Y(n_3120)
);

INVx1_ASAP7_75t_L g3121 ( 
.A(n_2854),
.Y(n_3121)
);

AND2x2_ASAP7_75t_L g3122 ( 
.A(n_2985),
.B(n_2537),
.Y(n_3122)
);

INVx1_ASAP7_75t_L g3123 ( 
.A(n_2879),
.Y(n_3123)
);

AND2x2_ASAP7_75t_L g3124 ( 
.A(n_2911),
.B(n_2537),
.Y(n_3124)
);

INVx1_ASAP7_75t_L g3125 ( 
.A(n_2905),
.Y(n_3125)
);

AND2x2_ASAP7_75t_L g3126 ( 
.A(n_2885),
.B(n_2616),
.Y(n_3126)
);

NAND2xp5_ASAP7_75t_L g3127 ( 
.A(n_2864),
.B(n_2587),
.Y(n_3127)
);

INVx1_ASAP7_75t_L g3128 ( 
.A(n_2908),
.Y(n_3128)
);

NAND2xp5_ASAP7_75t_L g3129 ( 
.A(n_2864),
.B(n_2693),
.Y(n_3129)
);

INVx1_ASAP7_75t_L g3130 ( 
.A(n_2910),
.Y(n_3130)
);

INVx1_ASAP7_75t_L g3131 ( 
.A(n_2924),
.Y(n_3131)
);

INVx1_ASAP7_75t_L g3132 ( 
.A(n_2932),
.Y(n_3132)
);

NAND2xp5_ASAP7_75t_L g3133 ( 
.A(n_2871),
.B(n_2695),
.Y(n_3133)
);

HB1xp67_ASAP7_75t_L g3134 ( 
.A(n_2829),
.Y(n_3134)
);

AND2x2_ASAP7_75t_L g3135 ( 
.A(n_2928),
.B(n_2617),
.Y(n_3135)
);

BUFx2_ASAP7_75t_L g3136 ( 
.A(n_3000),
.Y(n_3136)
);

AND2x2_ASAP7_75t_L g3137 ( 
.A(n_2844),
.B(n_2547),
.Y(n_3137)
);

AOI22xp33_ASAP7_75t_SL g3138 ( 
.A1(n_2942),
.A2(n_2202),
.B1(n_2200),
.B2(n_2240),
.Y(n_3138)
);

AND2x2_ASAP7_75t_L g3139 ( 
.A(n_2995),
.B(n_2774),
.Y(n_3139)
);

AND2x2_ASAP7_75t_L g3140 ( 
.A(n_2889),
.B(n_2918),
.Y(n_3140)
);

NAND2xp5_ASAP7_75t_L g3141 ( 
.A(n_2871),
.B(n_2704),
.Y(n_3141)
);

AND2x4_ASAP7_75t_L g3142 ( 
.A(n_2836),
.B(n_2548),
.Y(n_3142)
);

NAND2xp5_ASAP7_75t_L g3143 ( 
.A(n_2878),
.B(n_2705),
.Y(n_3143)
);

INVx1_ASAP7_75t_L g3144 ( 
.A(n_2935),
.Y(n_3144)
);

AO22x1_ASAP7_75t_L g3145 ( 
.A1(n_2997),
.A2(n_2636),
.B1(n_2604),
.B2(n_2758),
.Y(n_3145)
);

NAND2xp5_ASAP7_75t_L g3146 ( 
.A(n_2878),
.B(n_2707),
.Y(n_3146)
);

INVx1_ASAP7_75t_L g3147 ( 
.A(n_2992),
.Y(n_3147)
);

BUFx3_ASAP7_75t_L g3148 ( 
.A(n_2907),
.Y(n_3148)
);

AND2x2_ASAP7_75t_L g3149 ( 
.A(n_2889),
.B(n_2774),
.Y(n_3149)
);

AND2x2_ASAP7_75t_L g3150 ( 
.A(n_2829),
.B(n_2548),
.Y(n_3150)
);

AND2x2_ASAP7_75t_L g3151 ( 
.A(n_2838),
.B(n_2712),
.Y(n_3151)
);

INVx4_ASAP7_75t_L g3152 ( 
.A(n_3000),
.Y(n_3152)
);

AND2x2_ASAP7_75t_L g3153 ( 
.A(n_2838),
.B(n_2713),
.Y(n_3153)
);

NOR2xp33_ASAP7_75t_L g3154 ( 
.A(n_2975),
.B(n_2604),
.Y(n_3154)
);

NAND2x1p5_ASAP7_75t_L g3155 ( 
.A(n_3152),
.B(n_2801),
.Y(n_3155)
);

NAND2xp5_ASAP7_75t_L g3156 ( 
.A(n_3117),
.B(n_2787),
.Y(n_3156)
);

INVx1_ASAP7_75t_L g3157 ( 
.A(n_3034),
.Y(n_3157)
);

INVx2_ASAP7_75t_L g3158 ( 
.A(n_3030),
.Y(n_3158)
);

INVx2_ASAP7_75t_L g3159 ( 
.A(n_3030),
.Y(n_3159)
);

INVx1_ASAP7_75t_L g3160 ( 
.A(n_3039),
.Y(n_3160)
);

AND2x2_ASAP7_75t_L g3161 ( 
.A(n_3031),
.B(n_2913),
.Y(n_3161)
);

INVx1_ASAP7_75t_L g3162 ( 
.A(n_3007),
.Y(n_3162)
);

AND2x2_ASAP7_75t_L g3163 ( 
.A(n_3135),
.B(n_2929),
.Y(n_3163)
);

AND2x2_ASAP7_75t_L g3164 ( 
.A(n_3008),
.B(n_2917),
.Y(n_3164)
);

INVx2_ASAP7_75t_SL g3165 ( 
.A(n_3068),
.Y(n_3165)
);

OR2x2_ASAP7_75t_L g3166 ( 
.A(n_3035),
.B(n_3009),
.Y(n_3166)
);

BUFx3_ASAP7_75t_L g3167 ( 
.A(n_3068),
.Y(n_3167)
);

NAND2xp5_ASAP7_75t_L g3168 ( 
.A(n_3117),
.B(n_2787),
.Y(n_3168)
);

BUFx2_ASAP7_75t_L g3169 ( 
.A(n_3136),
.Y(n_3169)
);

NAND2xp5_ASAP7_75t_L g3170 ( 
.A(n_3121),
.B(n_2800),
.Y(n_3170)
);

INVx1_ASAP7_75t_L g3171 ( 
.A(n_3014),
.Y(n_3171)
);

AND2x2_ASAP7_75t_L g3172 ( 
.A(n_3079),
.B(n_2922),
.Y(n_3172)
);

INVx3_ASAP7_75t_L g3173 ( 
.A(n_3152),
.Y(n_3173)
);

AND2x2_ASAP7_75t_L g3174 ( 
.A(n_3025),
.B(n_2898),
.Y(n_3174)
);

OR2x2_ASAP7_75t_L g3175 ( 
.A(n_3035),
.B(n_3038),
.Y(n_3175)
);

INVx1_ASAP7_75t_L g3176 ( 
.A(n_3016),
.Y(n_3176)
);

OR2x2_ASAP7_75t_L g3177 ( 
.A(n_3038),
.B(n_2858),
.Y(n_3177)
);

AOI221xp5_ASAP7_75t_L g3178 ( 
.A1(n_3110),
.A2(n_2788),
.B1(n_2839),
.B2(n_2927),
.C(n_2976),
.Y(n_3178)
);

AND2x4_ASAP7_75t_L g3179 ( 
.A(n_3093),
.B(n_2987),
.Y(n_3179)
);

BUFx3_ASAP7_75t_L g3180 ( 
.A(n_3028),
.Y(n_3180)
);

OR2x2_ASAP7_75t_L g3181 ( 
.A(n_3123),
.B(n_2855),
.Y(n_3181)
);

HB1xp67_ASAP7_75t_L g3182 ( 
.A(n_3075),
.Y(n_3182)
);

INVx1_ASAP7_75t_L g3183 ( 
.A(n_3020),
.Y(n_3183)
);

BUFx2_ASAP7_75t_L g3184 ( 
.A(n_3102),
.Y(n_3184)
);

NAND2xp5_ASAP7_75t_L g3185 ( 
.A(n_3074),
.B(n_2800),
.Y(n_3185)
);

OR2x2_ASAP7_75t_L g3186 ( 
.A(n_3077),
.B(n_2855),
.Y(n_3186)
);

AND2x2_ASAP7_75t_L g3187 ( 
.A(n_3140),
.B(n_3011),
.Y(n_3187)
);

NAND2xp5_ASAP7_75t_L g3188 ( 
.A(n_3017),
.B(n_2978),
.Y(n_3188)
);

BUFx2_ASAP7_75t_L g3189 ( 
.A(n_3102),
.Y(n_3189)
);

NOR2xp33_ASAP7_75t_L g3190 ( 
.A(n_3154),
.B(n_2951),
.Y(n_3190)
);

AND2x4_ASAP7_75t_L g3191 ( 
.A(n_3093),
.B(n_2836),
.Y(n_3191)
);

HB1xp67_ASAP7_75t_L g3192 ( 
.A(n_3075),
.Y(n_3192)
);

INVx1_ASAP7_75t_L g3193 ( 
.A(n_3024),
.Y(n_3193)
);

NAND3xp33_ASAP7_75t_L g3194 ( 
.A(n_3110),
.B(n_2792),
.C(n_2784),
.Y(n_3194)
);

INVx1_ASAP7_75t_L g3195 ( 
.A(n_3027),
.Y(n_3195)
);

NAND2xp5_ASAP7_75t_L g3196 ( 
.A(n_3017),
.B(n_2831),
.Y(n_3196)
);

AND2x2_ASAP7_75t_L g3197 ( 
.A(n_3073),
.B(n_2893),
.Y(n_3197)
);

NAND2xp5_ASAP7_75t_L g3198 ( 
.A(n_3019),
.B(n_3049),
.Y(n_3198)
);

INVxp67_ASAP7_75t_L g3199 ( 
.A(n_3037),
.Y(n_3199)
);

NAND2xp5_ASAP7_75t_L g3200 ( 
.A(n_3019),
.B(n_2831),
.Y(n_3200)
);

INVx1_ASAP7_75t_L g3201 ( 
.A(n_3029),
.Y(n_3201)
);

INVx1_ASAP7_75t_L g3202 ( 
.A(n_3032),
.Y(n_3202)
);

INVx2_ASAP7_75t_L g3203 ( 
.A(n_3037),
.Y(n_3203)
);

AND2x4_ASAP7_75t_L g3204 ( 
.A(n_3106),
.B(n_2857),
.Y(n_3204)
);

INVx1_ASAP7_75t_L g3205 ( 
.A(n_3044),
.Y(n_3205)
);

INVx2_ASAP7_75t_L g3206 ( 
.A(n_3043),
.Y(n_3206)
);

AND2x2_ASAP7_75t_L g3207 ( 
.A(n_3085),
.B(n_3023),
.Y(n_3207)
);

OR2x2_ASAP7_75t_L g3208 ( 
.A(n_3026),
.B(n_2893),
.Y(n_3208)
);

AND2x2_ASAP7_75t_L g3209 ( 
.A(n_3137),
.B(n_2909),
.Y(n_3209)
);

INVx1_ASAP7_75t_L g3210 ( 
.A(n_3045),
.Y(n_3210)
);

AND2x2_ASAP7_75t_L g3211 ( 
.A(n_3015),
.B(n_2909),
.Y(n_3211)
);

INVx1_ASAP7_75t_L g3212 ( 
.A(n_3046),
.Y(n_3212)
);

INVx1_ASAP7_75t_L g3213 ( 
.A(n_3047),
.Y(n_3213)
);

INVx2_ASAP7_75t_L g3214 ( 
.A(n_3043),
.Y(n_3214)
);

INVx3_ASAP7_75t_R g3215 ( 
.A(n_3088),
.Y(n_3215)
);

AND2x2_ASAP7_75t_L g3216 ( 
.A(n_3059),
.B(n_2915),
.Y(n_3216)
);

NAND2xp5_ASAP7_75t_L g3217 ( 
.A(n_3010),
.B(n_2934),
.Y(n_3217)
);

OR2x2_ASAP7_75t_L g3218 ( 
.A(n_3026),
.B(n_3086),
.Y(n_3218)
);

INVx2_ASAP7_75t_L g3219 ( 
.A(n_3072),
.Y(n_3219)
);

NAND2xp5_ASAP7_75t_L g3220 ( 
.A(n_3010),
.B(n_2971),
.Y(n_3220)
);

BUFx6f_ASAP7_75t_L g3221 ( 
.A(n_3107),
.Y(n_3221)
);

AND2x2_ASAP7_75t_L g3222 ( 
.A(n_3065),
.B(n_2915),
.Y(n_3222)
);

AND2x2_ASAP7_75t_L g3223 ( 
.A(n_3069),
.B(n_2936),
.Y(n_3223)
);

HB1xp67_ASAP7_75t_L g3224 ( 
.A(n_3086),
.Y(n_3224)
);

AND2x4_ASAP7_75t_L g3225 ( 
.A(n_3106),
.B(n_3142),
.Y(n_3225)
);

INVx1_ASAP7_75t_L g3226 ( 
.A(n_3048),
.Y(n_3226)
);

AND2x2_ASAP7_75t_L g3227 ( 
.A(n_3069),
.B(n_3040),
.Y(n_3227)
);

INVx1_ASAP7_75t_L g3228 ( 
.A(n_3051),
.Y(n_3228)
);

NAND2xp5_ASAP7_75t_L g3229 ( 
.A(n_3012),
.B(n_2971),
.Y(n_3229)
);

AND2x2_ASAP7_75t_L g3230 ( 
.A(n_3101),
.B(n_2936),
.Y(n_3230)
);

INVx2_ASAP7_75t_L g3231 ( 
.A(n_3072),
.Y(n_3231)
);

NOR2xp33_ASAP7_75t_L g3232 ( 
.A(n_3154),
.B(n_2951),
.Y(n_3232)
);

OAI21xp5_ASAP7_75t_SL g3233 ( 
.A1(n_3006),
.A2(n_3041),
.B(n_3116),
.Y(n_3233)
);

NAND2xp5_ASAP7_75t_L g3234 ( 
.A(n_3012),
.B(n_2970),
.Y(n_3234)
);

OR2x2_ASAP7_75t_L g3235 ( 
.A(n_3087),
.B(n_2965),
.Y(n_3235)
);

INVx1_ASAP7_75t_L g3236 ( 
.A(n_3053),
.Y(n_3236)
);

INVx1_ASAP7_75t_L g3237 ( 
.A(n_3055),
.Y(n_3237)
);

OAI221xp5_ASAP7_75t_L g3238 ( 
.A1(n_3066),
.A2(n_2839),
.B1(n_2792),
.B2(n_2795),
.C(n_2942),
.Y(n_3238)
);

INVx1_ASAP7_75t_L g3239 ( 
.A(n_3082),
.Y(n_3239)
);

INVxp67_ASAP7_75t_L g3240 ( 
.A(n_3087),
.Y(n_3240)
);

INVx1_ASAP7_75t_L g3241 ( 
.A(n_3218),
.Y(n_3241)
);

AND2x2_ASAP7_75t_L g3242 ( 
.A(n_3227),
.B(n_3021),
.Y(n_3242)
);

OR2x2_ASAP7_75t_L g3243 ( 
.A(n_3175),
.B(n_3166),
.Y(n_3243)
);

NAND2xp5_ASAP7_75t_L g3244 ( 
.A(n_3198),
.B(n_3056),
.Y(n_3244)
);

AND2x4_ASAP7_75t_L g3245 ( 
.A(n_3225),
.B(n_3142),
.Y(n_3245)
);

INVx1_ASAP7_75t_L g3246 ( 
.A(n_3157),
.Y(n_3246)
);

INVx1_ASAP7_75t_L g3247 ( 
.A(n_3160),
.Y(n_3247)
);

INVx2_ASAP7_75t_L g3248 ( 
.A(n_3158),
.Y(n_3248)
);

AND2x2_ASAP7_75t_L g3249 ( 
.A(n_3187),
.B(n_3105),
.Y(n_3249)
);

AND2x2_ASAP7_75t_L g3250 ( 
.A(n_3161),
.B(n_3111),
.Y(n_3250)
);

INVxp67_ASAP7_75t_L g3251 ( 
.A(n_3169),
.Y(n_3251)
);

AND2x2_ASAP7_75t_L g3252 ( 
.A(n_3172),
.B(n_3124),
.Y(n_3252)
);

HB1xp67_ASAP7_75t_L g3253 ( 
.A(n_3199),
.Y(n_3253)
);

INVx1_ASAP7_75t_L g3254 ( 
.A(n_3162),
.Y(n_3254)
);

INVx1_ASAP7_75t_L g3255 ( 
.A(n_3171),
.Y(n_3255)
);

AND2x2_ASAP7_75t_L g3256 ( 
.A(n_3164),
.B(n_3067),
.Y(n_3256)
);

INVx1_ASAP7_75t_L g3257 ( 
.A(n_3176),
.Y(n_3257)
);

OAI221xp5_ASAP7_75t_SL g3258 ( 
.A1(n_3233),
.A2(n_3050),
.B1(n_3066),
.B2(n_3080),
.C(n_2976),
.Y(n_3258)
);

AOI32xp33_ASAP7_75t_L g3259 ( 
.A1(n_3184),
.A2(n_3006),
.A3(n_3058),
.B1(n_2852),
.B2(n_2964),
.Y(n_3259)
);

AND2x2_ASAP7_75t_L g3260 ( 
.A(n_3163),
.B(n_3223),
.Y(n_3260)
);

INVx2_ASAP7_75t_L g3261 ( 
.A(n_3159),
.Y(n_3261)
);

INVx1_ASAP7_75t_L g3262 ( 
.A(n_3183),
.Y(n_3262)
);

NAND2xp5_ASAP7_75t_L g3263 ( 
.A(n_3198),
.B(n_3057),
.Y(n_3263)
);

INVx1_ASAP7_75t_L g3264 ( 
.A(n_3193),
.Y(n_3264)
);

AND2x4_ASAP7_75t_L g3265 ( 
.A(n_3225),
.B(n_3204),
.Y(n_3265)
);

INVx1_ASAP7_75t_SL g3266 ( 
.A(n_3167),
.Y(n_3266)
);

INVx1_ASAP7_75t_L g3267 ( 
.A(n_3195),
.Y(n_3267)
);

NAND2xp5_ASAP7_75t_L g3268 ( 
.A(n_3211),
.B(n_3061),
.Y(n_3268)
);

BUFx3_ASAP7_75t_L g3269 ( 
.A(n_3189),
.Y(n_3269)
);

AND2x2_ASAP7_75t_L g3270 ( 
.A(n_3174),
.B(n_3071),
.Y(n_3270)
);

INVx1_ASAP7_75t_L g3271 ( 
.A(n_3201),
.Y(n_3271)
);

OAI21xp5_ASAP7_75t_L g3272 ( 
.A1(n_3233),
.A2(n_3054),
.B(n_3041),
.Y(n_3272)
);

AND2x2_ASAP7_75t_L g3273 ( 
.A(n_3207),
.B(n_3042),
.Y(n_3273)
);

NOR2xp33_ASAP7_75t_L g3274 ( 
.A(n_3215),
.B(n_3238),
.Y(n_3274)
);

OR2x2_ASAP7_75t_L g3275 ( 
.A(n_3177),
.B(n_3118),
.Y(n_3275)
);

INVxp67_ASAP7_75t_L g3276 ( 
.A(n_3182),
.Y(n_3276)
);

INVx3_ASAP7_75t_L g3277 ( 
.A(n_3173),
.Y(n_3277)
);

INVx1_ASAP7_75t_L g3278 ( 
.A(n_3202),
.Y(n_3278)
);

NOR2xp33_ASAP7_75t_L g3279 ( 
.A(n_3238),
.B(n_3080),
.Y(n_3279)
);

NOR2x1p5_ASAP7_75t_SL g3280 ( 
.A(n_3203),
.B(n_2853),
.Y(n_3280)
);

INVx2_ASAP7_75t_SL g3281 ( 
.A(n_3173),
.Y(n_3281)
);

INVx1_ASAP7_75t_L g3282 ( 
.A(n_3205),
.Y(n_3282)
);

AND2x4_ASAP7_75t_L g3283 ( 
.A(n_3204),
.B(n_3150),
.Y(n_3283)
);

AND2x2_ASAP7_75t_L g3284 ( 
.A(n_3230),
.B(n_3118),
.Y(n_3284)
);

AND2x2_ASAP7_75t_L g3285 ( 
.A(n_3209),
.B(n_3134),
.Y(n_3285)
);

INVx1_ASAP7_75t_L g3286 ( 
.A(n_3210),
.Y(n_3286)
);

AND2x2_ASAP7_75t_L g3287 ( 
.A(n_3216),
.B(n_3134),
.Y(n_3287)
);

INVx2_ASAP7_75t_L g3288 ( 
.A(n_3199),
.Y(n_3288)
);

INVx1_ASAP7_75t_L g3289 ( 
.A(n_3212),
.Y(n_3289)
);

INVxp67_ASAP7_75t_SL g3290 ( 
.A(n_3192),
.Y(n_3290)
);

AND2x4_ASAP7_75t_L g3291 ( 
.A(n_3179),
.B(n_3139),
.Y(n_3291)
);

INVx1_ASAP7_75t_SL g3292 ( 
.A(n_3180),
.Y(n_3292)
);

AOI22xp5_ASAP7_75t_L g3293 ( 
.A1(n_3194),
.A2(n_3013),
.B1(n_3145),
.B2(n_3050),
.Y(n_3293)
);

NAND2xp5_ASAP7_75t_L g3294 ( 
.A(n_3217),
.B(n_3064),
.Y(n_3294)
);

INVx1_ASAP7_75t_L g3295 ( 
.A(n_3213),
.Y(n_3295)
);

INVx1_ASAP7_75t_SL g3296 ( 
.A(n_3165),
.Y(n_3296)
);

INVx1_ASAP7_75t_L g3297 ( 
.A(n_3226),
.Y(n_3297)
);

BUFx3_ASAP7_75t_L g3298 ( 
.A(n_3155),
.Y(n_3298)
);

AND2x2_ASAP7_75t_L g3299 ( 
.A(n_3222),
.B(n_3090),
.Y(n_3299)
);

INVx1_ASAP7_75t_L g3300 ( 
.A(n_3228),
.Y(n_3300)
);

INVx2_ASAP7_75t_L g3301 ( 
.A(n_3236),
.Y(n_3301)
);

INVx1_ASAP7_75t_L g3302 ( 
.A(n_3237),
.Y(n_3302)
);

AND2x4_ASAP7_75t_L g3303 ( 
.A(n_3179),
.B(n_3033),
.Y(n_3303)
);

AND2x2_ASAP7_75t_L g3304 ( 
.A(n_3197),
.B(n_3191),
.Y(n_3304)
);

NAND2x1p5_ASAP7_75t_L g3305 ( 
.A(n_3191),
.B(n_3078),
.Y(n_3305)
);

HB1xp67_ASAP7_75t_L g3306 ( 
.A(n_3224),
.Y(n_3306)
);

INVx1_ASAP7_75t_L g3307 ( 
.A(n_3301),
.Y(n_3307)
);

OR2x2_ASAP7_75t_L g3308 ( 
.A(n_3243),
.B(n_3208),
.Y(n_3308)
);

OR2x2_ASAP7_75t_L g3309 ( 
.A(n_3275),
.B(n_3217),
.Y(n_3309)
);

INVx1_ASAP7_75t_L g3310 ( 
.A(n_3301),
.Y(n_3310)
);

INVx1_ASAP7_75t_L g3311 ( 
.A(n_3253),
.Y(n_3311)
);

OR2x2_ASAP7_75t_L g3312 ( 
.A(n_3241),
.B(n_3188),
.Y(n_3312)
);

INVx1_ASAP7_75t_L g3313 ( 
.A(n_3253),
.Y(n_3313)
);

OR2x2_ASAP7_75t_L g3314 ( 
.A(n_3268),
.B(n_3244),
.Y(n_3314)
);

INVx1_ASAP7_75t_L g3315 ( 
.A(n_3306),
.Y(n_3315)
);

INVx1_ASAP7_75t_L g3316 ( 
.A(n_3306),
.Y(n_3316)
);

INVx2_ASAP7_75t_L g3317 ( 
.A(n_3269),
.Y(n_3317)
);

AOI32xp33_ASAP7_75t_L g3318 ( 
.A1(n_3274),
.A2(n_3178),
.A3(n_3232),
.B1(n_3190),
.B2(n_3013),
.Y(n_3318)
);

NAND2x1_ASAP7_75t_L g3319 ( 
.A(n_3277),
.B(n_3109),
.Y(n_3319)
);

OAI21x1_ASAP7_75t_L g3320 ( 
.A1(n_3277),
.A2(n_3155),
.B(n_3109),
.Y(n_3320)
);

INVx1_ASAP7_75t_L g3321 ( 
.A(n_3246),
.Y(n_3321)
);

INVx1_ASAP7_75t_L g3322 ( 
.A(n_3247),
.Y(n_3322)
);

OAI22xp5_ASAP7_75t_L g3323 ( 
.A1(n_3258),
.A2(n_3178),
.B1(n_3194),
.B2(n_3081),
.Y(n_3323)
);

OAI22xp5_ASAP7_75t_L g3324 ( 
.A1(n_3258),
.A2(n_3081),
.B1(n_3138),
.B2(n_2795),
.Y(n_3324)
);

OR2x2_ASAP7_75t_L g3325 ( 
.A(n_3263),
.B(n_3188),
.Y(n_3325)
);

AOI22xp5_ASAP7_75t_L g3326 ( 
.A1(n_3279),
.A2(n_2788),
.B1(n_2963),
.B2(n_3062),
.Y(n_3326)
);

AOI32xp33_ASAP7_75t_L g3327 ( 
.A1(n_3274),
.A2(n_3062),
.A3(n_3138),
.B1(n_3148),
.B2(n_2798),
.Y(n_3327)
);

AND2x2_ASAP7_75t_L g3328 ( 
.A(n_3252),
.B(n_3240),
.Y(n_3328)
);

INVx1_ASAP7_75t_L g3329 ( 
.A(n_3254),
.Y(n_3329)
);

AND2x2_ASAP7_75t_L g3330 ( 
.A(n_3291),
.B(n_3240),
.Y(n_3330)
);

AND2x2_ASAP7_75t_L g3331 ( 
.A(n_3291),
.B(n_3206),
.Y(n_3331)
);

OAI22xp33_ASAP7_75t_L g3332 ( 
.A1(n_3272),
.A2(n_2798),
.B1(n_3148),
.B2(n_3018),
.Y(n_3332)
);

INVx2_ASAP7_75t_L g3333 ( 
.A(n_3269),
.Y(n_3333)
);

OAI211xp5_ASAP7_75t_L g3334 ( 
.A1(n_3259),
.A2(n_2732),
.B(n_2986),
.C(n_3220),
.Y(n_3334)
);

XOR2x2_ASAP7_75t_L g3335 ( 
.A(n_3279),
.B(n_2954),
.Y(n_3335)
);

NAND3xp33_ASAP7_75t_SL g3336 ( 
.A(n_3292),
.B(n_2906),
.C(n_2762),
.Y(n_3336)
);

INVxp67_ASAP7_75t_SL g3337 ( 
.A(n_3251),
.Y(n_3337)
);

INVx1_ASAP7_75t_SL g3338 ( 
.A(n_3266),
.Y(n_3338)
);

INVx2_ASAP7_75t_SL g3339 ( 
.A(n_3296),
.Y(n_3339)
);

INVx1_ASAP7_75t_L g3340 ( 
.A(n_3255),
.Y(n_3340)
);

NAND2xp5_ASAP7_75t_SL g3341 ( 
.A(n_3298),
.B(n_2783),
.Y(n_3341)
);

AND2x2_ASAP7_75t_L g3342 ( 
.A(n_3291),
.B(n_3214),
.Y(n_3342)
);

INVx2_ASAP7_75t_L g3343 ( 
.A(n_3288),
.Y(n_3343)
);

OR2x2_ASAP7_75t_L g3344 ( 
.A(n_3290),
.B(n_3170),
.Y(n_3344)
);

INVx1_ASAP7_75t_L g3345 ( 
.A(n_3257),
.Y(n_3345)
);

NAND2xp5_ASAP7_75t_L g3346 ( 
.A(n_3276),
.B(n_3156),
.Y(n_3346)
);

AOI22xp33_ASAP7_75t_L g3347 ( 
.A1(n_3293),
.A2(n_3229),
.B1(n_3220),
.B2(n_3156),
.Y(n_3347)
);

AND2x2_ASAP7_75t_L g3348 ( 
.A(n_3250),
.B(n_3219),
.Y(n_3348)
);

NAND2xp5_ASAP7_75t_SL g3349 ( 
.A(n_3298),
.B(n_2863),
.Y(n_3349)
);

INVx3_ASAP7_75t_L g3350 ( 
.A(n_3305),
.Y(n_3350)
);

AOI32xp33_ASAP7_75t_L g3351 ( 
.A1(n_3265),
.A2(n_3120),
.A3(n_3126),
.B1(n_2899),
.B2(n_2859),
.Y(n_3351)
);

INVx1_ASAP7_75t_L g3352 ( 
.A(n_3262),
.Y(n_3352)
);

INVxp67_ASAP7_75t_SL g3353 ( 
.A(n_3251),
.Y(n_3353)
);

NAND2xp5_ASAP7_75t_L g3354 ( 
.A(n_3276),
.B(n_3168),
.Y(n_3354)
);

AOI211xp5_ASAP7_75t_L g3355 ( 
.A1(n_3281),
.A2(n_2796),
.B(n_2805),
.C(n_2994),
.Y(n_3355)
);

NAND2xp5_ASAP7_75t_L g3356 ( 
.A(n_3284),
.B(n_3168),
.Y(n_3356)
);

CKINVDCx16_ASAP7_75t_R g3357 ( 
.A(n_3265),
.Y(n_3357)
);

INVx1_ASAP7_75t_L g3358 ( 
.A(n_3264),
.Y(n_3358)
);

INVx1_ASAP7_75t_L g3359 ( 
.A(n_3267),
.Y(n_3359)
);

AOI22xp5_ASAP7_75t_L g3360 ( 
.A1(n_3281),
.A2(n_3229),
.B1(n_2977),
.B2(n_3096),
.Y(n_3360)
);

AND2x2_ASAP7_75t_L g3361 ( 
.A(n_3249),
.B(n_3231),
.Y(n_3361)
);

AND2x2_ASAP7_75t_L g3362 ( 
.A(n_3283),
.B(n_3170),
.Y(n_3362)
);

NAND2xp5_ASAP7_75t_L g3363 ( 
.A(n_3288),
.B(n_3185),
.Y(n_3363)
);

OAI221xp5_ASAP7_75t_L g3364 ( 
.A1(n_3318),
.A2(n_3305),
.B1(n_3290),
.B2(n_3294),
.C(n_3278),
.Y(n_3364)
);

OAI22xp5_ASAP7_75t_L g3365 ( 
.A1(n_3357),
.A2(n_3265),
.B1(n_3283),
.B2(n_3245),
.Y(n_3365)
);

AOI22xp5_ASAP7_75t_L g3366 ( 
.A1(n_3323),
.A2(n_3283),
.B1(n_3303),
.B2(n_3285),
.Y(n_3366)
);

INVx1_ASAP7_75t_L g3367 ( 
.A(n_3337),
.Y(n_3367)
);

OAI21xp5_ASAP7_75t_L g3368 ( 
.A1(n_3323),
.A2(n_3084),
.B(n_2930),
.Y(n_3368)
);

INVx2_ASAP7_75t_SL g3369 ( 
.A(n_3338),
.Y(n_3369)
);

NOR2xp33_ASAP7_75t_SL g3370 ( 
.A(n_3338),
.B(n_2592),
.Y(n_3370)
);

AOI211xp5_ASAP7_75t_L g3371 ( 
.A1(n_3332),
.A2(n_2927),
.B(n_3084),
.C(n_3245),
.Y(n_3371)
);

INVx2_ASAP7_75t_SL g3372 ( 
.A(n_3339),
.Y(n_3372)
);

OAI22xp33_ASAP7_75t_L g3373 ( 
.A1(n_3350),
.A2(n_3303),
.B1(n_3245),
.B2(n_3304),
.Y(n_3373)
);

OAI22xp5_ASAP7_75t_L g3374 ( 
.A1(n_3355),
.A2(n_3303),
.B1(n_3114),
.B2(n_3273),
.Y(n_3374)
);

INVxp67_ASAP7_75t_L g3375 ( 
.A(n_3335),
.Y(n_3375)
);

NAND2xp5_ASAP7_75t_L g3376 ( 
.A(n_3347),
.B(n_3287),
.Y(n_3376)
);

AOI22xp33_ASAP7_75t_L g3377 ( 
.A1(n_3324),
.A2(n_3242),
.B1(n_3234),
.B2(n_3185),
.Y(n_3377)
);

NAND2xp5_ASAP7_75t_L g3378 ( 
.A(n_3315),
.B(n_3271),
.Y(n_3378)
);

HB1xp67_ASAP7_75t_L g3379 ( 
.A(n_3316),
.Y(n_3379)
);

OAI221xp5_ASAP7_75t_L g3380 ( 
.A1(n_3327),
.A2(n_3289),
.B1(n_3295),
.B2(n_3286),
.C(n_3282),
.Y(n_3380)
);

INVx1_ASAP7_75t_L g3381 ( 
.A(n_3353),
.Y(n_3381)
);

OAI21xp33_ASAP7_75t_L g3382 ( 
.A1(n_3334),
.A2(n_3234),
.B(n_3200),
.Y(n_3382)
);

AOI22xp33_ASAP7_75t_L g3383 ( 
.A1(n_3324),
.A2(n_3299),
.B1(n_3097),
.B2(n_3095),
.Y(n_3383)
);

INVx1_ASAP7_75t_L g3384 ( 
.A(n_3308),
.Y(n_3384)
);

AOI21xp5_ASAP7_75t_SL g3385 ( 
.A1(n_3341),
.A2(n_2809),
.B(n_2806),
.Y(n_3385)
);

AOI22xp33_ASAP7_75t_L g3386 ( 
.A1(n_3349),
.A2(n_3260),
.B1(n_3036),
.B2(n_3033),
.Y(n_3386)
);

OR2x2_ASAP7_75t_L g3387 ( 
.A(n_3344),
.B(n_3196),
.Y(n_3387)
);

AOI22xp5_ASAP7_75t_L g3388 ( 
.A1(n_3360),
.A2(n_3300),
.B1(n_3302),
.B2(n_3297),
.Y(n_3388)
);

OAI22xp5_ASAP7_75t_L g3389 ( 
.A1(n_3355),
.A2(n_3256),
.B1(n_3270),
.B2(n_3091),
.Y(n_3389)
);

INVx1_ASAP7_75t_L g3390 ( 
.A(n_3321),
.Y(n_3390)
);

INVx2_ASAP7_75t_L g3391 ( 
.A(n_3343),
.Y(n_3391)
);

OAI21xp33_ASAP7_75t_L g3392 ( 
.A1(n_3326),
.A2(n_3200),
.B(n_3196),
.Y(n_3392)
);

A2O1A1Ixp33_ASAP7_75t_L g3393 ( 
.A1(n_3351),
.A2(n_3280),
.B(n_2834),
.C(n_2886),
.Y(n_3393)
);

AO32x1_ASAP7_75t_L g3394 ( 
.A1(n_3317),
.A2(n_2941),
.A3(n_2961),
.B1(n_3100),
.B2(n_2990),
.Y(n_3394)
);

OAI221xp5_ASAP7_75t_L g3395 ( 
.A1(n_3360),
.A2(n_2895),
.B1(n_2863),
.B2(n_3181),
.C(n_3186),
.Y(n_3395)
);

INVx1_ASAP7_75t_L g3396 ( 
.A(n_3322),
.Y(n_3396)
);

NAND2xp33_ASAP7_75t_L g3397 ( 
.A(n_3350),
.B(n_2921),
.Y(n_3397)
);

OAI211xp5_ASAP7_75t_L g3398 ( 
.A1(n_3336),
.A2(n_2895),
.B(n_2926),
.C(n_3099),
.Y(n_3398)
);

AOI21xp5_ASAP7_75t_L g3399 ( 
.A1(n_3319),
.A2(n_3115),
.B(n_3108),
.Y(n_3399)
);

AOI21xp33_ASAP7_75t_SL g3400 ( 
.A1(n_3320),
.A2(n_3235),
.B(n_2990),
.Y(n_3400)
);

NAND2xp5_ASAP7_75t_SL g3401 ( 
.A(n_3333),
.B(n_3248),
.Y(n_3401)
);

A2O1A1Ixp33_ASAP7_75t_L g3402 ( 
.A1(n_3374),
.A2(n_3326),
.B(n_3330),
.C(n_3362),
.Y(n_3402)
);

AND2x4_ASAP7_75t_L g3403 ( 
.A(n_3369),
.B(n_3372),
.Y(n_3403)
);

NOR2xp33_ASAP7_75t_L g3404 ( 
.A(n_3375),
.B(n_3314),
.Y(n_3404)
);

AOI22xp5_ASAP7_75t_L g3405 ( 
.A1(n_3370),
.A2(n_3354),
.B1(n_3346),
.B2(n_3311),
.Y(n_3405)
);

INVx1_ASAP7_75t_L g3406 ( 
.A(n_3367),
.Y(n_3406)
);

INVx1_ASAP7_75t_L g3407 ( 
.A(n_3381),
.Y(n_3407)
);

AOI211x1_ASAP7_75t_L g3408 ( 
.A1(n_3380),
.A2(n_3313),
.B(n_3356),
.C(n_3328),
.Y(n_3408)
);

OA22x2_ASAP7_75t_L g3409 ( 
.A1(n_3366),
.A2(n_3331),
.B1(n_3342),
.B2(n_3340),
.Y(n_3409)
);

AOI22xp5_ASAP7_75t_L g3410 ( 
.A1(n_3370),
.A2(n_3329),
.B1(n_3352),
.B2(n_3345),
.Y(n_3410)
);

NOR4xp25_ASAP7_75t_SL g3411 ( 
.A(n_3364),
.B(n_3359),
.C(n_3358),
.D(n_2890),
.Y(n_3411)
);

OAI211xp5_ASAP7_75t_L g3412 ( 
.A1(n_3368),
.A2(n_2926),
.B(n_2890),
.C(n_3363),
.Y(n_3412)
);

A2O1A1Ixp33_ASAP7_75t_L g3413 ( 
.A1(n_3383),
.A2(n_3325),
.B(n_3309),
.C(n_3312),
.Y(n_3413)
);

NAND4xp25_ASAP7_75t_SL g3414 ( 
.A(n_3377),
.B(n_3363),
.C(n_3361),
.D(n_3348),
.Y(n_3414)
);

AOI22x1_ASAP7_75t_SL g3415 ( 
.A1(n_3385),
.A2(n_2592),
.B1(n_2877),
.B2(n_2834),
.Y(n_3415)
);

INVx1_ASAP7_75t_L g3416 ( 
.A(n_3384),
.Y(n_3416)
);

AOI21xp5_ASAP7_75t_L g3417 ( 
.A1(n_3394),
.A2(n_3310),
.B(n_3307),
.Y(n_3417)
);

OAI21xp5_ASAP7_75t_L g3418 ( 
.A1(n_3389),
.A2(n_2952),
.B(n_2912),
.Y(n_3418)
);

NOR2xp33_ASAP7_75t_L g3419 ( 
.A(n_3376),
.B(n_3239),
.Y(n_3419)
);

OAI22xp33_ASAP7_75t_SL g3420 ( 
.A1(n_3365),
.A2(n_2886),
.B1(n_2903),
.B2(n_2877),
.Y(n_3420)
);

AOI22x1_ASAP7_75t_L g3421 ( 
.A1(n_3399),
.A2(n_2801),
.B1(n_2991),
.B2(n_2959),
.Y(n_3421)
);

OAI221xp5_ASAP7_75t_L g3422 ( 
.A1(n_3371),
.A2(n_2979),
.B1(n_3119),
.B2(n_3113),
.C(n_3104),
.Y(n_3422)
);

NAND4xp25_ASAP7_75t_L g3423 ( 
.A(n_3386),
.B(n_2979),
.C(n_2887),
.D(n_2892),
.Y(n_3423)
);

INVx1_ASAP7_75t_SL g3424 ( 
.A(n_3401),
.Y(n_3424)
);

NAND2xp5_ASAP7_75t_L g3425 ( 
.A(n_3392),
.B(n_3261),
.Y(n_3425)
);

AND2x2_ASAP7_75t_L g3426 ( 
.A(n_3387),
.B(n_3248),
.Y(n_3426)
);

NOR2xp67_ASAP7_75t_L g3427 ( 
.A(n_3400),
.B(n_3261),
.Y(n_3427)
);

NAND3xp33_ASAP7_75t_L g3428 ( 
.A(n_3395),
.B(n_2952),
.C(n_3147),
.Y(n_3428)
);

OAI22xp33_ASAP7_75t_L g3429 ( 
.A1(n_3373),
.A2(n_3108),
.B1(n_3115),
.B2(n_2808),
.Y(n_3429)
);

NAND2xp33_ASAP7_75t_L g3430 ( 
.A(n_3393),
.B(n_3382),
.Y(n_3430)
);

AOI221x1_ASAP7_75t_L g3431 ( 
.A1(n_3390),
.A2(n_2944),
.B1(n_2794),
.B2(n_3089),
.C(n_3083),
.Y(n_3431)
);

AOI311xp33_ASAP7_75t_L g3432 ( 
.A1(n_3398),
.A2(n_3396),
.A3(n_3378),
.B(n_3070),
.C(n_3394),
.Y(n_3432)
);

INVx1_ASAP7_75t_L g3433 ( 
.A(n_3379),
.Y(n_3433)
);

OAI221xp5_ASAP7_75t_SL g3434 ( 
.A1(n_3388),
.A2(n_2912),
.B1(n_3094),
.B2(n_3063),
.C(n_2920),
.Y(n_3434)
);

OAI31xp33_ASAP7_75t_L g3435 ( 
.A1(n_3394),
.A2(n_3098),
.A3(n_2896),
.B(n_2903),
.Y(n_3435)
);

OAI221xp5_ASAP7_75t_L g3436 ( 
.A1(n_3397),
.A2(n_3103),
.B1(n_3112),
.B2(n_3127),
.C(n_2808),
.Y(n_3436)
);

NAND2xp5_ASAP7_75t_L g3437 ( 
.A(n_3391),
.B(n_3122),
.Y(n_3437)
);

INVx2_ASAP7_75t_L g3438 ( 
.A(n_3369),
.Y(n_3438)
);

AOI221xp5_ASAP7_75t_L g3439 ( 
.A1(n_3377),
.A2(n_3098),
.B1(n_3144),
.B2(n_3128),
.C(n_3131),
.Y(n_3439)
);

INVx1_ASAP7_75t_L g3440 ( 
.A(n_3367),
.Y(n_3440)
);

AOI211xp5_ASAP7_75t_L g3441 ( 
.A1(n_3430),
.A2(n_2921),
.B(n_2969),
.C(n_2968),
.Y(n_3441)
);

AOI221xp5_ASAP7_75t_L g3442 ( 
.A1(n_3408),
.A2(n_3125),
.B1(n_3130),
.B2(n_3132),
.C(n_3103),
.Y(n_3442)
);

AND4x1_ASAP7_75t_L g3443 ( 
.A(n_3432),
.B(n_2346),
.C(n_2999),
.D(n_2993),
.Y(n_3443)
);

AOI222xp33_ASAP7_75t_L g3444 ( 
.A1(n_3404),
.A2(n_3112),
.B1(n_3052),
.B2(n_3127),
.C1(n_3092),
.C2(n_2856),
.Y(n_3444)
);

NOR3xp33_ASAP7_75t_L g3445 ( 
.A(n_3422),
.B(n_2944),
.C(n_2305),
.Y(n_3445)
);

NOR2xp33_ASAP7_75t_L g3446 ( 
.A(n_3415),
.B(n_3060),
.Y(n_3446)
);

AOI211x1_ASAP7_75t_L g3447 ( 
.A1(n_3414),
.A2(n_2856),
.B(n_3092),
.C(n_2901),
.Y(n_3447)
);

NOR2xp33_ASAP7_75t_L g3448 ( 
.A(n_3403),
.B(n_3221),
.Y(n_3448)
);

AOI221xp5_ASAP7_75t_L g3449 ( 
.A1(n_3402),
.A2(n_3036),
.B1(n_3141),
.B2(n_3129),
.C(n_3133),
.Y(n_3449)
);

NAND2xp5_ASAP7_75t_SL g3450 ( 
.A(n_3420),
.B(n_3435),
.Y(n_3450)
);

NOR3x1_ASAP7_75t_L g3451 ( 
.A(n_3412),
.B(n_2940),
.C(n_2920),
.Y(n_3451)
);

NAND2xp5_ASAP7_75t_L g3452 ( 
.A(n_3419),
.B(n_3151),
.Y(n_3452)
);

OAI221xp5_ASAP7_75t_L g3453 ( 
.A1(n_3405),
.A2(n_2939),
.B1(n_2991),
.B2(n_2959),
.C(n_2940),
.Y(n_3453)
);

AOI221xp5_ASAP7_75t_SL g3454 ( 
.A1(n_3429),
.A2(n_2901),
.B1(n_3133),
.B2(n_3129),
.C(n_3141),
.Y(n_3454)
);

NOR4xp25_ASAP7_75t_L g3455 ( 
.A(n_3406),
.B(n_3440),
.C(n_3407),
.D(n_3433),
.Y(n_3455)
);

OAI21xp5_ASAP7_75t_L g3456 ( 
.A1(n_3427),
.A2(n_2984),
.B(n_2939),
.Y(n_3456)
);

AOI31xp33_ASAP7_75t_L g3457 ( 
.A1(n_3403),
.A2(n_2984),
.A3(n_2857),
.B(n_2802),
.Y(n_3457)
);

INVx3_ASAP7_75t_L g3458 ( 
.A(n_3438),
.Y(n_3458)
);

NAND2xp5_ASAP7_75t_L g3459 ( 
.A(n_3439),
.B(n_3153),
.Y(n_3459)
);

XOR2x2_ASAP7_75t_L g3460 ( 
.A(n_3409),
.B(n_2802),
.Y(n_3460)
);

NOR4xp25_ASAP7_75t_L g3461 ( 
.A(n_3424),
.B(n_2962),
.C(n_2974),
.D(n_3004),
.Y(n_3461)
);

INVx1_ASAP7_75t_L g3462 ( 
.A(n_3416),
.Y(n_3462)
);

NAND2xp5_ASAP7_75t_L g3463 ( 
.A(n_3413),
.B(n_3149),
.Y(n_3463)
);

NAND4xp25_ASAP7_75t_L g3464 ( 
.A(n_3418),
.B(n_2966),
.C(n_2888),
.D(n_2948),
.Y(n_3464)
);

NAND3xp33_ASAP7_75t_L g3465 ( 
.A(n_3411),
.B(n_2240),
.C(n_2949),
.Y(n_3465)
);

NAND2xp5_ASAP7_75t_L g3466 ( 
.A(n_3428),
.B(n_3143),
.Y(n_3466)
);

AOI211xp5_ASAP7_75t_L g3467 ( 
.A1(n_3420),
.A2(n_2888),
.B(n_2841),
.C(n_2953),
.Y(n_3467)
);

AND2x2_ASAP7_75t_L g3468 ( 
.A(n_3410),
.B(n_3221),
.Y(n_3468)
);

INVxp67_ASAP7_75t_L g3469 ( 
.A(n_3458),
.Y(n_3469)
);

NAND2xp5_ASAP7_75t_L g3470 ( 
.A(n_3455),
.B(n_3425),
.Y(n_3470)
);

NOR2xp33_ASAP7_75t_L g3471 ( 
.A(n_3458),
.B(n_3423),
.Y(n_3471)
);

NOR3xp33_ASAP7_75t_SL g3472 ( 
.A(n_3450),
.B(n_3434),
.C(n_3436),
.Y(n_3472)
);

OAI31xp33_ASAP7_75t_L g3473 ( 
.A1(n_3446),
.A2(n_3417),
.A3(n_3426),
.B(n_3421),
.Y(n_3473)
);

INVx2_ASAP7_75t_L g3474 ( 
.A(n_3462),
.Y(n_3474)
);

INVx1_ASAP7_75t_L g3475 ( 
.A(n_3466),
.Y(n_3475)
);

BUFx2_ASAP7_75t_L g3476 ( 
.A(n_3468),
.Y(n_3476)
);

INVx1_ASAP7_75t_L g3477 ( 
.A(n_3459),
.Y(n_3477)
);

NAND2xp5_ASAP7_75t_L g3478 ( 
.A(n_3442),
.B(n_3437),
.Y(n_3478)
);

NOR3xp33_ASAP7_75t_L g3479 ( 
.A(n_3445),
.B(n_2229),
.C(n_2219),
.Y(n_3479)
);

INVx2_ASAP7_75t_L g3480 ( 
.A(n_3448),
.Y(n_3480)
);

OAI322xp33_ASAP7_75t_L g3481 ( 
.A1(n_3463),
.A2(n_3453),
.A3(n_3465),
.B1(n_3451),
.B2(n_3443),
.C1(n_3447),
.C2(n_3452),
.Y(n_3481)
);

INVx2_ASAP7_75t_SL g3482 ( 
.A(n_3460),
.Y(n_3482)
);

INVx1_ASAP7_75t_L g3483 ( 
.A(n_3461),
.Y(n_3483)
);

NOR3xp33_ASAP7_75t_L g3484 ( 
.A(n_3464),
.B(n_2229),
.C(n_2219),
.Y(n_3484)
);

NOR2xp33_ASAP7_75t_SL g3485 ( 
.A(n_3456),
.B(n_3431),
.Y(n_3485)
);

OA22x2_ASAP7_75t_L g3486 ( 
.A1(n_3441),
.A2(n_2469),
.B1(n_2966),
.B2(n_2996),
.Y(n_3486)
);

HB1xp67_ASAP7_75t_L g3487 ( 
.A(n_3454),
.Y(n_3487)
);

INVx1_ASAP7_75t_L g3488 ( 
.A(n_3444),
.Y(n_3488)
);

INVx1_ASAP7_75t_L g3489 ( 
.A(n_3457),
.Y(n_3489)
);

AOI211x1_ASAP7_75t_L g3490 ( 
.A1(n_3449),
.A2(n_3146),
.B(n_3143),
.C(n_2998),
.Y(n_3490)
);

NOR2xp67_ASAP7_75t_L g3491 ( 
.A(n_3467),
.B(n_3146),
.Y(n_3491)
);

NAND3xp33_ASAP7_75t_L g3492 ( 
.A(n_3469),
.B(n_3472),
.C(n_3473),
.Y(n_3492)
);

NAND4xp25_ASAP7_75t_L g3493 ( 
.A(n_3488),
.B(n_2988),
.C(n_3002),
.D(n_3001),
.Y(n_3493)
);

AO22x2_ASAP7_75t_L g3494 ( 
.A1(n_3483),
.A2(n_2989),
.B1(n_2972),
.B2(n_2967),
.Y(n_3494)
);

OR2x2_ASAP7_75t_L g3495 ( 
.A(n_3487),
.B(n_3076),
.Y(n_3495)
);

NAND3xp33_ASAP7_75t_SL g3496 ( 
.A(n_3470),
.B(n_2874),
.C(n_2873),
.Y(n_3496)
);

NOR4xp25_ASAP7_75t_L g3497 ( 
.A(n_3477),
.B(n_2719),
.C(n_2727),
.D(n_2718),
.Y(n_3497)
);

HB1xp67_ASAP7_75t_L g3498 ( 
.A(n_3474),
.Y(n_3498)
);

NOR2x1p5_ASAP7_75t_L g3499 ( 
.A(n_3480),
.B(n_3489),
.Y(n_3499)
);

NOR2x1_ASAP7_75t_L g3500 ( 
.A(n_3481),
.B(n_2240),
.Y(n_3500)
);

NAND2x1p5_ASAP7_75t_L g3501 ( 
.A(n_3476),
.B(n_3107),
.Y(n_3501)
);

NAND2xp5_ASAP7_75t_L g3502 ( 
.A(n_3475),
.B(n_3022),
.Y(n_3502)
);

AOI22xp5_ASAP7_75t_L g3503 ( 
.A1(n_3471),
.A2(n_2469),
.B1(n_2982),
.B2(n_2989),
.Y(n_3503)
);

NOR2xp67_ASAP7_75t_L g3504 ( 
.A(n_3482),
.B(n_3478),
.Y(n_3504)
);

INVx1_ASAP7_75t_L g3505 ( 
.A(n_3478),
.Y(n_3505)
);

NAND4xp75_ASAP7_75t_L g3506 ( 
.A(n_3490),
.B(n_2431),
.C(n_2413),
.D(n_2698),
.Y(n_3506)
);

NOR2x1_ASAP7_75t_L g3507 ( 
.A(n_3491),
.B(n_3485),
.Y(n_3507)
);

INVxp67_ASAP7_75t_L g3508 ( 
.A(n_3485),
.Y(n_3508)
);

NAND4xp75_ASAP7_75t_L g3509 ( 
.A(n_3486),
.B(n_3479),
.C(n_3484),
.D(n_2431),
.Y(n_3509)
);

OR2x2_ASAP7_75t_L g3510 ( 
.A(n_3486),
.B(n_2845),
.Y(n_3510)
);

AOI211x1_ASAP7_75t_L g3511 ( 
.A1(n_3470),
.A2(n_2698),
.B(n_2730),
.C(n_2542),
.Y(n_3511)
);

NOR2x1_ASAP7_75t_L g3512 ( 
.A(n_3492),
.B(n_2491),
.Y(n_3512)
);

INVx1_ASAP7_75t_L g3513 ( 
.A(n_3498),
.Y(n_3513)
);

NOR2xp33_ASAP7_75t_L g3514 ( 
.A(n_3508),
.B(n_3221),
.Y(n_3514)
);

NOR3xp33_ASAP7_75t_L g3515 ( 
.A(n_3505),
.B(n_2416),
.C(n_2215),
.Y(n_3515)
);

NOR2x1_ASAP7_75t_L g3516 ( 
.A(n_3499),
.B(n_2469),
.Y(n_3516)
);

AOI21xp5_ASAP7_75t_L g3517 ( 
.A1(n_3504),
.A2(n_2487),
.B(n_2479),
.Y(n_3517)
);

INVx1_ASAP7_75t_L g3518 ( 
.A(n_3495),
.Y(n_3518)
);

INVx1_ASAP7_75t_L g3519 ( 
.A(n_3502),
.Y(n_3519)
);

NOR2x1_ASAP7_75t_L g3520 ( 
.A(n_3509),
.B(n_2310),
.Y(n_3520)
);

OR2x2_ASAP7_75t_L g3521 ( 
.A(n_3493),
.B(n_2845),
.Y(n_3521)
);

INVx1_ASAP7_75t_L g3522 ( 
.A(n_3494),
.Y(n_3522)
);

NOR3xp33_ASAP7_75t_L g3523 ( 
.A(n_3500),
.B(n_2416),
.C(n_2487),
.Y(n_3523)
);

XNOR2xp5_ASAP7_75t_L g3524 ( 
.A(n_3503),
.B(n_2967),
.Y(n_3524)
);

OA22x2_ASAP7_75t_L g3525 ( 
.A1(n_3513),
.A2(n_3507),
.B1(n_3494),
.B2(n_3501),
.Y(n_3525)
);

OR2x2_ASAP7_75t_L g3526 ( 
.A(n_3518),
.B(n_3496),
.Y(n_3526)
);

OR2x6_ASAP7_75t_L g3527 ( 
.A(n_3514),
.B(n_3511),
.Y(n_3527)
);

INVx2_ASAP7_75t_SL g3528 ( 
.A(n_3516),
.Y(n_3528)
);

NAND2x1p5_ASAP7_75t_L g3529 ( 
.A(n_3520),
.B(n_3519),
.Y(n_3529)
);

INVx1_ASAP7_75t_L g3530 ( 
.A(n_3522),
.Y(n_3530)
);

AND2x4_ASAP7_75t_L g3531 ( 
.A(n_3512),
.B(n_3510),
.Y(n_3531)
);

INVx1_ASAP7_75t_L g3532 ( 
.A(n_3521),
.Y(n_3532)
);

NOR2x1_ASAP7_75t_L g3533 ( 
.A(n_3524),
.B(n_3506),
.Y(n_3533)
);

XNOR2xp5_ASAP7_75t_L g3534 ( 
.A(n_3523),
.B(n_3497),
.Y(n_3534)
);

INVxp67_ASAP7_75t_L g3535 ( 
.A(n_3530),
.Y(n_3535)
);

OAI21xp5_ASAP7_75t_L g3536 ( 
.A1(n_3529),
.A2(n_3517),
.B(n_3515),
.Y(n_3536)
);

INVx1_ASAP7_75t_L g3537 ( 
.A(n_3526),
.Y(n_3537)
);

OAI211xp5_ASAP7_75t_L g3538 ( 
.A1(n_3532),
.A2(n_2352),
.B(n_2363),
.C(n_2357),
.Y(n_3538)
);

XNOR2xp5_ASAP7_75t_L g3539 ( 
.A(n_3525),
.B(n_2479),
.Y(n_3539)
);

NAND3xp33_ASAP7_75t_L g3540 ( 
.A(n_3535),
.B(n_3533),
.C(n_3527),
.Y(n_3540)
);

OAI21x1_ASAP7_75t_L g3541 ( 
.A1(n_3537),
.A2(n_3534),
.B(n_3528),
.Y(n_3541)
);

INVx2_ASAP7_75t_L g3542 ( 
.A(n_3539),
.Y(n_3542)
);

INVx3_ASAP7_75t_L g3543 ( 
.A(n_3538),
.Y(n_3543)
);

INVx1_ASAP7_75t_L g3544 ( 
.A(n_3536),
.Y(n_3544)
);

INVx1_ASAP7_75t_L g3545 ( 
.A(n_3544),
.Y(n_3545)
);

AOI22xp5_ASAP7_75t_SL g3546 ( 
.A1(n_3543),
.A2(n_3531),
.B1(n_3107),
.B2(n_2352),
.Y(n_3546)
);

INVx1_ASAP7_75t_L g3547 ( 
.A(n_3541),
.Y(n_3547)
);

INVxp33_ASAP7_75t_L g3548 ( 
.A(n_3540),
.Y(n_3548)
);

OAI21xp5_ASAP7_75t_L g3549 ( 
.A1(n_3548),
.A2(n_3540),
.B(n_3542),
.Y(n_3549)
);

INVx1_ASAP7_75t_L g3550 ( 
.A(n_3545),
.Y(n_3550)
);

NAND2xp33_ASAP7_75t_SL g3551 ( 
.A(n_3550),
.B(n_3543),
.Y(n_3551)
);

NAND2xp5_ASAP7_75t_SL g3552 ( 
.A(n_3551),
.B(n_3547),
.Y(n_3552)
);

OAI21xp5_ASAP7_75t_L g3553 ( 
.A1(n_3551),
.A2(n_3549),
.B(n_3546),
.Y(n_3553)
);

HB1xp67_ASAP7_75t_L g3554 ( 
.A(n_3553),
.Y(n_3554)
);

AOI22xp5_ASAP7_75t_L g3555 ( 
.A1(n_3554),
.A2(n_3552),
.B1(n_3107),
.B2(n_2982),
.Y(n_3555)
);


endmodule