module fake_jpeg_31756_n_364 (n_13, n_11, n_14, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_364);

input n_13;
input n_11;
input n_14;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_364;

wire n_253;
wire n_330;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_228;
wire n_134;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_340;
wire n_291;
wire n_236;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_148;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_17;
wire n_102;
wire n_196;
wire n_66;
wire n_142;
wire n_362;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_256;
wire n_221;
wire n_213;
wire n_292;
wire n_135;
wire n_189;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_225;
wire n_105;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_124;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_80;
wire n_204;
wire n_306;
wire n_298;
wire n_106;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_85;
wire n_163;
wire n_136;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_39;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_91;
wire n_305;
wire n_161;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_303;
wire n_259;
wire n_90;
wire n_344;
wire n_328;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_262;
wire n_240;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_275;
wire n_169;
wire n_153;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_114;
wire n_281;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_356;
wire n_119;
wire n_83;
wire n_125;
wire n_81;
wire n_224;
wire n_113;
wire n_248;
wire n_30;
wire n_307;
wire n_111;
wire n_197;
wire n_186;
wire n_202;
wire n_25;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_215;
wire n_212;
wire n_183;
wire n_249;
wire n_217;
wire n_53;
wire n_33;
wire n_54;
wire n_209;
wire n_22;
wire n_138;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

CKINVDCx20_ASAP7_75t_R g17 ( 
.A(n_14),
.Y(n_17)
);

INVx1_ASAP7_75t_L g18 ( 
.A(n_16),
.Y(n_18)
);

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_1),
.Y(n_19)
);

BUFx6f_ASAP7_75t_L g20 ( 
.A(n_5),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_2),
.Y(n_23)
);

BUFx16f_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx2_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

BUFx5_ASAP7_75t_L g26 ( 
.A(n_10),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_13),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_3),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_8),
.Y(n_29)
);

INVx1_ASAP7_75t_L g30 ( 
.A(n_1),
.Y(n_30)
);

CKINVDCx16_ASAP7_75t_R g31 ( 
.A(n_13),
.Y(n_31)
);

BUFx3_ASAP7_75t_L g32 ( 
.A(n_15),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_11),
.Y(n_33)
);

CKINVDCx20_ASAP7_75t_R g34 ( 
.A(n_16),
.Y(n_34)
);

INVx11_ASAP7_75t_L g35 ( 
.A(n_0),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_6),
.Y(n_36)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_14),
.Y(n_37)
);

CKINVDCx20_ASAP7_75t_R g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_8),
.Y(n_39)
);

INVx3_ASAP7_75t_L g40 ( 
.A(n_12),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx2_ASAP7_75t_L g42 ( 
.A(n_10),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_12),
.Y(n_43)
);

INVx6_ASAP7_75t_L g44 ( 
.A(n_19),
.Y(n_44)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_44),
.Y(n_95)
);

NOR2xp33_ASAP7_75t_L g45 ( 
.A(n_17),
.B(n_15),
.Y(n_45)
);

AND2x2_ASAP7_75t_L g100 ( 
.A(n_45),
.B(n_51),
.Y(n_100)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_25),
.Y(n_46)
);

INVx2_ASAP7_75t_L g89 ( 
.A(n_46),
.Y(n_89)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_25),
.Y(n_47)
);

INVx2_ASAP7_75t_L g93 ( 
.A(n_47),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_19),
.Y(n_48)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_48),
.Y(n_102)
);

AOI22xp33_ASAP7_75t_L g49 ( 
.A1(n_42),
.A2(n_0),
.B1(n_1),
.B2(n_2),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_49),
.A2(n_31),
.B1(n_23),
.B2(n_36),
.Y(n_83)
);

INVx13_ASAP7_75t_L g50 ( 
.A(n_24),
.Y(n_50)
);

INVx5_ASAP7_75t_L g109 ( 
.A(n_50),
.Y(n_109)
);

AND2x2_ASAP7_75t_L g51 ( 
.A(n_42),
.B(n_15),
.Y(n_51)
);

INVx6_ASAP7_75t_L g52 ( 
.A(n_19),
.Y(n_52)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_52),
.Y(n_103)
);

INVx5_ASAP7_75t_L g53 ( 
.A(n_26),
.Y(n_53)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_53),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g54 ( 
.A(n_19),
.Y(n_54)
);

INVx6_ASAP7_75t_L g81 ( 
.A(n_54),
.Y(n_81)
);

NOR2xp33_ASAP7_75t_L g55 ( 
.A(n_17),
.B(n_14),
.Y(n_55)
);

NOR2xp33_ASAP7_75t_L g85 ( 
.A(n_55),
.B(n_60),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_20),
.Y(n_56)
);

INVx6_ASAP7_75t_L g84 ( 
.A(n_56),
.Y(n_84)
);

BUFx12f_ASAP7_75t_L g57 ( 
.A(n_24),
.Y(n_57)
);

INVx3_ASAP7_75t_L g86 ( 
.A(n_57),
.Y(n_86)
);

BUFx6f_ASAP7_75t_L g58 ( 
.A(n_20),
.Y(n_58)
);

INVx6_ASAP7_75t_L g120 ( 
.A(n_58),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_24),
.Y(n_59)
);

INVx3_ASAP7_75t_L g105 ( 
.A(n_59),
.Y(n_105)
);

NOR2xp33_ASAP7_75t_L g60 ( 
.A(n_21),
.B(n_13),
.Y(n_60)
);

BUFx3_ASAP7_75t_L g61 ( 
.A(n_35),
.Y(n_61)
);

INVx4_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx5_ASAP7_75t_L g62 ( 
.A(n_26),
.Y(n_62)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_62),
.Y(n_118)
);

INVx8_ASAP7_75t_L g63 ( 
.A(n_26),
.Y(n_63)
);

INVx8_ASAP7_75t_L g94 ( 
.A(n_63),
.Y(n_94)
);

BUFx6f_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx8_ASAP7_75t_L g122 ( 
.A(n_64),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_20),
.Y(n_65)
);

INVx2_ASAP7_75t_L g99 ( 
.A(n_65),
.Y(n_99)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_40),
.Y(n_66)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_66),
.Y(n_107)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_21),
.B(n_12),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g87 ( 
.A(n_67),
.B(n_34),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx3_ASAP7_75t_L g119 ( 
.A(n_68),
.Y(n_119)
);

NOR2xp33_ASAP7_75t_L g69 ( 
.A(n_33),
.B(n_11),
.Y(n_69)
);

NOR2xp33_ASAP7_75t_L g90 ( 
.A(n_69),
.B(n_72),
.Y(n_90)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

INVx2_ASAP7_75t_SL g104 ( 
.A(n_70),
.Y(n_104)
);

INVx8_ASAP7_75t_L g71 ( 
.A(n_28),
.Y(n_71)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_71),
.Y(n_108)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_28),
.Y(n_72)
);

BUFx6f_ASAP7_75t_L g73 ( 
.A(n_28),
.Y(n_73)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_73),
.Y(n_113)
);

NOR2xp33_ASAP7_75t_L g74 ( 
.A(n_33),
.B(n_10),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_74),
.B(n_31),
.Y(n_98)
);

HB1xp67_ASAP7_75t_L g75 ( 
.A(n_40),
.Y(n_75)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_75),
.Y(n_88)
);

CKINVDCx20_ASAP7_75t_R g76 ( 
.A(n_61),
.Y(n_76)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_98),
.Y(n_130)
);

OAI22xp33_ASAP7_75t_SL g77 ( 
.A1(n_44),
.A2(n_43),
.B1(n_37),
.B2(n_39),
.Y(n_77)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_77),
.A2(n_101),
.B1(n_73),
.B2(n_65),
.Y(n_134)
);

NOR2x1_ASAP7_75t_L g78 ( 
.A(n_51),
.B(n_38),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_SL g159 ( 
.A(n_78),
.B(n_82),
.Y(n_159)
);

AOI22xp33_ASAP7_75t_SL g80 ( 
.A1(n_71),
.A2(n_40),
.B1(n_32),
.B2(n_39),
.Y(n_80)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_80),
.A2(n_115),
.B1(n_70),
.B2(n_41),
.Y(n_147)
);

NAND2xp5_ASAP7_75t_SL g82 ( 
.A(n_53),
.B(n_38),
.Y(n_82)
);

OA22x2_ASAP7_75t_L g126 ( 
.A1(n_83),
.A2(n_91),
.B1(n_43),
.B2(n_37),
.Y(n_126)
);

AND2x2_ASAP7_75t_L g125 ( 
.A(n_87),
.B(n_85),
.Y(n_125)
);

OA22x2_ASAP7_75t_L g91 ( 
.A1(n_49),
.A2(n_22),
.B1(n_30),
.B2(n_36),
.Y(n_91)
);

HB1xp67_ASAP7_75t_L g92 ( 
.A(n_68),
.Y(n_92)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_92),
.Y(n_124)
);

NAND2xp5_ASAP7_75t_L g96 ( 
.A(n_52),
.B(n_34),
.Y(n_96)
);

NAND2xp5_ASAP7_75t_L g155 ( 
.A(n_96),
.B(n_110),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g97 ( 
.A(n_62),
.B(n_27),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_97),
.B(n_109),
.Y(n_140)
);

OAI22xp33_ASAP7_75t_SL g101 ( 
.A1(n_48),
.A2(n_43),
.B1(n_37),
.B2(n_39),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g106 ( 
.A(n_57),
.B(n_27),
.Y(n_106)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_106),
.B(n_59),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_L g110 ( 
.A(n_54),
.B(n_23),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_SL g112 ( 
.A1(n_63),
.A2(n_18),
.B1(n_30),
.B2(n_22),
.Y(n_112)
);

OR2x2_ASAP7_75t_L g132 ( 
.A(n_112),
.B(n_114),
.Y(n_132)
);

OR2x2_ASAP7_75t_L g114 ( 
.A(n_50),
.B(n_18),
.Y(n_114)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_32),
.B1(n_41),
.B2(n_39),
.Y(n_115)
);

NOR2xp33_ASAP7_75t_SL g116 ( 
.A(n_57),
.B(n_9),
.Y(n_116)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_116),
.B(n_3),
.Y(n_164)
);

INVx2_ASAP7_75t_L g117 ( 
.A(n_56),
.Y(n_117)
);

INVx2_ASAP7_75t_L g157 ( 
.A(n_117),
.Y(n_157)
);

AND2x2_ASAP7_75t_SL g121 ( 
.A(n_58),
.B(n_41),
.Y(n_121)
);

XNOR2xp5_ASAP7_75t_L g128 ( 
.A(n_121),
.B(n_72),
.Y(n_128)
);

CKINVDCx20_ASAP7_75t_R g123 ( 
.A(n_114),
.Y(n_123)
);

NOR2xp33_ASAP7_75t_L g165 ( 
.A(n_123),
.B(n_135),
.Y(n_165)
);

NOR3xp33_ASAP7_75t_SL g185 ( 
.A(n_125),
.B(n_79),
.C(n_105),
.Y(n_185)
);

AOI22xp5_ASAP7_75t_L g169 ( 
.A1(n_126),
.A2(n_131),
.B1(n_134),
.B2(n_148),
.Y(n_169)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_102),
.Y(n_127)
);

INVx3_ASAP7_75t_L g192 ( 
.A(n_127),
.Y(n_192)
);

XNOR2xp5_ASAP7_75t_L g183 ( 
.A(n_128),
.B(n_94),
.Y(n_183)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_109),
.Y(n_129)
);

INVx2_ASAP7_75t_L g170 ( 
.A(n_129),
.Y(n_170)
);

OAI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_91),
.A2(n_78),
.B1(n_112),
.B2(n_95),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g133 ( 
.A(n_102),
.Y(n_133)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_133),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g136 ( 
.A(n_90),
.B(n_32),
.Y(n_136)
);

NOR2xp33_ASAP7_75t_L g178 ( 
.A(n_136),
.B(n_137),
.Y(n_178)
);

NOR2xp33_ASAP7_75t_L g137 ( 
.A(n_100),
.B(n_88),
.Y(n_137)
);

BUFx2_ASAP7_75t_L g138 ( 
.A(n_122),
.Y(n_138)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_138),
.Y(n_181)
);

AOI22xp33_ASAP7_75t_L g139 ( 
.A1(n_91),
.A2(n_64),
.B1(n_43),
.B2(n_37),
.Y(n_139)
);

OAI22xp5_ASAP7_75t_SL g171 ( 
.A1(n_139),
.A2(n_146),
.B1(n_158),
.B2(n_84),
.Y(n_171)
);

NOR2xp33_ASAP7_75t_L g191 ( 
.A(n_140),
.B(n_152),
.Y(n_191)
);

AND2x4_ASAP7_75t_L g141 ( 
.A(n_121),
.B(n_59),
.Y(n_141)
);

AND2x4_ASAP7_75t_SL g166 ( 
.A(n_141),
.B(n_118),
.Y(n_166)
);

INVx1_ASAP7_75t_L g142 ( 
.A(n_89),
.Y(n_142)
);

INVx1_ASAP7_75t_L g179 ( 
.A(n_142),
.Y(n_179)
);

INVx1_ASAP7_75t_L g143 ( 
.A(n_93),
.Y(n_143)
);

INVx1_ASAP7_75t_L g188 ( 
.A(n_143),
.Y(n_188)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_107),
.Y(n_144)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_144),
.Y(n_193)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_99),
.Y(n_145)
);

INVx1_ASAP7_75t_L g197 ( 
.A(n_145),
.Y(n_197)
);

AOI22xp33_ASAP7_75t_L g146 ( 
.A1(n_101),
.A2(n_41),
.B1(n_29),
.B2(n_72),
.Y(n_146)
);

OA22x2_ASAP7_75t_L g196 ( 
.A1(n_147),
.A2(n_4),
.B1(n_5),
.B2(n_6),
.Y(n_196)
);

OAI22xp5_ASAP7_75t_L g148 ( 
.A1(n_121),
.A2(n_29),
.B1(n_35),
.B2(n_9),
.Y(n_148)
);

INVx8_ASAP7_75t_L g149 ( 
.A(n_94),
.Y(n_149)
);

INVx1_ASAP7_75t_L g201 ( 
.A(n_149),
.Y(n_201)
);

OAI22xp5_ASAP7_75t_L g150 ( 
.A1(n_80),
.A2(n_29),
.B1(n_35),
.B2(n_9),
.Y(n_150)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_150),
.A2(n_103),
.B1(n_119),
.B2(n_86),
.Y(n_187)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_113),
.Y(n_151)
);

CKINVDCx16_ASAP7_75t_R g167 ( 
.A(n_151),
.Y(n_167)
);

CKINVDCx14_ASAP7_75t_R g152 ( 
.A(n_100),
.Y(n_152)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_111),
.Y(n_153)
);

NOR2xp33_ASAP7_75t_L g195 ( 
.A(n_153),
.B(n_154),
.Y(n_195)
);

CKINVDCx20_ASAP7_75t_R g154 ( 
.A(n_115),
.Y(n_154)
);

INVx1_ASAP7_75t_L g156 ( 
.A(n_108),
.Y(n_156)
);

CKINVDCx16_ASAP7_75t_R g176 ( 
.A(n_156),
.Y(n_176)
);

AOI22xp33_ASAP7_75t_L g158 ( 
.A1(n_77),
.A2(n_29),
.B1(n_1),
.B2(n_2),
.Y(n_158)
);

INVx1_ASAP7_75t_L g160 ( 
.A(n_95),
.Y(n_160)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_160),
.Y(n_184)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_118),
.B(n_0),
.Y(n_161)
);

NOR2xp33_ASAP7_75t_L g198 ( 
.A(n_161),
.B(n_162),
.Y(n_198)
);

CKINVDCx16_ASAP7_75t_R g162 ( 
.A(n_104),
.Y(n_162)
);

A2O1A1Ixp33_ASAP7_75t_L g163 ( 
.A1(n_104),
.A2(n_0),
.B(n_2),
.C(n_3),
.Y(n_163)
);

NOR3xp33_ASAP7_75t_L g177 ( 
.A(n_163),
.B(n_119),
.C(n_86),
.Y(n_177)
);

NOR2xp33_ASAP7_75t_L g200 ( 
.A(n_164),
.B(n_6),
.Y(n_200)
);

OAI21xp5_ASAP7_75t_L g211 ( 
.A1(n_166),
.A2(n_141),
.B(n_149),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_L g168 ( 
.A1(n_154),
.A2(n_84),
.B1(n_120),
.B2(n_81),
.Y(n_168)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_168),
.A2(n_171),
.B1(n_182),
.B2(n_199),
.Y(n_210)
);

CKINVDCx20_ASAP7_75t_R g173 ( 
.A(n_138),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g204 ( 
.A(n_173),
.B(n_200),
.Y(n_204)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_155),
.B(n_120),
.Y(n_174)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_174),
.B(n_175),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g175 ( 
.A(n_155),
.B(n_81),
.Y(n_175)
);

INVxp67_ASAP7_75t_L g232 ( 
.A(n_177),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g180 ( 
.A(n_128),
.B(n_79),
.C(n_105),
.Y(n_180)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_180),
.B(n_183),
.C(n_145),
.Y(n_234)
);

OAI22xp5_ASAP7_75t_SL g182 ( 
.A1(n_132),
.A2(n_103),
.B1(n_122),
.B2(n_111),
.Y(n_182)
);

NOR2xp33_ASAP7_75t_SL g214 ( 
.A(n_185),
.B(n_202),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g186 ( 
.A(n_132),
.B(n_140),
.Y(n_186)
);

NAND2xp5_ASAP7_75t_L g228 ( 
.A(n_186),
.B(n_190),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_L g212 ( 
.A1(n_187),
.A2(n_189),
.B1(n_196),
.B2(n_163),
.Y(n_212)
);

AOI22xp5_ASAP7_75t_L g189 ( 
.A1(n_134),
.A2(n_3),
.B1(n_4),
.B2(n_5),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_132),
.B(n_8),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g194 ( 
.A(n_141),
.B(n_8),
.Y(n_194)
);

NAND2xp5_ASAP7_75t_SL g216 ( 
.A(n_194),
.B(n_141),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_L g199 ( 
.A1(n_126),
.A2(n_7),
.B1(n_5),
.B2(n_6),
.Y(n_199)
);

NOR2xp33_ASAP7_75t_SL g202 ( 
.A(n_123),
.B(n_7),
.Y(n_202)
);

CKINVDCx20_ASAP7_75t_R g203 ( 
.A(n_165),
.Y(n_203)
);

NOR2xp33_ASAP7_75t_L g242 ( 
.A(n_203),
.B(n_209),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_L g205 ( 
.A1(n_199),
.A2(n_150),
.B1(n_126),
.B2(n_148),
.Y(n_205)
);

AOI22xp5_ASAP7_75t_L g264 ( 
.A1(n_205),
.A2(n_212),
.B1(n_229),
.B2(n_127),
.Y(n_264)
);

INVx2_ASAP7_75t_L g206 ( 
.A(n_172),
.Y(n_206)
);

INVx1_ASAP7_75t_L g243 ( 
.A(n_206),
.Y(n_243)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_179),
.Y(n_207)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_207),
.Y(n_250)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_179),
.Y(n_208)
);

INVx1_ASAP7_75t_L g263 ( 
.A(n_208),
.Y(n_263)
);

CKINVDCx20_ASAP7_75t_R g209 ( 
.A(n_174),
.Y(n_209)
);

AND2x2_ASAP7_75t_L g244 ( 
.A(n_211),
.B(n_223),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g213 ( 
.A(n_202),
.B(n_130),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_L g241 ( 
.A(n_213),
.B(n_218),
.Y(n_241)
);

INVx1_ASAP7_75t_L g215 ( 
.A(n_188),
.Y(n_215)
);

CKINVDCx16_ASAP7_75t_R g239 ( 
.A(n_215),
.Y(n_239)
);

XNOR2xp5_ASAP7_75t_SL g254 ( 
.A(n_216),
.B(n_234),
.Y(n_254)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_171),
.A2(n_126),
.B1(n_125),
.B2(n_142),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g247 ( 
.A1(n_217),
.A2(n_235),
.B1(n_176),
.B2(n_184),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_L g218 ( 
.A(n_175),
.B(n_198),
.Y(n_218)
);

NOR2xp33_ASAP7_75t_L g219 ( 
.A(n_186),
.B(n_178),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_219),
.B(n_224),
.Y(n_248)
);

INVx1_ASAP7_75t_L g220 ( 
.A(n_188),
.Y(n_220)
);

NOR2xp33_ASAP7_75t_L g252 ( 
.A(n_220),
.B(n_226),
.Y(n_252)
);

OAI21xp5_ASAP7_75t_L g222 ( 
.A1(n_190),
.A2(n_159),
.B(n_125),
.Y(n_222)
);

OAI21xp5_ASAP7_75t_L g245 ( 
.A1(n_222),
.A2(n_166),
.B(n_189),
.Y(n_245)
);

OA21x2_ASAP7_75t_L g223 ( 
.A1(n_195),
.A2(n_124),
.B(n_156),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_183),
.B(n_143),
.Y(n_224)
);

NOR2xp33_ASAP7_75t_L g225 ( 
.A(n_191),
.B(n_124),
.Y(n_225)
);

NAND2xp5_ASAP7_75t_L g257 ( 
.A(n_225),
.B(n_170),
.Y(n_257)
);

INVx1_ASAP7_75t_L g226 ( 
.A(n_193),
.Y(n_226)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_193),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_227),
.B(n_230),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_169),
.A2(n_160),
.B1(n_144),
.B2(n_133),
.Y(n_229)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_197),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g231 ( 
.A(n_185),
.Y(n_231)
);

NOR2xp33_ASAP7_75t_L g261 ( 
.A(n_231),
.B(n_233),
.Y(n_261)
);

INVxp33_ASAP7_75t_L g233 ( 
.A(n_182),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_L g235 ( 
.A1(n_169),
.A2(n_151),
.B1(n_157),
.B2(n_133),
.Y(n_235)
);

CKINVDCx20_ASAP7_75t_R g236 ( 
.A(n_167),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_236),
.Y(n_237)
);

OAI22x1_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_196),
.B1(n_166),
.B2(n_187),
.Y(n_238)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_238),
.A2(n_247),
.B1(n_229),
.B2(n_209),
.Y(n_268)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_232),
.A2(n_180),
.B(n_194),
.Y(n_240)
);

AOI21xp5_ASAP7_75t_L g273 ( 
.A1(n_240),
.A2(n_255),
.B(n_262),
.Y(n_273)
);

XOR2xp5_ASAP7_75t_L g266 ( 
.A(n_245),
.B(n_211),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g246 ( 
.A(n_228),
.B(n_197),
.Y(n_246)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_246),
.B(n_257),
.Y(n_277)
);

MAJIxp5_ASAP7_75t_L g249 ( 
.A(n_234),
.B(n_166),
.C(n_201),
.Y(n_249)
);

MAJIxp5_ASAP7_75t_L g269 ( 
.A(n_249),
.B(n_265),
.C(n_216),
.Y(n_269)
);

NOR2xp33_ASAP7_75t_SL g251 ( 
.A(n_219),
.B(n_168),
.Y(n_251)
);

NOR2xp33_ASAP7_75t_SL g278 ( 
.A(n_251),
.B(n_253),
.Y(n_278)
);

NOR2xp33_ASAP7_75t_SL g253 ( 
.A(n_213),
.B(n_201),
.Y(n_253)
);

OAI21xp5_ASAP7_75t_SL g255 ( 
.A1(n_212),
.A2(n_196),
.B(n_170),
.Y(n_255)
);

NOR2xp33_ASAP7_75t_SL g256 ( 
.A(n_203),
.B(n_173),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_256),
.B(n_258),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_SL g258 ( 
.A(n_225),
.B(n_196),
.Y(n_258)
);

CKINVDCx20_ASAP7_75t_R g260 ( 
.A(n_204),
.Y(n_260)
);

NOR2xp33_ASAP7_75t_L g270 ( 
.A(n_260),
.B(n_236),
.Y(n_270)
);

OAI21xp5_ASAP7_75t_SL g262 ( 
.A1(n_228),
.A2(n_153),
.B(n_181),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g283 ( 
.A1(n_264),
.A2(n_223),
.B1(n_227),
.B2(n_226),
.Y(n_283)
);

XOR2xp5_ASAP7_75t_L g265 ( 
.A(n_224),
.B(n_162),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_SL g291 ( 
.A(n_266),
.B(n_244),
.Y(n_291)
);

INVx1_ASAP7_75t_L g267 ( 
.A(n_252),
.Y(n_267)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_267),
.Y(n_297)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_268),
.A2(n_276),
.B1(n_245),
.B2(n_261),
.Y(n_293)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_269),
.B(n_271),
.Y(n_292)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_270),
.Y(n_302)
);

MAJIxp5_ASAP7_75t_L g271 ( 
.A(n_254),
.B(n_221),
.C(n_218),
.Y(n_271)
);

INVxp67_ASAP7_75t_L g272 ( 
.A(n_256),
.Y(n_272)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_272),
.B(n_274),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_L g274 ( 
.A(n_237),
.B(n_204),
.Y(n_274)
);

NOR3xp33_ASAP7_75t_L g275 ( 
.A(n_237),
.B(n_231),
.C(n_214),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_SL g300 ( 
.A(n_275),
.B(n_241),
.Y(n_300)
);

AOI22xp5_ASAP7_75t_L g276 ( 
.A1(n_238),
.A2(n_210),
.B1(n_235),
.B2(n_217),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_242),
.B(n_246),
.Y(n_279)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_279),
.Y(n_299)
);

OAI22xp5_ASAP7_75t_L g280 ( 
.A1(n_264),
.A2(n_210),
.B1(n_221),
.B2(n_214),
.Y(n_280)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_280),
.B(n_281),
.Y(n_290)
);

INVxp67_ASAP7_75t_L g281 ( 
.A(n_244),
.Y(n_281)
);

MAJIxp5_ASAP7_75t_L g282 ( 
.A(n_254),
.B(n_222),
.C(n_230),
.Y(n_282)
);

XNOR2xp5_ASAP7_75t_L g304 ( 
.A(n_282),
.B(n_265),
.Y(n_304)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_283),
.B(n_284),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g284 ( 
.A(n_253),
.B(n_223),
.Y(n_284)
);

AO21x1_ASAP7_75t_L g285 ( 
.A1(n_244),
.A2(n_223),
.B(n_220),
.Y(n_285)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_285),
.B(n_288),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_L g287 ( 
.A(n_242),
.B(n_215),
.Y(n_287)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_287),
.Y(n_307)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_260),
.B(n_208),
.Y(n_288)
);

XNOR2xp5_ASAP7_75t_SL g313 ( 
.A(n_291),
.B(n_266),
.Y(n_313)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_293),
.A2(n_301),
.B1(n_305),
.B2(n_284),
.Y(n_309)
);

CKINVDCx16_ASAP7_75t_R g295 ( 
.A(n_270),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_SL g319 ( 
.A(n_295),
.B(n_296),
.Y(n_319)
);

AOI322xp5_ASAP7_75t_L g296 ( 
.A1(n_280),
.A2(n_255),
.A3(n_261),
.B1(n_240),
.B2(n_262),
.C1(n_247),
.C2(n_248),
.Y(n_296)
);

OAI22xp5_ASAP7_75t_L g298 ( 
.A1(n_276),
.A2(n_241),
.B1(n_251),
.B2(n_258),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g317 ( 
.A1(n_298),
.A2(n_278),
.B1(n_287),
.B2(n_277),
.Y(n_317)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_300),
.B(n_303),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g301 ( 
.A1(n_268),
.A2(n_249),
.B1(n_248),
.B2(n_257),
.Y(n_301)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_278),
.B(n_239),
.Y(n_303)
);

XOR2xp5_ASAP7_75t_L g312 ( 
.A(n_304),
.B(n_271),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g305 ( 
.A1(n_286),
.A2(n_259),
.B1(n_252),
.B2(n_239),
.Y(n_305)
);

MAJIxp5_ASAP7_75t_L g308 ( 
.A(n_292),
.B(n_282),
.C(n_269),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g325 ( 
.A(n_308),
.B(n_315),
.C(n_304),
.Y(n_325)
);

XOR2xp5_ASAP7_75t_L g331 ( 
.A(n_309),
.B(n_312),
.Y(n_331)
);

NAND2x1_ASAP7_75t_SL g310 ( 
.A(n_302),
.B(n_286),
.Y(n_310)
);

OR2x2_ASAP7_75t_L g334 ( 
.A(n_310),
.B(n_323),
.Y(n_334)
);

XNOR2xp5_ASAP7_75t_L g328 ( 
.A(n_313),
.B(n_314),
.Y(n_328)
);

OAI21xp5_ASAP7_75t_SL g314 ( 
.A1(n_306),
.A2(n_273),
.B(n_285),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g315 ( 
.A(n_292),
.B(n_273),
.Y(n_315)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_290),
.A2(n_279),
.B1(n_267),
.B2(n_288),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g330 ( 
.A1(n_316),
.A2(n_317),
.B1(n_318),
.B2(n_305),
.Y(n_330)
);

AOI22xp5_ASAP7_75t_SL g318 ( 
.A1(n_293),
.A2(n_283),
.B1(n_285),
.B2(n_274),
.Y(n_318)
);

INVx1_ASAP7_75t_L g320 ( 
.A(n_289),
.Y(n_320)
);

INVx1_ASAP7_75t_L g326 ( 
.A(n_320),
.Y(n_326)
);

AOI21xp5_ASAP7_75t_SL g321 ( 
.A1(n_306),
.A2(n_277),
.B(n_259),
.Y(n_321)
);

INVx1_ASAP7_75t_L g335 ( 
.A(n_321),
.Y(n_335)
);

NAND4xp25_ASAP7_75t_SL g322 ( 
.A(n_302),
.B(n_138),
.C(n_129),
.D(n_181),
.Y(n_322)
);

NOR2xp33_ASAP7_75t_SL g324 ( 
.A(n_322),
.B(n_297),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_L g323 ( 
.A1(n_294),
.A2(n_263),
.B(n_250),
.Y(n_323)
);

NAND2xp5_ASAP7_75t_L g339 ( 
.A(n_324),
.B(n_329),
.Y(n_339)
);

XOR2xp5_ASAP7_75t_L g342 ( 
.A(n_325),
.B(n_314),
.Y(n_342)
);

MAJIxp5_ASAP7_75t_L g327 ( 
.A(n_308),
.B(n_301),
.C(n_291),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g345 ( 
.A(n_327),
.B(n_332),
.C(n_333),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g329 ( 
.A(n_319),
.B(n_289),
.C(n_290),
.Y(n_329)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_330),
.A2(n_334),
.B1(n_323),
.B2(n_321),
.Y(n_341)
);

MAJIxp5_ASAP7_75t_L g332 ( 
.A(n_312),
.B(n_297),
.C(n_294),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g333 ( 
.A(n_315),
.B(n_299),
.C(n_307),
.Y(n_333)
);

AOI22xp5_ASAP7_75t_SL g336 ( 
.A1(n_335),
.A2(n_320),
.B1(n_316),
.B2(n_313),
.Y(n_336)
);

AND2x2_ASAP7_75t_L g351 ( 
.A(n_336),
.B(n_343),
.Y(n_351)
);

AOI22xp5_ASAP7_75t_L g337 ( 
.A1(n_326),
.A2(n_311),
.B1(n_299),
.B2(n_307),
.Y(n_337)
);

OAI22xp5_ASAP7_75t_L g349 ( 
.A1(n_337),
.A2(n_340),
.B1(n_243),
.B2(n_206),
.Y(n_349)
);

NAND4xp25_ASAP7_75t_SL g338 ( 
.A(n_334),
.B(n_322),
.C(n_310),
.D(n_309),
.Y(n_338)
);

NAND2xp5_ASAP7_75t_L g353 ( 
.A(n_338),
.B(n_344),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_328),
.A2(n_331),
.B1(n_318),
.B2(n_263),
.Y(n_340)
);

INVxp67_ASAP7_75t_L g347 ( 
.A(n_341),
.Y(n_347)
);

MAJIxp5_ASAP7_75t_L g352 ( 
.A(n_342),
.B(n_192),
.C(n_157),
.Y(n_352)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_331),
.B(n_250),
.Y(n_343)
);

XOR2xp5_ASAP7_75t_L g346 ( 
.A(n_343),
.B(n_327),
.Y(n_346)
);

BUFx24_ASAP7_75t_SL g344 ( 
.A(n_325),
.Y(n_344)
);

XOR2xp5_ASAP7_75t_L g354 ( 
.A(n_346),
.B(n_349),
.Y(n_354)
);

AOI21xp33_ASAP7_75t_L g348 ( 
.A1(n_339),
.A2(n_243),
.B(n_207),
.Y(n_348)
);

OR2x2_ASAP7_75t_L g356 ( 
.A(n_348),
.B(n_350),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_L g350 ( 
.A1(n_338),
.A2(n_192),
.B1(n_172),
.B2(n_127),
.Y(n_350)
);

AND2x2_ASAP7_75t_L g355 ( 
.A(n_351),
.B(n_352),
.Y(n_355)
);

NOR2xp33_ASAP7_75t_L g357 ( 
.A(n_353),
.B(n_342),
.Y(n_357)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_357),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g358 ( 
.A1(n_347),
.A2(n_345),
.B1(n_351),
.B2(n_346),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g361 ( 
.A(n_358),
.B(n_345),
.Y(n_361)
);

NOR2xp67_ASAP7_75t_SL g359 ( 
.A(n_357),
.B(n_347),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g362 ( 
.A(n_359),
.B(n_361),
.C(n_355),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_362),
.A2(n_360),
.B1(n_355),
.B2(n_356),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_SL g364 ( 
.A(n_363),
.B(n_354),
.Y(n_364)
);


endmodule