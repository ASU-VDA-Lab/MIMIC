module fake_jpeg_22706_n_79 (n_3, n_2, n_1, n_0, n_4, n_8, n_6, n_5, n_7, n_79);

input n_3;
input n_2;
input n_1;
input n_0;
input n_4;
input n_8;
input n_6;
input n_5;
input n_7;

output n_79;

wire n_10;
wire n_55;
wire n_64;
wire n_47;
wire n_51;
wire n_14;
wire n_73;
wire n_19;
wire n_59;
wire n_65;
wire n_42;
wire n_16;
wire n_49;
wire n_76;
wire n_28;
wire n_38;
wire n_26;
wire n_74;
wire n_31;
wire n_29;
wire n_50;
wire n_15;
wire n_13;
wire n_21;
wire n_57;
wire n_23;
wire n_69;
wire n_27;
wire n_40;
wire n_71;
wire n_30;
wire n_24;
wire n_44;
wire n_17;
wire n_25;
wire n_75;
wire n_37;
wire n_70;
wire n_66;
wire n_77;
wire n_61;
wire n_45;
wire n_78;
wire n_18;
wire n_20;
wire n_68;
wire n_52;
wire n_58;
wire n_41;
wire n_60;
wire n_63;
wire n_34;
wire n_39;
wire n_72;
wire n_11;
wire n_56;
wire n_12;
wire n_67;
wire n_53;
wire n_33;
wire n_54;
wire n_22;
wire n_35;
wire n_48;
wire n_46;
wire n_9;
wire n_36;
wire n_62;
wire n_43;
wire n_32;

BUFx16f_ASAP7_75t_L g9 ( 
.A(n_7),
.Y(n_9)
);

INVx6_ASAP7_75t_L g10 ( 
.A(n_5),
.Y(n_10)
);

BUFx6f_ASAP7_75t_L g11 ( 
.A(n_5),
.Y(n_11)
);

BUFx16f_ASAP7_75t_L g12 ( 
.A(n_7),
.Y(n_12)
);

INVx1_ASAP7_75t_L g13 ( 
.A(n_4),
.Y(n_13)
);

INVx1_ASAP7_75t_L g14 ( 
.A(n_1),
.Y(n_14)
);

CKINVDCx20_ASAP7_75t_R g15 ( 
.A(n_4),
.Y(n_15)
);

BUFx16f_ASAP7_75t_L g16 ( 
.A(n_0),
.Y(n_16)
);

BUFx3_ASAP7_75t_L g17 ( 
.A(n_0),
.Y(n_17)
);

INVx5_ASAP7_75t_L g18 ( 
.A(n_10),
.Y(n_18)
);

NOR2xp33_ASAP7_75t_L g24 ( 
.A(n_18),
.B(n_20),
.Y(n_24)
);

INVx2_ASAP7_75t_L g19 ( 
.A(n_9),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g26 ( 
.A(n_19),
.B(n_9),
.Y(n_26)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_15),
.Y(n_20)
);

INVx5_ASAP7_75t_L g21 ( 
.A(n_10),
.Y(n_21)
);

NOR2xp33_ASAP7_75t_L g25 ( 
.A(n_21),
.B(n_22),
.Y(n_25)
);

NOR2xp33_ASAP7_75t_L g22 ( 
.A(n_9),
.B(n_0),
.Y(n_22)
);

BUFx6f_ASAP7_75t_L g23 ( 
.A(n_17),
.Y(n_23)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_23),
.Y(n_27)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_26),
.Y(n_32)
);

OAI22xp5_ASAP7_75t_L g28 ( 
.A1(n_18),
.A2(n_10),
.B1(n_17),
.B2(n_14),
.Y(n_28)
);

AOI22xp5_ASAP7_75t_SL g35 ( 
.A1(n_28),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_35)
);

NOR2xp33_ASAP7_75t_L g29 ( 
.A(n_20),
.B(n_9),
.Y(n_29)
);

NAND2xp5_ASAP7_75t_L g33 ( 
.A(n_29),
.B(n_9),
.Y(n_33)
);

MAJIxp5_ASAP7_75t_SL g30 ( 
.A(n_28),
.B(n_17),
.C(n_12),
.Y(n_30)
);

CKINVDCx14_ASAP7_75t_R g38 ( 
.A(n_30),
.Y(n_38)
);

AND2x6_ASAP7_75t_L g31 ( 
.A(n_25),
.B(n_1),
.Y(n_31)
);

OAI22xp5_ASAP7_75t_SL g46 ( 
.A1(n_31),
.A2(n_35),
.B1(n_13),
.B2(n_14),
.Y(n_46)
);

NAND2xp5_ASAP7_75t_SL g39 ( 
.A(n_33),
.B(n_24),
.Y(n_39)
);

INVx13_ASAP7_75t_L g34 ( 
.A(n_27),
.Y(n_34)
);

NOR2xp33_ASAP7_75t_L g42 ( 
.A(n_34),
.B(n_12),
.Y(n_42)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_27),
.Y(n_36)
);

INVxp67_ASAP7_75t_L g41 ( 
.A(n_36),
.Y(n_41)
);

MAJIxp5_ASAP7_75t_L g37 ( 
.A(n_25),
.B(n_22),
.C(n_19),
.Y(n_37)
);

NAND2xp5_ASAP7_75t_L g45 ( 
.A(n_37),
.B(n_16),
.Y(n_45)
);

NAND2xp5_ASAP7_75t_L g54 ( 
.A(n_39),
.B(n_42),
.Y(n_54)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_36),
.Y(n_40)
);

NOR2xp33_ASAP7_75t_L g49 ( 
.A(n_40),
.B(n_44),
.Y(n_49)
);

NAND2xp5_ASAP7_75t_SL g43 ( 
.A(n_37),
.B(n_24),
.Y(n_43)
);

XNOR2xp5_ASAP7_75t_L g53 ( 
.A(n_43),
.B(n_21),
.Y(n_53)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_35),
.Y(n_44)
);

MAJIxp5_ASAP7_75t_L g51 ( 
.A(n_45),
.B(n_13),
.C(n_21),
.Y(n_51)
);

AND2x2_ASAP7_75t_L g50 ( 
.A(n_46),
.B(n_8),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_L g47 ( 
.A1(n_44),
.A2(n_30),
.B1(n_31),
.B2(n_32),
.Y(n_47)
);

OAI22xp5_ASAP7_75t_L g61 ( 
.A1(n_47),
.A2(n_48),
.B1(n_55),
.B2(n_23),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_SL g48 ( 
.A1(n_38),
.A2(n_31),
.B1(n_32),
.B2(n_33),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g62 ( 
.A(n_50),
.B(n_52),
.Y(n_62)
);

MAJIxp5_ASAP7_75t_L g57 ( 
.A(n_51),
.B(n_42),
.C(n_11),
.Y(n_57)
);

NOR2xp33_ASAP7_75t_L g52 ( 
.A(n_40),
.B(n_34),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g59 ( 
.A(n_53),
.B(n_23),
.Y(n_59)
);

OAI22xp5_ASAP7_75t_SL g55 ( 
.A1(n_43),
.A2(n_45),
.B1(n_46),
.B2(n_18),
.Y(n_55)
);

AOI322xp5_ASAP7_75t_SL g56 ( 
.A1(n_50),
.A2(n_39),
.A3(n_8),
.B1(n_41),
.B2(n_4),
.C1(n_5),
.C2(n_1),
.Y(n_56)
);

XNOR2xp5_ASAP7_75t_L g65 ( 
.A(n_56),
.B(n_58),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g63 ( 
.A(n_57),
.B(n_60),
.C(n_51),
.Y(n_63)
);

AOI21xp5_ASAP7_75t_L g58 ( 
.A1(n_49),
.A2(n_16),
.B(n_12),
.Y(n_58)
);

XNOR2xp5_ASAP7_75t_L g67 ( 
.A(n_59),
.B(n_61),
.Y(n_67)
);

MAJIxp5_ASAP7_75t_L g60 ( 
.A(n_55),
.B(n_23),
.C(n_34),
.Y(n_60)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_63),
.B(n_64),
.C(n_66),
.Y(n_69)
);

MAJIxp5_ASAP7_75t_L g64 ( 
.A(n_57),
.B(n_54),
.C(n_53),
.Y(n_64)
);

NAND2xp5_ASAP7_75t_SL g66 ( 
.A(n_62),
.B(n_60),
.Y(n_66)
);

OAI321xp33_ASAP7_75t_L g68 ( 
.A1(n_67),
.A2(n_48),
.A3(n_11),
.B1(n_12),
.B2(n_16),
.C(n_3),
.Y(n_68)
);

NAND2xp5_ASAP7_75t_L g73 ( 
.A(n_68),
.B(n_70),
.Y(n_73)
);

AOI21xp5_ASAP7_75t_SL g70 ( 
.A1(n_66),
.A2(n_12),
.B(n_16),
.Y(n_70)
);

OAI22xp5_ASAP7_75t_SL g71 ( 
.A1(n_69),
.A2(n_65),
.B1(n_11),
.B2(n_6),
.Y(n_71)
);

XNOR2xp5_ASAP7_75t_SL g75 ( 
.A(n_71),
.B(n_72),
.Y(n_75)
);

OAI22xp5_ASAP7_75t_L g72 ( 
.A1(n_68),
.A2(n_11),
.B1(n_3),
.B2(n_6),
.Y(n_72)
);

NOR2x1_ASAP7_75t_L g74 ( 
.A(n_73),
.B(n_16),
.Y(n_74)
);

OAI21xp5_ASAP7_75t_L g76 ( 
.A1(n_74),
.A2(n_73),
.B(n_71),
.Y(n_76)
);

INVx1_ASAP7_75t_L g77 ( 
.A(n_76),
.Y(n_77)
);

AOI21xp5_ASAP7_75t_L g78 ( 
.A1(n_77),
.A2(n_75),
.B(n_3),
.Y(n_78)
);

AOI221xp5_ASAP7_75t_L g79 ( 
.A1(n_78),
.A2(n_2),
.B1(n_6),
.B2(n_7),
.C(n_72),
.Y(n_79)
);


endmodule