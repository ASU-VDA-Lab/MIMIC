module fake_jpeg_12821_n_524 (n_13, n_11, n_14, n_17, n_16, n_3, n_2, n_1, n_0, n_10, n_12, n_4, n_8, n_9, n_15, n_6, n_5, n_7, n_524);

input n_13;
input n_11;
input n_14;
input n_17;
input n_16;
input n_3;
input n_2;
input n_1;
input n_0;
input n_10;
input n_12;
input n_4;
input n_8;
input n_9;
input n_15;
input n_6;
input n_5;
input n_7;

output n_524;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_415;
wire n_479;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_465;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_393;
wire n_349;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_486;
wire n_511;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_296;
wire n_384;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_491;
wire n_24;
wire n_467;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_18;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_494;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_492;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_472;
wire n_279;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_482;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_471;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVx1_ASAP7_75t_L g18 ( 
.A(n_3),
.Y(n_18)
);

INVx1_ASAP7_75t_L g19 ( 
.A(n_16),
.Y(n_19)
);

CKINVDCx20_ASAP7_75t_R g20 ( 
.A(n_9),
.Y(n_20)
);

BUFx6f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_1),
.Y(n_22)
);

CKINVDCx20_ASAP7_75t_R g23 ( 
.A(n_0),
.Y(n_23)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_2),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_12),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_15),
.Y(n_26)
);

NAND2xp5_ASAP7_75t_L g27 ( 
.A(n_11),
.B(n_4),
.Y(n_27)
);

INVx1_ASAP7_75t_L g28 ( 
.A(n_12),
.Y(n_28)
);

BUFx6f_ASAP7_75t_L g29 ( 
.A(n_10),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_11),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g31 ( 
.A(n_1),
.Y(n_31)
);

INVx1_ASAP7_75t_L g32 ( 
.A(n_2),
.Y(n_32)
);

INVx4_ASAP7_75t_L g33 ( 
.A(n_12),
.Y(n_33)
);

BUFx3_ASAP7_75t_L g34 ( 
.A(n_12),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_9),
.Y(n_35)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_14),
.Y(n_37)
);

INVx6_ASAP7_75t_L g38 ( 
.A(n_2),
.Y(n_38)
);

INVx6_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_11),
.Y(n_40)
);

BUFx5_ASAP7_75t_L g41 ( 
.A(n_3),
.Y(n_41)
);

BUFx12f_ASAP7_75t_L g42 ( 
.A(n_9),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_11),
.Y(n_43)
);

INVx2_ASAP7_75t_L g44 ( 
.A(n_4),
.Y(n_44)
);

CKINVDCx20_ASAP7_75t_R g45 ( 
.A(n_1),
.Y(n_45)
);

NOR2xp33_ASAP7_75t_L g46 ( 
.A(n_7),
.B(n_8),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

BUFx6f_ASAP7_75t_L g48 ( 
.A(n_2),
.Y(n_48)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_17),
.Y(n_50)
);

NOR2xp33_ASAP7_75t_L g51 ( 
.A(n_46),
.B(n_17),
.Y(n_51)
);

NOR2xp33_ASAP7_75t_SL g132 ( 
.A(n_51),
.B(n_76),
.Y(n_132)
);

INVx4_ASAP7_75t_SL g52 ( 
.A(n_21),
.Y(n_52)
);

INVx2_ASAP7_75t_SL g119 ( 
.A(n_52),
.Y(n_119)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_21),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_53),
.Y(n_111)
);

INVx1_ASAP7_75t_L g54 ( 
.A(n_35),
.Y(n_54)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_54),
.Y(n_118)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_33),
.Y(n_55)
);

INVx3_ASAP7_75t_L g104 ( 
.A(n_55),
.Y(n_104)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_35),
.Y(n_56)
);

NOR2xp33_ASAP7_75t_L g108 ( 
.A(n_56),
.B(n_59),
.Y(n_108)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_21),
.Y(n_57)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_57),
.Y(n_120)
);

NAND2xp5_ASAP7_75t_L g58 ( 
.A(n_27),
.B(n_16),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_L g121 ( 
.A(n_58),
.B(n_61),
.Y(n_121)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_44),
.Y(n_59)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_41),
.Y(n_60)
);

INVx3_ASAP7_75t_L g136 ( 
.A(n_60),
.Y(n_136)
);

NAND2xp5_ASAP7_75t_L g61 ( 
.A(n_27),
.B(n_16),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g62 ( 
.A(n_21),
.Y(n_62)
);

BUFx6f_ASAP7_75t_L g145 ( 
.A(n_62),
.Y(n_145)
);

BUFx24_ASAP7_75t_L g63 ( 
.A(n_41),
.Y(n_63)
);

BUFx5_ASAP7_75t_L g157 ( 
.A(n_63),
.Y(n_157)
);

INVx4_ASAP7_75t_L g64 ( 
.A(n_41),
.Y(n_64)
);

INVx3_ASAP7_75t_L g143 ( 
.A(n_64),
.Y(n_143)
);

INVx5_ASAP7_75t_L g65 ( 
.A(n_33),
.Y(n_65)
);

BUFx2_ASAP7_75t_L g161 ( 
.A(n_65),
.Y(n_161)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_29),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g148 ( 
.A(n_66),
.Y(n_148)
);

INVx8_ASAP7_75t_L g67 ( 
.A(n_29),
.Y(n_67)
);

INVx5_ASAP7_75t_L g105 ( 
.A(n_67),
.Y(n_105)
);

INVx11_ASAP7_75t_L g68 ( 
.A(n_42),
.Y(n_68)
);

INVx8_ASAP7_75t_L g126 ( 
.A(n_68),
.Y(n_126)
);

INVx2_ASAP7_75t_L g69 ( 
.A(n_44),
.Y(n_69)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_69),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g70 ( 
.A(n_29),
.Y(n_70)
);

BUFx6f_ASAP7_75t_L g153 ( 
.A(n_70),
.Y(n_153)
);

BUFx3_ASAP7_75t_L g71 ( 
.A(n_30),
.Y(n_71)
);

BUFx3_ASAP7_75t_L g159 ( 
.A(n_71),
.Y(n_159)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_30),
.Y(n_72)
);

INVx5_ASAP7_75t_L g107 ( 
.A(n_72),
.Y(n_107)
);

BUFx3_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_73),
.Y(n_125)
);

NOR2xp33_ASAP7_75t_SL g74 ( 
.A(n_36),
.B(n_0),
.Y(n_74)
);

NOR2xp33_ASAP7_75t_L g123 ( 
.A(n_74),
.B(n_83),
.Y(n_123)
);

INVx8_ASAP7_75t_L g75 ( 
.A(n_29),
.Y(n_75)
);

INVx5_ASAP7_75t_L g149 ( 
.A(n_75),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g76 ( 
.A(n_46),
.B(n_0),
.Y(n_76)
);

INVx5_ASAP7_75t_L g77 ( 
.A(n_33),
.Y(n_77)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_77),
.Y(n_160)
);

INVx2_ASAP7_75t_L g78 ( 
.A(n_44),
.Y(n_78)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_78),
.Y(n_106)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_42),
.Y(n_79)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_79),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g80 ( 
.A(n_34),
.Y(n_80)
);

INVx4_ASAP7_75t_L g110 ( 
.A(n_80),
.Y(n_110)
);

NOR2xp33_ASAP7_75t_L g81 ( 
.A(n_27),
.B(n_1),
.Y(n_81)
);

NAND2xp5_ASAP7_75t_SL g112 ( 
.A(n_81),
.B(n_87),
.Y(n_112)
);

BUFx8_ASAP7_75t_L g82 ( 
.A(n_34),
.Y(n_82)
);

INVx2_ASAP7_75t_SL g140 ( 
.A(n_82),
.Y(n_140)
);

INVx1_ASAP7_75t_L g83 ( 
.A(n_42),
.Y(n_83)
);

BUFx12_ASAP7_75t_L g84 ( 
.A(n_42),
.Y(n_84)
);

INVx8_ASAP7_75t_L g133 ( 
.A(n_84),
.Y(n_133)
);

INVx6_ASAP7_75t_L g85 ( 
.A(n_40),
.Y(n_85)
);

INVx6_ASAP7_75t_L g102 ( 
.A(n_85),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g86 ( 
.A(n_42),
.Y(n_86)
);

HB1xp67_ASAP7_75t_L g139 ( 
.A(n_86),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_36),
.B(n_3),
.Y(n_87)
);

BUFx5_ASAP7_75t_L g88 ( 
.A(n_40),
.Y(n_88)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_88),
.Y(n_124)
);

INVx4_ASAP7_75t_L g89 ( 
.A(n_42),
.Y(n_89)
);

INVx4_ASAP7_75t_L g137 ( 
.A(n_89),
.Y(n_137)
);

INVx1_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

NOR2xp33_ASAP7_75t_L g128 ( 
.A(n_90),
.B(n_50),
.Y(n_128)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_91),
.Y(n_114)
);

BUFx12f_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx4_ASAP7_75t_L g150 ( 
.A(n_92),
.Y(n_150)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_40),
.Y(n_93)
);

INVx6_ASAP7_75t_L g117 ( 
.A(n_93),
.Y(n_117)
);

INVx2_ASAP7_75t_L g94 ( 
.A(n_38),
.Y(n_94)
);

INVx2_ASAP7_75t_L g116 ( 
.A(n_94),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_40),
.Y(n_95)
);

INVx6_ASAP7_75t_L g127 ( 
.A(n_95),
.Y(n_127)
);

BUFx6f_ASAP7_75t_L g96 ( 
.A(n_48),
.Y(n_96)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_96),
.Y(n_141)
);

NAND2xp5_ASAP7_75t_L g97 ( 
.A(n_50),
.B(n_16),
.Y(n_97)
);

NAND2xp5_ASAP7_75t_L g144 ( 
.A(n_97),
.B(n_3),
.Y(n_144)
);

BUFx6f_ASAP7_75t_L g98 ( 
.A(n_48),
.Y(n_98)
);

INVx6_ASAP7_75t_L g146 ( 
.A(n_98),
.Y(n_146)
);

INVx3_ASAP7_75t_L g99 ( 
.A(n_39),
.Y(n_99)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_99),
.Y(n_122)
);

BUFx6f_ASAP7_75t_L g100 ( 
.A(n_48),
.Y(n_100)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_100),
.Y(n_151)
);

BUFx6f_ASAP7_75t_L g101 ( 
.A(n_48),
.Y(n_101)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_101),
.Y(n_142)
);

AND2x2_ASAP7_75t_SL g113 ( 
.A(n_81),
.B(n_39),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g170 ( 
.A(n_113),
.B(n_92),
.Y(n_170)
);

AOI22xp33_ASAP7_75t_SL g115 ( 
.A1(n_63),
.A2(n_39),
.B1(n_86),
.B2(n_67),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_L g176 ( 
.A1(n_115),
.A2(n_131),
.B1(n_134),
.B2(n_152),
.Y(n_176)
);

NOR2xp33_ASAP7_75t_L g164 ( 
.A(n_128),
.B(n_23),
.Y(n_164)
);

AND2x2_ASAP7_75t_L g129 ( 
.A(n_51),
.B(n_45),
.Y(n_129)
);

AOI21xp33_ASAP7_75t_L g196 ( 
.A1(n_129),
.A2(n_138),
.B(n_155),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_76),
.B(n_45),
.Y(n_130)
);

NAND2xp5_ASAP7_75t_SL g194 ( 
.A(n_130),
.B(n_135),
.Y(n_194)
);

AOI22xp33_ASAP7_75t_SL g131 ( 
.A1(n_75),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_131)
);

AO22x1_ASAP7_75t_SL g134 ( 
.A1(n_82),
.A2(n_49),
.B1(n_47),
.B2(n_43),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g135 ( 
.A(n_87),
.B(n_20),
.Y(n_135)
);

AND2x2_ASAP7_75t_L g138 ( 
.A(n_52),
.B(n_20),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g197 ( 
.A(n_144),
.B(n_162),
.Y(n_197)
);

AOI22xp5_ASAP7_75t_SL g147 ( 
.A1(n_73),
.A2(n_37),
.B1(n_31),
.B2(n_25),
.Y(n_147)
);

AOI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_147),
.A2(n_163),
.B1(n_93),
.B2(n_70),
.Y(n_222)
);

AOI22xp33_ASAP7_75t_SL g152 ( 
.A1(n_72),
.A2(n_22),
.B1(n_47),
.B2(n_43),
.Y(n_152)
);

AOI22xp33_ASAP7_75t_SL g154 ( 
.A1(n_72),
.A2(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g186 ( 
.A1(n_154),
.A2(n_156),
.B1(n_24),
.B2(n_49),
.Y(n_186)
);

AND2x2_ASAP7_75t_L g155 ( 
.A(n_80),
.B(n_23),
.Y(n_155)
);

AOI22xp33_ASAP7_75t_SL g156 ( 
.A1(n_80),
.A2(n_19),
.B1(n_32),
.B2(n_28),
.Y(n_156)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_85),
.Y(n_158)
);

INVx1_ASAP7_75t_L g167 ( 
.A(n_158),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_L g162 ( 
.A(n_53),
.B(n_25),
.Y(n_162)
);

OAI22xp5_ASAP7_75t_L g163 ( 
.A1(n_57),
.A2(n_101),
.B1(n_100),
.B2(n_98),
.Y(n_163)
);

NOR2xp33_ASAP7_75t_SL g254 ( 
.A(n_164),
.B(n_173),
.Y(n_254)
);

CKINVDCx16_ASAP7_75t_R g165 ( 
.A(n_139),
.Y(n_165)
);

NAND2xp5_ASAP7_75t_SL g248 ( 
.A(n_165),
.B(n_207),
.Y(n_248)
);

INVx1_ASAP7_75t_L g166 ( 
.A(n_139),
.Y(n_166)
);

INVx1_ASAP7_75t_L g224 ( 
.A(n_166),
.Y(n_224)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_142),
.Y(n_168)
);

INVx2_ASAP7_75t_L g247 ( 
.A(n_168),
.Y(n_247)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_119),
.Y(n_169)
);

INVx1_ASAP7_75t_SL g226 ( 
.A(n_169),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g231 ( 
.A1(n_170),
.A2(n_202),
.B(n_115),
.Y(n_231)
);

INVx3_ASAP7_75t_L g171 ( 
.A(n_105),
.Y(n_171)
);

INVx4_ASAP7_75t_L g229 ( 
.A(n_171),
.Y(n_229)
);

INVx6_ASAP7_75t_L g172 ( 
.A(n_111),
.Y(n_172)
);

BUFx6f_ASAP7_75t_L g230 ( 
.A(n_172),
.Y(n_230)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_123),
.B(n_92),
.Y(n_173)
);

INVx5_ASAP7_75t_L g174 ( 
.A(n_125),
.Y(n_174)
);

INVx3_ASAP7_75t_L g246 ( 
.A(n_174),
.Y(n_246)
);

INVx1_ASAP7_75t_L g175 ( 
.A(n_118),
.Y(n_175)
);

INVx2_ASAP7_75t_SL g275 ( 
.A(n_175),
.Y(n_275)
);

MAJIxp5_ASAP7_75t_L g177 ( 
.A(n_113),
.B(n_84),
.C(n_95),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_177),
.B(n_126),
.Y(n_266)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_114),
.Y(n_178)
);

INVx2_ASAP7_75t_L g264 ( 
.A(n_178),
.Y(n_264)
);

BUFx3_ASAP7_75t_L g179 ( 
.A(n_140),
.Y(n_179)
);

INVx5_ASAP7_75t_L g234 ( 
.A(n_179),
.Y(n_234)
);

INVx1_ASAP7_75t_L g180 ( 
.A(n_108),
.Y(n_180)
);

INVx1_ASAP7_75t_L g227 ( 
.A(n_180),
.Y(n_227)
);

INVx1_ASAP7_75t_L g181 ( 
.A(n_116),
.Y(n_181)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_181),
.Y(n_228)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_103),
.Y(n_182)
);

INVx1_ASAP7_75t_L g232 ( 
.A(n_182),
.Y(n_232)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_119),
.Y(n_183)
);

INVx1_ASAP7_75t_L g236 ( 
.A(n_183),
.Y(n_236)
);

INVx2_ASAP7_75t_SL g184 ( 
.A(n_157),
.Y(n_184)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_184),
.Y(n_253)
);

INVx2_ASAP7_75t_L g185 ( 
.A(n_106),
.Y(n_185)
);

INVx1_ASAP7_75t_L g257 ( 
.A(n_185),
.Y(n_257)
);

INVxp67_ASAP7_75t_L g263 ( 
.A(n_186),
.Y(n_263)
);

BUFx6f_ASAP7_75t_L g187 ( 
.A(n_111),
.Y(n_187)
);

INVx3_ASAP7_75t_L g252 ( 
.A(n_187),
.Y(n_252)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_155),
.Y(n_188)
);

NOR2xp33_ASAP7_75t_L g241 ( 
.A(n_188),
.B(n_193),
.Y(n_241)
);

INVx1_ASAP7_75t_L g189 ( 
.A(n_122),
.Y(n_189)
);

INVx1_ASAP7_75t_L g270 ( 
.A(n_189),
.Y(n_270)
);

INVx2_ASAP7_75t_L g190 ( 
.A(n_109),
.Y(n_190)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_190),
.Y(n_262)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_102),
.Y(n_191)
);

INVx3_ASAP7_75t_L g271 ( 
.A(n_191),
.Y(n_271)
);

HB1xp67_ASAP7_75t_L g192 ( 
.A(n_137),
.Y(n_192)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_192),
.Y(n_258)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_104),
.Y(n_193)
);

INVx1_ASAP7_75t_SL g195 ( 
.A(n_133),
.Y(n_195)
);

CKINVDCx14_ASAP7_75t_R g255 ( 
.A(n_195),
.Y(n_255)
);

AND2x2_ASAP7_75t_SL g198 ( 
.A(n_121),
.B(n_96),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_SL g249 ( 
.A(n_198),
.B(n_146),
.Y(n_249)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_120),
.Y(n_199)
);

INVx3_ASAP7_75t_L g273 ( 
.A(n_199),
.Y(n_273)
);

INVx3_ASAP7_75t_L g200 ( 
.A(n_149),
.Y(n_200)
);

CKINVDCx20_ASAP7_75t_R g237 ( 
.A(n_200),
.Y(n_237)
);

BUFx12f_ASAP7_75t_L g201 ( 
.A(n_159),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_201),
.B(n_203),
.Y(n_245)
);

OAI21xp33_ASAP7_75t_SL g202 ( 
.A1(n_129),
.A2(n_134),
.B(n_132),
.Y(n_202)
);

INVx1_ASAP7_75t_L g203 ( 
.A(n_138),
.Y(n_203)
);

INVx5_ASAP7_75t_L g204 ( 
.A(n_110),
.Y(n_204)
);

INVxp33_ASAP7_75t_L g242 ( 
.A(n_204),
.Y(n_242)
);

AOI22xp33_ASAP7_75t_SL g205 ( 
.A1(n_161),
.A2(n_18),
.B1(n_24),
.B2(n_22),
.Y(n_205)
);

AOI22xp33_ASAP7_75t_SL g238 ( 
.A1(n_205),
.A2(n_206),
.B1(n_210),
.B2(n_215),
.Y(n_238)
);

AOI22xp33_ASAP7_75t_SL g206 ( 
.A1(n_161),
.A2(n_22),
.B1(n_18),
.B2(n_32),
.Y(n_206)
);

INVx1_ASAP7_75t_L g207 ( 
.A(n_137),
.Y(n_207)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_160),
.Y(n_208)
);

NOR2xp33_ASAP7_75t_L g259 ( 
.A(n_208),
.B(n_211),
.Y(n_259)
);

HB1xp67_ASAP7_75t_L g209 ( 
.A(n_110),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g240 ( 
.A(n_209),
.Y(n_240)
);

AOI22xp33_ASAP7_75t_SL g210 ( 
.A1(n_136),
.A2(n_19),
.B1(n_28),
.B2(n_26),
.Y(n_210)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_102),
.Y(n_211)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_143),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_SL g256 ( 
.A(n_212),
.B(n_213),
.Y(n_256)
);

INVx4_ASAP7_75t_L g213 ( 
.A(n_150),
.Y(n_213)
);

INVx1_ASAP7_75t_L g214 ( 
.A(n_140),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_SL g260 ( 
.A(n_214),
.B(n_216),
.Y(n_260)
);

INVx5_ASAP7_75t_L g215 ( 
.A(n_150),
.Y(n_215)
);

INVx2_ASAP7_75t_L g216 ( 
.A(n_117),
.Y(n_216)
);

AOI22xp33_ASAP7_75t_SL g217 ( 
.A1(n_159),
.A2(n_18),
.B1(n_26),
.B2(n_24),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_L g272 ( 
.A1(n_217),
.A2(n_220),
.B1(n_222),
.B2(n_5),
.Y(n_272)
);

INVx5_ASAP7_75t_L g218 ( 
.A(n_124),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_219),
.Y(n_267)
);

INVx1_ASAP7_75t_L g219 ( 
.A(n_117),
.Y(n_219)
);

AOI22xp33_ASAP7_75t_SL g220 ( 
.A1(n_124),
.A2(n_26),
.B1(n_37),
.B2(n_31),
.Y(n_220)
);

INVx2_ASAP7_75t_L g221 ( 
.A(n_127),
.Y(n_221)
);

NAND2xp5_ASAP7_75t_L g225 ( 
.A(n_221),
.B(n_141),
.Y(n_225)
);

NOR2xp33_ASAP7_75t_L g223 ( 
.A(n_112),
.B(n_4),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_SL g268 ( 
.A(n_223),
.B(n_4),
.Y(n_268)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_225),
.Y(n_297)
);

AND2x2_ASAP7_75t_L g293 ( 
.A(n_231),
.B(n_272),
.Y(n_293)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_198),
.B(n_131),
.Y(n_233)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_233),
.B(n_274),
.Y(n_306)
);

OAI21xp5_ASAP7_75t_SL g235 ( 
.A1(n_170),
.A2(n_154),
.B(n_152),
.Y(n_235)
);

AOI21xp5_ASAP7_75t_SL g283 ( 
.A1(n_235),
.A2(n_263),
.B(n_231),
.Y(n_283)
);

AOI22xp33_ASAP7_75t_L g239 ( 
.A1(n_222),
.A2(n_141),
.B1(n_127),
.B2(n_151),
.Y(n_239)
);

OAI22xp5_ASAP7_75t_L g311 ( 
.A1(n_239),
.A2(n_244),
.B1(n_250),
.B2(n_251),
.Y(n_311)
);

OAI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_177),
.A2(n_156),
.B1(n_66),
.B2(n_62),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_243),
.A2(n_184),
.B1(n_204),
.B2(n_201),
.Y(n_295)
);

AOI22xp5_ASAP7_75t_L g244 ( 
.A1(n_176),
.A2(n_151),
.B1(n_146),
.B2(n_148),
.Y(n_244)
);

XNOR2xp5_ASAP7_75t_L g278 ( 
.A(n_249),
.B(n_266),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g250 ( 
.A1(n_170),
.A2(n_153),
.B1(n_148),
.B2(n_145),
.Y(n_250)
);

AOI22xp33_ASAP7_75t_L g251 ( 
.A1(n_197),
.A2(n_153),
.B1(n_145),
.B2(n_120),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g261 ( 
.A1(n_198),
.A2(n_126),
.B1(n_107),
.B2(n_133),
.Y(n_261)
);

OAI22xp5_ASAP7_75t_SL g277 ( 
.A1(n_261),
.A2(n_265),
.B1(n_274),
.B2(n_238),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g265 ( 
.A1(n_191),
.A2(n_211),
.B1(n_196),
.B2(n_182),
.Y(n_265)
);

NAND2xp5_ASAP7_75t_SL g310 ( 
.A(n_268),
.B(n_10),
.Y(n_310)
);

AOI22xp33_ASAP7_75t_L g269 ( 
.A1(n_178),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_269)
);

OAI22xp33_ASAP7_75t_L g276 ( 
.A1(n_269),
.A2(n_172),
.B1(n_199),
.B2(n_187),
.Y(n_276)
);

AOI22xp5_ASAP7_75t_L g274 ( 
.A1(n_185),
.A2(n_5),
.B1(n_6),
.B2(n_7),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g361 ( 
.A(n_276),
.B(n_307),
.Y(n_361)
);

AOI22xp5_ASAP7_75t_L g327 ( 
.A1(n_277),
.A2(n_292),
.B1(n_255),
.B2(n_237),
.Y(n_327)
);

AOI22xp33_ASAP7_75t_L g279 ( 
.A1(n_263),
.A2(n_171),
.B1(n_200),
.B2(n_221),
.Y(n_279)
);

CKINVDCx16_ASAP7_75t_R g342 ( 
.A(n_279),
.Y(n_342)
);

INVx2_ASAP7_75t_SL g280 ( 
.A(n_253),
.Y(n_280)
);

INVx1_ASAP7_75t_L g332 ( 
.A(n_280),
.Y(n_332)
);

INVx2_ASAP7_75t_L g281 ( 
.A(n_271),
.Y(n_281)
);

INVx1_ASAP7_75t_L g333 ( 
.A(n_281),
.Y(n_333)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_249),
.B(n_167),
.Y(n_282)
);

NAND2xp5_ASAP7_75t_L g323 ( 
.A(n_282),
.B(n_288),
.Y(n_323)
);

OAI21xp5_ASAP7_75t_SL g329 ( 
.A1(n_283),
.A2(n_306),
.B(n_320),
.Y(n_329)
);

XNOR2xp5_ASAP7_75t_L g284 ( 
.A(n_266),
.B(n_194),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_284),
.B(n_286),
.C(n_316),
.Y(n_358)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_271),
.Y(n_285)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_285),
.Y(n_352)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_265),
.B(n_166),
.C(n_190),
.Y(n_286)
);

INVx2_ASAP7_75t_L g287 ( 
.A(n_247),
.Y(n_287)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_287),
.Y(n_353)
);

NAND2xp5_ASAP7_75t_L g288 ( 
.A(n_233),
.B(n_168),
.Y(n_288)
);

OAI21xp5_ASAP7_75t_SL g289 ( 
.A1(n_261),
.A2(n_207),
.B(n_195),
.Y(n_289)
);

AOI21xp5_ASAP7_75t_L g350 ( 
.A1(n_289),
.A2(n_234),
.B(n_246),
.Y(n_350)
);

NOR2xp33_ASAP7_75t_L g290 ( 
.A(n_254),
.B(n_179),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g336 ( 
.A(n_290),
.B(n_303),
.Y(n_336)
);

NOR2x1_ASAP7_75t_L g291 ( 
.A(n_275),
.B(n_213),
.Y(n_291)
);

NAND2xp5_ASAP7_75t_SL g360 ( 
.A(n_291),
.B(n_314),
.Y(n_360)
);

OAI22xp5_ASAP7_75t_SL g292 ( 
.A1(n_244),
.A2(n_216),
.B1(n_174),
.B2(n_218),
.Y(n_292)
);

NAND2xp5_ASAP7_75t_L g294 ( 
.A(n_243),
.B(n_215),
.Y(n_294)
);

NAND2xp5_ASAP7_75t_L g338 ( 
.A(n_294),
.B(n_308),
.Y(n_338)
);

OAI22xp5_ASAP7_75t_SL g344 ( 
.A1(n_295),
.A2(n_294),
.B1(n_296),
.B2(n_283),
.Y(n_344)
);

OAI21xp5_ASAP7_75t_L g296 ( 
.A1(n_235),
.A2(n_201),
.B(n_6),
.Y(n_296)
);

OAI21xp5_ASAP7_75t_L g328 ( 
.A1(n_296),
.A2(n_242),
.B(n_226),
.Y(n_328)
);

AOI22xp5_ASAP7_75t_L g298 ( 
.A1(n_225),
.A2(n_5),
.B1(n_7),
.B2(n_8),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_298),
.A2(n_317),
.B1(n_252),
.B2(n_273),
.Y(n_346)
);

INVx1_ASAP7_75t_L g299 ( 
.A(n_224),
.Y(n_299)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_299),
.Y(n_355)
);

INVx2_ASAP7_75t_L g300 ( 
.A(n_247),
.Y(n_300)
);

BUFx3_ASAP7_75t_L g325 ( 
.A(n_300),
.Y(n_325)
);

AND2x2_ASAP7_75t_L g301 ( 
.A(n_241),
.B(n_8),
.Y(n_301)
);

OAI21xp33_ASAP7_75t_L g326 ( 
.A1(n_301),
.A2(n_15),
.B(n_240),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g302 ( 
.A(n_245),
.Y(n_302)
);

NOR2xp33_ASAP7_75t_L g331 ( 
.A(n_302),
.B(n_305),
.Y(n_331)
);

NOR2xp33_ASAP7_75t_L g303 ( 
.A(n_227),
.B(n_268),
.Y(n_303)
);

INVxp67_ASAP7_75t_L g304 ( 
.A(n_267),
.Y(n_304)
);

INVx13_ASAP7_75t_L g348 ( 
.A(n_304),
.Y(n_348)
);

BUFx24_ASAP7_75t_SL g305 ( 
.A(n_227),
.Y(n_305)
);

INVx1_ASAP7_75t_SL g307 ( 
.A(n_253),
.Y(n_307)
);

OA22x2_ASAP7_75t_L g308 ( 
.A1(n_237),
.A2(n_8),
.B1(n_10),
.B2(n_13),
.Y(n_308)
);

NOR2xp33_ASAP7_75t_L g309 ( 
.A(n_236),
.B(n_10),
.Y(n_309)
);

NOR2xp33_ASAP7_75t_L g347 ( 
.A(n_309),
.B(n_310),
.Y(n_347)
);

CKINVDCx20_ASAP7_75t_R g312 ( 
.A(n_259),
.Y(n_312)
);

NOR2xp33_ASAP7_75t_L g356 ( 
.A(n_312),
.B(n_313),
.Y(n_356)
);

INVxp67_ASAP7_75t_L g313 ( 
.A(n_256),
.Y(n_313)
);

NAND2xp5_ASAP7_75t_L g314 ( 
.A(n_240),
.B(n_13),
.Y(n_314)
);

A2O1A1Ixp33_ASAP7_75t_L g315 ( 
.A1(n_236),
.A2(n_224),
.B(n_228),
.C(n_270),
.Y(n_315)
);

O2A1O1Ixp33_ASAP7_75t_L g351 ( 
.A1(n_315),
.A2(n_258),
.B(n_262),
.C(n_264),
.Y(n_351)
);

MAJIxp5_ASAP7_75t_L g316 ( 
.A(n_248),
.B(n_13),
.C(n_14),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_L g317 ( 
.A1(n_275),
.A2(n_13),
.B1(n_14),
.B2(n_15),
.Y(n_317)
);

INVx1_ASAP7_75t_L g318 ( 
.A(n_275),
.Y(n_318)
);

BUFx3_ASAP7_75t_L g349 ( 
.A(n_318),
.Y(n_349)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_228),
.Y(n_319)
);

BUFx5_ASAP7_75t_L g334 ( 
.A(n_319),
.Y(n_334)
);

AO22x1_ASAP7_75t_L g320 ( 
.A1(n_270),
.A2(n_15),
.B1(n_229),
.B2(n_232),
.Y(n_320)
);

CKINVDCx20_ASAP7_75t_R g321 ( 
.A(n_260),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g330 ( 
.A(n_321),
.Y(n_330)
);

INVx2_ASAP7_75t_L g322 ( 
.A(n_229),
.Y(n_322)
);

CKINVDCx20_ASAP7_75t_R g337 ( 
.A(n_322),
.Y(n_337)
);

OA21x2_ASAP7_75t_L g324 ( 
.A1(n_293),
.A2(n_226),
.B(n_246),
.Y(n_324)
);

OAI21xp5_ASAP7_75t_SL g370 ( 
.A1(n_324),
.A2(n_350),
.B(n_280),
.Y(n_370)
);

XOR2xp5_ASAP7_75t_SL g376 ( 
.A(n_326),
.B(n_317),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_L g368 ( 
.A1(n_327),
.A2(n_280),
.B1(n_292),
.B2(n_298),
.Y(n_368)
);

INVxp67_ASAP7_75t_L g385 ( 
.A(n_328),
.Y(n_385)
);

XNOR2xp5_ASAP7_75t_L g335 ( 
.A(n_278),
.B(n_232),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_335),
.B(n_339),
.C(n_359),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g339 ( 
.A(n_278),
.B(n_257),
.Y(n_339)
);

AOI22xp5_ASAP7_75t_L g340 ( 
.A1(n_277),
.A2(n_273),
.B1(n_252),
.B2(n_230),
.Y(n_340)
);

OAI22xp5_ASAP7_75t_SL g378 ( 
.A1(n_340),
.A2(n_342),
.B1(n_327),
.B2(n_350),
.Y(n_378)
);

CKINVDCx20_ASAP7_75t_R g341 ( 
.A(n_315),
.Y(n_341)
);

NOR2xp33_ASAP7_75t_L g371 ( 
.A(n_341),
.B(n_354),
.Y(n_371)
);

OAI32xp33_ASAP7_75t_L g343 ( 
.A1(n_288),
.A2(n_242),
.A3(n_257),
.B1(n_264),
.B2(n_230),
.Y(n_343)
);

NAND2xp5_ASAP7_75t_L g377 ( 
.A(n_343),
.B(n_308),
.Y(n_377)
);

AOI22xp5_ASAP7_75t_L g372 ( 
.A1(n_344),
.A2(n_346),
.B1(n_357),
.B2(n_363),
.Y(n_372)
);

OAI21xp5_ASAP7_75t_SL g345 ( 
.A1(n_293),
.A2(n_282),
.B(n_286),
.Y(n_345)
);

AOI21xp5_ASAP7_75t_L g364 ( 
.A1(n_345),
.A2(n_289),
.B(n_301),
.Y(n_364)
);

AND2x2_ASAP7_75t_L g365 ( 
.A(n_351),
.B(n_291),
.Y(n_365)
);

CKINVDCx16_ASAP7_75t_R g354 ( 
.A(n_301),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g357 ( 
.A1(n_297),
.A2(n_293),
.B1(n_295),
.B2(n_304),
.Y(n_357)
);

XNOR2xp5_ASAP7_75t_L g359 ( 
.A(n_284),
.B(n_262),
.Y(n_359)
);

CKINVDCx20_ASAP7_75t_R g362 ( 
.A(n_287),
.Y(n_362)
);

NOR2xp33_ASAP7_75t_L g380 ( 
.A(n_362),
.B(n_332),
.Y(n_380)
);

OAI22xp5_ASAP7_75t_L g363 ( 
.A1(n_313),
.A2(n_234),
.B1(n_311),
.B2(n_307),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g421 ( 
.A(n_364),
.B(n_392),
.Y(n_421)
);

INVx1_ASAP7_75t_L g411 ( 
.A(n_365),
.Y(n_411)
);

CKINVDCx20_ASAP7_75t_R g366 ( 
.A(n_356),
.Y(n_366)
);

INVx13_ASAP7_75t_L g413 ( 
.A(n_366),
.Y(n_413)
);

XOR2x1_ASAP7_75t_SL g367 ( 
.A(n_344),
.B(n_320),
.Y(n_367)
);

NAND2x1_ASAP7_75t_SL g426 ( 
.A(n_367),
.B(n_392),
.Y(n_426)
);

AOI22xp5_ASAP7_75t_L g402 ( 
.A1(n_368),
.A2(n_378),
.B1(n_393),
.B2(n_346),
.Y(n_402)
);

OAI32xp33_ASAP7_75t_L g369 ( 
.A1(n_338),
.A2(n_320),
.A3(n_322),
.B1(n_308),
.B2(n_285),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g404 ( 
.A(n_369),
.B(n_384),
.Y(n_404)
);

OAI21xp5_ASAP7_75t_L g415 ( 
.A1(n_370),
.A2(n_375),
.B(n_379),
.Y(n_415)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_355),
.Y(n_373)
);

INVx1_ASAP7_75t_L g417 ( 
.A(n_373),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g374 ( 
.A1(n_357),
.A2(n_281),
.B1(n_300),
.B2(n_276),
.Y(n_374)
);

OAI22xp5_ASAP7_75t_L g401 ( 
.A1(n_374),
.A2(n_377),
.B1(n_337),
.B2(n_349),
.Y(n_401)
);

OAI21xp5_ASAP7_75t_SL g375 ( 
.A1(n_324),
.A2(n_316),
.B(n_308),
.Y(n_375)
);

NAND2xp5_ASAP7_75t_SL g428 ( 
.A(n_376),
.B(n_381),
.Y(n_428)
);

AOI21xp5_ASAP7_75t_L g379 ( 
.A1(n_329),
.A2(n_341),
.B(n_328),
.Y(n_379)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_380),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_L g381 ( 
.A(n_336),
.B(n_330),
.Y(n_381)
);

NAND2xp5_ASAP7_75t_L g382 ( 
.A(n_330),
.B(n_332),
.Y(n_382)
);

INVx1_ASAP7_75t_L g427 ( 
.A(n_382),
.Y(n_427)
);

INVx2_ASAP7_75t_L g383 ( 
.A(n_325),
.Y(n_383)
);

HB1xp67_ASAP7_75t_L g416 ( 
.A(n_383),
.Y(n_416)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_355),
.Y(n_384)
);

XOR2xp5_ASAP7_75t_L g386 ( 
.A(n_335),
.B(n_339),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g407 ( 
.A(n_386),
.B(n_347),
.C(n_333),
.Y(n_407)
);

CKINVDCx20_ASAP7_75t_R g387 ( 
.A(n_360),
.Y(n_387)
);

NAND2xp5_ASAP7_75t_L g408 ( 
.A(n_387),
.B(n_390),
.Y(n_408)
);

OAI21xp5_ASAP7_75t_SL g388 ( 
.A1(n_324),
.A2(n_338),
.B(n_360),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g418 ( 
.A(n_388),
.B(n_397),
.Y(n_418)
);

INVx6_ASAP7_75t_L g389 ( 
.A(n_348),
.Y(n_389)
);

BUFx6f_ASAP7_75t_L g406 ( 
.A(n_389),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g390 ( 
.A(n_336),
.B(n_331),
.Y(n_390)
);

BUFx3_ASAP7_75t_L g391 ( 
.A(n_349),
.Y(n_391)
);

AOI22xp33_ASAP7_75t_SL g412 ( 
.A1(n_391),
.A2(n_394),
.B1(n_396),
.B2(n_352),
.Y(n_412)
);

AOI21xp5_ASAP7_75t_L g392 ( 
.A1(n_329),
.A2(n_345),
.B(n_361),
.Y(n_392)
);

OAI22xp5_ASAP7_75t_SL g393 ( 
.A1(n_340),
.A2(n_323),
.B1(n_342),
.B2(n_358),
.Y(n_393)
);

INVx1_ASAP7_75t_L g394 ( 
.A(n_353),
.Y(n_394)
);

INVx1_ASAP7_75t_L g396 ( 
.A(n_353),
.Y(n_396)
);

CKINVDCx20_ASAP7_75t_R g397 ( 
.A(n_363),
.Y(n_397)
);

CKINVDCx20_ASAP7_75t_R g398 ( 
.A(n_361),
.Y(n_398)
);

CKINVDCx20_ASAP7_75t_R g403 ( 
.A(n_398),
.Y(n_403)
);

OAI22xp5_ASAP7_75t_SL g399 ( 
.A1(n_372),
.A2(n_323),
.B1(n_358),
.B2(n_354),
.Y(n_399)
);

AOI22xp5_ASAP7_75t_L g444 ( 
.A1(n_399),
.A2(n_400),
.B1(n_401),
.B2(n_405),
.Y(n_444)
);

OAI22x1_ASAP7_75t_SL g400 ( 
.A1(n_372),
.A2(n_351),
.B1(n_361),
.B2(n_348),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_402),
.B(n_422),
.Y(n_429)
);

OAI22xp5_ASAP7_75t_SL g405 ( 
.A1(n_377),
.A2(n_343),
.B1(n_359),
.B2(n_337),
.Y(n_405)
);

XOR2xp5_ASAP7_75t_L g452 ( 
.A(n_407),
.B(n_409),
.Y(n_452)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_395),
.B(n_333),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g410 ( 
.A1(n_387),
.A2(n_362),
.B1(n_352),
.B2(n_325),
.Y(n_410)
);

INVx1_ASAP7_75t_L g433 ( 
.A(n_410),
.Y(n_433)
);

INVxp67_ASAP7_75t_L g445 ( 
.A(n_412),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_382),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_414),
.B(n_381),
.Y(n_431)
);

XOR2xp5_ASAP7_75t_L g419 ( 
.A(n_395),
.B(n_334),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g434 ( 
.A(n_419),
.B(n_420),
.C(n_425),
.Y(n_434)
);

MAJIxp5_ASAP7_75t_L g420 ( 
.A(n_386),
.B(n_334),
.C(n_393),
.Y(n_420)
);

AND2x2_ASAP7_75t_SL g430 ( 
.A(n_421),
.B(n_370),
.Y(n_430)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_397),
.A2(n_379),
.B1(n_398),
.B2(n_371),
.Y(n_422)
);

AOI22xp5_ASAP7_75t_L g423 ( 
.A1(n_378),
.A2(n_368),
.B1(n_385),
.B2(n_365),
.Y(n_423)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_423),
.B(n_369),
.Y(n_438)
);

XNOR2xp5_ASAP7_75t_L g425 ( 
.A(n_371),
.B(n_388),
.Y(n_425)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_430),
.B(n_453),
.Y(n_455)
);

INVx1_ASAP7_75t_L g462 ( 
.A(n_431),
.Y(n_462)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_406),
.Y(n_432)
);

INVx1_ASAP7_75t_L g466 ( 
.A(n_432),
.Y(n_466)
);

XNOR2xp5_ASAP7_75t_L g435 ( 
.A(n_409),
.B(n_419),
.Y(n_435)
);

XNOR2xp5_ASAP7_75t_L g454 ( 
.A(n_435),
.B(n_415),
.Y(n_454)
);

A2O1A1Ixp33_ASAP7_75t_SL g436 ( 
.A1(n_411),
.A2(n_367),
.B(n_365),
.C(n_364),
.Y(n_436)
);

OAI22xp5_ASAP7_75t_SL g457 ( 
.A1(n_436),
.A2(n_438),
.B1(n_415),
.B2(n_423),
.Y(n_457)
);

OAI21xp5_ASAP7_75t_SL g437 ( 
.A1(n_418),
.A2(n_367),
.B(n_366),
.Y(n_437)
);

AOI21xp5_ASAP7_75t_L g465 ( 
.A1(n_437),
.A2(n_451),
.B(n_404),
.Y(n_465)
);

MAJIxp5_ASAP7_75t_L g439 ( 
.A(n_420),
.B(n_380),
.C(n_394),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g456 ( 
.A(n_439),
.B(n_448),
.C(n_450),
.Y(n_456)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_424),
.Y(n_440)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_440),
.Y(n_470)
);

CKINVDCx20_ASAP7_75t_R g441 ( 
.A(n_416),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_L g459 ( 
.A(n_441),
.B(n_443),
.Y(n_459)
);

NOR2xp33_ASAP7_75t_L g442 ( 
.A(n_408),
.B(n_390),
.Y(n_442)
);

NOR2xp33_ASAP7_75t_SL g468 ( 
.A(n_442),
.B(n_389),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g443 ( 
.A(n_408),
.Y(n_443)
);

INVx1_ASAP7_75t_L g446 ( 
.A(n_424),
.Y(n_446)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_446),
.B(n_447),
.Y(n_461)
);

INVxp67_ASAP7_75t_L g447 ( 
.A(n_422),
.Y(n_447)
);

MAJIxp5_ASAP7_75t_L g448 ( 
.A(n_407),
.B(n_399),
.C(n_421),
.Y(n_448)
);

CKINVDCx14_ASAP7_75t_R g449 ( 
.A(n_428),
.Y(n_449)
);

NAND2xp5_ASAP7_75t_SL g471 ( 
.A(n_449),
.B(n_413),
.Y(n_471)
);

MAJIxp5_ASAP7_75t_L g450 ( 
.A(n_425),
.B(n_396),
.C(n_375),
.Y(n_450)
);

OAI21xp5_ASAP7_75t_SL g451 ( 
.A1(n_403),
.A2(n_376),
.B(n_373),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_SL g453 ( 
.A(n_405),
.B(n_384),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_SL g487 ( 
.A(n_454),
.B(n_463),
.Y(n_487)
);

INVxp67_ASAP7_75t_L g479 ( 
.A(n_457),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g458 ( 
.A(n_452),
.B(n_427),
.C(n_411),
.Y(n_458)
);

NAND2xp5_ASAP7_75t_L g475 ( 
.A(n_458),
.B(n_460),
.Y(n_475)
);

MAJIxp5_ASAP7_75t_L g460 ( 
.A(n_452),
.B(n_427),
.C(n_402),
.Y(n_460)
);

XOR2xp5_ASAP7_75t_L g463 ( 
.A(n_435),
.B(n_434),
.Y(n_463)
);

XNOR2xp5_ASAP7_75t_L g464 ( 
.A(n_434),
.B(n_426),
.Y(n_464)
);

XNOR2xp5_ASAP7_75t_L g480 ( 
.A(n_464),
.B(n_465),
.Y(n_480)
);

XNOR2xp5_ASAP7_75t_L g467 ( 
.A(n_448),
.B(n_426),
.Y(n_467)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_467),
.B(n_469),
.Y(n_476)
);

INVx1_ASAP7_75t_L g474 ( 
.A(n_468),
.Y(n_474)
);

MAJIxp5_ASAP7_75t_L g469 ( 
.A(n_439),
.B(n_404),
.C(n_400),
.Y(n_469)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_471),
.Y(n_482)
);

AOI22xp5_ASAP7_75t_L g472 ( 
.A1(n_447),
.A2(n_417),
.B1(n_413),
.B2(n_389),
.Y(n_472)
);

OAI22xp5_ASAP7_75t_SL g484 ( 
.A1(n_472),
.A2(n_445),
.B1(n_429),
.B2(n_444),
.Y(n_484)
);

OAI22xp5_ASAP7_75t_SL g473 ( 
.A1(n_444),
.A2(n_417),
.B1(n_406),
.B2(n_391),
.Y(n_473)
);

AOI22xp5_ASAP7_75t_L g486 ( 
.A1(n_473),
.A2(n_445),
.B1(n_432),
.B2(n_453),
.Y(n_486)
);

NAND2xp5_ASAP7_75t_L g477 ( 
.A(n_462),
.B(n_470),
.Y(n_477)
);

INVx1_ASAP7_75t_L g500 ( 
.A(n_477),
.Y(n_500)
);

FAx1_ASAP7_75t_L g478 ( 
.A(n_457),
.B(n_436),
.CI(n_430),
.CON(n_478),
.SN(n_478)
);

OAI21xp5_ASAP7_75t_L g494 ( 
.A1(n_478),
.A2(n_436),
.B(n_455),
.Y(n_494)
);

AOI22xp5_ASAP7_75t_L g481 ( 
.A1(n_473),
.A2(n_433),
.B1(n_438),
.B2(n_469),
.Y(n_481)
);

INVx1_ASAP7_75t_L g493 ( 
.A(n_481),
.Y(n_493)
);

MAJIxp5_ASAP7_75t_L g483 ( 
.A(n_456),
.B(n_450),
.C(n_429),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_SL g498 ( 
.A(n_483),
.B(n_485),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g490 ( 
.A1(n_484),
.A2(n_460),
.B1(n_458),
.B2(n_436),
.Y(n_490)
);

NOR2xp67_ASAP7_75t_SL g485 ( 
.A(n_467),
.B(n_430),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_L g495 ( 
.A(n_486),
.B(n_488),
.Y(n_495)
);

OAI22xp33_ASAP7_75t_L g488 ( 
.A1(n_461),
.A2(n_436),
.B1(n_451),
.B2(n_437),
.Y(n_488)
);

INVx1_ASAP7_75t_L g489 ( 
.A(n_459),
.Y(n_489)
);

NOR2xp33_ASAP7_75t_L g491 ( 
.A(n_489),
.B(n_456),
.Y(n_491)
);

INVx1_ASAP7_75t_L g505 ( 
.A(n_490),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_L g502 ( 
.A(n_491),
.B(n_492),
.Y(n_502)
);

NOR2xp33_ASAP7_75t_L g492 ( 
.A(n_483),
.B(n_466),
.Y(n_492)
);

NAND2xp5_ASAP7_75t_L g506 ( 
.A(n_494),
.B(n_496),
.Y(n_506)
);

NOR2xp33_ASAP7_75t_L g496 ( 
.A(n_482),
.B(n_391),
.Y(n_496)
);

XOR2xp5_ASAP7_75t_L g497 ( 
.A(n_480),
.B(n_454),
.Y(n_497)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_497),
.B(n_501),
.C(n_487),
.Y(n_503)
);

NOR2xp33_ASAP7_75t_L g499 ( 
.A(n_474),
.B(n_463),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_SL g504 ( 
.A(n_499),
.B(n_475),
.Y(n_504)
);

MAJIxp5_ASAP7_75t_L g501 ( 
.A(n_487),
.B(n_464),
.C(n_472),
.Y(n_501)
);

INVxp67_ASAP7_75t_L g510 ( 
.A(n_503),
.Y(n_510)
);

CKINVDCx14_ASAP7_75t_R g511 ( 
.A(n_504),
.Y(n_511)
);

AOI22xp5_ASAP7_75t_L g507 ( 
.A1(n_493),
.A2(n_479),
.B1(n_488),
.B2(n_476),
.Y(n_507)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_507),
.B(n_495),
.C(n_481),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_SL g508 ( 
.A(n_498),
.B(n_480),
.Y(n_508)
);

NOR2xp33_ASAP7_75t_SL g514 ( 
.A(n_508),
.B(n_501),
.Y(n_514)
);

OAI21xp5_ASAP7_75t_SL g509 ( 
.A1(n_490),
.A2(n_479),
.B(n_478),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_SL g512 ( 
.A(n_509),
.B(n_495),
.Y(n_512)
);

INVx1_ASAP7_75t_L g516 ( 
.A(n_512),
.Y(n_516)
);

INVxp67_ASAP7_75t_L g515 ( 
.A(n_513),
.Y(n_515)
);

NOR3xp33_ASAP7_75t_L g517 ( 
.A(n_514),
.B(n_502),
.C(n_503),
.Y(n_517)
);

NOR2xp33_ASAP7_75t_L g518 ( 
.A(n_517),
.B(n_510),
.Y(n_518)
);

NAND2xp5_ASAP7_75t_L g520 ( 
.A(n_518),
.B(n_519),
.Y(n_520)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_515),
.B(n_505),
.C(n_506),
.Y(n_519)
);

MAJIxp5_ASAP7_75t_L g521 ( 
.A(n_520),
.B(n_516),
.C(n_511),
.Y(n_521)
);

OAI321xp33_ASAP7_75t_L g522 ( 
.A1(n_521),
.A2(n_500),
.A3(n_493),
.B1(n_507),
.B2(n_478),
.C(n_494),
.Y(n_522)
);

AOI21xp5_ASAP7_75t_L g523 ( 
.A1(n_522),
.A2(n_497),
.B(n_455),
.Y(n_523)
);

OR2x2_ASAP7_75t_L g524 ( 
.A(n_523),
.B(n_383),
.Y(n_524)
);


endmodule