module real_jpeg_11670_n_17 (n_5, n_4, n_8, n_0, n_12, n_1, n_11, n_14, n_2, n_13, n_15, n_6, n_7, n_16, n_3, n_10, n_9, n_330, n_17);

input n_5;
input n_4;
input n_8;
input n_0;
input n_12;
input n_1;
input n_11;
input n_14;
input n_2;
input n_13;
input n_15;
input n_6;
input n_7;
input n_16;
input n_3;
input n_10;
input n_9;
input n_330;

output n_17;

wire n_37;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_300;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_47;
wire n_271;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_199;
wire n_95;
wire n_238;
wire n_67;
wire n_235;
wire n_107;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_123;
wire n_50;
wire n_186;
wire n_137;
wire n_72;
wire n_171;
wire n_151;
wire n_272;
wire n_198;
wire n_203;
wire n_23;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_80;
wire n_30;
wire n_149;
wire n_259;
wire n_57;
wire n_157;
wire n_84;
wire n_55;
wire n_58;
wire n_52;
wire n_230;
wire n_128;
wire n_202;
wire n_216;
wire n_127;
wire n_36;
wire n_102;
wire n_81;
wire n_101;
wire n_317;
wire n_108;
wire n_233;
wire n_73;
wire n_252;
wire n_310;
wire n_83;
wire n_78;
wire n_288;
wire n_221;
wire n_104;
wire n_153;
wire n_131;
wire n_322;
wire n_87;
wire n_40;
wire n_98;
wire n_200;
wire n_214;
wire n_113;
wire n_251;
wire n_139;
wire n_33;
wire n_175;
wire n_156;
wire n_66;
wire n_305;
wire n_62;
wire n_254;
wire n_250;
wire n_304;
wire n_77;
wire n_219;
wire n_122;
wire n_19;
wire n_262;
wire n_246;
wire n_21;
wire n_69;
wire n_31;
wire n_154;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_110;
wire n_195;
wire n_289;
wire n_117;
wire n_193;
wire n_20;
wire n_314;
wire n_278;
wire n_103;
wire n_232;
wire n_212;
wire n_284;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_213;
wire n_25;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_89;
wire n_49;
wire n_68;
wire n_146;
wire n_323;
wire n_166;
wire n_215;
wire n_286;
wire n_176;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_237;
wire n_173;
wire n_115;
wire n_184;
wire n_164;
wire n_140;
wire n_126;
wire n_120;
wire n_155;
wire n_319;
wire n_93;
wire n_242;
wire n_142;
wire n_76;
wire n_79;
wire n_282;
wire n_147;
wire n_265;
wire n_231;
wire n_44;
wire n_208;
wire n_162;
wire n_106;
wire n_172;
wire n_285;
wire n_112;
wire n_18;
wire n_145;
wire n_266;
wire n_109;
wire n_148;
wire n_196;
wire n_298;
wire n_152;
wire n_270;
wire n_159;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_90;
wire n_258;
wire n_150;
wire n_41;
wire n_74;
wire n_158;
wire n_204;
wire n_241;
wire n_111;
wire n_226;
wire n_125;
wire n_297;
wire n_75;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_119;
wire n_283;
wire n_181;
wire n_256;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_201;
wire n_260;
wire n_247;
wire n_249;
wire n_292;
wire n_64;
wire n_291;
wire n_236;
wire n_276;
wire n_287;
wire n_174;
wire n_255;
wire n_243;
wire n_299;
wire n_56;
wire n_293;
wire n_275;
wire n_227;
wire n_229;
wire n_141;
wire n_65;
wire n_188;
wire n_178;
wire n_189;
wire n_170;
wire n_28;
wire n_245;
wire n_45;
wire n_313;
wire n_42;
wire n_268;
wire n_94;
wire n_309;
wire n_294;
wire n_116;
wire n_143;
wire n_129;
wire n_135;
wire n_306;
wire n_218;
wire n_165;
wire n_303;
wire n_321;
wire n_100;
wire n_51;
wire n_205;
wire n_261;
wire n_86;
wire n_324;
wire n_70;
wire n_32;
wire n_228;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_191;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_133;
wire n_257;
wire n_210;
wire n_206;
wire n_85;
wire n_96;
wire n_308;

BUFx2_ASAP7_75t_L g32 ( 
.A(n_0),
.Y(n_32)
);

BUFx16f_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

BUFx12_ASAP7_75t_L g54 ( 
.A(n_2),
.Y(n_54)
);

INVx1_ASAP7_75t_L g144 ( 
.A(n_3),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g146 ( 
.A(n_3),
.B(n_53),
.Y(n_146)
);

NAND2xp5_ASAP7_75t_L g172 ( 
.A(n_3),
.B(n_173),
.Y(n_172)
);

O2A1O1Ixp33_ASAP7_75t_L g218 ( 
.A1(n_3),
.A2(n_57),
.B(n_74),
.C(n_219),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_L g232 ( 
.A1(n_3),
.A2(n_40),
.B1(n_41),
.B2(n_144),
.Y(n_232)
);

MAJIxp5_ASAP7_75t_L g234 ( 
.A(n_3),
.B(n_30),
.C(n_44),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_3),
.B(n_75),
.Y(n_238)
);

OAI21xp33_ASAP7_75t_L g258 ( 
.A1(n_3),
.A2(n_110),
.B(n_244),
.Y(n_258)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_3),
.A2(n_57),
.B1(n_58),
.B2(n_144),
.Y(n_270)
);

BUFx12f_ASAP7_75t_L g40 ( 
.A(n_4),
.Y(n_40)
);

AOI22xp33_ASAP7_75t_SL g149 ( 
.A1(n_5),
.A2(n_57),
.B1(n_58),
.B2(n_150),
.Y(n_149)
);

CKINVDCx20_ASAP7_75t_R g150 ( 
.A(n_5),
.Y(n_150)
);

AOI22xp33_ASAP7_75t_SL g190 ( 
.A1(n_5),
.A2(n_53),
.B1(n_54),
.B2(n_150),
.Y(n_190)
);

AOI22xp5_ASAP7_75t_SL g241 ( 
.A1(n_5),
.A2(n_40),
.B1(n_41),
.B2(n_150),
.Y(n_241)
);

AOI22xp33_ASAP7_75t_L g249 ( 
.A1(n_5),
.A2(n_29),
.B1(n_30),
.B2(n_150),
.Y(n_249)
);

AOI22xp33_ASAP7_75t_L g66 ( 
.A1(n_6),
.A2(n_53),
.B1(n_54),
.B2(n_67),
.Y(n_66)
);

CKINVDCx20_ASAP7_75t_R g67 ( 
.A(n_6),
.Y(n_67)
);

OAI22xp5_ASAP7_75t_SL g156 ( 
.A1(n_6),
.A2(n_40),
.B1(n_41),
.B2(n_67),
.Y(n_156)
);

OAI22xp33_ASAP7_75t_SL g170 ( 
.A1(n_6),
.A2(n_57),
.B1(n_58),
.B2(n_67),
.Y(n_170)
);

OAI22xp5_ASAP7_75t_SL g222 ( 
.A1(n_6),
.A2(n_29),
.B1(n_30),
.B2(n_67),
.Y(n_222)
);

OAI22xp5_ASAP7_75t_L g38 ( 
.A1(n_7),
.A2(n_39),
.B1(n_40),
.B2(n_41),
.Y(n_38)
);

INVx1_ASAP7_75t_L g39 ( 
.A(n_7),
.Y(n_39)
);

AOI22xp33_ASAP7_75t_SL g79 ( 
.A1(n_7),
.A2(n_39),
.B1(n_57),
.B2(n_58),
.Y(n_79)
);

AOI22xp33_ASAP7_75t_SL g128 ( 
.A1(n_7),
.A2(n_39),
.B1(n_53),
.B2(n_54),
.Y(n_128)
);

OAI22xp33_ASAP7_75t_SL g166 ( 
.A1(n_7),
.A2(n_29),
.B1(n_30),
.B2(n_39),
.Y(n_166)
);

BUFx12f_ASAP7_75t_L g59 ( 
.A(n_8),
.Y(n_59)
);

AOI22xp33_ASAP7_75t_SL g76 ( 
.A1(n_9),
.A2(n_57),
.B1(n_58),
.B2(n_77),
.Y(n_76)
);

CKINVDCx16_ASAP7_75t_R g77 ( 
.A(n_9),
.Y(n_77)
);

AOI22xp33_ASAP7_75t_SL g95 ( 
.A1(n_9),
.A2(n_53),
.B1(n_54),
.B2(n_77),
.Y(n_95)
);

OAI22xp5_ASAP7_75t_L g114 ( 
.A1(n_9),
.A2(n_40),
.B1(n_41),
.B2(n_77),
.Y(n_114)
);

AOI22xp5_ASAP7_75t_SL g164 ( 
.A1(n_9),
.A2(n_29),
.B1(n_30),
.B2(n_77),
.Y(n_164)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_10),
.Y(n_73)
);

AOI22xp5_ASAP7_75t_L g56 ( 
.A1(n_11),
.A2(n_57),
.B1(n_58),
.B2(n_60),
.Y(n_56)
);

INVx4_ASAP7_75t_L g60 ( 
.A(n_11),
.Y(n_60)
);

OAI22xp5_ASAP7_75t_SL g64 ( 
.A1(n_11),
.A2(n_53),
.B1(n_54),
.B2(n_60),
.Y(n_64)
);

NAND2xp33_ASAP7_75t_SL g161 ( 
.A(n_11),
.B(n_58),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_SL g34 ( 
.A1(n_12),
.A2(n_29),
.B1(n_30),
.B2(n_35),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_12),
.Y(n_35)
);

AOI22xp33_ASAP7_75t_SL g82 ( 
.A1(n_12),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_82)
);

AOI22xp33_ASAP7_75t_SL g132 ( 
.A1(n_12),
.A2(n_35),
.B1(n_57),
.B2(n_58),
.Y(n_132)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_12),
.A2(n_35),
.B1(n_53),
.B2(n_54),
.Y(n_323)
);

AOI22xp33_ASAP7_75t_SL g118 ( 
.A1(n_13),
.A2(n_53),
.B1(n_54),
.B2(n_119),
.Y(n_118)
);

CKINVDCx20_ASAP7_75t_R g119 ( 
.A(n_13),
.Y(n_119)
);

AOI22xp33_ASAP7_75t_SL g151 ( 
.A1(n_13),
.A2(n_57),
.B1(n_58),
.B2(n_119),
.Y(n_151)
);

OAI22xp5_ASAP7_75t_L g214 ( 
.A1(n_13),
.A2(n_40),
.B1(n_41),
.B2(n_119),
.Y(n_214)
);

AOI22xp5_ASAP7_75t_SL g243 ( 
.A1(n_13),
.A2(n_29),
.B1(n_30),
.B2(n_119),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g52 ( 
.A1(n_14),
.A2(n_53),
.B1(n_54),
.B2(n_55),
.Y(n_52)
);

CKINVDCx20_ASAP7_75t_R g55 ( 
.A(n_14),
.Y(n_55)
);

AOI22xp33_ASAP7_75t_SL g116 ( 
.A1(n_14),
.A2(n_55),
.B1(n_57),
.B2(n_58),
.Y(n_116)
);

OAI22xp5_ASAP7_75t_L g154 ( 
.A1(n_14),
.A2(n_40),
.B1(n_41),
.B2(n_55),
.Y(n_154)
);

AOI22xp33_ASAP7_75t_SL g175 ( 
.A1(n_14),
.A2(n_29),
.B1(n_30),
.B2(n_55),
.Y(n_175)
);

AOI22xp33_ASAP7_75t_SL g48 ( 
.A1(n_15),
.A2(n_40),
.B1(n_41),
.B2(n_49),
.Y(n_48)
);

CKINVDCx16_ASAP7_75t_R g49 ( 
.A(n_15),
.Y(n_49)
);

AOI22xp5_ASAP7_75t_L g88 ( 
.A1(n_15),
.A2(n_49),
.B1(n_57),
.B2(n_58),
.Y(n_88)
);

OAI22xp5_ASAP7_75t_L g109 ( 
.A1(n_15),
.A2(n_29),
.B1(n_30),
.B2(n_49),
.Y(n_109)
);

OAI22xp5_ASAP7_75t_L g314 ( 
.A1(n_15),
.A2(n_49),
.B1(n_53),
.B2(n_54),
.Y(n_314)
);

INVx11_ASAP7_75t_L g31 ( 
.A(n_16),
.Y(n_31)
);

XOR2xp5_ASAP7_75t_L g17 ( 
.A(n_18),
.B(n_320),
.Y(n_17)
);

AOI21xp5_ASAP7_75t_L g18 ( 
.A1(n_19),
.A2(n_307),
.B(n_319),
.Y(n_18)
);

AO21x1_ASAP7_75t_L g19 ( 
.A1(n_20),
.A2(n_135),
.B(n_304),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_122),
.Y(n_20)
);

NOR2xp33_ASAP7_75t_L g21 ( 
.A(n_22),
.B(n_97),
.Y(n_21)
);

NAND2xp5_ASAP7_75t_L g305 ( 
.A(n_22),
.B(n_97),
.Y(n_305)
);

BUFx24_ASAP7_75t_SL g328 ( 
.A(n_22),
.Y(n_328)
);

FAx1_ASAP7_75t_L g22 ( 
.A(n_23),
.B(n_68),
.CI(n_83),
.CON(n_22),
.SN(n_22)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_23),
.B(n_68),
.C(n_83),
.Y(n_134)
);

OAI21xp5_ASAP7_75t_L g23 ( 
.A1(n_24),
.A2(n_27),
.B(n_51),
.Y(n_23)
);

OAI22xp5_ASAP7_75t_SL g99 ( 
.A1(n_24),
.A2(n_25),
.B1(n_100),
.B2(n_101),
.Y(n_99)
);

INVx1_ASAP7_75t_L g24 ( 
.A(n_25),
.Y(n_24)
);

NAND2xp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g101 ( 
.A1(n_26),
.A2(n_27),
.B1(n_51),
.B2(n_102),
.Y(n_101)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_26),
.A2(n_27),
.B1(n_36),
.B2(n_37),
.Y(n_291)
);

CKINVDCx20_ASAP7_75t_R g26 ( 
.A(n_27),
.Y(n_26)
);

OAI21xp5_ASAP7_75t_SL g27 ( 
.A1(n_28),
.A2(n_32),
.B(n_33),
.Y(n_27)
);

INVx1_ASAP7_75t_L g110 ( 
.A(n_28),
.Y(n_110)
);

AOI22xp5_ASAP7_75t_L g180 ( 
.A1(n_28),
.A2(n_32),
.B1(n_109),
.B2(n_166),
.Y(n_180)
);

NAND2xp5_ASAP7_75t_L g221 ( 
.A(n_28),
.B(n_222),
.Y(n_221)
);

AOI22xp5_ASAP7_75t_SL g247 ( 
.A1(n_28),
.A2(n_32),
.B1(n_248),
.B2(n_250),
.Y(n_247)
);

NOR2xp33_ASAP7_75t_SL g28 ( 
.A(n_29),
.B(n_32),
.Y(n_28)
);

OA22x2_ASAP7_75t_L g46 ( 
.A1(n_29),
.A2(n_30),
.B1(n_44),
.B2(n_45),
.Y(n_46)
);

NOR2xp33_ASAP7_75t_SL g259 ( 
.A(n_29),
.B(n_260),
.Y(n_259)
);

INVx5_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

CKINVDCx20_ASAP7_75t_R g111 ( 
.A(n_32),
.Y(n_111)
);

NAND2xp5_ASAP7_75t_SL g244 ( 
.A(n_32),
.B(n_222),
.Y(n_244)
);

INVxp67_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

OAI22xp5_ASAP7_75t_SL g107 ( 
.A1(n_34),
.A2(n_108),
.B1(n_110),
.B2(n_111),
.Y(n_107)
);

CKINVDCx20_ASAP7_75t_R g36 ( 
.A(n_37),
.Y(n_36)
);

AOI22xp5_ASAP7_75t_L g37 ( 
.A1(n_38),
.A2(n_42),
.B1(n_47),
.B2(n_50),
.Y(n_37)
);

AOI22xp5_ASAP7_75t_L g113 ( 
.A1(n_38),
.A2(n_42),
.B1(n_50),
.B2(n_114),
.Y(n_113)
);

INVx4_ASAP7_75t_SL g41 ( 
.A(n_40),
.Y(n_41)
);

OAI22xp33_ASAP7_75t_L g43 ( 
.A1(n_40),
.A2(n_41),
.B1(n_44),
.B2(n_45),
.Y(n_43)
);

AO22x1_ASAP7_75t_SL g75 ( 
.A1(n_40),
.A2(n_41),
.B1(n_73),
.B2(n_74),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_SL g233 ( 
.A(n_40),
.B(n_234),
.Y(n_233)
);

OAI21xp33_ASAP7_75t_L g219 ( 
.A1(n_41),
.A2(n_73),
.B(n_144),
.Y(n_219)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_42),
.Y(n_81)
);

OAI21xp5_ASAP7_75t_L g90 ( 
.A1(n_42),
.A2(n_50),
.B(n_91),
.Y(n_90)
);

NAND2xp5_ASAP7_75t_SL g155 ( 
.A(n_42),
.B(n_156),
.Y(n_155)
);

AOI22xp5_ASAP7_75t_L g181 ( 
.A1(n_42),
.A2(n_50),
.B1(n_114),
.B2(n_154),
.Y(n_181)
);

AOI22xp5_ASAP7_75t_L g271 ( 
.A1(n_42),
.A2(n_50),
.B1(n_214),
.B2(n_272),
.Y(n_271)
);

AND2x2_ASAP7_75t_L g42 ( 
.A(n_43),
.B(n_46),
.Y(n_42)
);

INVx6_ASAP7_75t_L g45 ( 
.A(n_44),
.Y(n_45)
);

INVx1_ASAP7_75t_L g50 ( 
.A(n_46),
.Y(n_50)
);

OAI22xp5_ASAP7_75t_SL g80 ( 
.A1(n_46),
.A2(n_48),
.B1(n_81),
.B2(n_82),
.Y(n_80)
);

OAI21xp5_ASAP7_75t_L g152 ( 
.A1(n_46),
.A2(n_153),
.B(n_155),
.Y(n_152)
);

OAI21xp5_ASAP7_75t_L g240 ( 
.A1(n_46),
.A2(n_155),
.B(n_241),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_SL g255 ( 
.A(n_46),
.B(n_144),
.Y(n_255)
);

INVxp67_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

NAND2xp5_ASAP7_75t_L g215 ( 
.A(n_50),
.B(n_156),
.Y(n_215)
);

INVx1_ASAP7_75t_L g102 ( 
.A(n_51),
.Y(n_102)
);

OAI21xp5_ASAP7_75t_L g51 ( 
.A1(n_52),
.A2(n_56),
.B(n_61),
.Y(n_51)
);

OAI22xp5_ASAP7_75t_L g94 ( 
.A1(n_52),
.A2(n_56),
.B1(n_63),
.B2(n_95),
.Y(n_94)
);

INVx4_ASAP7_75t_L g53 ( 
.A(n_54),
.Y(n_53)
);

O2A1O1Ixp33_ASAP7_75t_L g143 ( 
.A1(n_54),
.A2(n_63),
.B(n_144),
.C(n_145),
.Y(n_143)
);

AOI32xp33_ASAP7_75t_L g160 ( 
.A1(n_54),
.A2(n_57),
.A3(n_60),
.B1(n_146),
.B2(n_161),
.Y(n_160)
);

NAND2xp5_ASAP7_75t_SL g63 ( 
.A(n_56),
.B(n_64),
.Y(n_63)
);

NOR2xp33_ASAP7_75t_L g121 ( 
.A(n_56),
.B(n_66),
.Y(n_121)
);

OAI22xp5_ASAP7_75t_SL g127 ( 
.A1(n_56),
.A2(n_63),
.B1(n_95),
.B2(n_128),
.Y(n_127)
);

INVx1_ASAP7_75t_L g173 ( 
.A(n_56),
.Y(n_173)
);

OAI21xp5_ASAP7_75t_L g189 ( 
.A1(n_56),
.A2(n_61),
.B(n_190),
.Y(n_189)
);

OAI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_56),
.A2(n_63),
.B1(n_118),
.B2(n_190),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_L g72 ( 
.A1(n_57),
.A2(n_58),
.B1(n_73),
.B2(n_74),
.Y(n_72)
);

INVx8_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

BUFx12f_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

NAND2xp5_ASAP7_75t_SL g61 ( 
.A(n_62),
.B(n_65),
.Y(n_61)
);

AOI22xp5_ASAP7_75t_L g312 ( 
.A1(n_62),
.A2(n_173),
.B1(n_313),
.B2(n_314),
.Y(n_312)
);

AOI22xp5_ASAP7_75t_L g322 ( 
.A1(n_62),
.A2(n_173),
.B1(n_314),
.B2(n_323),
.Y(n_322)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

OAI21xp5_ASAP7_75t_L g117 ( 
.A1(n_63),
.A2(n_118),
.B(n_120),
.Y(n_117)
);

INVxp67_ASAP7_75t_L g65 ( 
.A(n_66),
.Y(n_65)
);

AOI21xp5_ASAP7_75t_L g103 ( 
.A1(n_68),
.A2(n_69),
.B(n_80),
.Y(n_103)
);

NOR2xp33_ASAP7_75t_L g68 ( 
.A(n_69),
.B(n_80),
.Y(n_68)
);

OAI22xp5_ASAP7_75t_SL g69 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_79),
.Y(n_69)
);

OAI22xp5_ASAP7_75t_SL g115 ( 
.A1(n_70),
.A2(n_76),
.B1(n_78),
.B2(n_116),
.Y(n_115)
);

OAI22xp5_ASAP7_75t_SL g131 ( 
.A1(n_70),
.A2(n_78),
.B1(n_88),
.B2(n_132),
.Y(n_131)
);

OAI22xp5_ASAP7_75t_SL g148 ( 
.A1(n_70),
.A2(n_78),
.B1(n_149),
.B2(n_151),
.Y(n_148)
);

OAI21xp5_ASAP7_75t_L g187 ( 
.A1(n_70),
.A2(n_151),
.B(n_188),
.Y(n_187)
);

OAI21xp5_ASAP7_75t_SL g269 ( 
.A1(n_70),
.A2(n_188),
.B(n_270),
.Y(n_269)
);

INVx1_ASAP7_75t_L g70 ( 
.A(n_71),
.Y(n_70)
);

AOI22xp5_ASAP7_75t_L g85 ( 
.A1(n_71),
.A2(n_75),
.B1(n_86),
.B2(n_87),
.Y(n_85)
);

NAND2xp5_ASAP7_75t_L g169 ( 
.A(n_71),
.B(n_170),
.Y(n_169)
);

OAI21xp5_ASAP7_75t_SL g310 ( 
.A1(n_71),
.A2(n_75),
.B(n_311),
.Y(n_310)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_72),
.B(n_75),
.Y(n_71)
);

INVx8_ASAP7_75t_L g74 ( 
.A(n_73),
.Y(n_74)
);

INVx1_ASAP7_75t_L g78 ( 
.A(n_75),
.Y(n_78)
);

NAND2xp5_ASAP7_75t_L g188 ( 
.A(n_75),
.B(n_170),
.Y(n_188)
);

OAI21xp5_ASAP7_75t_SL g168 ( 
.A1(n_78),
.A2(n_149),
.B(n_169),
.Y(n_168)
);

OAI21xp5_ASAP7_75t_SL g202 ( 
.A1(n_78),
.A2(n_116),
.B(n_169),
.Y(n_202)
);

INVxp67_ASAP7_75t_L g86 ( 
.A(n_79),
.Y(n_86)
);

OAI21xp5_ASAP7_75t_SL g212 ( 
.A1(n_81),
.A2(n_213),
.B(n_215),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g231 ( 
.A1(n_81),
.A2(n_215),
.B(n_232),
.Y(n_231)
);

CKINVDCx14_ASAP7_75t_R g91 ( 
.A(n_82),
.Y(n_91)
);

AOI22xp5_ASAP7_75t_L g83 ( 
.A1(n_84),
.A2(n_93),
.B1(n_94),
.B2(n_96),
.Y(n_83)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_84),
.Y(n_96)
);

AOI22xp5_ASAP7_75t_L g84 ( 
.A1(n_85),
.A2(n_89),
.B1(n_90),
.B2(n_92),
.Y(n_84)
);

CKINVDCx16_ASAP7_75t_R g92 ( 
.A(n_85),
.Y(n_92)
);

MAJIxp5_ASAP7_75t_SL g133 ( 
.A(n_85),
.B(n_90),
.C(n_94),
.Y(n_133)
);

INVx1_ASAP7_75t_L g87 ( 
.A(n_88),
.Y(n_87)
);

AOI22xp5_ASAP7_75t_L g129 ( 
.A1(n_89),
.A2(n_90),
.B1(n_130),
.B2(n_131),
.Y(n_129)
);

CKINVDCx16_ASAP7_75t_R g89 ( 
.A(n_90),
.Y(n_89)
);

MAJIxp5_ASAP7_75t_L g317 ( 
.A(n_90),
.B(n_127),
.C(n_131),
.Y(n_317)
);

AOI22xp5_ASAP7_75t_L g124 ( 
.A1(n_93),
.A2(n_94),
.B1(n_125),
.B2(n_126),
.Y(n_124)
);

CKINVDCx16_ASAP7_75t_R g93 ( 
.A(n_94),
.Y(n_93)
);

MAJIxp5_ASAP7_75t_L g318 ( 
.A(n_94),
.B(n_126),
.C(n_133),
.Y(n_318)
);

MAJIxp5_ASAP7_75t_L g97 ( 
.A(n_98),
.B(n_103),
.C(n_104),
.Y(n_97)
);

AOI22xp5_ASAP7_75t_L g301 ( 
.A1(n_98),
.A2(n_99),
.B1(n_103),
.B2(n_302),
.Y(n_301)
);

INVx1_ASAP7_75t_L g98 ( 
.A(n_99),
.Y(n_98)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx1_ASAP7_75t_L g302 ( 
.A(n_103),
.Y(n_302)
);

XOR2xp5_ASAP7_75t_L g300 ( 
.A(n_104),
.B(n_301),
.Y(n_300)
);

MAJIxp5_ASAP7_75t_L g104 ( 
.A(n_105),
.B(n_115),
.C(n_117),
.Y(n_104)
);

OAI22xp5_ASAP7_75t_SL g293 ( 
.A1(n_105),
.A2(n_106),
.B1(n_294),
.B2(n_295),
.Y(n_293)
);

INVx1_ASAP7_75t_L g105 ( 
.A(n_106),
.Y(n_105)
);

NAND2xp5_ASAP7_75t_L g106 ( 
.A(n_107),
.B(n_112),
.Y(n_106)
);

OAI22xp5_ASAP7_75t_SL g197 ( 
.A1(n_107),
.A2(n_112),
.B1(n_113),
.B2(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

INVxp67_ASAP7_75t_L g108 ( 
.A(n_109),
.Y(n_108)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_110),
.A2(n_111),
.B1(n_164),
.B2(n_165),
.Y(n_163)
);

OAI22xp5_ASAP7_75t_SL g174 ( 
.A1(n_110),
.A2(n_111),
.B1(n_164),
.B2(n_175),
.Y(n_174)
);

OAI21xp5_ASAP7_75t_L g242 ( 
.A1(n_110),
.A2(n_243),
.B(n_244),
.Y(n_242)
);

OAI21xp5_ASAP7_75t_L g220 ( 
.A1(n_111),
.A2(n_175),
.B(n_221),
.Y(n_220)
);

OAI21xp5_ASAP7_75t_SL g256 ( 
.A1(n_111),
.A2(n_221),
.B(n_249),
.Y(n_256)
);

NOR2xp33_ASAP7_75t_L g260 ( 
.A(n_111),
.B(n_144),
.Y(n_260)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_113),
.Y(n_112)
);

XNOR2xp5_ASAP7_75t_SL g295 ( 
.A(n_115),
.B(n_117),
.Y(n_295)
);

INVxp67_ASAP7_75t_L g120 ( 
.A(n_121),
.Y(n_120)
);

NOR2xp33_ASAP7_75t_SL g142 ( 
.A(n_121),
.B(n_143),
.Y(n_142)
);

OAI21xp33_ASAP7_75t_L g304 ( 
.A1(n_122),
.A2(n_305),
.B(n_306),
.Y(n_304)
);

NOR2xp33_ASAP7_75t_SL g122 ( 
.A(n_123),
.B(n_134),
.Y(n_122)
);

NAND2xp5_ASAP7_75t_L g306 ( 
.A(n_123),
.B(n_134),
.Y(n_306)
);

XNOR2xp5_ASAP7_75t_L g123 ( 
.A(n_124),
.B(n_133),
.Y(n_123)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_126),
.Y(n_125)
);

XNOR2xp5_ASAP7_75t_L g126 ( 
.A(n_127),
.B(n_129),
.Y(n_126)
);

CKINVDCx20_ASAP7_75t_R g313 ( 
.A(n_128),
.Y(n_313)
);

INVx1_ASAP7_75t_L g130 ( 
.A(n_131),
.Y(n_130)
);

CKINVDCx16_ASAP7_75t_R g311 ( 
.A(n_132),
.Y(n_311)
);

OAI21xp5_ASAP7_75t_SL g135 ( 
.A1(n_136),
.A2(n_298),
.B(n_303),
.Y(n_135)
);

AOI21xp5_ASAP7_75t_SL g136 ( 
.A1(n_137),
.A2(n_286),
.B(n_297),
.Y(n_136)
);

OAI321xp33_ASAP7_75t_L g137 ( 
.A1(n_138),
.A2(n_193),
.A3(n_205),
.B1(n_284),
.B2(n_285),
.C(n_330),
.Y(n_137)
);

NOR2xp33_ASAP7_75t_L g138 ( 
.A(n_139),
.B(n_176),
.Y(n_138)
);

NAND2xp5_ASAP7_75t_SL g284 ( 
.A(n_139),
.B(n_176),
.Y(n_284)
);

MAJIxp5_ASAP7_75t_L g139 ( 
.A(n_140),
.B(n_158),
.C(n_167),
.Y(n_139)
);

XNOR2xp5_ASAP7_75t_L g223 ( 
.A(n_140),
.B(n_224),
.Y(n_223)
);

AOI22xp5_ASAP7_75t_L g140 ( 
.A1(n_141),
.A2(n_142),
.B1(n_147),
.B2(n_157),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g182 ( 
.A(n_141),
.B(n_148),
.C(n_152),
.Y(n_182)
);

INVx1_ASAP7_75t_L g141 ( 
.A(n_142),
.Y(n_141)
);

INVxp67_ASAP7_75t_L g145 ( 
.A(n_146),
.Y(n_145)
);

INVx1_ASAP7_75t_L g157 ( 
.A(n_147),
.Y(n_157)
);

XNOR2xp5_ASAP7_75t_SL g147 ( 
.A(n_148),
.B(n_152),
.Y(n_147)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_154),
.Y(n_153)
);

XNOR2xp5_ASAP7_75t_L g224 ( 
.A(n_158),
.B(n_167),
.Y(n_224)
);

AOI22xp5_ASAP7_75t_L g158 ( 
.A1(n_159),
.A2(n_160),
.B1(n_162),
.B2(n_163),
.Y(n_158)
);

NAND2xp5_ASAP7_75t_L g192 ( 
.A(n_159),
.B(n_163),
.Y(n_192)
);

INVx1_ASAP7_75t_L g159 ( 
.A(n_160),
.Y(n_159)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_163),
.Y(n_162)
);

INVxp67_ASAP7_75t_L g165 ( 
.A(n_166),
.Y(n_165)
);

MAJIxp5_ASAP7_75t_L g167 ( 
.A(n_168),
.B(n_171),
.C(n_174),
.Y(n_167)
);

XOR2xp5_ASAP7_75t_L g209 ( 
.A(n_168),
.B(n_210),
.Y(n_209)
);

AOI22xp5_ASAP7_75t_L g210 ( 
.A1(n_171),
.A2(n_172),
.B1(n_174),
.B2(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g171 ( 
.A(n_172),
.Y(n_171)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_174),
.Y(n_211)
);

OAI22xp5_ASAP7_75t_SL g176 ( 
.A1(n_177),
.A2(n_178),
.B1(n_183),
.B2(n_184),
.Y(n_176)
);

INVx1_ASAP7_75t_L g177 ( 
.A(n_178),
.Y(n_177)
);

XNOR2xp5_ASAP7_75t_SL g178 ( 
.A(n_179),
.B(n_182),
.Y(n_178)
);

MAJIxp5_ASAP7_75t_L g194 ( 
.A(n_179),
.B(n_182),
.C(n_183),
.Y(n_194)
);

XNOR2xp5_ASAP7_75t_L g179 ( 
.A(n_180),
.B(n_181),
.Y(n_179)
);

NOR2xp33_ASAP7_75t_L g203 ( 
.A(n_180),
.B(n_181),
.Y(n_203)
);

INVx1_ASAP7_75t_L g183 ( 
.A(n_184),
.Y(n_183)
);

XOR2xp5_ASAP7_75t_L g184 ( 
.A(n_185),
.B(n_192),
.Y(n_184)
);

AOI22xp5_ASAP7_75t_L g185 ( 
.A1(n_186),
.A2(n_187),
.B1(n_189),
.B2(n_191),
.Y(n_185)
);

MAJIxp5_ASAP7_75t_L g204 ( 
.A(n_186),
.B(n_191),
.C(n_192),
.Y(n_204)
);

INVx1_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_189),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g193 ( 
.A(n_194),
.B(n_195),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g285 ( 
.A(n_194),
.B(n_195),
.Y(n_285)
);

XNOR2xp5_ASAP7_75t_L g195 ( 
.A(n_196),
.B(n_204),
.Y(n_195)
);

XNOR2xp5_ASAP7_75t_L g196 ( 
.A(n_197),
.B(n_199),
.Y(n_196)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_197),
.B(n_199),
.C(n_204),
.Y(n_296)
);

XNOR2xp5_ASAP7_75t_SL g199 ( 
.A(n_200),
.B(n_203),
.Y(n_199)
);

XNOR2xp5_ASAP7_75t_L g200 ( 
.A(n_201),
.B(n_202),
.Y(n_200)
);

MAJIxp5_ASAP7_75t_L g288 ( 
.A(n_201),
.B(n_202),
.C(n_203),
.Y(n_288)
);

AOI21xp5_ASAP7_75t_SL g205 ( 
.A1(n_206),
.A2(n_225),
.B(n_283),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g206 ( 
.A(n_207),
.B(n_223),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_SL g283 ( 
.A(n_207),
.B(n_223),
.Y(n_283)
);

MAJIxp5_ASAP7_75t_L g207 ( 
.A(n_208),
.B(n_212),
.C(n_216),
.Y(n_207)
);

OAI22xp5_ASAP7_75t_SL g278 ( 
.A1(n_208),
.A2(n_209),
.B1(n_279),
.B2(n_280),
.Y(n_278)
);

INVx1_ASAP7_75t_L g208 ( 
.A(n_209),
.Y(n_208)
);

OAI22xp5_ASAP7_75t_SL g280 ( 
.A1(n_212),
.A2(n_216),
.B1(n_217),
.B2(n_281),
.Y(n_280)
);

INVx1_ASAP7_75t_L g281 ( 
.A(n_212),
.Y(n_281)
);

INVxp67_ASAP7_75t_L g213 ( 
.A(n_214),
.Y(n_213)
);

INVx1_ASAP7_75t_L g216 ( 
.A(n_217),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_220),
.Y(n_217)
);

XNOR2xp5_ASAP7_75t_SL g267 ( 
.A(n_218),
.B(n_220),
.Y(n_267)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_226),
.A2(n_276),
.B(n_282),
.Y(n_225)
);

AOI21xp5_ASAP7_75t_L g226 ( 
.A1(n_227),
.A2(n_264),
.B(n_275),
.Y(n_226)
);

OAI21xp5_ASAP7_75t_SL g227 ( 
.A1(n_228),
.A2(n_245),
.B(n_263),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_229),
.B(n_235),
.Y(n_228)
);

NAND2xp5_ASAP7_75t_SL g263 ( 
.A(n_229),
.B(n_235),
.Y(n_263)
);

NOR2xp33_ASAP7_75t_SL g229 ( 
.A(n_230),
.B(n_233),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_SL g251 ( 
.A1(n_230),
.A2(n_231),
.B1(n_233),
.B2(n_252),
.Y(n_251)
);

INVx1_ASAP7_75t_L g230 ( 
.A(n_231),
.Y(n_230)
);

CKINVDCx20_ASAP7_75t_R g252 ( 
.A(n_233),
.Y(n_252)
);

XNOR2xp5_ASAP7_75t_L g235 ( 
.A(n_236),
.B(n_242),
.Y(n_235)
);

AOI22xp5_ASAP7_75t_L g236 ( 
.A1(n_237),
.A2(n_238),
.B1(n_239),
.B2(n_240),
.Y(n_236)
);

MAJIxp5_ASAP7_75t_L g265 ( 
.A(n_237),
.B(n_240),
.C(n_242),
.Y(n_265)
);

CKINVDCx14_ASAP7_75t_R g237 ( 
.A(n_238),
.Y(n_237)
);

INVx1_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

CKINVDCx14_ASAP7_75t_R g272 ( 
.A(n_241),
.Y(n_272)
);

INVxp67_ASAP7_75t_L g250 ( 
.A(n_243),
.Y(n_250)
);

AOI21xp5_ASAP7_75t_L g245 ( 
.A1(n_246),
.A2(n_253),
.B(n_262),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_L g246 ( 
.A(n_247),
.B(n_251),
.Y(n_246)
);

NOR2xp33_ASAP7_75t_SL g262 ( 
.A(n_247),
.B(n_251),
.Y(n_262)
);

INVxp67_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

OAI21xp5_ASAP7_75t_SL g253 ( 
.A1(n_254),
.A2(n_257),
.B(n_261),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g254 ( 
.A(n_255),
.B(n_256),
.Y(n_254)
);

NAND2xp5_ASAP7_75t_SL g261 ( 
.A(n_255),
.B(n_256),
.Y(n_261)
);

NAND2xp5_ASAP7_75t_SL g257 ( 
.A(n_258),
.B(n_259),
.Y(n_257)
);

NAND2xp5_ASAP7_75t_L g264 ( 
.A(n_265),
.B(n_266),
.Y(n_264)
);

NOR2xp33_ASAP7_75t_SL g275 ( 
.A(n_265),
.B(n_266),
.Y(n_275)
);

XNOR2xp5_ASAP7_75t_L g266 ( 
.A(n_267),
.B(n_268),
.Y(n_266)
);

MAJIxp5_ASAP7_75t_L g277 ( 
.A(n_267),
.B(n_271),
.C(n_274),
.Y(n_277)
);

AOI22xp5_ASAP7_75t_L g268 ( 
.A1(n_269),
.A2(n_271),
.B1(n_273),
.B2(n_274),
.Y(n_268)
);

INVx1_ASAP7_75t_L g274 ( 
.A(n_269),
.Y(n_274)
);

INVx1_ASAP7_75t_L g273 ( 
.A(n_271),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_277),
.B(n_278),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_SL g282 ( 
.A(n_277),
.B(n_278),
.Y(n_282)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_SL g286 ( 
.A(n_287),
.B(n_296),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g297 ( 
.A(n_287),
.B(n_296),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g287 ( 
.A(n_288),
.B(n_289),
.Y(n_287)
);

MAJIxp5_ASAP7_75t_L g299 ( 
.A(n_288),
.B(n_291),
.C(n_292),
.Y(n_299)
);

AOI22xp5_ASAP7_75t_L g289 ( 
.A1(n_290),
.A2(n_291),
.B1(n_292),
.B2(n_293),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_291),
.Y(n_290)
);

INVx1_ASAP7_75t_L g292 ( 
.A(n_293),
.Y(n_292)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_295),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g298 ( 
.A(n_299),
.B(n_300),
.Y(n_298)
);

NAND2xp5_ASAP7_75t_L g303 ( 
.A(n_299),
.B(n_300),
.Y(n_303)
);

NAND2xp5_ASAP7_75t_L g307 ( 
.A(n_308),
.B(n_318),
.Y(n_307)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_308),
.B(n_318),
.Y(n_319)
);

XNOR2xp5_ASAP7_75t_L g308 ( 
.A(n_309),
.B(n_317),
.Y(n_308)
);

AOI22xp5_ASAP7_75t_L g309 ( 
.A1(n_310),
.A2(n_312),
.B1(n_315),
.B2(n_316),
.Y(n_309)
);

CKINVDCx20_ASAP7_75t_R g315 ( 
.A(n_310),
.Y(n_315)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_312),
.Y(n_316)
);

MAJIxp5_ASAP7_75t_L g324 ( 
.A(n_312),
.B(n_315),
.C(n_317),
.Y(n_324)
);

NOR2xp33_ASAP7_75t_L g320 ( 
.A(n_321),
.B(n_325),
.Y(n_320)
);

NOR2xp33_ASAP7_75t_L g321 ( 
.A(n_322),
.B(n_324),
.Y(n_321)
);

CKINVDCx20_ASAP7_75t_R g326 ( 
.A(n_322),
.Y(n_326)
);

CKINVDCx16_ASAP7_75t_R g327 ( 
.A(n_324),
.Y(n_327)
);

NOR2xp33_ASAP7_75t_L g325 ( 
.A(n_326),
.B(n_327),
.Y(n_325)
);


endmodule