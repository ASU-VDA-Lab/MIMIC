module real_jpeg_18559_n_19 (n_17, n_8, n_0, n_2, n_10, n_9, n_12, n_6, n_11, n_14, n_7, n_18, n_3, n_5, n_4, n_1, n_16, n_15, n_13, n_19);

input n_17;
input n_8;
input n_0;
input n_2;
input n_10;
input n_9;
input n_12;
input n_6;
input n_11;
input n_14;
input n_7;
input n_18;
input n_3;
input n_5;
input n_4;
input n_1;
input n_16;
input n_15;
input n_13;

output n_19;

wire n_384;
wire n_37;
wire n_430;
wire n_35;
wire n_29;
wire n_91;
wire n_114;
wire n_460;
wire n_300;
wire n_415;
wire n_194;
wire n_301;
wire n_280;
wire n_177;
wire n_271;
wire n_47;
wire n_281;
wire n_311;
wire n_163;
wire n_22;
wire n_320;
wire n_197;
wire n_105;
wire n_27;
wire n_48;
wire n_518;
wire n_446;
wire n_199;
wire n_535;
wire n_95;
wire n_541;
wire n_441;
wire n_557;
wire n_238;
wire n_67;
wire n_350;
wire n_235;
wire n_107;
wire n_369;
wire n_498;
wire n_471;
wire n_376;
wire n_354;
wire n_136;
wire n_267;
wire n_239;
wire n_290;
wire n_553;
wire n_121;
wire n_234;
wire n_160;
wire n_211;
wire n_574;
wire n_490;
wire n_39;
wire n_302;
wire n_26;
wire n_222;
wire n_118;
wire n_220;
wire n_355;
wire n_123;
wire n_463;
wire n_425;
wire n_455;
wire n_462;
wire n_50;
wire n_409;
wire n_485;
wire n_186;
wire n_137;
wire n_491;
wire n_72;
wire n_440;
wire n_171;
wire n_151;
wire n_272;
wire n_461;
wire n_198;
wire n_203;
wire n_500;
wire n_562;
wire n_23;
wire n_362;
wire n_71;
wire n_61;
wire n_99;
wire n_327;
wire n_326;
wire n_339;
wire n_80;
wire n_30;
wire n_328;
wire n_149;
wire n_366;
wire n_332;
wire n_578;
wire n_456;
wire n_259;
wire n_556;
wire n_57;
wire n_507;
wire n_157;
wire n_84;
wire n_560;
wire n_538;
wire n_527;
wire n_55;
wire n_499;
wire n_58;
wire n_52;
wire n_565;
wire n_466;
wire n_353;
wire n_453;
wire n_551;
wire n_230;
wire n_417;
wire n_428;
wire n_128;
wire n_202;
wire n_216;
wire n_483;
wire n_367;
wire n_127;
wire n_356;
wire n_365;
wire n_423;
wire n_464;
wire n_36;
wire n_81;
wire n_102;
wire n_101;
wire n_422;
wire n_317;
wire n_506;
wire n_108;
wire n_550;
wire n_233;
wire n_73;
wire n_532;
wire n_348;
wire n_516;
wire n_473;
wire n_252;
wire n_363;
wire n_310;
wire n_345;
wire n_78;
wire n_83;
wire n_288;
wire n_525;
wire n_221;
wire n_393;
wire n_489;
wire n_104;
wire n_153;
wire n_443;
wire n_337;
wire n_544;
wire n_131;
wire n_439;
wire n_517;
wire n_322;
wire n_87;
wire n_40;
wire n_561;
wire n_98;
wire n_378;
wire n_469;
wire n_200;
wire n_432;
wire n_465;
wire n_569;
wire n_335;
wire n_214;
wire n_113;
wire n_566;
wire n_543;
wire n_251;
wire n_459;
wire n_576;
wire n_139;
wire n_33;
wire n_175;
wire n_338;
wire n_488;
wire n_156;
wire n_387;
wire n_434;
wire n_66;
wire n_577;
wire n_305;
wire n_505;
wire n_62;
wire n_254;
wire n_250;
wire n_564;
wire n_304;
wire n_390;
wire n_77;
wire n_399;
wire n_219;
wire n_470;
wire n_372;
wire n_122;
wire n_262;
wire n_334;
wire n_383;
wire n_246;
wire n_523;
wire n_21;
wire n_476;
wire n_529;
wire n_69;
wire n_31;
wire n_426;
wire n_590;
wire n_154;
wire n_495;
wire n_315;
wire n_296;
wire n_134;
wire n_223;
wire n_371;
wire n_410;
wire n_421;
wire n_110;
wire n_195;
wire n_592;
wire n_533;
wire n_289;
wire n_117;
wire n_193;
wire n_382;
wire n_411;
wire n_20;
wire n_278;
wire n_314;
wire n_103;
wire n_559;
wire n_232;
wire n_582;
wire n_448;
wire n_212;
wire n_579;
wire n_284;
wire n_402;
wire n_478;
wire n_180;
wire n_124;
wire n_264;
wire n_97;
wire n_34;
wire n_190;
wire n_583;
wire n_60;
wire n_263;
wire n_46;
wire n_59;
wire n_452;
wire n_213;
wire n_511;
wire n_524;
wire n_589;
wire n_25;
wire n_480;
wire n_542;
wire n_329;
wire n_224;
wire n_274;
wire n_182;
wire n_269;
wire n_515;
wire n_89;
wire n_407;
wire n_419;
wire n_386;
wire n_521;
wire n_341;
wire n_331;
wire n_49;
wire n_514;
wire n_68;
wire n_497;
wire n_395;
wire n_146;
wire n_496;
wire n_286;
wire n_166;
wire n_176;
wire n_215;
wire n_323;
wire n_312;
wire n_325;
wire n_307;
wire n_316;
wire n_161;
wire n_207;
wire n_526;
wire n_431;
wire n_420;
wire n_357;
wire n_237;
wire n_445;
wire n_173;
wire n_115;
wire n_474;
wire n_184;
wire n_164;
wire n_380;
wire n_414;
wire n_140;
wire n_126;
wire n_342;
wire n_586;
wire n_155;
wire n_120;
wire n_405;
wire n_412;
wire n_572;
wire n_548;
wire n_319;
wire n_93;
wire n_493;
wire n_242;
wire n_487;
wire n_142;
wire n_522;
wire n_397;
wire n_76;
wire n_403;
wire n_79;
wire n_282;
wire n_147;
wire n_359;
wire n_265;
wire n_231;
wire n_44;
wire n_482;
wire n_208;
wire n_162;
wire n_449;
wire n_106;
wire n_172;
wire n_285;
wire n_531;
wire n_546;
wire n_112;
wire n_554;
wire n_508;
wire n_145;
wire n_266;
wire n_377;
wire n_109;
wire n_503;
wire n_391;
wire n_427;
wire n_401;
wire n_536;
wire n_148;
wire n_373;
wire n_563;
wire n_558;
wire n_510;
wire n_396;
wire n_501;
wire n_392;
wire n_575;
wire n_375;
wire n_196;
wire n_298;
wire n_330;
wire n_333;
wire n_450;
wire n_492;
wire n_152;
wire n_584;
wire n_270;
wire n_159;
wire n_429;
wire n_347;
wire n_183;
wire n_248;
wire n_192;
wire n_318;
wire n_537;
wire n_90;
wire n_336;
wire n_258;
wire n_458;
wire n_150;
wire n_41;
wire n_74;
wire n_475;
wire n_404;
wire n_158;
wire n_204;
wire n_241;
wire n_504;
wire n_111;
wire n_479;
wire n_226;
wire n_125;
wire n_297;
wire n_413;
wire n_585;
wire n_494;
wire n_539;
wire n_512;
wire n_75;
wire n_581;
wire n_346;
wire n_340;
wire n_279;
wire n_244;
wire n_179;
wire n_138;
wire n_217;
wire n_53;
wire n_457;
wire n_119;
wire n_283;
wire n_181;
wire n_358;
wire n_534;
wire n_256;
wire n_520;
wire n_253;
wire n_273;
wire n_54;
wire n_168;
wire n_38;
wire n_442;
wire n_385;
wire n_545;
wire n_201;
wire n_484;
wire n_587;
wire n_260;
wire n_247;
wire n_249;
wire n_349;
wire n_418;
wire n_502;
wire n_472;
wire n_292;
wire n_343;
wire n_486;
wire n_64;
wire n_291;
wire n_236;
wire n_370;
wire n_276;
wire n_374;
wire n_287;
wire n_388;
wire n_174;
wire n_400;
wire n_255;
wire n_299;
wire n_243;
wire n_352;
wire n_477;
wire n_56;
wire n_293;
wire n_275;
wire n_381;
wire n_227;
wire n_229;
wire n_454;
wire n_571;
wire n_573;
wire n_379;
wire n_141;
wire n_555;
wire n_65;
wire n_188;
wire n_444;
wire n_178;
wire n_360;
wire n_398;
wire n_189;
wire n_170;
wire n_570;
wire n_28;
wire n_245;
wire n_451;
wire n_45;
wire n_437;
wire n_268;
wire n_42;
wire n_313;
wire n_94;
wire n_547;
wire n_309;
wire n_294;
wire n_116;
wire n_416;
wire n_513;
wire n_143;
wire n_588;
wire n_351;
wire n_467;
wire n_129;
wire n_135;
wire n_306;
wire n_540;
wire n_218;
wire n_528;
wire n_165;
wire n_406;
wire n_303;
wire n_321;
wire n_100;
wire n_368;
wire n_567;
wire n_51;
wire n_509;
wire n_205;
wire n_519;
wire n_530;
wire n_361;
wire n_261;
wire n_86;
wire n_324;
wire n_549;
wire n_70;
wire n_568;
wire n_435;
wire n_32;
wire n_228;
wire n_389;
wire n_580;
wire n_144;
wire n_130;
wire n_225;
wire n_43;
wire n_438;
wire n_82;
wire n_132;
wire n_277;
wire n_185;
wire n_240;
wire n_209;
wire n_481;
wire n_191;
wire n_394;
wire n_63;
wire n_24;
wire n_92;
wire n_187;
wire n_436;
wire n_88;
wire n_169;
wire n_167;
wire n_295;
wire n_424;
wire n_133;
wire n_468;
wire n_447;
wire n_257;
wire n_344;
wire n_210;
wire n_206;
wire n_552;
wire n_408;
wire n_85;
wire n_591;
wire n_96;
wire n_308;
wire n_433;
wire n_364;

AOI21xp5_ASAP7_75t_L g19 ( 
.A1(n_0),
.A2(n_20),
.B(n_591),
.Y(n_19)
);

NOR2xp33_ASAP7_75t_L g591 ( 
.A(n_0),
.B(n_592),
.Y(n_591)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_1),
.B(n_96),
.Y(n_95)
);

AND2x2_ASAP7_75t_L g172 ( 
.A(n_1),
.B(n_173),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_SL g218 ( 
.A(n_1),
.B(n_219),
.Y(n_218)
);

NAND2xp5_ASAP7_75t_SL g237 ( 
.A(n_1),
.B(n_238),
.Y(n_237)
);

AND2x2_ASAP7_75t_L g249 ( 
.A(n_1),
.B(n_250),
.Y(n_249)
);

INVx1_ASAP7_75t_L g305 ( 
.A(n_1),
.Y(n_305)
);

NAND2xp5_ASAP7_75t_L g344 ( 
.A(n_1),
.B(n_46),
.Y(n_344)
);

AND2x2_ASAP7_75t_L g370 ( 
.A(n_1),
.B(n_371),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_L g36 ( 
.A(n_2),
.B(n_37),
.Y(n_36)
);

NAND2xp5_ASAP7_75t_L g53 ( 
.A(n_2),
.B(n_54),
.Y(n_53)
);

NAND2xp5_ASAP7_75t_L g89 ( 
.A(n_2),
.B(n_90),
.Y(n_89)
);

NAND2xp5_ASAP7_75t_L g103 ( 
.A(n_2),
.B(n_104),
.Y(n_103)
);

AND2x2_ASAP7_75t_L g146 ( 
.A(n_2),
.B(n_147),
.Y(n_146)
);

AND2x2_ASAP7_75t_L g213 ( 
.A(n_2),
.B(n_214),
.Y(n_213)
);

NAND2xp5_ASAP7_75t_SL g270 ( 
.A(n_2),
.B(n_271),
.Y(n_270)
);

NAND2xp5_ASAP7_75t_L g347 ( 
.A(n_2),
.B(n_348),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g70 ( 
.A(n_3),
.B(n_71),
.Y(n_70)
);

CKINVDCx16_ASAP7_75t_R g110 ( 
.A(n_3),
.Y(n_110)
);

AND2x2_ASAP7_75t_L g165 ( 
.A(n_3),
.B(n_166),
.Y(n_165)
);

AND2x4_ASAP7_75t_L g185 ( 
.A(n_3),
.B(n_186),
.Y(n_185)
);

NAND2xp5_ASAP7_75t_L g232 ( 
.A(n_3),
.B(n_180),
.Y(n_232)
);

NAND2xp5_ASAP7_75t_L g275 ( 
.A(n_3),
.B(n_276),
.Y(n_275)
);

AND2x2_ASAP7_75t_SL g306 ( 
.A(n_3),
.B(n_307),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g334 ( 
.A(n_3),
.B(n_335),
.Y(n_334)
);

INVx2_ASAP7_75t_L g150 ( 
.A(n_4),
.Y(n_150)
);

BUFx5_ASAP7_75t_L g154 ( 
.A(n_4),
.Y(n_154)
);

BUFx5_ASAP7_75t_L g372 ( 
.A(n_4),
.Y(n_372)
);

BUFx3_ASAP7_75t_L g441 ( 
.A(n_4),
.Y(n_441)
);

AOI22xp5_ASAP7_75t_SL g152 ( 
.A1(n_5),
.A2(n_9),
.B1(n_153),
.B2(n_155),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_SL g205 ( 
.A(n_5),
.B(n_206),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_SL g223 ( 
.A(n_5),
.B(n_224),
.Y(n_223)
);

AND2x2_ASAP7_75t_L g311 ( 
.A(n_5),
.B(n_312),
.Y(n_311)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_5),
.B(n_379),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g400 ( 
.A(n_5),
.B(n_401),
.Y(n_400)
);

NAND2xp5_ASAP7_75t_L g433 ( 
.A(n_5),
.B(n_434),
.Y(n_433)
);

AND2x2_ASAP7_75t_L g437 ( 
.A(n_5),
.B(n_438),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g471 ( 
.A(n_5),
.B(n_472),
.Y(n_471)
);

INVx6_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

INVx1_ASAP7_75t_L g49 ( 
.A(n_6),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_6),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g113 ( 
.A(n_6),
.Y(n_113)
);

AND2x2_ASAP7_75t_L g162 ( 
.A(n_7),
.B(n_163),
.Y(n_162)
);

NAND2xp33_ASAP7_75t_SL g189 ( 
.A(n_7),
.B(n_190),
.Y(n_189)
);

NAND2xp5_ASAP7_75t_SL g234 ( 
.A(n_7),
.B(n_235),
.Y(n_234)
);

NAND2xp5_ASAP7_75t_SL g254 ( 
.A(n_7),
.B(n_255),
.Y(n_254)
);

AND2x2_ASAP7_75t_L g316 ( 
.A(n_7),
.B(n_317),
.Y(n_316)
);

AND2x2_ASAP7_75t_L g439 ( 
.A(n_7),
.B(n_440),
.Y(n_439)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_7),
.B(n_444),
.Y(n_443)
);

NAND2xp5_ASAP7_75t_L g461 ( 
.A(n_7),
.B(n_462),
.Y(n_461)
);

NAND2xp5_ASAP7_75t_SL g177 ( 
.A(n_8),
.B(n_178),
.Y(n_177)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_8),
.B(n_375),
.Y(n_374)
);

NAND2xp5_ASAP7_75t_SL g396 ( 
.A(n_8),
.B(n_397),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_L g429 ( 
.A(n_8),
.B(n_430),
.Y(n_429)
);

NAND2xp5_ASAP7_75t_L g480 ( 
.A(n_8),
.B(n_481),
.Y(n_480)
);

NAND2xp5_ASAP7_75t_SL g485 ( 
.A(n_8),
.B(n_486),
.Y(n_485)
);

NAND2xp5_ASAP7_75t_SL g494 ( 
.A(n_8),
.B(n_495),
.Y(n_494)
);

NAND2xp5_ASAP7_75t_L g67 ( 
.A(n_9),
.B(n_68),
.Y(n_67)
);

NAND2xp5_ASAP7_75t_L g83 ( 
.A(n_9),
.B(n_84),
.Y(n_83)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_9),
.B(n_100),
.Y(n_99)
);

AND2x2_ASAP7_75t_L g142 ( 
.A(n_9),
.B(n_143),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_9),
.B(n_186),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g279 ( 
.A(n_9),
.B(n_280),
.Y(n_279)
);

NAND2xp5_ASAP7_75t_L g346 ( 
.A(n_9),
.B(n_312),
.Y(n_346)
);

CKINVDCx14_ASAP7_75t_R g383 ( 
.A(n_9),
.Y(n_383)
);

NAND2xp5_ASAP7_75t_L g26 ( 
.A(n_10),
.B(n_27),
.Y(n_26)
);

AND2x2_ASAP7_75t_SL g32 ( 
.A(n_10),
.B(n_33),
.Y(n_32)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_10),
.Y(n_50)
);

AND2x2_ASAP7_75t_L g74 ( 
.A(n_10),
.B(n_75),
.Y(n_74)
);

AND2x2_ASAP7_75t_L g209 ( 
.A(n_10),
.B(n_210),
.Y(n_209)
);

NAND2xp5_ASAP7_75t_L g585 ( 
.A(n_10),
.B(n_586),
.Y(n_585)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_11),
.Y(n_118)
);

BUFx6f_ASAP7_75t_L g176 ( 
.A(n_11),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_11),
.Y(n_188)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_11),
.Y(n_273)
);

BUFx5_ASAP7_75t_L g490 ( 
.A(n_11),
.Y(n_490)
);

BUFx4f_ASAP7_75t_L g145 ( 
.A(n_12),
.Y(n_145)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_12),
.Y(n_168)
);

BUFx12f_ASAP7_75t_L g215 ( 
.A(n_12),
.Y(n_215)
);

BUFx6f_ASAP7_75t_L g265 ( 
.A(n_12),
.Y(n_265)
);

CKINVDCx20_ASAP7_75t_R g592 ( 
.A(n_13),
.Y(n_592)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_14),
.Y(n_35)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_14),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g164 ( 
.A(n_14),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g241 ( 
.A(n_14),
.Y(n_241)
);

NAND2xp5_ASAP7_75t_L g138 ( 
.A(n_15),
.B(n_139),
.Y(n_138)
);

CKINVDCx16_ASAP7_75t_R g160 ( 
.A(n_15),
.Y(n_160)
);

AND2x4_ASAP7_75t_SL g179 ( 
.A(n_15),
.B(n_180),
.Y(n_179)
);

AND2x2_ASAP7_75t_SL g196 ( 
.A(n_15),
.B(n_197),
.Y(n_196)
);

AND2x2_ASAP7_75t_L g226 ( 
.A(n_15),
.B(n_227),
.Y(n_226)
);

AND2x2_ASAP7_75t_L g314 ( 
.A(n_15),
.B(n_315),
.Y(n_314)
);

AND2x2_ASAP7_75t_L g367 ( 
.A(n_15),
.B(n_368),
.Y(n_367)
);

AND2x2_ASAP7_75t_L g446 ( 
.A(n_15),
.B(n_447),
.Y(n_446)
);

BUFx6f_ASAP7_75t_L g77 ( 
.A(n_16),
.Y(n_77)
);

INVx3_ASAP7_75t_L g183 ( 
.A(n_16),
.Y(n_183)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_16),
.Y(n_222)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_16),
.Y(n_283)
);

BUFx3_ASAP7_75t_L g319 ( 
.A(n_16),
.Y(n_319)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g107 ( 
.A(n_17),
.Y(n_107)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_18),
.Y(n_60)
);

BUFx5_ASAP7_75t_L g68 ( 
.A(n_18),
.Y(n_68)
);

BUFx8_ASAP7_75t_L g72 ( 
.A(n_18),
.Y(n_72)
);

BUFx3_ASAP7_75t_L g256 ( 
.A(n_18),
.Y(n_256)
);

XOR2x2_ASAP7_75t_L g20 ( 
.A(n_21),
.B(n_580),
.Y(n_20)
);

OAI21x1_ASAP7_75t_L g21 ( 
.A1(n_22),
.A2(n_127),
.B(n_579),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_23),
.Y(n_22)
);

NAND2xp5_ASAP7_75t_L g23 ( 
.A(n_24),
.B(n_78),
.Y(n_23)
);

OR2x2_ASAP7_75t_L g579 ( 
.A(n_24),
.B(n_78),
.Y(n_579)
);

BUFx24_ASAP7_75t_SL g594 ( 
.A(n_24),
.Y(n_594)
);

FAx1_ASAP7_75t_SL g24 ( 
.A(n_25),
.B(n_41),
.CI(n_61),
.CON(n_24),
.SN(n_24)
);

MAJIxp5_ASAP7_75t_L g589 ( 
.A(n_25),
.B(n_41),
.C(n_61),
.Y(n_589)
);

MAJIxp5_ASAP7_75t_L g25 ( 
.A(n_26),
.B(n_32),
.C(n_36),
.Y(n_25)
);

AOI22xp5_ASAP7_75t_L g42 ( 
.A1(n_26),
.A2(n_43),
.B1(n_51),
.B2(n_52),
.Y(n_42)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_26),
.Y(n_51)
);

AOI22xp5_ASAP7_75t_L g64 ( 
.A1(n_26),
.A2(n_32),
.B1(n_51),
.B2(n_65),
.Y(n_64)
);

MAJIxp5_ASAP7_75t_SL g583 ( 
.A(n_26),
.B(n_43),
.C(n_53),
.Y(n_583)
);

HB1xp67_ASAP7_75t_L g27 ( 
.A(n_28),
.Y(n_27)
);

INVx2_ASAP7_75t_L g28 ( 
.A(n_29),
.Y(n_28)
);

INVx2_ASAP7_75t_L g29 ( 
.A(n_30),
.Y(n_29)
);

BUFx6f_ASAP7_75t_L g30 ( 
.A(n_31),
.Y(n_30)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_31),
.Y(n_87)
);

BUFx6f_ASAP7_75t_L g252 ( 
.A(n_31),
.Y(n_252)
);

BUFx6f_ASAP7_75t_L g399 ( 
.A(n_31),
.Y(n_399)
);

INVx1_ASAP7_75t_SL g65 ( 
.A(n_32),
.Y(n_65)
);

MAJIxp5_ASAP7_75t_L g69 ( 
.A(n_32),
.B(n_70),
.C(n_73),
.Y(n_69)
);

AOI22xp5_ASAP7_75t_L g121 ( 
.A1(n_32),
.A2(n_65),
.B1(n_73),
.B2(n_74),
.Y(n_121)
);

INVx3_ASAP7_75t_L g33 ( 
.A(n_34),
.Y(n_33)
);

INVx5_ASAP7_75t_L g278 ( 
.A(n_34),
.Y(n_278)
);

BUFx6f_ASAP7_75t_L g34 ( 
.A(n_35),
.Y(n_34)
);

XOR2xp5_ASAP7_75t_L g63 ( 
.A(n_36),
.B(n_64),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g37 ( 
.A(n_38),
.Y(n_37)
);

INVx4_ASAP7_75t_L g38 ( 
.A(n_39),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_40),
.Y(n_39)
);

INVx4_ASAP7_75t_L g375 ( 
.A(n_40),
.Y(n_375)
);

XNOR2xp5_ASAP7_75t_L g41 ( 
.A(n_42),
.B(n_53),
.Y(n_41)
);

INVx1_ASAP7_75t_L g52 ( 
.A(n_43),
.Y(n_52)
);

AOI22xp5_ASAP7_75t_L g584 ( 
.A1(n_43),
.A2(n_52),
.B1(n_585),
.B2(n_588),
.Y(n_584)
);

NOR2xp33_ASAP7_75t_SL g43 ( 
.A(n_44),
.B(n_50),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_45),
.Y(n_44)
);

HB1xp67_ASAP7_75t_L g45 ( 
.A(n_46),
.Y(n_45)
);

INVx2_ASAP7_75t_L g46 ( 
.A(n_47),
.Y(n_46)
);

INVx2_ASAP7_75t_L g47 ( 
.A(n_48),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_49),
.Y(n_48)
);

OR2x2_ASAP7_75t_SL g114 ( 
.A(n_50),
.B(n_115),
.Y(n_114)
);

OR2x2_ASAP7_75t_L g261 ( 
.A(n_50),
.B(n_262),
.Y(n_261)
);

BUFx2_ASAP7_75t_L g54 ( 
.A(n_55),
.Y(n_54)
);

INVx3_ASAP7_75t_L g55 ( 
.A(n_56),
.Y(n_55)
);

INVx2_ASAP7_75t_L g56 ( 
.A(n_57),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g57 ( 
.A(n_58),
.Y(n_57)
);

INVx4_ASAP7_75t_L g58 ( 
.A(n_59),
.Y(n_58)
);

INVx8_ASAP7_75t_L g207 ( 
.A(n_59),
.Y(n_207)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_60),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

MAJIxp5_ASAP7_75t_L g61 ( 
.A(n_62),
.B(n_66),
.C(n_69),
.Y(n_61)
);

OAI22xp5_ASAP7_75t_L g123 ( 
.A1(n_62),
.A2(n_63),
.B1(n_124),
.B2(n_125),
.Y(n_123)
);

INVx1_ASAP7_75t_L g62 ( 
.A(n_63),
.Y(n_62)
);

AOI22xp5_ASAP7_75t_L g125 ( 
.A1(n_66),
.A2(n_67),
.B1(n_69),
.B2(n_126),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g66 ( 
.A(n_67),
.Y(n_66)
);

INVx1_ASAP7_75t_L g126 ( 
.A(n_69),
.Y(n_126)
);

XOR2xp5_ASAP7_75t_L g120 ( 
.A(n_70),
.B(n_121),
.Y(n_120)
);

BUFx12f_ASAP7_75t_L g71 ( 
.A(n_72),
.Y(n_71)
);

INVx3_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

INVx1_ASAP7_75t_L g587 ( 
.A(n_72),
.Y(n_587)
);

AOI22xp5_ASAP7_75t_L g545 ( 
.A1(n_73),
.A2(n_74),
.B1(n_114),
.B2(n_340),
.Y(n_545)
);

INVx2_ASAP7_75t_L g73 ( 
.A(n_74),
.Y(n_73)
);

MAJIxp5_ASAP7_75t_SL g108 ( 
.A(n_74),
.B(n_109),
.C(n_114),
.Y(n_108)
);

INVx3_ASAP7_75t_L g75 ( 
.A(n_76),
.Y(n_75)
);

INVx4_ASAP7_75t_L g76 ( 
.A(n_77),
.Y(n_76)
);

MAJIxp5_ASAP7_75t_L g78 ( 
.A(n_79),
.B(n_122),
.C(n_123),
.Y(n_78)
);

XNOR2xp5_ASAP7_75t_L g551 ( 
.A(n_79),
.B(n_552),
.Y(n_551)
);

MAJIxp5_ASAP7_75t_L g79 ( 
.A(n_80),
.B(n_108),
.C(n_119),
.Y(n_79)
);

XOR2xp5_ASAP7_75t_L g549 ( 
.A(n_80),
.B(n_550),
.Y(n_549)
);

XNOR2xp5_ASAP7_75t_L g80 ( 
.A(n_81),
.B(n_98),
.Y(n_80)
);

MAJIxp5_ASAP7_75t_L g122 ( 
.A(n_81),
.B(n_99),
.C(n_103),
.Y(n_122)
);

MAJIxp5_ASAP7_75t_L g81 ( 
.A(n_82),
.B(n_88),
.C(n_95),
.Y(n_81)
);

AOI22xp5_ASAP7_75t_L g541 ( 
.A1(n_82),
.A2(n_83),
.B1(n_88),
.B2(n_89),
.Y(n_541)
);

INVx1_ASAP7_75t_L g82 ( 
.A(n_83),
.Y(n_82)
);

HB1xp67_ASAP7_75t_L g84 ( 
.A(n_85),
.Y(n_84)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_86),
.Y(n_85)
);

BUFx6f_ASAP7_75t_L g156 ( 
.A(n_86),
.Y(n_156)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_87),
.Y(n_86)
);

INVx1_ASAP7_75t_L g88 ( 
.A(n_89),
.Y(n_88)
);

INVx2_ASAP7_75t_L g90 ( 
.A(n_91),
.Y(n_90)
);

INVx2_ASAP7_75t_L g91 ( 
.A(n_92),
.Y(n_91)
);

INVx4_ASAP7_75t_L g92 ( 
.A(n_93),
.Y(n_92)
);

INVx2_ASAP7_75t_L g432 ( 
.A(n_93),
.Y(n_432)
);

BUFx3_ASAP7_75t_L g93 ( 
.A(n_94),
.Y(n_93)
);

INVx2_ASAP7_75t_L g229 ( 
.A(n_94),
.Y(n_229)
);

XNOR2xp5_ASAP7_75t_L g540 ( 
.A(n_95),
.B(n_541),
.Y(n_540)
);

INVx1_ASAP7_75t_L g96 ( 
.A(n_97),
.Y(n_96)
);

XNOR2xp5_ASAP7_75t_L g98 ( 
.A(n_99),
.B(n_103),
.Y(n_98)
);

INVx2_ASAP7_75t_L g100 ( 
.A(n_101),
.Y(n_100)
);

INVx4_ASAP7_75t_L g101 ( 
.A(n_102),
.Y(n_101)
);

INVx2_ASAP7_75t_L g161 ( 
.A(n_102),
.Y(n_161)
);

INVx6_ASAP7_75t_L g236 ( 
.A(n_102),
.Y(n_236)
);

BUFx3_ASAP7_75t_L g104 ( 
.A(n_105),
.Y(n_104)
);

INVx2_ASAP7_75t_SL g105 ( 
.A(n_106),
.Y(n_105)
);

INVx1_ASAP7_75t_L g106 ( 
.A(n_107),
.Y(n_106)
);

BUFx6f_ASAP7_75t_L g190 ( 
.A(n_107),
.Y(n_190)
);

INVx4_ASAP7_75t_L g198 ( 
.A(n_107),
.Y(n_198)
);

XNOR2xp5_ASAP7_75t_L g550 ( 
.A(n_108),
.B(n_120),
.Y(n_550)
);

XNOR2xp5_ASAP7_75t_SL g544 ( 
.A(n_109),
.B(n_545),
.Y(n_544)
);

NOR2xp33_ASAP7_75t_L g109 ( 
.A(n_110),
.B(n_111),
.Y(n_109)
);

HB1xp67_ASAP7_75t_L g111 ( 
.A(n_112),
.Y(n_111)
);

INVx2_ASAP7_75t_L g224 ( 
.A(n_112),
.Y(n_224)
);

INVx3_ASAP7_75t_L g112 ( 
.A(n_113),
.Y(n_112)
);

AOI22xp33_ASAP7_75t_L g339 ( 
.A1(n_114),
.A2(n_261),
.B1(n_266),
.B2(n_340),
.Y(n_339)
);

INVx1_ASAP7_75t_L g340 ( 
.A(n_114),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_114),
.B(n_266),
.C(n_334),
.Y(n_546)
);

INVx3_ASAP7_75t_L g115 ( 
.A(n_116),
.Y(n_115)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_117),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g117 ( 
.A(n_118),
.Y(n_117)
);

HB1xp67_ASAP7_75t_L g119 ( 
.A(n_120),
.Y(n_119)
);

XNOR2xp5_ASAP7_75t_L g552 ( 
.A(n_122),
.B(n_123),
.Y(n_552)
);

INVx1_ASAP7_75t_L g124 ( 
.A(n_125),
.Y(n_124)
);

AOI21x1_ASAP7_75t_L g127 ( 
.A1(n_128),
.A2(n_533),
.B(n_574),
.Y(n_127)
);

AO21x2_ASAP7_75t_L g128 ( 
.A1(n_129),
.A2(n_360),
.B(n_530),
.Y(n_128)
);

NOR2xp33_ASAP7_75t_L g129 ( 
.A(n_130),
.B(n_326),
.Y(n_129)
);

AND2x2_ASAP7_75t_L g130 ( 
.A(n_131),
.B(n_286),
.Y(n_130)
);

OR2x2_ASAP7_75t_L g531 ( 
.A(n_131),
.B(n_286),
.Y(n_531)
);

XNOR2xp5_ASAP7_75t_L g131 ( 
.A(n_132),
.B(n_201),
.Y(n_131)
);

INVxp67_ASAP7_75t_SL g359 ( 
.A(n_132),
.Y(n_359)
);

MAJIxp5_ASAP7_75t_L g132 ( 
.A(n_133),
.B(n_169),
.C(n_191),
.Y(n_132)
);

INVxp33_ASAP7_75t_SL g133 ( 
.A(n_134),
.Y(n_133)
);

XNOR2xp5_ASAP7_75t_L g288 ( 
.A(n_134),
.B(n_289),
.Y(n_288)
);

MAJIxp5_ASAP7_75t_L g134 ( 
.A(n_135),
.B(n_151),
.C(n_157),
.Y(n_134)
);

XNOR2xp5_ASAP7_75t_L g412 ( 
.A(n_135),
.B(n_413),
.Y(n_412)
);

XNOR2xp5_ASAP7_75t_L g135 ( 
.A(n_136),
.B(n_141),
.Y(n_135)
);

MAJx2_ASAP7_75t_L g542 ( 
.A(n_136),
.B(n_249),
.C(n_356),
.Y(n_542)
);

INVx1_ASAP7_75t_L g136 ( 
.A(n_137),
.Y(n_136)
);

XNOR2xp5_ASAP7_75t_L g353 ( 
.A(n_137),
.B(n_249),
.Y(n_353)
);

INVx1_ASAP7_75t_L g137 ( 
.A(n_138),
.Y(n_137)
);

MAJIxp5_ASAP7_75t_L g193 ( 
.A(n_138),
.B(n_142),
.C(n_146),
.Y(n_193)
);

INVx4_ASAP7_75t_L g139 ( 
.A(n_140),
.Y(n_139)
);

INVx6_ASAP7_75t_L g178 ( 
.A(n_140),
.Y(n_178)
);

XNOR2xp5_ASAP7_75t_L g141 ( 
.A(n_142),
.B(n_146),
.Y(n_141)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_144),
.Y(n_143)
);

INVx2_ASAP7_75t_L g144 ( 
.A(n_145),
.Y(n_144)
);

INVx2_ASAP7_75t_L g147 ( 
.A(n_148),
.Y(n_147)
);

INVx1_ASAP7_75t_L g148 ( 
.A(n_149),
.Y(n_148)
);

INVx1_ASAP7_75t_L g211 ( 
.A(n_149),
.Y(n_211)
);

BUFx6f_ASAP7_75t_L g309 ( 
.A(n_149),
.Y(n_309)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_150),
.Y(n_149)
);

AOI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_151),
.A2(n_152),
.B1(n_157),
.B2(n_414),
.Y(n_413)
);

INVx1_ASAP7_75t_L g151 ( 
.A(n_152),
.Y(n_151)
);

AOI21xp5_ASAP7_75t_L g377 ( 
.A1(n_152),
.A2(n_378),
.B(n_382),
.Y(n_377)
);

BUFx12f_ASAP7_75t_L g153 ( 
.A(n_154),
.Y(n_153)
);

INVx3_ASAP7_75t_L g155 ( 
.A(n_156),
.Y(n_155)
);

INVx1_ASAP7_75t_L g414 ( 
.A(n_157),
.Y(n_414)
);

MAJx2_ASAP7_75t_L g157 ( 
.A(n_158),
.B(n_162),
.C(n_165),
.Y(n_157)
);

AOI22xp5_ASAP7_75t_L g258 ( 
.A1(n_158),
.A2(n_159),
.B1(n_259),
.B2(n_260),
.Y(n_258)
);

AOI22xp5_ASAP7_75t_L g299 ( 
.A1(n_158),
.A2(n_159),
.B1(n_165),
.B2(n_300),
.Y(n_299)
);

INVx1_ASAP7_75t_SL g158 ( 
.A(n_159),
.Y(n_158)
);

MAJx2_ASAP7_75t_L g354 ( 
.A(n_159),
.B(n_209),
.C(n_261),
.Y(n_354)
);

OR2x2_ASAP7_75t_L g159 ( 
.A(n_160),
.B(n_161),
.Y(n_159)
);

XNOR2xp5_ASAP7_75t_L g298 ( 
.A(n_162),
.B(n_299),
.Y(n_298)
);

BUFx3_ASAP7_75t_L g163 ( 
.A(n_164),
.Y(n_163)
);

INVx2_ASAP7_75t_L g313 ( 
.A(n_164),
.Y(n_313)
);

INVx1_ASAP7_75t_L g300 ( 
.A(n_165),
.Y(n_300)
);

INVx2_ASAP7_75t_L g166 ( 
.A(n_167),
.Y(n_166)
);

BUFx6f_ASAP7_75t_L g167 ( 
.A(n_168),
.Y(n_167)
);

HB1xp67_ASAP7_75t_L g169 ( 
.A(n_170),
.Y(n_169)
);

AOI22xp5_ASAP7_75t_SL g289 ( 
.A1(n_170),
.A2(n_191),
.B1(n_192),
.B2(n_290),
.Y(n_289)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_170),
.Y(n_290)
);

MAJIxp5_ASAP7_75t_L g170 ( 
.A(n_171),
.B(n_184),
.C(n_189),
.Y(n_170)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_171),
.B(n_321),
.Y(n_320)
);

MAJIxp5_ASAP7_75t_L g171 ( 
.A(n_172),
.B(n_177),
.C(n_179),
.Y(n_171)
);

AOI22xp5_ASAP7_75t_L g388 ( 
.A1(n_172),
.A2(n_179),
.B1(n_389),
.B2(n_390),
.Y(n_388)
);

INVxp67_ASAP7_75t_L g390 ( 
.A(n_172),
.Y(n_390)
);

INVx2_ASAP7_75t_L g173 ( 
.A(n_174),
.Y(n_173)
);

INVx3_ASAP7_75t_L g174 ( 
.A(n_175),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g175 ( 
.A(n_176),
.Y(n_175)
);

INVx6_ASAP7_75t_L g465 ( 
.A(n_176),
.Y(n_465)
);

XOR2xp5_ASAP7_75t_SL g387 ( 
.A(n_177),
.B(n_388),
.Y(n_387)
);

INVx1_ASAP7_75t_L g389 ( 
.A(n_179),
.Y(n_389)
);

XNOR2xp5_ASAP7_75t_L g427 ( 
.A(n_179),
.B(n_428),
.Y(n_427)
);

INVx2_ASAP7_75t_L g180 ( 
.A(n_181),
.Y(n_180)
);

INVx2_ASAP7_75t_L g181 ( 
.A(n_182),
.Y(n_181)
);

INVx1_ASAP7_75t_L g182 ( 
.A(n_183),
.Y(n_182)
);

AOI22xp5_ASAP7_75t_L g321 ( 
.A1(n_184),
.A2(n_185),
.B1(n_189),
.B2(n_322),
.Y(n_321)
);

CKINVDCx16_ASAP7_75t_R g184 ( 
.A(n_185),
.Y(n_184)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_187),
.Y(n_186)
);

INVx8_ASAP7_75t_L g187 ( 
.A(n_188),
.Y(n_187)
);

INVx1_ASAP7_75t_L g322 ( 
.A(n_189),
.Y(n_322)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_192),
.Y(n_191)
);

XNOR2x1_ASAP7_75t_L g192 ( 
.A(n_193),
.B(n_194),
.Y(n_192)
);

MAJx2_ASAP7_75t_L g243 ( 
.A(n_193),
.B(n_195),
.C(n_244),
.Y(n_243)
);

AOI22xp5_ASAP7_75t_L g194 ( 
.A1(n_195),
.A2(n_196),
.B1(n_199),
.B2(n_200),
.Y(n_194)
);

AOI22xp5_ASAP7_75t_L g516 ( 
.A1(n_195),
.A2(n_196),
.B1(n_373),
.B2(n_374),
.Y(n_516)
);

INVx2_ASAP7_75t_SL g195 ( 
.A(n_196),
.Y(n_195)
);

MAJIxp5_ASAP7_75t_L g365 ( 
.A(n_196),
.B(n_366),
.C(n_373),
.Y(n_365)
);

INVx6_ASAP7_75t_L g197 ( 
.A(n_198),
.Y(n_197)
);

INVx1_ASAP7_75t_L g199 ( 
.A(n_200),
.Y(n_199)
);

HB1xp67_ASAP7_75t_L g244 ( 
.A(n_200),
.Y(n_244)
);

AOI22xp5_ASAP7_75t_SL g201 ( 
.A1(n_202),
.A2(n_257),
.B1(n_284),
.B2(n_285),
.Y(n_201)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_202),
.Y(n_284)
);

XNOR2x1_ASAP7_75t_SL g202 ( 
.A(n_203),
.B(n_242),
.Y(n_202)
);

MAJIxp5_ASAP7_75t_L g328 ( 
.A(n_203),
.B(n_243),
.C(n_329),
.Y(n_328)
);

MAJIxp5_ASAP7_75t_L g203 ( 
.A(n_204),
.B(n_217),
.C(n_230),
.Y(n_203)
);

XNOR2xp5_ASAP7_75t_L g292 ( 
.A(n_204),
.B(n_217),
.Y(n_292)
);

XNOR2x1_ASAP7_75t_L g204 ( 
.A(n_205),
.B(n_208),
.Y(n_204)
);

MAJIxp5_ASAP7_75t_L g268 ( 
.A(n_205),
.B(n_209),
.C(n_213),
.Y(n_268)
);

BUFx2_ASAP7_75t_L g206 ( 
.A(n_207),
.Y(n_206)
);

AOI22xp5_ASAP7_75t_SL g208 ( 
.A1(n_209),
.A2(n_212),
.B1(n_213),
.B2(n_216),
.Y(n_208)
);

INVx1_ASAP7_75t_SL g216 ( 
.A(n_209),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_209),
.A2(n_216),
.B1(n_261),
.B2(n_266),
.Y(n_260)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_211),
.Y(n_210)
);

INVx1_ASAP7_75t_L g212 ( 
.A(n_213),
.Y(n_212)
);

BUFx6f_ASAP7_75t_L g214 ( 
.A(n_215),
.Y(n_214)
);

INVx2_ASAP7_75t_L g369 ( 
.A(n_215),
.Y(n_369)
);

INVx2_ASAP7_75t_L g445 ( 
.A(n_215),
.Y(n_445)
);

INVx3_ASAP7_75t_L g496 ( 
.A(n_215),
.Y(n_496)
);

MAJIxp5_ASAP7_75t_L g217 ( 
.A(n_218),
.B(n_223),
.C(n_225),
.Y(n_217)
);

XOR2xp5_ASAP7_75t_L g323 ( 
.A(n_218),
.B(n_324),
.Y(n_323)
);

INVx5_ASAP7_75t_L g219 ( 
.A(n_220),
.Y(n_219)
);

BUFx6f_ASAP7_75t_L g220 ( 
.A(n_221),
.Y(n_220)
);

BUFx6f_ASAP7_75t_L g221 ( 
.A(n_222),
.Y(n_221)
);

AOI22xp33_ASAP7_75t_L g324 ( 
.A1(n_223),
.A2(n_225),
.B1(n_226),
.B2(n_325),
.Y(n_324)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_223),
.Y(n_325)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_225),
.B(n_396),
.C(n_400),
.Y(n_395)
);

AOI22xp5_ASAP7_75t_L g455 ( 
.A1(n_225),
.A2(n_226),
.B1(n_396),
.B2(n_456),
.Y(n_455)
);

INVx1_ASAP7_75t_L g225 ( 
.A(n_226),
.Y(n_225)
);

INVx2_ASAP7_75t_L g227 ( 
.A(n_228),
.Y(n_227)
);

INVx2_ASAP7_75t_L g228 ( 
.A(n_229),
.Y(n_228)
);

INVx1_ASAP7_75t_L g293 ( 
.A(n_230),
.Y(n_293)
);

XOR2xp5_ASAP7_75t_L g230 ( 
.A(n_231),
.B(n_233),
.Y(n_230)
);

HB1xp67_ASAP7_75t_L g231 ( 
.A(n_232),
.Y(n_231)
);

MAJIxp5_ASAP7_75t_L g246 ( 
.A(n_232),
.B(n_234),
.C(n_237),
.Y(n_246)
);

XNOR2xp5_ASAP7_75t_L g233 ( 
.A(n_234),
.B(n_237),
.Y(n_233)
);

INVx4_ASAP7_75t_L g235 ( 
.A(n_236),
.Y(n_235)
);

INVx8_ASAP7_75t_L g238 ( 
.A(n_239),
.Y(n_238)
);

INVx6_ASAP7_75t_L g239 ( 
.A(n_240),
.Y(n_239)
);

BUFx6f_ASAP7_75t_L g240 ( 
.A(n_241),
.Y(n_240)
);

XNOR2x1_ASAP7_75t_L g242 ( 
.A(n_243),
.B(n_245),
.Y(n_242)
);

HB1xp67_ASAP7_75t_L g329 ( 
.A(n_245),
.Y(n_329)
);

XNOR2x1_ASAP7_75t_L g245 ( 
.A(n_246),
.B(n_247),
.Y(n_245)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_246),
.B(n_248),
.C(n_254),
.Y(n_357)
);

OAI22x1_ASAP7_75t_SL g247 ( 
.A1(n_248),
.A2(n_249),
.B1(n_253),
.B2(n_254),
.Y(n_247)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_249),
.Y(n_248)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_250),
.Y(n_381)
);

INVx2_ASAP7_75t_L g250 ( 
.A(n_251),
.Y(n_250)
);

INVx3_ASAP7_75t_L g251 ( 
.A(n_252),
.Y(n_251)
);

INVx3_ASAP7_75t_L g338 ( 
.A(n_252),
.Y(n_338)
);

INVx1_ASAP7_75t_L g253 ( 
.A(n_254),
.Y(n_253)
);

BUFx6f_ASAP7_75t_L g255 ( 
.A(n_256),
.Y(n_255)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_257),
.Y(n_285)
);

MAJIxp5_ASAP7_75t_L g358 ( 
.A(n_257),
.B(n_284),
.C(n_359),
.Y(n_358)
);

XOR2x2_ASAP7_75t_L g257 ( 
.A(n_258),
.B(n_267),
.Y(n_257)
);

MAJIxp5_ASAP7_75t_L g350 ( 
.A(n_258),
.B(n_268),
.C(n_269),
.Y(n_350)
);

INVx1_ASAP7_75t_L g259 ( 
.A(n_260),
.Y(n_259)
);

INVx2_ASAP7_75t_SL g266 ( 
.A(n_261),
.Y(n_266)
);

INVx3_ASAP7_75t_L g438 ( 
.A(n_262),
.Y(n_438)
);

INVx2_ASAP7_75t_L g262 ( 
.A(n_263),
.Y(n_262)
);

INVx2_ASAP7_75t_L g263 ( 
.A(n_264),
.Y(n_263)
);

INVx2_ASAP7_75t_L g304 ( 
.A(n_264),
.Y(n_304)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_265),
.Y(n_264)
);

XNOR2x1_ASAP7_75t_L g267 ( 
.A(n_268),
.B(n_269),
.Y(n_267)
);

XNOR2x1_ASAP7_75t_L g269 ( 
.A(n_270),
.B(n_274),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g342 ( 
.A(n_270),
.B(n_275),
.C(n_279),
.Y(n_342)
);

INVx4_ASAP7_75t_L g271 ( 
.A(n_272),
.Y(n_271)
);

INVx6_ASAP7_75t_L g272 ( 
.A(n_273),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g315 ( 
.A(n_273),
.Y(n_315)
);

BUFx2_ASAP7_75t_L g434 ( 
.A(n_273),
.Y(n_434)
);

XNOR2x1_ASAP7_75t_L g274 ( 
.A(n_275),
.B(n_279),
.Y(n_274)
);

INVx2_ASAP7_75t_L g276 ( 
.A(n_277),
.Y(n_276)
);

INVx4_ASAP7_75t_L g277 ( 
.A(n_278),
.Y(n_277)
);

BUFx6f_ASAP7_75t_L g280 ( 
.A(n_281),
.Y(n_280)
);

INVx2_ASAP7_75t_L g482 ( 
.A(n_281),
.Y(n_482)
);

INVx4_ASAP7_75t_L g281 ( 
.A(n_282),
.Y(n_281)
);

INVx6_ASAP7_75t_L g282 ( 
.A(n_283),
.Y(n_282)
);

BUFx6f_ASAP7_75t_L g348 ( 
.A(n_283),
.Y(n_348)
);

INVx2_ASAP7_75t_L g403 ( 
.A(n_283),
.Y(n_403)
);

MAJIxp5_ASAP7_75t_L g286 ( 
.A(n_287),
.B(n_291),
.C(n_294),
.Y(n_286)
);

AOI22xp5_ASAP7_75t_SL g420 ( 
.A1(n_287),
.A2(n_288),
.B1(n_291),
.B2(n_421),
.Y(n_420)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_288),
.Y(n_287)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_291),
.Y(n_421)
);

XOR2x2_ASAP7_75t_L g291 ( 
.A(n_292),
.B(n_293),
.Y(n_291)
);

INVxp67_ASAP7_75t_SL g294 ( 
.A(n_295),
.Y(n_294)
);

XNOR2xp5_ASAP7_75t_L g419 ( 
.A(n_295),
.B(n_420),
.Y(n_419)
);

MAJIxp5_ASAP7_75t_L g295 ( 
.A(n_296),
.B(n_320),
.C(n_323),
.Y(n_295)
);

XNOR2xp5_ASAP7_75t_SL g415 ( 
.A(n_296),
.B(n_416),
.Y(n_415)
);

MAJIxp5_ASAP7_75t_L g296 ( 
.A(n_297),
.B(n_301),
.C(n_310),
.Y(n_296)
);

INVx1_ASAP7_75t_L g297 ( 
.A(n_298),
.Y(n_297)
);

XNOR2xp5_ASAP7_75t_L g407 ( 
.A(n_298),
.B(n_408),
.Y(n_407)
);

XNOR2xp5_ASAP7_75t_L g408 ( 
.A(n_301),
.B(n_310),
.Y(n_408)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_302),
.B(n_306),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g405 ( 
.A(n_302),
.B(n_306),
.Y(n_405)
);

NOR2xp33_ASAP7_75t_L g302 ( 
.A(n_303),
.B(n_305),
.Y(n_302)
);

INVx2_ASAP7_75t_L g303 ( 
.A(n_304),
.Y(n_303)
);

INVx2_ASAP7_75t_L g307 ( 
.A(n_308),
.Y(n_307)
);

INVx2_ASAP7_75t_L g308 ( 
.A(n_309),
.Y(n_308)
);

MAJIxp5_ASAP7_75t_L g310 ( 
.A(n_311),
.B(n_314),
.C(n_316),
.Y(n_310)
);

XNOR2xp5_ASAP7_75t_SL g393 ( 
.A(n_311),
.B(n_314),
.Y(n_393)
);

INVx3_ASAP7_75t_L g312 ( 
.A(n_313),
.Y(n_312)
);

XNOR2xp5_ASAP7_75t_SL g479 ( 
.A(n_314),
.B(n_480),
.Y(n_479)
);

MAJIxp5_ASAP7_75t_L g503 ( 
.A(n_314),
.B(n_476),
.C(n_504),
.Y(n_503)
);

XOR2x1_ASAP7_75t_SL g392 ( 
.A(n_316),
.B(n_393),
.Y(n_392)
);

INVx3_ASAP7_75t_L g317 ( 
.A(n_318),
.Y(n_317)
);

INVx5_ASAP7_75t_L g318 ( 
.A(n_319),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g416 ( 
.A(n_320),
.B(n_323),
.Y(n_416)
);

OAI21xp5_ASAP7_75t_L g530 ( 
.A1(n_326),
.A2(n_531),
.B(n_532),
.Y(n_530)
);

AND2x2_ASAP7_75t_SL g326 ( 
.A(n_327),
.B(n_358),
.Y(n_326)
);

OR2x2_ASAP7_75t_L g532 ( 
.A(n_327),
.B(n_358),
.Y(n_532)
);

XOR2xp5_ASAP7_75t_L g327 ( 
.A(n_328),
.B(n_330),
.Y(n_327)
);

MAJIxp5_ASAP7_75t_L g568 ( 
.A(n_328),
.B(n_569),
.C(n_570),
.Y(n_568)
);

XNOR2x1_ASAP7_75t_L g330 ( 
.A(n_331),
.B(n_349),
.Y(n_330)
);

HB1xp67_ASAP7_75t_L g570 ( 
.A(n_331),
.Y(n_570)
);

XNOR2xp5_ASAP7_75t_L g331 ( 
.A(n_332),
.B(n_341),
.Y(n_331)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_333),
.Y(n_332)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_333),
.B(n_342),
.C(n_343),
.Y(n_538)
);

XOR2xp5_ASAP7_75t_L g333 ( 
.A(n_334),
.B(n_339),
.Y(n_333)
);

INVx4_ASAP7_75t_L g335 ( 
.A(n_336),
.Y(n_335)
);

INVx2_ASAP7_75t_L g336 ( 
.A(n_337),
.Y(n_336)
);

INVx1_ASAP7_75t_L g337 ( 
.A(n_338),
.Y(n_337)
);

XNOR2xp5_ASAP7_75t_L g341 ( 
.A(n_342),
.B(n_343),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g343 ( 
.A(n_344),
.B(n_345),
.Y(n_343)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_344),
.B(n_346),
.C(n_347),
.Y(n_547)
);

XNOR2xp5_ASAP7_75t_L g345 ( 
.A(n_346),
.B(n_347),
.Y(n_345)
);

HB1xp67_ASAP7_75t_L g569 ( 
.A(n_349),
.Y(n_569)
);

XNOR2x1_ASAP7_75t_L g349 ( 
.A(n_350),
.B(n_351),
.Y(n_349)
);

INVxp33_ASAP7_75t_SL g565 ( 
.A(n_350),
.Y(n_565)
);

XNOR2xp5_ASAP7_75t_L g351 ( 
.A(n_352),
.B(n_357),
.Y(n_351)
);

HB1xp67_ASAP7_75t_L g566 ( 
.A(n_352),
.Y(n_566)
);

AOI22xp5_ASAP7_75t_L g352 ( 
.A1(n_353),
.A2(n_354),
.B1(n_355),
.B2(n_356),
.Y(n_352)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_353),
.Y(n_355)
);

INVx1_ASAP7_75t_SL g356 ( 
.A(n_354),
.Y(n_356)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_357),
.B(n_565),
.C(n_566),
.Y(n_564)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_361),
.B(n_526),
.Y(n_360)
);

NAND3xp33_ASAP7_75t_SL g361 ( 
.A(n_362),
.B(n_417),
.C(n_422),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_L g362 ( 
.A(n_363),
.B(n_409),
.Y(n_362)
);

NOR2xp67_ASAP7_75t_L g529 ( 
.A(n_363),
.B(n_409),
.Y(n_529)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_364),
.B(n_391),
.C(n_406),
.Y(n_363)
);

XNOR2xp5_ASAP7_75t_L g523 ( 
.A(n_364),
.B(n_524),
.Y(n_523)
);

XOR2xp5_ASAP7_75t_L g364 ( 
.A(n_365),
.B(n_376),
.Y(n_364)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_365),
.B(n_377),
.C(n_387),
.Y(n_411)
);

XNOR2xp5_ASAP7_75t_SL g515 ( 
.A(n_366),
.B(n_516),
.Y(n_515)
);

AND2x2_ASAP7_75t_L g366 ( 
.A(n_367),
.B(n_370),
.Y(n_366)
);

XNOR2x1_ASAP7_75t_SL g460 ( 
.A(n_367),
.B(n_370),
.Y(n_460)
);

INVx1_ASAP7_75t_L g470 ( 
.A(n_367),
.Y(n_470)
);

AOI22xp5_ASAP7_75t_L g491 ( 
.A1(n_367),
.A2(n_470),
.B1(n_471),
.B2(n_492),
.Y(n_491)
);

INVx2_ASAP7_75t_L g368 ( 
.A(n_369),
.Y(n_368)
);

BUFx3_ASAP7_75t_L g371 ( 
.A(n_372),
.Y(n_371)
);

INVx3_ASAP7_75t_L g386 ( 
.A(n_372),
.Y(n_386)
);

INVx1_ASAP7_75t_L g373 ( 
.A(n_374),
.Y(n_373)
);

XNOR2xp5_ASAP7_75t_L g376 ( 
.A(n_377),
.B(n_387),
.Y(n_376)
);

INVx1_ASAP7_75t_L g379 ( 
.A(n_380),
.Y(n_379)
);

HB1xp67_ASAP7_75t_L g380 ( 
.A(n_381),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_383),
.B(n_384),
.Y(n_382)
);

INVx1_ASAP7_75t_L g384 ( 
.A(n_385),
.Y(n_384)
);

INVx1_ASAP7_75t_L g385 ( 
.A(n_386),
.Y(n_385)
);

MAJIxp5_ASAP7_75t_L g453 ( 
.A(n_389),
.B(n_429),
.C(n_433),
.Y(n_453)
);

XNOR2xp5_ASAP7_75t_L g524 ( 
.A(n_391),
.B(n_407),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g391 ( 
.A(n_392),
.B(n_394),
.C(n_404),
.Y(n_391)
);

XOR2xp5_ASAP7_75t_L g510 ( 
.A(n_392),
.B(n_511),
.Y(n_510)
);

INVxp67_ASAP7_75t_SL g394 ( 
.A(n_395),
.Y(n_394)
);

XNOR2xp5_ASAP7_75t_L g511 ( 
.A(n_395),
.B(n_405),
.Y(n_511)
);

INVx1_ASAP7_75t_L g456 ( 
.A(n_396),
.Y(n_456)
);

INVx2_ASAP7_75t_L g397 ( 
.A(n_398),
.Y(n_397)
);

INVx1_ASAP7_75t_L g398 ( 
.A(n_399),
.Y(n_398)
);

XOR2x2_ASAP7_75t_L g454 ( 
.A(n_400),
.B(n_455),
.Y(n_454)
);

BUFx2_ASAP7_75t_L g401 ( 
.A(n_402),
.Y(n_401)
);

INVx5_ASAP7_75t_L g402 ( 
.A(n_403),
.Y(n_402)
);

INVx1_ASAP7_75t_L g404 ( 
.A(n_405),
.Y(n_404)
);

HB1xp67_ASAP7_75t_L g406 ( 
.A(n_407),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g409 ( 
.A(n_410),
.B(n_415),
.Y(n_409)
);

XNOR2xp5_ASAP7_75t_L g410 ( 
.A(n_411),
.B(n_412),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g418 ( 
.A(n_411),
.B(n_412),
.C(n_415),
.Y(n_418)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_418),
.B(n_419),
.Y(n_417)
);

INVx1_ASAP7_75t_L g528 ( 
.A(n_418),
.Y(n_528)
);

INVx1_ASAP7_75t_L g527 ( 
.A(n_419),
.Y(n_527)
);

OAI21xp5_ASAP7_75t_SL g422 ( 
.A1(n_423),
.A2(n_521),
.B(n_525),
.Y(n_422)
);

AOI21xp5_ASAP7_75t_L g423 ( 
.A1(n_424),
.A2(n_507),
.B(n_520),
.Y(n_423)
);

OAI21x1_ASAP7_75t_SL g424 ( 
.A1(n_425),
.A2(n_466),
.B(n_506),
.Y(n_424)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_426),
.B(n_451),
.Y(n_425)
);

OR2x2_ASAP7_75t_L g506 ( 
.A(n_426),
.B(n_451),
.Y(n_506)
);

MAJIxp5_ASAP7_75t_L g426 ( 
.A(n_427),
.B(n_435),
.C(n_442),
.Y(n_426)
);

XOR2xp5_ASAP7_75t_L g500 ( 
.A(n_427),
.B(n_501),
.Y(n_500)
);

XNOR2xp5_ASAP7_75t_L g428 ( 
.A(n_429),
.B(n_433),
.Y(n_428)
);

INVx1_ASAP7_75t_L g430 ( 
.A(n_431),
.Y(n_430)
);

INVx1_ASAP7_75t_L g431 ( 
.A(n_432),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g501 ( 
.A1(n_435),
.A2(n_436),
.B1(n_442),
.B2(n_502),
.Y(n_501)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_436),
.Y(n_435)
);

NAND2xp5_ASAP7_75t_L g436 ( 
.A(n_437),
.B(n_439),
.Y(n_436)
);

XNOR2xp5_ASAP7_75t_SL g477 ( 
.A(n_437),
.B(n_439),
.Y(n_477)
);

BUFx3_ASAP7_75t_L g440 ( 
.A(n_441),
.Y(n_440)
);

INVx3_ASAP7_75t_L g448 ( 
.A(n_441),
.Y(n_448)
);

INVx1_ASAP7_75t_L g502 ( 
.A(n_442),
.Y(n_502)
);

AO22x1_ASAP7_75t_SL g442 ( 
.A1(n_443),
.A2(n_446),
.B1(n_449),
.B2(n_450),
.Y(n_442)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_443),
.Y(n_449)
);

INVx2_ASAP7_75t_L g444 ( 
.A(n_445),
.Y(n_444)
);

INVx1_ASAP7_75t_SL g450 ( 
.A(n_446),
.Y(n_450)
);

NAND2xp5_ASAP7_75t_SL g458 ( 
.A(n_446),
.B(n_449),
.Y(n_458)
);

INVx4_ASAP7_75t_L g447 ( 
.A(n_448),
.Y(n_447)
);

INVx5_ASAP7_75t_L g474 ( 
.A(n_448),
.Y(n_474)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_450),
.B(n_494),
.Y(n_493)
);

XOR2xp5_ASAP7_75t_L g451 ( 
.A(n_452),
.B(n_457),
.Y(n_451)
);

XNOR2xp5_ASAP7_75t_L g452 ( 
.A(n_453),
.B(n_454),
.Y(n_452)
);

MAJIxp5_ASAP7_75t_L g519 ( 
.A(n_453),
.B(n_454),
.C(n_457),
.Y(n_519)
);

XOR2xp5_ASAP7_75t_L g457 ( 
.A(n_458),
.B(n_459),
.Y(n_457)
);

MAJx2_ASAP7_75t_L g518 ( 
.A(n_458),
.B(n_460),
.C(n_461),
.Y(n_518)
);

XNOR2xp5_ASAP7_75t_L g459 ( 
.A(n_460),
.B(n_461),
.Y(n_459)
);

INVx2_ASAP7_75t_L g462 ( 
.A(n_463),
.Y(n_462)
);

INVx4_ASAP7_75t_L g463 ( 
.A(n_464),
.Y(n_463)
);

INVx3_ASAP7_75t_L g464 ( 
.A(n_465),
.Y(n_464)
);

AOI21xp5_ASAP7_75t_L g466 ( 
.A1(n_467),
.A2(n_499),
.B(n_505),
.Y(n_466)
);

OAI21xp5_ASAP7_75t_SL g467 ( 
.A1(n_468),
.A2(n_483),
.B(n_498),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g468 ( 
.A(n_469),
.B(n_475),
.Y(n_468)
);

NAND2xp33_ASAP7_75t_SL g498 ( 
.A(n_469),
.B(n_475),
.Y(n_498)
);

NOR2xp33_ASAP7_75t_SL g469 ( 
.A(n_470),
.B(n_471),
.Y(n_469)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_471),
.Y(n_492)
);

INVx5_ASAP7_75t_L g472 ( 
.A(n_473),
.Y(n_472)
);

INVx6_ASAP7_75t_L g473 ( 
.A(n_474),
.Y(n_473)
);

OAI22xp5_ASAP7_75t_SL g475 ( 
.A1(n_476),
.A2(n_477),
.B1(n_478),
.B2(n_479),
.Y(n_475)
);

INVx1_ASAP7_75t_L g476 ( 
.A(n_477),
.Y(n_476)
);

INVx1_ASAP7_75t_L g478 ( 
.A(n_479),
.Y(n_478)
);

INVx1_ASAP7_75t_L g504 ( 
.A(n_480),
.Y(n_504)
);

INVx2_ASAP7_75t_L g481 ( 
.A(n_482),
.Y(n_481)
);

AOI21xp5_ASAP7_75t_L g483 ( 
.A1(n_484),
.A2(n_493),
.B(n_497),
.Y(n_483)
);

NAND2xp5_ASAP7_75t_L g484 ( 
.A(n_485),
.B(n_491),
.Y(n_484)
);

NOR2xp33_ASAP7_75t_L g497 ( 
.A(n_485),
.B(n_491),
.Y(n_497)
);

INVx1_ASAP7_75t_SL g486 ( 
.A(n_487),
.Y(n_486)
);

INVx1_ASAP7_75t_L g487 ( 
.A(n_488),
.Y(n_487)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_489),
.Y(n_488)
);

INVx2_ASAP7_75t_L g489 ( 
.A(n_490),
.Y(n_489)
);

INVx4_ASAP7_75t_L g495 ( 
.A(n_496),
.Y(n_495)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_500),
.B(n_503),
.Y(n_499)
);

NOR2xp33_ASAP7_75t_L g505 ( 
.A(n_500),
.B(n_503),
.Y(n_505)
);

NAND2xp5_ASAP7_75t_SL g507 ( 
.A(n_508),
.B(n_519),
.Y(n_507)
);

NOR2xp67_ASAP7_75t_L g520 ( 
.A(n_508),
.B(n_519),
.Y(n_520)
);

AOI22xp5_ASAP7_75t_L g508 ( 
.A1(n_509),
.A2(n_510),
.B1(n_512),
.B2(n_513),
.Y(n_508)
);

MAJIxp5_ASAP7_75t_L g522 ( 
.A(n_509),
.B(n_514),
.C(n_518),
.Y(n_522)
);

INVx1_ASAP7_75t_L g509 ( 
.A(n_510),
.Y(n_509)
);

INVx1_ASAP7_75t_L g512 ( 
.A(n_513),
.Y(n_512)
);

AOI22xp5_ASAP7_75t_L g513 ( 
.A1(n_514),
.A2(n_515),
.B1(n_517),
.B2(n_518),
.Y(n_513)
);

INVx1_ASAP7_75t_L g514 ( 
.A(n_515),
.Y(n_514)
);

INVx1_ASAP7_75t_L g517 ( 
.A(n_518),
.Y(n_517)
);

NOR2xp67_ASAP7_75t_SL g521 ( 
.A(n_522),
.B(n_523),
.Y(n_521)
);

NAND2xp5_ASAP7_75t_L g525 ( 
.A(n_522),
.B(n_523),
.Y(n_525)
);

MAJIxp5_ASAP7_75t_L g526 ( 
.A(n_527),
.B(n_528),
.C(n_529),
.Y(n_526)
);

NOR3xp33_ASAP7_75t_SL g533 ( 
.A(n_534),
.B(n_553),
.C(n_567),
.Y(n_533)
);

OAI21xp5_ASAP7_75t_SL g574 ( 
.A1(n_534),
.A2(n_575),
.B(n_578),
.Y(n_574)
);

NOR2xp67_ASAP7_75t_SL g534 ( 
.A(n_535),
.B(n_551),
.Y(n_534)
);

NAND2xp5_ASAP7_75t_L g578 ( 
.A(n_535),
.B(n_551),
.Y(n_578)
);

MAJIxp5_ASAP7_75t_L g535 ( 
.A(n_536),
.B(n_543),
.C(n_548),
.Y(n_535)
);

XNOR2xp5_ASAP7_75t_L g555 ( 
.A(n_536),
.B(n_556),
.Y(n_555)
);

MAJIxp5_ASAP7_75t_L g536 ( 
.A(n_537),
.B(n_539),
.C(n_542),
.Y(n_536)
);

INVxp33_ASAP7_75t_L g537 ( 
.A(n_538),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g560 ( 
.A(n_538),
.B(n_561),
.Y(n_560)
);

HB1xp67_ASAP7_75t_L g539 ( 
.A(n_540),
.Y(n_539)
);

XNOR2xp5_ASAP7_75t_L g561 ( 
.A(n_540),
.B(n_542),
.Y(n_561)
);

AOI22xp5_ASAP7_75t_L g556 ( 
.A1(n_543),
.A2(n_548),
.B1(n_549),
.B2(n_557),
.Y(n_556)
);

INVxp67_ASAP7_75t_SL g557 ( 
.A(n_543),
.Y(n_557)
);

MAJIxp5_ASAP7_75t_L g543 ( 
.A(n_544),
.B(n_546),
.C(n_547),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_544),
.B(n_563),
.Y(n_562)
);

XNOR2xp5_ASAP7_75t_L g563 ( 
.A(n_546),
.B(n_547),
.Y(n_563)
);

INVx1_ASAP7_75t_L g548 ( 
.A(n_549),
.Y(n_548)
);

INVx1_ASAP7_75t_L g553 ( 
.A(n_554),
.Y(n_553)
);

AOI21xp5_ASAP7_75t_L g575 ( 
.A1(n_554),
.A2(n_576),
.B(n_577),
.Y(n_575)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_555),
.B(n_558),
.Y(n_554)
);

NOR2xp33_ASAP7_75t_L g577 ( 
.A(n_555),
.B(n_558),
.Y(n_577)
);

MAJIxp5_ASAP7_75t_L g558 ( 
.A(n_559),
.B(n_562),
.C(n_564),
.Y(n_558)
);

AOI22xp5_ASAP7_75t_L g572 ( 
.A1(n_559),
.A2(n_560),
.B1(n_562),
.B2(n_573),
.Y(n_572)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_560),
.Y(n_559)
);

INVx1_ASAP7_75t_L g573 ( 
.A(n_562),
.Y(n_573)
);

XOR2xp5_ASAP7_75t_L g571 ( 
.A(n_564),
.B(n_572),
.Y(n_571)
);

AND2x2_ASAP7_75t_L g567 ( 
.A(n_568),
.B(n_571),
.Y(n_567)
);

NOR2xp33_ASAP7_75t_L g576 ( 
.A(n_568),
.B(n_571),
.Y(n_576)
);

NOR2xp33_ASAP7_75t_SL g580 ( 
.A(n_581),
.B(n_590),
.Y(n_580)
);

NOR2xp67_ASAP7_75t_R g581 ( 
.A(n_582),
.B(n_589),
.Y(n_581)
);

AND2x2_ASAP7_75t_L g590 ( 
.A(n_582),
.B(n_589),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_583),
.B(n_584),
.Y(n_582)
);

CKINVDCx20_ASAP7_75t_R g588 ( 
.A(n_585),
.Y(n_588)
);

INVx2_ASAP7_75t_L g586 ( 
.A(n_587),
.Y(n_586)
);


endmodule