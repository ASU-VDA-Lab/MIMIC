module fake_jpeg_29075_n_455 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_455);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_455;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_265;
wire n_192;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_84;
wire n_59;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_378;
wire n_132;
wire n_133;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_412;
wire n_249;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx6f_ASAP7_75t_L g19 ( 
.A(n_5),
.Y(n_19)
);

BUFx5_ASAP7_75t_L g20 ( 
.A(n_10),
.Y(n_20)
);

BUFx12f_ASAP7_75t_L g21 ( 
.A(n_14),
.Y(n_21)
);

BUFx6f_ASAP7_75t_L g22 ( 
.A(n_4),
.Y(n_22)
);

INVx4_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx1_ASAP7_75t_L g25 ( 
.A(n_18),
.Y(n_25)
);

INVx1_ASAP7_75t_L g26 ( 
.A(n_9),
.Y(n_26)
);

INVx1_ASAP7_75t_L g27 ( 
.A(n_5),
.Y(n_27)
);

INVx4_ASAP7_75t_L g28 ( 
.A(n_6),
.Y(n_28)
);

INVx11_ASAP7_75t_SL g29 ( 
.A(n_14),
.Y(n_29)
);

INVx8_ASAP7_75t_L g30 ( 
.A(n_10),
.Y(n_30)
);

INVx1_ASAP7_75t_L g31 ( 
.A(n_3),
.Y(n_31)
);

BUFx6f_ASAP7_75t_L g32 ( 
.A(n_9),
.Y(n_32)
);

INVx6_ASAP7_75t_L g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_1),
.Y(n_34)
);

INVx6_ASAP7_75t_SL g35 ( 
.A(n_6),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_17),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_18),
.Y(n_37)
);

BUFx4f_ASAP7_75t_L g38 ( 
.A(n_16),
.Y(n_38)
);

BUFx12f_ASAP7_75t_L g39 ( 
.A(n_18),
.Y(n_39)
);

INVx2_ASAP7_75t_L g40 ( 
.A(n_16),
.Y(n_40)
);

BUFx6f_ASAP7_75t_L g41 ( 
.A(n_7),
.Y(n_41)
);

INVx1_ASAP7_75t_L g42 ( 
.A(n_2),
.Y(n_42)
);

INVx1_ASAP7_75t_L g43 ( 
.A(n_7),
.Y(n_43)
);

BUFx6f_ASAP7_75t_L g44 ( 
.A(n_16),
.Y(n_44)
);

CKINVDCx16_ASAP7_75t_R g45 ( 
.A(n_14),
.Y(n_45)
);

BUFx10_ASAP7_75t_L g46 ( 
.A(n_5),
.Y(n_46)
);

INVx6_ASAP7_75t_SL g47 ( 
.A(n_29),
.Y(n_47)
);

INVx13_ASAP7_75t_L g110 ( 
.A(n_47),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_29),
.Y(n_48)
);

NAND2xp5_ASAP7_75t_SL g93 ( 
.A(n_48),
.B(n_54),
.Y(n_93)
);

INVx2_ASAP7_75t_SL g49 ( 
.A(n_38),
.Y(n_49)
);

INVxp67_ASAP7_75t_L g133 ( 
.A(n_49),
.Y(n_133)
);

INVx2_ASAP7_75t_L g50 ( 
.A(n_40),
.Y(n_50)
);

INVx2_ASAP7_75t_L g96 ( 
.A(n_50),
.Y(n_96)
);

INVx1_ASAP7_75t_L g51 ( 
.A(n_40),
.Y(n_51)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_51),
.Y(n_100)
);

INVx8_ASAP7_75t_L g52 ( 
.A(n_20),
.Y(n_52)
);

INVx11_ASAP7_75t_L g130 ( 
.A(n_52),
.Y(n_130)
);

BUFx6f_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

BUFx6f_ASAP7_75t_L g94 ( 
.A(n_53),
.Y(n_94)
);

CKINVDCx20_ASAP7_75t_R g54 ( 
.A(n_38),
.Y(n_54)
);

INVx11_ASAP7_75t_L g55 ( 
.A(n_30),
.Y(n_55)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_55),
.Y(n_95)
);

INVx1_ASAP7_75t_L g56 ( 
.A(n_25),
.Y(n_56)
);

INVx1_ASAP7_75t_L g125 ( 
.A(n_56),
.Y(n_125)
);

INVx4_ASAP7_75t_L g57 ( 
.A(n_23),
.Y(n_57)
);

INVx4_ASAP7_75t_L g116 ( 
.A(n_57),
.Y(n_116)
);

BUFx24_ASAP7_75t_L g58 ( 
.A(n_38),
.Y(n_58)
);

BUFx12f_ASAP7_75t_L g103 ( 
.A(n_58),
.Y(n_103)
);

BUFx6f_ASAP7_75t_L g59 ( 
.A(n_19),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g97 ( 
.A(n_59),
.Y(n_97)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_23),
.Y(n_60)
);

INVx2_ASAP7_75t_L g104 ( 
.A(n_60),
.Y(n_104)
);

INVx13_ASAP7_75t_L g61 ( 
.A(n_30),
.Y(n_61)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_61),
.Y(n_131)
);

NOR2xp33_ASAP7_75t_SL g62 ( 
.A(n_37),
.B(n_17),
.Y(n_62)
);

NOR2xp33_ASAP7_75t_SL g140 ( 
.A(n_62),
.B(n_13),
.Y(n_140)
);

INVx3_ASAP7_75t_L g63 ( 
.A(n_21),
.Y(n_63)
);

INVx3_ASAP7_75t_L g101 ( 
.A(n_63),
.Y(n_101)
);

BUFx4f_ASAP7_75t_SL g64 ( 
.A(n_38),
.Y(n_64)
);

BUFx12f_ASAP7_75t_L g137 ( 
.A(n_64),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_19),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_65),
.Y(n_111)
);

BUFx6f_ASAP7_75t_L g66 ( 
.A(n_19),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g118 ( 
.A(n_66),
.Y(n_118)
);

INVx2_ASAP7_75t_L g67 ( 
.A(n_23),
.Y(n_67)
);

INVx2_ASAP7_75t_L g107 ( 
.A(n_67),
.Y(n_107)
);

INVx2_ASAP7_75t_L g68 ( 
.A(n_24),
.Y(n_68)
);

INVx2_ASAP7_75t_L g109 ( 
.A(n_68),
.Y(n_109)
);

BUFx12f_ASAP7_75t_L g69 ( 
.A(n_22),
.Y(n_69)
);

INVx3_ASAP7_75t_L g117 ( 
.A(n_69),
.Y(n_117)
);

INVx3_ASAP7_75t_L g70 ( 
.A(n_21),
.Y(n_70)
);

INVx3_ASAP7_75t_L g129 ( 
.A(n_70),
.Y(n_129)
);

NOR2xp33_ASAP7_75t_L g71 ( 
.A(n_37),
.B(n_17),
.Y(n_71)
);

AND2x2_ASAP7_75t_L g106 ( 
.A(n_71),
.B(n_87),
.Y(n_106)
);

INVx4_ASAP7_75t_L g72 ( 
.A(n_24),
.Y(n_72)
);

INVx4_ASAP7_75t_L g126 ( 
.A(n_72),
.Y(n_126)
);

INVx11_ASAP7_75t_L g73 ( 
.A(n_30),
.Y(n_73)
);

INVx5_ASAP7_75t_L g128 ( 
.A(n_73),
.Y(n_128)
);

INVx3_ASAP7_75t_L g74 ( 
.A(n_21),
.Y(n_74)
);

INVx5_ASAP7_75t_L g135 ( 
.A(n_74),
.Y(n_135)
);

NAND2xp5_ASAP7_75t_SL g75 ( 
.A(n_45),
.B(n_15),
.Y(n_75)
);

NAND2xp5_ASAP7_75t_L g105 ( 
.A(n_75),
.B(n_15),
.Y(n_105)
);

INVx3_ASAP7_75t_L g76 ( 
.A(n_21),
.Y(n_76)
);

INVx4_ASAP7_75t_L g98 ( 
.A(n_76),
.Y(n_98)
);

INVx4_ASAP7_75t_L g77 ( 
.A(n_24),
.Y(n_77)
);

INVx4_ASAP7_75t_L g119 ( 
.A(n_77),
.Y(n_119)
);

BUFx3_ASAP7_75t_L g78 ( 
.A(n_20),
.Y(n_78)
);

BUFx3_ASAP7_75t_L g120 ( 
.A(n_78),
.Y(n_120)
);

INVx4_ASAP7_75t_L g79 ( 
.A(n_28),
.Y(n_79)
);

INVx2_ASAP7_75t_L g112 ( 
.A(n_79),
.Y(n_112)
);

BUFx6f_ASAP7_75t_L g80 ( 
.A(n_22),
.Y(n_80)
);

INVx8_ASAP7_75t_L g142 ( 
.A(n_80),
.Y(n_142)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_25),
.Y(n_81)
);

INVx1_ASAP7_75t_L g138 ( 
.A(n_81),
.Y(n_138)
);

INVx13_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g139 ( 
.A(n_82),
.Y(n_139)
);

BUFx12f_ASAP7_75t_L g83 ( 
.A(n_22),
.Y(n_83)
);

BUFx3_ASAP7_75t_L g123 ( 
.A(n_83),
.Y(n_123)
);

BUFx12f_ASAP7_75t_L g84 ( 
.A(n_22),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g127 ( 
.A(n_84),
.Y(n_127)
);

INVx2_ASAP7_75t_L g85 ( 
.A(n_28),
.Y(n_85)
);

INVx2_ASAP7_75t_L g113 ( 
.A(n_85),
.Y(n_113)
);

INVx1_ASAP7_75t_L g86 ( 
.A(n_36),
.Y(n_86)
);

CKINVDCx16_ASAP7_75t_R g121 ( 
.A(n_86),
.Y(n_121)
);

NOR2xp33_ASAP7_75t_L g87 ( 
.A(n_45),
.B(n_15),
.Y(n_87)
);

INVx8_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

BUFx3_ASAP7_75t_L g136 ( 
.A(n_88),
.Y(n_136)
);

INVx6_ASAP7_75t_L g89 ( 
.A(n_32),
.Y(n_89)
);

INVx2_ASAP7_75t_L g114 ( 
.A(n_89),
.Y(n_114)
);

BUFx3_ASAP7_75t_L g90 ( 
.A(n_32),
.Y(n_90)
);

INVx2_ASAP7_75t_L g115 ( 
.A(n_90),
.Y(n_115)
);

AND2x2_ASAP7_75t_SL g91 ( 
.A(n_28),
.B(n_0),
.Y(n_91)
);

A2O1A1Ixp33_ASAP7_75t_L g132 ( 
.A1(n_91),
.A2(n_34),
.B(n_43),
.C(n_42),
.Y(n_132)
);

BUFx6f_ASAP7_75t_L g92 ( 
.A(n_32),
.Y(n_92)
);

INVx2_ASAP7_75t_L g122 ( 
.A(n_92),
.Y(n_122)
);

OAI22xp5_ASAP7_75t_L g99 ( 
.A1(n_91),
.A2(n_44),
.B1(n_33),
.B2(n_36),
.Y(n_99)
);

AOI22xp5_ASAP7_75t_L g161 ( 
.A1(n_99),
.A2(n_108),
.B1(n_41),
.B2(n_65),
.Y(n_161)
);

BUFx4f_ASAP7_75t_L g102 ( 
.A(n_58),
.Y(n_102)
);

INVx2_ASAP7_75t_SL g173 ( 
.A(n_102),
.Y(n_173)
);

NOR2xp33_ASAP7_75t_L g144 ( 
.A(n_105),
.B(n_134),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_L g108 ( 
.A1(n_53),
.A2(n_44),
.B1(n_33),
.B2(n_32),
.Y(n_108)
);

AOI22xp33_ASAP7_75t_L g124 ( 
.A1(n_89),
.A2(n_33),
.B1(n_44),
.B2(n_41),
.Y(n_124)
);

OAI22xp5_ASAP7_75t_SL g163 ( 
.A1(n_124),
.A2(n_92),
.B1(n_59),
.B2(n_66),
.Y(n_163)
);

A2O1A1Ixp33_ASAP7_75t_L g176 ( 
.A1(n_132),
.A2(n_27),
.B(n_31),
.C(n_43),
.Y(n_176)
);

NAND2xp5_ASAP7_75t_SL g134 ( 
.A(n_63),
.B(n_34),
.Y(n_134)
);

NOR2xp33_ASAP7_75t_L g154 ( 
.A(n_140),
.B(n_13),
.Y(n_154)
);

AOI21xp5_ASAP7_75t_L g141 ( 
.A1(n_78),
.A2(n_13),
.B(n_1),
.Y(n_141)
);

OAI21xp5_ASAP7_75t_L g157 ( 
.A1(n_141),
.A2(n_21),
.B(n_39),
.Y(n_157)
);

BUFx6f_ASAP7_75t_L g143 ( 
.A(n_94),
.Y(n_143)
);

INVx8_ASAP7_75t_L g186 ( 
.A(n_143),
.Y(n_186)
);

INVx1_ASAP7_75t_L g145 ( 
.A(n_100),
.Y(n_145)
);

INVx1_ASAP7_75t_L g187 ( 
.A(n_145),
.Y(n_187)
);

INVx2_ASAP7_75t_L g146 ( 
.A(n_101),
.Y(n_146)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_146),
.Y(n_204)
);

AOI22xp33_ASAP7_75t_SL g147 ( 
.A1(n_125),
.A2(n_35),
.B1(n_57),
.B2(n_77),
.Y(n_147)
);

INVxp67_ASAP7_75t_L g185 ( 
.A(n_147),
.Y(n_185)
);

CKINVDCx9p33_ASAP7_75t_R g148 ( 
.A(n_102),
.Y(n_148)
);

INVxp67_ASAP7_75t_SL g192 ( 
.A(n_148),
.Y(n_192)
);

INVx2_ASAP7_75t_L g149 ( 
.A(n_129),
.Y(n_149)
);

INVx2_ASAP7_75t_L g207 ( 
.A(n_149),
.Y(n_207)
);

BUFx10_ASAP7_75t_L g150 ( 
.A(n_131),
.Y(n_150)
);

CKINVDCx20_ASAP7_75t_R g183 ( 
.A(n_150),
.Y(n_183)
);

BUFx6f_ASAP7_75t_L g151 ( 
.A(n_94),
.Y(n_151)
);

INVx6_ASAP7_75t_L g180 ( 
.A(n_151),
.Y(n_180)
);

INVx8_ASAP7_75t_L g152 ( 
.A(n_95),
.Y(n_152)
);

INVx3_ASAP7_75t_L g196 ( 
.A(n_152),
.Y(n_196)
);

INVx1_ASAP7_75t_L g153 ( 
.A(n_138),
.Y(n_153)
);

INVx1_ASAP7_75t_L g191 ( 
.A(n_153),
.Y(n_191)
);

NOR2xp33_ASAP7_75t_L g181 ( 
.A(n_154),
.B(n_162),
.Y(n_181)
);

INVx2_ASAP7_75t_L g155 ( 
.A(n_112),
.Y(n_155)
);

CKINVDCx14_ASAP7_75t_R g184 ( 
.A(n_155),
.Y(n_184)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_114),
.Y(n_156)
);

INVx1_ASAP7_75t_L g198 ( 
.A(n_156),
.Y(n_198)
);

AND2x2_ASAP7_75t_L g199 ( 
.A(n_157),
.B(n_161),
.Y(n_199)
);

MAJIxp5_ASAP7_75t_L g158 ( 
.A(n_96),
.B(n_72),
.C(n_79),
.Y(n_158)
);

AND2x2_ASAP7_75t_L g189 ( 
.A(n_158),
.B(n_163),
.Y(n_189)
);

AOI22xp33_ASAP7_75t_SL g159 ( 
.A1(n_142),
.A2(n_35),
.B1(n_39),
.B2(n_90),
.Y(n_159)
);

OAI22xp5_ASAP7_75t_L g201 ( 
.A1(n_159),
.A2(n_160),
.B1(n_166),
.B2(n_175),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g160 ( 
.A1(n_142),
.A2(n_35),
.B1(n_39),
.B2(n_70),
.Y(n_160)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_131),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g164 ( 
.A(n_121),
.B(n_106),
.Y(n_164)
);

NAND2xp5_ASAP7_75t_L g182 ( 
.A(n_164),
.B(n_170),
.Y(n_182)
);

INVx1_ASAP7_75t_L g165 ( 
.A(n_93),
.Y(n_165)
);

NOR2xp33_ASAP7_75t_L g206 ( 
.A(n_165),
.B(n_167),
.Y(n_206)
);

OAI22xp5_ASAP7_75t_L g166 ( 
.A1(n_106),
.A2(n_80),
.B1(n_44),
.B2(n_41),
.Y(n_166)
);

INVx3_ASAP7_75t_L g167 ( 
.A(n_131),
.Y(n_167)
);

INVx4_ASAP7_75t_L g168 ( 
.A(n_117),
.Y(n_168)
);

CKINVDCx20_ASAP7_75t_R g188 ( 
.A(n_168),
.Y(n_188)
);

INVx1_ASAP7_75t_L g169 ( 
.A(n_104),
.Y(n_169)
);

CKINVDCx20_ASAP7_75t_R g193 ( 
.A(n_169),
.Y(n_193)
);

NAND2xp5_ASAP7_75t_L g170 ( 
.A(n_107),
.B(n_26),
.Y(n_170)
);

INVx4_ASAP7_75t_L g171 ( 
.A(n_115),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g202 ( 
.A(n_171),
.Y(n_202)
);

INVx2_ASAP7_75t_L g172 ( 
.A(n_122),
.Y(n_172)
);

AND2x2_ASAP7_75t_L g208 ( 
.A(n_172),
.B(n_174),
.Y(n_208)
);

INVx2_ASAP7_75t_L g174 ( 
.A(n_119),
.Y(n_174)
);

OAI22xp5_ASAP7_75t_L g175 ( 
.A1(n_97),
.A2(n_41),
.B1(n_26),
.B2(n_42),
.Y(n_175)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_176),
.B(n_133),
.Y(n_195)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_139),
.Y(n_177)
);

AND2x2_ASAP7_75t_L g194 ( 
.A(n_177),
.B(n_178),
.Y(n_194)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_97),
.Y(n_178)
);

OAI22xp5_ASAP7_75t_SL g179 ( 
.A1(n_124),
.A2(n_49),
.B1(n_73),
.B2(n_55),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g197 ( 
.A(n_179),
.B(n_64),
.Y(n_197)
);

AOI32xp33_ASAP7_75t_L g190 ( 
.A1(n_157),
.A2(n_126),
.A3(n_116),
.B1(n_98),
.B2(n_119),
.Y(n_190)
);

NOR2xp33_ASAP7_75t_L g210 ( 
.A(n_190),
.B(n_195),
.Y(n_210)
);

AND2x2_ASAP7_75t_L g219 ( 
.A(n_197),
.B(n_88),
.Y(n_219)
);

NAND2xp5_ASAP7_75t_L g200 ( 
.A(n_170),
.B(n_109),
.Y(n_200)
);

NAND2xp5_ASAP7_75t_L g211 ( 
.A(n_200),
.B(n_203),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g203 ( 
.A(n_144),
.B(n_113),
.Y(n_203)
);

NAND2xp5_ASAP7_75t_L g205 ( 
.A(n_145),
.B(n_133),
.Y(n_205)
);

NAND2xp5_ASAP7_75t_L g226 ( 
.A(n_205),
.B(n_150),
.Y(n_226)
);

INVx2_ASAP7_75t_L g209 ( 
.A(n_204),
.Y(n_209)
);

INVx2_ASAP7_75t_L g237 ( 
.A(n_209),
.Y(n_237)
);

NOR2xp33_ASAP7_75t_L g212 ( 
.A(n_205),
.B(n_203),
.Y(n_212)
);

NAND2xp5_ASAP7_75t_L g236 ( 
.A(n_212),
.B(n_214),
.Y(n_236)
);

CKINVDCx20_ASAP7_75t_R g213 ( 
.A(n_208),
.Y(n_213)
);

NOR2xp33_ASAP7_75t_L g235 ( 
.A(n_213),
.B(n_222),
.Y(n_235)
);

NAND2xp5_ASAP7_75t_SL g214 ( 
.A(n_200),
.B(n_176),
.Y(n_214)
);

INVx13_ASAP7_75t_L g215 ( 
.A(n_186),
.Y(n_215)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_215),
.Y(n_252)
);

AOI22xp5_ASAP7_75t_SL g216 ( 
.A1(n_185),
.A2(n_179),
.B1(n_153),
.B2(n_163),
.Y(n_216)
);

AOI21xp5_ASAP7_75t_L g251 ( 
.A1(n_216),
.A2(n_194),
.B(n_120),
.Y(n_251)
);

AOI22xp5_ASAP7_75t_L g217 ( 
.A1(n_199),
.A2(n_161),
.B1(n_156),
.B2(n_111),
.Y(n_217)
);

OAI22xp5_ASAP7_75t_SL g246 ( 
.A1(n_217),
.A2(n_184),
.B1(n_191),
.B2(n_188),
.Y(n_246)
);

OAI22xp5_ASAP7_75t_SL g218 ( 
.A1(n_199),
.A2(n_158),
.B1(n_164),
.B2(n_118),
.Y(n_218)
);

AOI22xp5_ASAP7_75t_L g240 ( 
.A1(n_218),
.A2(n_230),
.B1(n_189),
.B2(n_201),
.Y(n_240)
);

NAND2xp5_ASAP7_75t_L g247 ( 
.A(n_219),
.B(n_224),
.Y(n_247)
);

INVx2_ASAP7_75t_L g220 ( 
.A(n_204),
.Y(n_220)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_220),
.Y(n_248)
);

MAJIxp5_ASAP7_75t_L g221 ( 
.A(n_182),
.B(n_155),
.C(n_171),
.Y(n_221)
);

MAJIxp5_ASAP7_75t_L g239 ( 
.A(n_221),
.B(n_189),
.C(n_218),
.Y(n_239)
);

AND2x6_ASAP7_75t_L g222 ( 
.A(n_199),
.B(n_110),
.Y(n_222)
);

INVx13_ASAP7_75t_L g223 ( 
.A(n_186),
.Y(n_223)
);

NOR2xp33_ASAP7_75t_L g256 ( 
.A(n_223),
.B(n_227),
.Y(n_256)
);

NAND2xp5_ASAP7_75t_SL g224 ( 
.A(n_182),
.B(n_172),
.Y(n_224)
);

AO21x2_ASAP7_75t_SL g225 ( 
.A1(n_197),
.A2(n_64),
.B(n_137),
.Y(n_225)
);

AO22x1_ASAP7_75t_L g244 ( 
.A1(n_225),
.A2(n_194),
.B1(n_137),
.B2(n_208),
.Y(n_244)
);

NAND2xp5_ASAP7_75t_SL g238 ( 
.A(n_226),
.B(n_228),
.Y(n_238)
);

INVx13_ASAP7_75t_L g227 ( 
.A(n_186),
.Y(n_227)
);

NOR2xp33_ASAP7_75t_L g228 ( 
.A(n_206),
.B(n_146),
.Y(n_228)
);

BUFx4f_ASAP7_75t_SL g229 ( 
.A(n_183),
.Y(n_229)
);

INVx1_ASAP7_75t_L g250 ( 
.A(n_229),
.Y(n_250)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_189),
.A2(n_111),
.B1(n_118),
.B2(n_151),
.Y(n_230)
);

INVx5_ASAP7_75t_L g231 ( 
.A(n_180),
.Y(n_231)
);

INVx1_ASAP7_75t_L g258 ( 
.A(n_231),
.Y(n_258)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_206),
.B(n_149),
.Y(n_232)
);

XOR2xp5_ASAP7_75t_L g243 ( 
.A(n_232),
.B(n_208),
.Y(n_243)
);

INVx1_ASAP7_75t_L g233 ( 
.A(n_187),
.Y(n_233)
);

AOI22xp5_ASAP7_75t_SL g245 ( 
.A1(n_233),
.A2(n_208),
.B1(n_184),
.B2(n_193),
.Y(n_245)
);

OAI32xp33_ASAP7_75t_L g234 ( 
.A1(n_210),
.A2(n_195),
.A3(n_189),
.B1(n_201),
.B2(n_190),
.Y(n_234)
);

INVx1_ASAP7_75t_L g265 ( 
.A(n_234),
.Y(n_265)
);

XNOR2xp5_ASAP7_75t_L g277 ( 
.A(n_239),
.B(n_241),
.Y(n_277)
);

OAI22xp5_ASAP7_75t_SL g270 ( 
.A1(n_240),
.A2(n_242),
.B1(n_255),
.B2(n_257),
.Y(n_270)
);

XNOR2x1_ASAP7_75t_L g241 ( 
.A(n_221),
.B(n_181),
.Y(n_241)
);

AOI22xp5_ASAP7_75t_L g242 ( 
.A1(n_230),
.A2(n_191),
.B1(n_187),
.B2(n_194),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g276 ( 
.A(n_243),
.B(n_245),
.Y(n_276)
);

AO22x1_ASAP7_75t_L g278 ( 
.A1(n_244),
.A2(n_137),
.B1(n_103),
.B2(n_139),
.Y(n_278)
);

AOI22xp33_ASAP7_75t_L g263 ( 
.A1(n_246),
.A2(n_213),
.B1(n_216),
.B2(n_233),
.Y(n_263)
);

XOR2xp5_ASAP7_75t_L g249 ( 
.A(n_221),
.B(n_181),
.Y(n_249)
);

INVxp67_ASAP7_75t_L g285 ( 
.A(n_249),
.Y(n_285)
);

OAI21xp5_ASAP7_75t_SL g260 ( 
.A1(n_251),
.A2(n_219),
.B(n_226),
.Y(n_260)
);

MAJIxp5_ASAP7_75t_L g253 ( 
.A(n_210),
.B(n_224),
.C(n_211),
.Y(n_253)
);

NOR2xp33_ASAP7_75t_L g279 ( 
.A(n_253),
.B(n_254),
.Y(n_279)
);

MAJIxp5_ASAP7_75t_L g254 ( 
.A(n_211),
.B(n_202),
.C(n_188),
.Y(n_254)
);

OAI22xp5_ASAP7_75t_SL g255 ( 
.A1(n_217),
.A2(n_193),
.B1(n_202),
.B2(n_178),
.Y(n_255)
);

AOI22xp5_ASAP7_75t_L g257 ( 
.A1(n_219),
.A2(n_194),
.B1(n_198),
.B2(n_180),
.Y(n_257)
);

OAI21xp5_ASAP7_75t_L g259 ( 
.A1(n_235),
.A2(n_222),
.B(n_214),
.Y(n_259)
);

OAI21xp5_ASAP7_75t_L g291 ( 
.A1(n_259),
.A2(n_262),
.B(n_247),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g306 ( 
.A1(n_260),
.A2(n_120),
.B(n_177),
.Y(n_306)
);

AND2x6_ASAP7_75t_L g261 ( 
.A(n_244),
.B(n_222),
.Y(n_261)
);

NOR3xp33_ASAP7_75t_L g301 ( 
.A(n_261),
.B(n_162),
.C(n_167),
.Y(n_301)
);

OAI21xp5_ASAP7_75t_L g262 ( 
.A1(n_251),
.A2(n_219),
.B(n_229),
.Y(n_262)
);

OAI22xp5_ASAP7_75t_SL g307 ( 
.A1(n_263),
.A2(n_267),
.B1(n_173),
.B2(n_174),
.Y(n_307)
);

OAI22xp5_ASAP7_75t_L g264 ( 
.A1(n_240),
.A2(n_225),
.B1(n_212),
.B2(n_232),
.Y(n_264)
);

AOI22xp5_ASAP7_75t_L g297 ( 
.A1(n_264),
.A2(n_272),
.B1(n_282),
.B2(n_283),
.Y(n_297)
);

NOR2x1_ASAP7_75t_L g266 ( 
.A(n_244),
.B(n_225),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_L g292 ( 
.A(n_266),
.B(n_274),
.Y(n_292)
);

AOI22xp33_ASAP7_75t_L g267 ( 
.A1(n_255),
.A2(n_228),
.B1(n_225),
.B2(n_231),
.Y(n_267)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_248),
.Y(n_268)
);

INVx1_ASAP7_75t_L g290 ( 
.A(n_268),
.Y(n_290)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_248),
.Y(n_269)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_269),
.Y(n_310)
);

CKINVDCx16_ASAP7_75t_R g271 ( 
.A(n_250),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g298 ( 
.A(n_271),
.B(n_280),
.Y(n_298)
);

OAI22xp5_ASAP7_75t_SL g272 ( 
.A1(n_239),
.A2(n_225),
.B1(n_229),
.B2(n_231),
.Y(n_272)
);

HB1xp67_ASAP7_75t_L g273 ( 
.A(n_250),
.Y(n_273)
);

NOR2xp33_ASAP7_75t_L g308 ( 
.A(n_273),
.B(n_281),
.Y(n_308)
);

NOR2x1_ASAP7_75t_L g274 ( 
.A(n_257),
.B(n_229),
.Y(n_274)
);

NOR2xp33_ASAP7_75t_L g275 ( 
.A(n_238),
.B(n_183),
.Y(n_275)
);

CKINVDCx14_ASAP7_75t_R g293 ( 
.A(n_275),
.Y(n_293)
);

AND2x2_ASAP7_75t_L g313 ( 
.A(n_278),
.B(n_136),
.Y(n_313)
);

NOR2xp33_ASAP7_75t_L g280 ( 
.A(n_236),
.B(n_220),
.Y(n_280)
);

CKINVDCx20_ASAP7_75t_R g281 ( 
.A(n_256),
.Y(n_281)
);

OAI22xp5_ASAP7_75t_L g282 ( 
.A1(n_242),
.A2(n_180),
.B1(n_143),
.B2(n_196),
.Y(n_282)
);

OAI22xp5_ASAP7_75t_L g283 ( 
.A1(n_247),
.A2(n_196),
.B1(n_152),
.B2(n_198),
.Y(n_283)
);

INVx1_ASAP7_75t_L g284 ( 
.A(n_237),
.Y(n_284)
);

INVx1_ASAP7_75t_SL g299 ( 
.A(n_284),
.Y(n_299)
);

INVxp67_ASAP7_75t_SL g286 ( 
.A(n_246),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g312 ( 
.A(n_286),
.B(n_227),
.Y(n_312)
);

OAI22xp5_ASAP7_75t_SL g287 ( 
.A1(n_234),
.A2(n_209),
.B1(n_207),
.B2(n_136),
.Y(n_287)
);

AOI22xp5_ASAP7_75t_L g300 ( 
.A1(n_287),
.A2(n_243),
.B1(n_258),
.B2(n_252),
.Y(n_300)
);

NOR2xp33_ASAP7_75t_SL g288 ( 
.A(n_281),
.B(n_236),
.Y(n_288)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_288),
.B(n_311),
.Y(n_319)
);

MAJIxp5_ASAP7_75t_L g289 ( 
.A(n_277),
.B(n_249),
.C(n_241),
.Y(n_289)
);

MAJIxp5_ASAP7_75t_L g323 ( 
.A(n_289),
.B(n_285),
.C(n_260),
.Y(n_323)
);

XNOR2xp5_ASAP7_75t_L g321 ( 
.A(n_291),
.B(n_302),
.Y(n_321)
);

AOI22xp5_ASAP7_75t_SL g294 ( 
.A1(n_287),
.A2(n_258),
.B1(n_254),
.B2(n_245),
.Y(n_294)
);

OAI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_294),
.A2(n_315),
.B1(n_300),
.B2(n_297),
.Y(n_329)
);

XOR2xp5_ASAP7_75t_L g295 ( 
.A(n_277),
.B(n_253),
.Y(n_295)
);

XOR2xp5_ASAP7_75t_L g320 ( 
.A(n_295),
.B(n_305),
.Y(n_320)
);

NAND2xp5_ASAP7_75t_L g296 ( 
.A(n_275),
.B(n_238),
.Y(n_296)
);

INVx1_ASAP7_75t_L g325 ( 
.A(n_296),
.Y(n_325)
);

OAI22xp5_ASAP7_75t_L g324 ( 
.A1(n_300),
.A2(n_312),
.B1(n_294),
.B2(n_313),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g318 ( 
.A(n_301),
.B(n_307),
.Y(n_318)
);

XNOR2xp5_ASAP7_75t_L g302 ( 
.A(n_279),
.B(n_207),
.Y(n_302)
);

XNOR2xp5_ASAP7_75t_L g303 ( 
.A(n_276),
.B(n_168),
.Y(n_303)
);

XNOR2xp5_ASAP7_75t_L g327 ( 
.A(n_303),
.B(n_262),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_L g304 ( 
.A(n_274),
.B(n_237),
.Y(n_304)
);

INVx1_ASAP7_75t_L g342 ( 
.A(n_304),
.Y(n_342)
);

A2O1A1O1Ixp25_ASAP7_75t_L g305 ( 
.A1(n_259),
.A2(n_31),
.B(n_27),
.C(n_150),
.D(n_252),
.Y(n_305)
);

OAI21xp5_ASAP7_75t_SL g326 ( 
.A1(n_306),
.A2(n_313),
.B(n_283),
.Y(n_326)
);

XNOR2xp5_ASAP7_75t_SL g309 ( 
.A(n_276),
.B(n_58),
.Y(n_309)
);

XOR2xp5_ASAP7_75t_L g330 ( 
.A(n_309),
.B(n_303),
.Y(n_330)
);

INVxp67_ASAP7_75t_SL g311 ( 
.A(n_278),
.Y(n_311)
);

NOR2xp33_ASAP7_75t_SL g314 ( 
.A(n_271),
.B(n_265),
.Y(n_314)
);

NOR2xp33_ASAP7_75t_SL g340 ( 
.A(n_314),
.B(n_316),
.Y(n_340)
);

AOI22xp5_ASAP7_75t_L g315 ( 
.A1(n_264),
.A2(n_223),
.B1(n_215),
.B2(n_227),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g316 ( 
.A(n_265),
.B(n_272),
.Y(n_316)
);

NAND3xp33_ASAP7_75t_L g317 ( 
.A(n_278),
.B(n_150),
.C(n_110),
.Y(n_317)
);

CKINVDCx20_ASAP7_75t_R g334 ( 
.A(n_317),
.Y(n_334)
);

BUFx2_ASAP7_75t_L g322 ( 
.A(n_315),
.Y(n_322)
);

INVx2_ASAP7_75t_L g355 ( 
.A(n_322),
.Y(n_355)
);

XOR2xp5_ASAP7_75t_L g344 ( 
.A(n_323),
.B(n_327),
.Y(n_344)
);

AOI22xp5_ASAP7_75t_L g350 ( 
.A1(n_324),
.A2(n_329),
.B1(n_333),
.B2(n_339),
.Y(n_350)
);

INVxp67_ASAP7_75t_L g352 ( 
.A(n_326),
.Y(n_352)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_292),
.Y(n_328)
);

INVx1_ASAP7_75t_L g348 ( 
.A(n_328),
.Y(n_348)
);

XOR2xp5_ASAP7_75t_L g349 ( 
.A(n_330),
.B(n_309),
.Y(n_349)
);

NAND2xp5_ASAP7_75t_L g331 ( 
.A(n_293),
.B(n_274),
.Y(n_331)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_331),
.Y(n_360)
);

OAI21xp5_ASAP7_75t_SL g332 ( 
.A1(n_292),
.A2(n_261),
.B(n_266),
.Y(n_332)
);

NOR2xp33_ASAP7_75t_L g354 ( 
.A(n_332),
.B(n_299),
.Y(n_354)
);

OAI22xp5_ASAP7_75t_SL g333 ( 
.A1(n_297),
.A2(n_270),
.B1(n_266),
.B2(n_285),
.Y(n_333)
);

MAJIxp5_ASAP7_75t_L g335 ( 
.A(n_295),
.B(n_270),
.C(n_268),
.Y(n_335)
);

MAJIxp5_ASAP7_75t_L g353 ( 
.A(n_335),
.B(n_336),
.C(n_337),
.Y(n_353)
);

MAJIxp5_ASAP7_75t_L g336 ( 
.A(n_289),
.B(n_269),
.C(n_282),
.Y(n_336)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_302),
.B(n_284),
.C(n_98),
.Y(n_337)
);

INVx1_ASAP7_75t_L g338 ( 
.A(n_304),
.Y(n_338)
);

INVx1_ASAP7_75t_L g366 ( 
.A(n_338),
.Y(n_366)
);

OAI22xp5_ASAP7_75t_SL g339 ( 
.A1(n_291),
.A2(n_223),
.B1(n_215),
.B2(n_130),
.Y(n_339)
);

INVx2_ASAP7_75t_L g341 ( 
.A(n_290),
.Y(n_341)
);

NAND2xp5_ASAP7_75t_L g343 ( 
.A(n_341),
.B(n_296),
.Y(n_343)
);

INVx1_ASAP7_75t_L g368 ( 
.A(n_343),
.Y(n_368)
);

OAI22xp5_ASAP7_75t_L g345 ( 
.A1(n_334),
.A2(n_340),
.B1(n_319),
.B2(n_322),
.Y(n_345)
);

INVx1_ASAP7_75t_L g369 ( 
.A(n_345),
.Y(n_369)
);

OAI21xp5_ASAP7_75t_L g346 ( 
.A1(n_331),
.A2(n_306),
.B(n_313),
.Y(n_346)
);

OAI21xp5_ASAP7_75t_L g367 ( 
.A1(n_346),
.A2(n_338),
.B(n_342),
.Y(n_367)
);

OAI22xp5_ASAP7_75t_SL g347 ( 
.A1(n_318),
.A2(n_298),
.B1(n_308),
.B2(n_310),
.Y(n_347)
);

NAND2xp5_ASAP7_75t_L g371 ( 
.A(n_347),
.B(n_356),
.Y(n_371)
);

XNOR2x1_ASAP7_75t_L g381 ( 
.A(n_349),
.B(n_362),
.Y(n_381)
);

XOR2xp5_ASAP7_75t_L g351 ( 
.A(n_323),
.B(n_307),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g373 ( 
.A(n_351),
.B(n_359),
.Y(n_373)
);

INVxp67_ASAP7_75t_L g374 ( 
.A(n_354),
.Y(n_374)
);

FAx1_ASAP7_75t_SL g356 ( 
.A(n_321),
.B(n_305),
.CI(n_299),
.CON(n_356),
.SN(n_356)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_335),
.B(n_123),
.C(n_127),
.Y(n_357)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_357),
.B(n_363),
.C(n_52),
.Y(n_383)
);

INVxp33_ASAP7_75t_L g358 ( 
.A(n_318),
.Y(n_358)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_358),
.Y(n_382)
);

XOR2xp5_ASAP7_75t_L g359 ( 
.A(n_321),
.B(n_61),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g361 ( 
.A(n_336),
.B(n_320),
.Y(n_361)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_361),
.B(n_135),
.Y(n_385)
);

XOR2xp5_ASAP7_75t_L g362 ( 
.A(n_330),
.B(n_123),
.Y(n_362)
);

MAJIxp5_ASAP7_75t_L g363 ( 
.A(n_337),
.B(n_127),
.C(n_95),
.Y(n_363)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_325),
.B(n_0),
.Y(n_364)
);

INVx1_ASAP7_75t_L g387 ( 
.A(n_364),
.Y(n_387)
);

CKINVDCx16_ASAP7_75t_R g365 ( 
.A(n_328),
.Y(n_365)
);

NAND2xp5_ASAP7_75t_L g378 ( 
.A(n_365),
.B(n_348),
.Y(n_378)
);

AOI21xp5_ASAP7_75t_L g399 ( 
.A1(n_367),
.A2(n_366),
.B(n_355),
.Y(n_399)
);

FAx1_ASAP7_75t_L g370 ( 
.A(n_346),
.B(n_332),
.CI(n_327),
.CON(n_370),
.SN(n_370)
);

NAND2xp5_ASAP7_75t_L g389 ( 
.A(n_370),
.B(n_376),
.Y(n_389)
);

OAI22xp5_ASAP7_75t_SL g372 ( 
.A1(n_350),
.A2(n_329),
.B1(n_333),
.B2(n_326),
.Y(n_372)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_372),
.Y(n_388)
);

OAI22xp5_ASAP7_75t_L g375 ( 
.A1(n_350),
.A2(n_341),
.B1(n_320),
.B2(n_339),
.Y(n_375)
);

INVx1_ASAP7_75t_L g391 ( 
.A(n_375),
.Y(n_391)
);

NOR2xp33_ASAP7_75t_SL g376 ( 
.A(n_356),
.B(n_173),
.Y(n_376)
);

OAI22xp5_ASAP7_75t_SL g377 ( 
.A1(n_360),
.A2(n_173),
.B1(n_128),
.B2(n_69),
.Y(n_377)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_377),
.Y(n_400)
);

NOR2xp33_ASAP7_75t_L g393 ( 
.A(n_378),
.B(n_380),
.Y(n_393)
);

OAI22xp5_ASAP7_75t_SL g379 ( 
.A1(n_352),
.A2(n_84),
.B1(n_69),
.B2(n_83),
.Y(n_379)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_379),
.B(n_383),
.Y(n_392)
);

BUFx12_ASAP7_75t_L g380 ( 
.A(n_358),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g384 ( 
.A(n_353),
.B(n_83),
.C(n_84),
.Y(n_384)
);

MAJIxp5_ASAP7_75t_L g390 ( 
.A(n_384),
.B(n_344),
.C(n_353),
.Y(n_390)
);

XOR2xp5_ASAP7_75t_L g401 ( 
.A(n_385),
.B(n_386),
.Y(n_401)
);

XNOR2x1_ASAP7_75t_L g386 ( 
.A(n_351),
.B(n_0),
.Y(n_386)
);

NAND2xp5_ASAP7_75t_SL g405 ( 
.A(n_390),
.B(n_384),
.Y(n_405)
);

INVx3_ASAP7_75t_L g394 ( 
.A(n_387),
.Y(n_394)
);

NAND2xp5_ASAP7_75t_L g416 ( 
.A(n_394),
.B(n_1),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g395 ( 
.A(n_383),
.B(n_344),
.C(n_361),
.Y(n_395)
);

MAJIxp5_ASAP7_75t_L g413 ( 
.A(n_395),
.B(n_396),
.C(n_398),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g396 ( 
.A(n_373),
.B(n_357),
.C(n_363),
.Y(n_396)
);

NOR2xp33_ASAP7_75t_SL g397 ( 
.A(n_374),
.B(n_356),
.Y(n_397)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_397),
.B(n_381),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g398 ( 
.A(n_373),
.B(n_362),
.C(n_352),
.Y(n_398)
);

OAI21xp5_ASAP7_75t_L g409 ( 
.A1(n_399),
.A2(n_367),
.B(n_382),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_L g402 ( 
.A1(n_369),
.A2(n_359),
.B1(n_349),
.B2(n_192),
.Y(n_402)
);

AOI22xp5_ASAP7_75t_L g404 ( 
.A1(n_402),
.A2(n_403),
.B1(n_377),
.B2(n_368),
.Y(n_404)
);

OAI22xp5_ASAP7_75t_SL g403 ( 
.A1(n_371),
.A2(n_39),
.B1(n_103),
.B2(n_139),
.Y(n_403)
);

INVxp67_ASAP7_75t_L g422 ( 
.A(n_404),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_405),
.B(n_406),
.Y(n_420)
);

NOR2xp33_ASAP7_75t_SL g406 ( 
.A(n_394),
.B(n_374),
.Y(n_406)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_395),
.B(n_372),
.Y(n_407)
);

NAND2xp5_ASAP7_75t_L g421 ( 
.A(n_407),
.B(n_408),
.Y(n_421)
);

NOR2xp33_ASAP7_75t_L g408 ( 
.A(n_389),
.B(n_393),
.Y(n_408)
);

AO21x1_ASAP7_75t_SL g428 ( 
.A1(n_409),
.A2(n_416),
.B(n_1),
.Y(n_428)
);

FAx1_ASAP7_75t_L g410 ( 
.A(n_388),
.B(n_370),
.CI(n_371),
.CON(n_410),
.SN(n_410)
);

OR2x2_ASAP7_75t_L g423 ( 
.A(n_410),
.B(n_392),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_L g411 ( 
.A1(n_391),
.A2(n_370),
.B1(n_380),
.B2(n_386),
.Y(n_411)
);

NAND2xp5_ASAP7_75t_L g425 ( 
.A(n_411),
.B(n_414),
.Y(n_425)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_412),
.Y(n_424)
);

NOR2xp33_ASAP7_75t_SL g414 ( 
.A(n_390),
.B(n_379),
.Y(n_414)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_399),
.B(n_380),
.Y(n_415)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_415),
.B(n_39),
.Y(n_427)
);

FAx1_ASAP7_75t_SL g417 ( 
.A(n_409),
.B(n_401),
.CI(n_398),
.CON(n_417),
.SN(n_417)
);

INVx1_ASAP7_75t_L g429 ( 
.A(n_417),
.Y(n_429)
);

AOI21xp5_ASAP7_75t_L g418 ( 
.A1(n_413),
.A2(n_396),
.B(n_400),
.Y(n_418)
);

OAI21xp5_ASAP7_75t_SL g436 ( 
.A1(n_418),
.A2(n_4),
.B(n_6),
.Y(n_436)
);

AOI21xp33_ASAP7_75t_L g419 ( 
.A1(n_410),
.A2(n_403),
.B(n_392),
.Y(n_419)
);

AO22x1_ASAP7_75t_L g433 ( 
.A1(n_419),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_433)
);

NAND2xp5_ASAP7_75t_SL g437 ( 
.A(n_423),
.B(n_8),
.Y(n_437)
);

AOI31xp67_ASAP7_75t_L g426 ( 
.A1(n_410),
.A2(n_401),
.A3(n_381),
.B(n_3),
.Y(n_426)
);

OR2x2_ASAP7_75t_L g434 ( 
.A(n_426),
.B(n_2),
.Y(n_434)
);

NAND2xp5_ASAP7_75t_L g438 ( 
.A(n_427),
.B(n_46),
.Y(n_438)
);

XOR2xp5_ASAP7_75t_L g432 ( 
.A(n_428),
.B(n_2),
.Y(n_432)
);

AOI322xp5_ASAP7_75t_L g430 ( 
.A1(n_422),
.A2(n_407),
.A3(n_413),
.B1(n_103),
.B2(n_82),
.C1(n_6),
.C2(n_7),
.Y(n_430)
);

AOI22xp5_ASAP7_75t_SL g441 ( 
.A1(n_430),
.A2(n_433),
.B1(n_435),
.B2(n_424),
.Y(n_441)
);

NAND4xp25_ASAP7_75t_SL g431 ( 
.A(n_420),
.B(n_46),
.C(n_3),
.D(n_4),
.Y(n_431)
);

AOI21xp5_ASAP7_75t_L g439 ( 
.A1(n_431),
.A2(n_8),
.B(n_9),
.Y(n_439)
);

MAJIxp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_436),
.C(n_438),
.Y(n_443)
);

INVx1_ASAP7_75t_SL g440 ( 
.A(n_434),
.Y(n_440)
);

AND2x2_ASAP7_75t_L g435 ( 
.A(n_421),
.B(n_46),
.Y(n_435)
);

OAI21xp5_ASAP7_75t_L g444 ( 
.A1(n_437),
.A2(n_423),
.B(n_9),
.Y(n_444)
);

AOI21xp5_ASAP7_75t_SL g447 ( 
.A1(n_439),
.A2(n_442),
.B(n_445),
.Y(n_447)
);

AO21x1_ASAP7_75t_L g446 ( 
.A1(n_441),
.A2(n_444),
.B(n_430),
.Y(n_446)
);

MAJx2_ASAP7_75t_L g442 ( 
.A(n_429),
.B(n_425),
.C(n_417),
.Y(n_442)
);

OAI21xp5_ASAP7_75t_L g445 ( 
.A1(n_437),
.A2(n_8),
.B(n_10),
.Y(n_445)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_446),
.B(n_11),
.Y(n_451)
);

AOI322xp5_ASAP7_75t_L g448 ( 
.A1(n_440),
.A2(n_8),
.A3(n_10),
.B1(n_11),
.B2(n_12),
.C1(n_46),
.C2(n_443),
.Y(n_448)
);

OAI21xp33_ASAP7_75t_L g450 ( 
.A1(n_448),
.A2(n_449),
.B(n_447),
.Y(n_450)
);

AO21x1_ASAP7_75t_L g449 ( 
.A1(n_444),
.A2(n_11),
.B(n_12),
.Y(n_449)
);

AOI21xp5_ASAP7_75t_SL g452 ( 
.A1(n_450),
.A2(n_451),
.B(n_11),
.Y(n_452)
);

CKINVDCx20_ASAP7_75t_R g453 ( 
.A(n_452),
.Y(n_453)
);

AOI21xp5_ASAP7_75t_L g454 ( 
.A1(n_453),
.A2(n_12),
.B(n_46),
.Y(n_454)
);

XOR2xp5_ASAP7_75t_L g455 ( 
.A(n_454),
.B(n_12),
.Y(n_455)
);


endmodule