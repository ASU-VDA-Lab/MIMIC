module fake_jpeg_29338_n_452 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_452);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_452;

wire n_390;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_182;
wire n_19;
wire n_252;
wire n_385;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_377;
wire n_291;
wire n_236;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_44;
wire n_355;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_196;
wire n_66;
wire n_374;
wire n_142;
wire n_362;
wire n_417;
wire n_172;
wire n_345;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_304;
wire n_60;
wire n_283;
wire n_107;
wire n_415;
wire n_357;
wire n_89;
wire n_131;
wire n_294;
wire n_230;
wire n_170;
wire n_313;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_48;
wire n_200;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_416;
wire n_221;
wire n_256;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_82;
wire n_155;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_42;
wire n_49;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_31;
wire n_277;
wire n_255;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_408;
wire n_80;
wire n_204;
wire n_306;
wire n_429;
wire n_368;
wire n_298;
wire n_106;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_254;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_268;
wire n_404;
wire n_91;
wire n_305;
wire n_161;
wire n_441;
wire n_342;
wire n_101;
wire n_226;
wire n_149;
wire n_87;
wire n_46;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_97;
wire n_382;
wire n_237;
wire n_188;
wire n_174;
wire n_198;
wire n_422;
wire n_190;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_110;
wire n_76;
wire n_278;
wire n_343;
wire n_26;
wire n_88;
wire n_397;
wire n_363;
wire n_238;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_301;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_389;
wire n_339;
wire n_109;
wire n_267;
wire n_296;
wire n_384;
wire n_168;
wire n_274;
wire n_24;
wire n_269;
wire n_287;
wire n_219;
wire n_433;
wire n_77;
wire n_45;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_239;
wire n_243;
wire n_348;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_333;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_302;
wire n_216;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_199;
wire n_260;
wire n_413;
wire n_275;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_36;
wire n_62;
wire n_118;
wire n_140;
wire n_361;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_347;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_279;
wire n_154;
wire n_205;
wire n_379;
wire n_114;
wire n_444;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_257;
wire n_61;
wire n_173;
wire n_244;
wire n_232;
wire n_58;
wire n_41;
wire n_266;
wire n_72;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_183;
wire n_409;
wire n_249;
wire n_412;
wire n_217;
wire n_53;
wire n_372;
wire n_33;
wire n_54;
wire n_391;
wire n_209;
wire n_22;
wire n_138;
wire n_402;
wire n_438;
wire n_247;
wire n_157;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_151;
wire n_341;
wire n_426;
wire n_290;
wire n_242;
wire n_351;
wire n_325;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_282;
wire n_181;

BUFx3_ASAP7_75t_L g19 ( 
.A(n_3),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_7),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_13),
.Y(n_21)
);

INVx1_ASAP7_75t_L g22 ( 
.A(n_8),
.Y(n_22)
);

BUFx10_ASAP7_75t_L g23 ( 
.A(n_0),
.Y(n_23)
);

INVx4_ASAP7_75t_L g24 ( 
.A(n_7),
.Y(n_24)
);

INVx6_ASAP7_75t_L g25 ( 
.A(n_4),
.Y(n_25)
);

INVx2_ASAP7_75t_L g26 ( 
.A(n_1),
.Y(n_26)
);

INVx8_ASAP7_75t_L g27 ( 
.A(n_10),
.Y(n_27)
);

BUFx10_ASAP7_75t_L g28 ( 
.A(n_10),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_16),
.Y(n_29)
);

BUFx12f_ASAP7_75t_L g30 ( 
.A(n_5),
.Y(n_30)
);

BUFx12f_ASAP7_75t_L g31 ( 
.A(n_2),
.Y(n_31)
);

CKINVDCx20_ASAP7_75t_R g32 ( 
.A(n_6),
.Y(n_32)
);

CKINVDCx20_ASAP7_75t_R g33 ( 
.A(n_3),
.Y(n_33)
);

INVx1_ASAP7_75t_L g34 ( 
.A(n_4),
.Y(n_34)
);

INVx1_ASAP7_75t_L g35 ( 
.A(n_7),
.Y(n_35)
);

INVx1_ASAP7_75t_L g36 ( 
.A(n_2),
.Y(n_36)
);

CKINVDCx20_ASAP7_75t_R g37 ( 
.A(n_15),
.Y(n_37)
);

BUFx10_ASAP7_75t_L g38 ( 
.A(n_15),
.Y(n_38)
);

BUFx6f_ASAP7_75t_L g39 ( 
.A(n_0),
.Y(n_39)
);

INVx1_ASAP7_75t_L g40 ( 
.A(n_10),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_6),
.Y(n_41)
);

INVx4_ASAP7_75t_L g42 ( 
.A(n_1),
.Y(n_42)
);

BUFx6f_ASAP7_75t_L g43 ( 
.A(n_17),
.Y(n_43)
);

INVx1_ASAP7_75t_L g44 ( 
.A(n_1),
.Y(n_44)
);

INVx2_ASAP7_75t_SL g45 ( 
.A(n_2),
.Y(n_45)
);

BUFx5_ASAP7_75t_L g46 ( 
.A(n_20),
.Y(n_46)
);

INVx3_ASAP7_75t_SL g105 ( 
.A(n_46),
.Y(n_105)
);

INVx8_ASAP7_75t_L g47 ( 
.A(n_42),
.Y(n_47)
);

INVx8_ASAP7_75t_L g145 ( 
.A(n_47),
.Y(n_145)
);

CKINVDCx20_ASAP7_75t_R g48 ( 
.A(n_28),
.Y(n_48)
);

NOR2xp33_ASAP7_75t_L g96 ( 
.A(n_48),
.B(n_58),
.Y(n_96)
);

BUFx6f_ASAP7_75t_L g49 ( 
.A(n_39),
.Y(n_49)
);

BUFx6f_ASAP7_75t_L g103 ( 
.A(n_49),
.Y(n_103)
);

BUFx12f_ASAP7_75t_L g50 ( 
.A(n_39),
.Y(n_50)
);

BUFx5_ASAP7_75t_L g113 ( 
.A(n_50),
.Y(n_113)
);

INVx3_ASAP7_75t_L g51 ( 
.A(n_24),
.Y(n_51)
);

INVx3_ASAP7_75t_L g118 ( 
.A(n_51),
.Y(n_118)
);

NAND2xp5_ASAP7_75t_L g52 ( 
.A(n_21),
.B(n_9),
.Y(n_52)
);

NAND2xp5_ASAP7_75t_L g116 ( 
.A(n_52),
.B(n_32),
.Y(n_116)
);

BUFx3_ASAP7_75t_L g53 ( 
.A(n_19),
.Y(n_53)
);

INVx4_ASAP7_75t_L g130 ( 
.A(n_53),
.Y(n_130)
);

INVx3_ASAP7_75t_L g54 ( 
.A(n_24),
.Y(n_54)
);

INVx3_ASAP7_75t_L g132 ( 
.A(n_54),
.Y(n_132)
);

BUFx3_ASAP7_75t_L g55 ( 
.A(n_19),
.Y(n_55)
);

INVx4_ASAP7_75t_L g135 ( 
.A(n_55),
.Y(n_135)
);

BUFx6f_ASAP7_75t_L g56 ( 
.A(n_39),
.Y(n_56)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_56),
.Y(n_109)
);

BUFx8_ASAP7_75t_L g57 ( 
.A(n_20),
.Y(n_57)
);

BUFx2_ASAP7_75t_L g140 ( 
.A(n_57),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g58 ( 
.A(n_28),
.Y(n_58)
);

INVx6_ASAP7_75t_L g59 ( 
.A(n_39),
.Y(n_59)
);

BUFx6f_ASAP7_75t_L g110 ( 
.A(n_59),
.Y(n_110)
);

CKINVDCx20_ASAP7_75t_R g60 ( 
.A(n_28),
.Y(n_60)
);

NOR2xp33_ASAP7_75t_L g98 ( 
.A(n_60),
.B(n_63),
.Y(n_98)
);

BUFx6f_ASAP7_75t_L g61 ( 
.A(n_43),
.Y(n_61)
);

BUFx6f_ASAP7_75t_L g111 ( 
.A(n_61),
.Y(n_111)
);

INVx3_ASAP7_75t_L g62 ( 
.A(n_24),
.Y(n_62)
);

INVx5_ASAP7_75t_L g125 ( 
.A(n_62),
.Y(n_125)
);

CKINVDCx20_ASAP7_75t_R g63 ( 
.A(n_28),
.Y(n_63)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_20),
.Y(n_64)
);

INVx5_ASAP7_75t_L g131 ( 
.A(n_64),
.Y(n_131)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_43),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g115 ( 
.A(n_65),
.Y(n_115)
);

INVx6_ASAP7_75t_L g66 ( 
.A(n_43),
.Y(n_66)
);

BUFx6f_ASAP7_75t_L g120 ( 
.A(n_66),
.Y(n_120)
);

INVx1_ASAP7_75t_L g67 ( 
.A(n_22),
.Y(n_67)
);

INVx1_ASAP7_75t_L g94 ( 
.A(n_67),
.Y(n_94)
);

BUFx3_ASAP7_75t_L g68 ( 
.A(n_19),
.Y(n_68)
);

BUFx3_ASAP7_75t_L g102 ( 
.A(n_68),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g69 ( 
.A(n_43),
.Y(n_69)
);

BUFx6f_ASAP7_75t_L g124 ( 
.A(n_69),
.Y(n_124)
);

BUFx12f_ASAP7_75t_L g70 ( 
.A(n_28),
.Y(n_70)
);

NOR2xp33_ASAP7_75t_L g99 ( 
.A(n_70),
.B(n_73),
.Y(n_99)
);

BUFx6f_ASAP7_75t_L g71 ( 
.A(n_25),
.Y(n_71)
);

BUFx6f_ASAP7_75t_L g127 ( 
.A(n_71),
.Y(n_127)
);

INVx1_ASAP7_75t_L g72 ( 
.A(n_22),
.Y(n_72)
);

INVx1_ASAP7_75t_L g97 ( 
.A(n_72),
.Y(n_97)
);

NOR2xp33_ASAP7_75t_L g73 ( 
.A(n_21),
.B(n_18),
.Y(n_73)
);

INVx2_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

INVx2_ASAP7_75t_L g101 ( 
.A(n_74),
.Y(n_101)
);

INVx4_ASAP7_75t_L g75 ( 
.A(n_42),
.Y(n_75)
);

INVx3_ASAP7_75t_SL g107 ( 
.A(n_75),
.Y(n_107)
);

INVx1_ASAP7_75t_L g76 ( 
.A(n_29),
.Y(n_76)
);

INVx1_ASAP7_75t_L g100 ( 
.A(n_76),
.Y(n_100)
);

CKINVDCx20_ASAP7_75t_R g77 ( 
.A(n_28),
.Y(n_77)
);

NOR2xp33_ASAP7_75t_L g122 ( 
.A(n_77),
.B(n_84),
.Y(n_122)
);

INVx4_ASAP7_75t_L g78 ( 
.A(n_42),
.Y(n_78)
);

INVx4_ASAP7_75t_SL g146 ( 
.A(n_78),
.Y(n_146)
);

BUFx6f_ASAP7_75t_L g79 ( 
.A(n_25),
.Y(n_79)
);

BUFx6f_ASAP7_75t_L g136 ( 
.A(n_79),
.Y(n_136)
);

INVx5_ASAP7_75t_L g80 ( 
.A(n_27),
.Y(n_80)
);

BUFx3_ASAP7_75t_L g114 ( 
.A(n_80),
.Y(n_114)
);

INVx1_ASAP7_75t_L g81 ( 
.A(n_29),
.Y(n_81)
);

INVx1_ASAP7_75t_L g121 ( 
.A(n_81),
.Y(n_121)
);

BUFx16f_ASAP7_75t_L g82 ( 
.A(n_38),
.Y(n_82)
);

BUFx12f_ASAP7_75t_L g117 ( 
.A(n_82),
.Y(n_117)
);

INVx3_ASAP7_75t_L g83 ( 
.A(n_20),
.Y(n_83)
);

INVx2_ASAP7_75t_L g106 ( 
.A(n_83),
.Y(n_106)
);

CKINVDCx20_ASAP7_75t_R g84 ( 
.A(n_38),
.Y(n_84)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_25),
.Y(n_85)
);

CKINVDCx14_ASAP7_75t_R g137 ( 
.A(n_85),
.Y(n_137)
);

BUFx6f_ASAP7_75t_L g86 ( 
.A(n_26),
.Y(n_86)
);

INVx6_ASAP7_75t_L g141 ( 
.A(n_86),
.Y(n_141)
);

INVx2_ASAP7_75t_L g87 ( 
.A(n_26),
.Y(n_87)
);

INVx2_ASAP7_75t_L g108 ( 
.A(n_87),
.Y(n_108)
);

INVx2_ASAP7_75t_L g88 ( 
.A(n_27),
.Y(n_88)
);

INVx2_ASAP7_75t_L g133 ( 
.A(n_88),
.Y(n_133)
);

INVx13_ASAP7_75t_L g89 ( 
.A(n_27),
.Y(n_89)
);

BUFx12f_ASAP7_75t_L g123 ( 
.A(n_89),
.Y(n_123)
);

BUFx6f_ASAP7_75t_L g90 ( 
.A(n_38),
.Y(n_90)
);

INVx2_ASAP7_75t_L g138 ( 
.A(n_90),
.Y(n_138)
);

BUFx12f_ASAP7_75t_L g91 ( 
.A(n_38),
.Y(n_91)
);

CKINVDCx16_ASAP7_75t_R g143 ( 
.A(n_91),
.Y(n_143)
);

INVx2_ASAP7_75t_L g92 ( 
.A(n_34),
.Y(n_92)
);

INVx2_ASAP7_75t_L g142 ( 
.A(n_92),
.Y(n_142)
);

INVx13_ASAP7_75t_L g93 ( 
.A(n_38),
.Y(n_93)
);

BUFx12_ASAP7_75t_L g112 ( 
.A(n_93),
.Y(n_112)
);

NAND2xp5_ASAP7_75t_SL g95 ( 
.A(n_75),
.B(n_37),
.Y(n_95)
);

NAND2xp5_ASAP7_75t_SL g167 ( 
.A(n_95),
.B(n_104),
.Y(n_167)
);

NAND2xp5_ASAP7_75t_SL g104 ( 
.A(n_78),
.B(n_37),
.Y(n_104)
);

AND2x2_ASAP7_75t_L g147 ( 
.A(n_116),
.B(n_35),
.Y(n_147)
);

BUFx12_ASAP7_75t_L g119 ( 
.A(n_82),
.Y(n_119)
);

BUFx12f_ASAP7_75t_L g181 ( 
.A(n_119),
.Y(n_181)
);

OR2x2_ASAP7_75t_L g126 ( 
.A(n_93),
.B(n_32),
.Y(n_126)
);

NOR2xp33_ASAP7_75t_L g152 ( 
.A(n_126),
.B(n_129),
.Y(n_152)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_86),
.B(n_33),
.Y(n_128)
);

NAND2xp5_ASAP7_75t_L g148 ( 
.A(n_128),
.B(n_33),
.Y(n_148)
);

INVx1_ASAP7_75t_L g129 ( 
.A(n_47),
.Y(n_129)
);

OAI22xp5_ASAP7_75t_L g134 ( 
.A1(n_71),
.A2(n_35),
.B1(n_40),
.B2(n_41),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_L g166 ( 
.A1(n_134),
.A2(n_34),
.B1(n_36),
.B2(n_44),
.Y(n_166)
);

NOR2xp33_ASAP7_75t_SL g139 ( 
.A(n_57),
.B(n_40),
.Y(n_139)
);

NOR2xp33_ASAP7_75t_L g161 ( 
.A(n_139),
.B(n_41),
.Y(n_161)
);

AOI22xp33_ASAP7_75t_L g144 ( 
.A1(n_66),
.A2(n_20),
.B1(n_30),
.B2(n_31),
.Y(n_144)
);

OAI22xp5_ASAP7_75t_SL g165 ( 
.A1(n_144),
.A2(n_45),
.B1(n_70),
.B2(n_91),
.Y(n_165)
);

AND2x2_ASAP7_75t_L g206 ( 
.A(n_147),
.B(n_148),
.Y(n_206)
);

CKINVDCx16_ASAP7_75t_R g149 ( 
.A(n_126),
.Y(n_149)
);

NOR2xp33_ASAP7_75t_L g205 ( 
.A(n_149),
.B(n_151),
.Y(n_205)
);

INVx1_ASAP7_75t_L g150 ( 
.A(n_142),
.Y(n_150)
);

INVx1_ASAP7_75t_L g190 ( 
.A(n_150),
.Y(n_190)
);

CKINVDCx16_ASAP7_75t_R g151 ( 
.A(n_96),
.Y(n_151)
);

CKINVDCx20_ASAP7_75t_R g153 ( 
.A(n_96),
.Y(n_153)
);

NAND3xp33_ASAP7_75t_L g199 ( 
.A(n_153),
.B(n_159),
.C(n_169),
.Y(n_199)
);

NAND2xp5_ASAP7_75t_L g154 ( 
.A(n_94),
.B(n_97),
.Y(n_154)
);

NAND2xp5_ASAP7_75t_L g195 ( 
.A(n_154),
.B(n_157),
.Y(n_195)
);

INVx5_ASAP7_75t_L g155 ( 
.A(n_113),
.Y(n_155)
);

INVx11_ASAP7_75t_L g188 ( 
.A(n_155),
.Y(n_188)
);

INVx2_ASAP7_75t_L g156 ( 
.A(n_101),
.Y(n_156)
);

INVx2_ASAP7_75t_L g191 ( 
.A(n_156),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_L g157 ( 
.A(n_100),
.B(n_36),
.Y(n_157)
);

AOI22xp33_ASAP7_75t_SL g158 ( 
.A1(n_146),
.A2(n_80),
.B1(n_45),
.B2(n_55),
.Y(n_158)
);

AOI22xp33_ASAP7_75t_SL g189 ( 
.A1(n_158),
.A2(n_171),
.B1(n_179),
.B2(n_140),
.Y(n_189)
);

CKINVDCx16_ASAP7_75t_R g159 ( 
.A(n_121),
.Y(n_159)
);

INVx2_ASAP7_75t_L g160 ( 
.A(n_108),
.Y(n_160)
);

INVx2_ASAP7_75t_L g192 ( 
.A(n_160),
.Y(n_192)
);

NOR2xp33_ASAP7_75t_SL g203 ( 
.A(n_161),
.B(n_168),
.Y(n_203)
);

INVx1_ASAP7_75t_L g162 ( 
.A(n_133),
.Y(n_162)
);

INVx1_ASAP7_75t_L g213 ( 
.A(n_162),
.Y(n_213)
);

INVx2_ASAP7_75t_L g163 ( 
.A(n_138),
.Y(n_163)
);

INVx2_ASAP7_75t_L g204 ( 
.A(n_163),
.Y(n_204)
);

BUFx6f_ASAP7_75t_L g164 ( 
.A(n_111),
.Y(n_164)
);

INVx11_ASAP7_75t_L g198 ( 
.A(n_164),
.Y(n_198)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_165),
.A2(n_166),
.B1(n_176),
.B2(n_149),
.Y(n_187)
);

NOR2xp33_ASAP7_75t_L g168 ( 
.A(n_99),
.B(n_44),
.Y(n_168)
);

NOR2xp33_ASAP7_75t_L g169 ( 
.A(n_99),
.B(n_89),
.Y(n_169)
);

NOR2xp33_ASAP7_75t_L g170 ( 
.A(n_98),
.B(n_30),
.Y(n_170)
);

NAND2xp5_ASAP7_75t_L g201 ( 
.A(n_170),
.B(n_172),
.Y(n_201)
);

AOI22xp33_ASAP7_75t_SL g171 ( 
.A1(n_146),
.A2(n_45),
.B1(n_68),
.B2(n_53),
.Y(n_171)
);

CKINVDCx20_ASAP7_75t_R g172 ( 
.A(n_98),
.Y(n_172)
);

NOR2xp33_ASAP7_75t_L g173 ( 
.A(n_122),
.B(n_31),
.Y(n_173)
);

XNOR2xp5_ASAP7_75t_L g193 ( 
.A(n_173),
.B(n_175),
.Y(n_193)
);

INVx6_ASAP7_75t_L g174 ( 
.A(n_111),
.Y(n_174)
);

BUFx6f_ASAP7_75t_L g196 ( 
.A(n_174),
.Y(n_196)
);

NOR2xp33_ASAP7_75t_L g175 ( 
.A(n_122),
.B(n_31),
.Y(n_175)
);

AOI21xp5_ASAP7_75t_L g176 ( 
.A1(n_105),
.A2(n_45),
.B(n_85),
.Y(n_176)
);

AOI21xp5_ASAP7_75t_L g186 ( 
.A1(n_176),
.A2(n_105),
.B(n_107),
.Y(n_186)
);

INVx3_ASAP7_75t_L g177 ( 
.A(n_123),
.Y(n_177)
);

INVx3_ASAP7_75t_L g197 ( 
.A(n_177),
.Y(n_197)
);

INVx2_ASAP7_75t_L g178 ( 
.A(n_106),
.Y(n_178)
);

INVx2_ASAP7_75t_L g210 ( 
.A(n_178),
.Y(n_210)
);

INVx3_ASAP7_75t_SL g179 ( 
.A(n_130),
.Y(n_179)
);

BUFx6f_ASAP7_75t_L g180 ( 
.A(n_115),
.Y(n_180)
);

INVx6_ASAP7_75t_L g202 ( 
.A(n_180),
.Y(n_202)
);

INVx2_ASAP7_75t_L g182 ( 
.A(n_141),
.Y(n_182)
);

INVx2_ASAP7_75t_L g211 ( 
.A(n_182),
.Y(n_211)
);

NAND2xp5_ASAP7_75t_L g183 ( 
.A(n_110),
.B(n_38),
.Y(n_183)
);

MAJIxp5_ASAP7_75t_L g200 ( 
.A(n_183),
.B(n_165),
.C(n_137),
.Y(n_200)
);

INVx1_ASAP7_75t_L g184 ( 
.A(n_107),
.Y(n_184)
);

BUFx3_ASAP7_75t_L g207 ( 
.A(n_184),
.Y(n_207)
);

INVx6_ASAP7_75t_L g185 ( 
.A(n_115),
.Y(n_185)
);

INVx6_ASAP7_75t_L g209 ( 
.A(n_185),
.Y(n_209)
);

AOI21xp5_ASAP7_75t_L g236 ( 
.A1(n_186),
.A2(n_194),
.B(n_135),
.Y(n_236)
);

OAI22xp5_ASAP7_75t_L g230 ( 
.A1(n_187),
.A2(n_79),
.B1(n_125),
.B2(n_114),
.Y(n_230)
);

OAI21xp33_ASAP7_75t_SL g234 ( 
.A1(n_189),
.A2(n_202),
.B(n_209),
.Y(n_234)
);

OAI21xp5_ASAP7_75t_SL g194 ( 
.A1(n_152),
.A2(n_144),
.B(n_118),
.Y(n_194)
);

MAJIxp5_ASAP7_75t_L g218 ( 
.A(n_200),
.B(n_150),
.C(n_162),
.Y(n_218)
);

AOI22xp33_ASAP7_75t_SL g208 ( 
.A1(n_153),
.A2(n_137),
.B1(n_140),
.B2(n_172),
.Y(n_208)
);

BUFx24_ASAP7_75t_L g221 ( 
.A(n_208),
.Y(n_221)
);

O2A1O1Ixp33_ASAP7_75t_L g212 ( 
.A1(n_157),
.A2(n_112),
.B(n_123),
.C(n_143),
.Y(n_212)
);

OAI21xp5_ASAP7_75t_L g225 ( 
.A1(n_212),
.A2(n_184),
.B(n_132),
.Y(n_225)
);

INVx6_ASAP7_75t_L g214 ( 
.A(n_198),
.Y(n_214)
);

INVx1_ASAP7_75t_L g248 ( 
.A(n_214),
.Y(n_248)
);

NOR2xp33_ASAP7_75t_L g215 ( 
.A(n_203),
.B(n_154),
.Y(n_215)
);

NAND2xp5_ASAP7_75t_L g242 ( 
.A(n_215),
.B(n_216),
.Y(n_242)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_195),
.B(n_148),
.Y(n_216)
);

OAI22xp5_ASAP7_75t_SL g217 ( 
.A1(n_187),
.A2(n_183),
.B1(n_167),
.B2(n_127),
.Y(n_217)
);

AOI22xp5_ASAP7_75t_L g249 ( 
.A1(n_217),
.A2(n_223),
.B1(n_228),
.B2(n_229),
.Y(n_249)
);

XNOR2xp5_ASAP7_75t_L g243 ( 
.A(n_218),
.B(n_224),
.Y(n_243)
);

CKINVDCx14_ASAP7_75t_R g219 ( 
.A(n_207),
.Y(n_219)
);

NOR2xp33_ASAP7_75t_L g245 ( 
.A(n_219),
.B(n_222),
.Y(n_245)
);

NAND2xp5_ASAP7_75t_SL g220 ( 
.A(n_195),
.B(n_147),
.Y(n_220)
);

NAND2xp5_ASAP7_75t_L g255 ( 
.A(n_220),
.B(n_226),
.Y(n_255)
);

INVx2_ASAP7_75t_L g222 ( 
.A(n_211),
.Y(n_222)
);

OAI22xp33_ASAP7_75t_SL g223 ( 
.A1(n_186),
.A2(n_159),
.B1(n_182),
.B2(n_179),
.Y(n_223)
);

MAJIxp5_ASAP7_75t_L g224 ( 
.A(n_193),
.B(n_147),
.C(n_156),
.Y(n_224)
);

INVxp67_ASAP7_75t_L g253 ( 
.A(n_225),
.Y(n_253)
);

NAND2xp5_ASAP7_75t_SL g226 ( 
.A(n_206),
.B(n_160),
.Y(n_226)
);

NOR2xp33_ASAP7_75t_L g227 ( 
.A(n_201),
.B(n_205),
.Y(n_227)
);

CKINVDCx16_ASAP7_75t_R g258 ( 
.A(n_227),
.Y(n_258)
);

OAI22xp33_ASAP7_75t_SL g228 ( 
.A1(n_194),
.A2(n_179),
.B1(n_178),
.B2(n_185),
.Y(n_228)
);

OAI22xp5_ASAP7_75t_SL g229 ( 
.A1(n_200),
.A2(n_127),
.B1(n_136),
.B2(n_110),
.Y(n_229)
);

AOI22xp5_ASAP7_75t_L g254 ( 
.A1(n_230),
.A2(n_234),
.B1(n_236),
.B2(n_221),
.Y(n_254)
);

AND2x2_ASAP7_75t_SL g231 ( 
.A(n_201),
.B(n_163),
.Y(n_231)
);

AND2x4_ASAP7_75t_L g244 ( 
.A(n_231),
.B(n_191),
.Y(n_244)
);

NOR2xp33_ASAP7_75t_L g232 ( 
.A(n_199),
.B(n_112),
.Y(n_232)
);

NOR2xp33_ASAP7_75t_L g247 ( 
.A(n_232),
.B(n_233),
.Y(n_247)
);

FAx1_ASAP7_75t_SL g233 ( 
.A(n_206),
.B(n_57),
.CI(n_91),
.CON(n_233),
.SN(n_233)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_190),
.Y(n_235)
);

AOI22xp33_ASAP7_75t_SL g239 ( 
.A1(n_235),
.A2(n_207),
.B1(n_213),
.B2(n_202),
.Y(n_239)
);

OAI21xp5_ASAP7_75t_SL g240 ( 
.A1(n_236),
.A2(n_211),
.B(n_210),
.Y(n_240)
);

NOR2xp33_ASAP7_75t_L g237 ( 
.A(n_193),
.B(n_177),
.Y(n_237)
);

CKINVDCx20_ASAP7_75t_R g250 ( 
.A(n_237),
.Y(n_250)
);

AO22x1_ASAP7_75t_SL g238 ( 
.A1(n_190),
.A2(n_213),
.B1(n_212),
.B2(n_206),
.Y(n_238)
);

OA21x2_ASAP7_75t_L g241 ( 
.A1(n_238),
.A2(n_50),
.B(n_70),
.Y(n_241)
);

INVxp67_ASAP7_75t_L g290 ( 
.A(n_239),
.Y(n_290)
);

AOI21xp5_ASAP7_75t_L g275 ( 
.A1(n_240),
.A2(n_238),
.B(n_233),
.Y(n_275)
);

NAND2xp5_ASAP7_75t_L g270 ( 
.A(n_241),
.B(n_244),
.Y(n_270)
);

OAI32xp33_ASAP7_75t_L g246 ( 
.A1(n_220),
.A2(n_191),
.A3(n_192),
.B1(n_204),
.B2(n_210),
.Y(n_246)
);

INVx1_ASAP7_75t_L g268 ( 
.A(n_246),
.Y(n_268)
);

XOR2xp5_ASAP7_75t_L g251 ( 
.A(n_218),
.B(n_192),
.Y(n_251)
);

MAJIxp5_ASAP7_75t_L g273 ( 
.A(n_251),
.B(n_229),
.C(n_233),
.Y(n_273)
);

AOI22xp33_ASAP7_75t_SL g252 ( 
.A1(n_221),
.A2(n_197),
.B1(n_155),
.B2(n_209),
.Y(n_252)
);

MAJIxp5_ASAP7_75t_SL g278 ( 
.A(n_252),
.B(n_257),
.C(n_188),
.Y(n_278)
);

OAI22xp5_ASAP7_75t_SL g284 ( 
.A1(n_254),
.A2(n_188),
.B1(n_214),
.B2(n_102),
.Y(n_284)
);

OAI22xp5_ASAP7_75t_SL g256 ( 
.A1(n_216),
.A2(n_136),
.B1(n_103),
.B2(n_109),
.Y(n_256)
);

AOI22xp5_ASAP7_75t_L g282 ( 
.A1(n_256),
.A2(n_259),
.B1(n_260),
.B2(n_262),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_SL g257 ( 
.A1(n_221),
.A2(n_234),
.B1(n_219),
.B2(n_214),
.Y(n_257)
);

OAI22xp5_ASAP7_75t_SL g259 ( 
.A1(n_217),
.A2(n_109),
.B1(n_103),
.B2(n_124),
.Y(n_259)
);

OAI22xp5_ASAP7_75t_SL g260 ( 
.A1(n_226),
.A2(n_237),
.B1(n_225),
.B2(n_221),
.Y(n_260)
);

CKINVDCx20_ASAP7_75t_R g261 ( 
.A(n_231),
.Y(n_261)
);

OR2x2_ASAP7_75t_L g265 ( 
.A(n_261),
.B(n_263),
.Y(n_265)
);

OAI22xp5_ASAP7_75t_L g262 ( 
.A1(n_231),
.A2(n_174),
.B1(n_180),
.B2(n_164),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g263 ( 
.A(n_231),
.Y(n_263)
);

OAI21xp5_ASAP7_75t_L g264 ( 
.A1(n_253),
.A2(n_232),
.B(n_227),
.Y(n_264)
);

OAI21xp5_ASAP7_75t_L g299 ( 
.A1(n_264),
.A2(n_275),
.B(n_288),
.Y(n_299)
);

CKINVDCx20_ASAP7_75t_R g266 ( 
.A(n_245),
.Y(n_266)
);

NAND2xp5_ASAP7_75t_SL g293 ( 
.A(n_266),
.B(n_281),
.Y(n_293)
);

AO22x2_ASAP7_75t_L g267 ( 
.A1(n_241),
.A2(n_238),
.B1(n_230),
.B2(n_235),
.Y(n_267)
);

NAND2xp5_ASAP7_75t_L g301 ( 
.A(n_267),
.B(n_283),
.Y(n_301)
);

XOR2xp5_ASAP7_75t_L g269 ( 
.A(n_243),
.B(n_224),
.Y(n_269)
);

MAJIxp5_ASAP7_75t_L g307 ( 
.A(n_269),
.B(n_273),
.C(n_274),
.Y(n_307)
);

INVx1_ASAP7_75t_L g271 ( 
.A(n_245),
.Y(n_271)
);

INVx1_ASAP7_75t_L g294 ( 
.A(n_271),
.Y(n_294)
);

NOR2xp33_ASAP7_75t_L g272 ( 
.A(n_258),
.B(n_215),
.Y(n_272)
);

INVx1_ASAP7_75t_L g316 ( 
.A(n_272),
.Y(n_316)
);

XOR2xp5_ASAP7_75t_L g274 ( 
.A(n_243),
.B(n_238),
.Y(n_274)
);

INVx1_ASAP7_75t_L g276 ( 
.A(n_246),
.Y(n_276)
);

INVx1_ASAP7_75t_L g319 ( 
.A(n_276),
.Y(n_319)
);

NAND2xp5_ASAP7_75t_L g277 ( 
.A(n_242),
.B(n_233),
.Y(n_277)
);

INVx1_ASAP7_75t_L g304 ( 
.A(n_277),
.Y(n_304)
);

HAxp5_ASAP7_75t_SL g309 ( 
.A(n_278),
.B(n_198),
.CON(n_309),
.SN(n_309)
);

INVx1_ASAP7_75t_L g279 ( 
.A(n_262),
.Y(n_279)
);

INVx1_ASAP7_75t_L g310 ( 
.A(n_279),
.Y(n_310)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_256),
.Y(n_280)
);

INVx1_ASAP7_75t_L g315 ( 
.A(n_280),
.Y(n_315)
);

NOR2xp33_ASAP7_75t_L g281 ( 
.A(n_258),
.B(n_197),
.Y(n_281)
);

AOI22xp5_ASAP7_75t_L g283 ( 
.A1(n_260),
.A2(n_259),
.B1(n_249),
.B2(n_250),
.Y(n_283)
);

AOI22xp5_ASAP7_75t_L g295 ( 
.A1(n_284),
.A2(n_291),
.B1(n_244),
.B2(n_251),
.Y(n_295)
);

INVx1_ASAP7_75t_L g285 ( 
.A(n_248),
.Y(n_285)
);

CKINVDCx16_ASAP7_75t_R g308 ( 
.A(n_285),
.Y(n_308)
);

INVx8_ASAP7_75t_L g286 ( 
.A(n_248),
.Y(n_286)
);

NOR2xp33_ASAP7_75t_L g296 ( 
.A(n_286),
.B(n_287),
.Y(n_296)
);

INVx1_ASAP7_75t_L g287 ( 
.A(n_240),
.Y(n_287)
);

OAI21xp5_ASAP7_75t_L g288 ( 
.A1(n_241),
.A2(n_222),
.B(n_181),
.Y(n_288)
);

CKINVDCx20_ASAP7_75t_R g289 ( 
.A(n_241),
.Y(n_289)
);

NOR2xp33_ASAP7_75t_SL g302 ( 
.A(n_289),
.B(n_255),
.Y(n_302)
);

AOI22xp5_ASAP7_75t_L g291 ( 
.A1(n_249),
.A2(n_250),
.B1(n_254),
.B2(n_263),
.Y(n_291)
);

AOI21xp5_ASAP7_75t_L g292 ( 
.A1(n_270),
.A2(n_261),
.B(n_247),
.Y(n_292)
);

INVxp67_ASAP7_75t_L g324 ( 
.A(n_292),
.Y(n_324)
);

OAI22xp5_ASAP7_75t_SL g323 ( 
.A1(n_295),
.A2(n_276),
.B1(n_268),
.B2(n_282),
.Y(n_323)
);

XOR2xp5_ASAP7_75t_L g297 ( 
.A(n_269),
.B(n_274),
.Y(n_297)
);

MAJIxp5_ASAP7_75t_L g321 ( 
.A(n_297),
.B(n_298),
.C(n_306),
.Y(n_321)
);

XOR2xp5_ASAP7_75t_L g298 ( 
.A(n_273),
.B(n_255),
.Y(n_298)
);

AOI21xp5_ASAP7_75t_L g300 ( 
.A1(n_270),
.A2(n_288),
.B(n_275),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g338 ( 
.A(n_300),
.Y(n_338)
);

INVx1_ASAP7_75t_L g329 ( 
.A(n_302),
.Y(n_329)
);

AND2x2_ASAP7_75t_L g303 ( 
.A(n_271),
.B(n_244),
.Y(n_303)
);

INVx1_ASAP7_75t_SL g320 ( 
.A(n_303),
.Y(n_320)
);

AOI21xp5_ASAP7_75t_L g305 ( 
.A1(n_290),
.A2(n_244),
.B(n_242),
.Y(n_305)
);

NOR2xp33_ASAP7_75t_L g341 ( 
.A(n_305),
.B(n_31),
.Y(n_341)
);

XOR2xp5_ASAP7_75t_L g306 ( 
.A(n_277),
.B(n_244),
.Y(n_306)
);

OAI22xp5_ASAP7_75t_L g322 ( 
.A1(n_309),
.A2(n_278),
.B1(n_290),
.B2(n_279),
.Y(n_322)
);

XOR2xp5_ASAP7_75t_L g311 ( 
.A(n_291),
.B(n_204),
.Y(n_311)
);

MAJIxp5_ASAP7_75t_L g326 ( 
.A(n_311),
.B(n_313),
.C(n_284),
.Y(n_326)
);

OAI21xp5_ASAP7_75t_L g312 ( 
.A1(n_265),
.A2(n_181),
.B(n_117),
.Y(n_312)
);

NAND2xp5_ASAP7_75t_SL g340 ( 
.A(n_312),
.B(n_314),
.Y(n_340)
);

MAJIxp5_ASAP7_75t_L g313 ( 
.A(n_265),
.B(n_196),
.C(n_145),
.Y(n_313)
);

OAI21xp5_ASAP7_75t_L g314 ( 
.A1(n_268),
.A2(n_181),
.B(n_117),
.Y(n_314)
);

XNOR2xp5_ASAP7_75t_L g317 ( 
.A(n_283),
.B(n_181),
.Y(n_317)
);

XNOR2xp5_ASAP7_75t_L g332 ( 
.A(n_317),
.B(n_267),
.Y(n_332)
);

OAI31xp33_ASAP7_75t_L g318 ( 
.A1(n_267),
.A2(n_50),
.A3(n_23),
.B(n_196),
.Y(n_318)
);

NAND2xp5_ASAP7_75t_L g328 ( 
.A(n_318),
.B(n_312),
.Y(n_328)
);

CKINVDCx16_ASAP7_75t_R g353 ( 
.A(n_322),
.Y(n_353)
);

AOI22xp5_ASAP7_75t_L g347 ( 
.A1(n_323),
.A2(n_335),
.B1(n_317),
.B2(n_305),
.Y(n_347)
);

INVx2_ASAP7_75t_L g325 ( 
.A(n_294),
.Y(n_325)
);

INVx1_ASAP7_75t_L g359 ( 
.A(n_325),
.Y(n_359)
);

XNOR2xp5_ASAP7_75t_L g354 ( 
.A(n_326),
.B(n_332),
.Y(n_354)
);

INVx1_ASAP7_75t_L g327 ( 
.A(n_293),
.Y(n_327)
);

INVx1_ASAP7_75t_L g360 ( 
.A(n_327),
.Y(n_360)
);

INVx1_ASAP7_75t_L g352 ( 
.A(n_328),
.Y(n_352)
);

AOI22xp5_ASAP7_75t_L g330 ( 
.A1(n_311),
.A2(n_280),
.B1(n_282),
.B2(n_267),
.Y(n_330)
);

OAI22xp5_ASAP7_75t_SL g350 ( 
.A1(n_330),
.A2(n_310),
.B1(n_314),
.B2(n_315),
.Y(n_350)
);

OAI22xp5_ASAP7_75t_L g331 ( 
.A1(n_319),
.A2(n_264),
.B1(n_286),
.B2(n_267),
.Y(n_331)
);

INVx1_ASAP7_75t_L g361 ( 
.A(n_331),
.Y(n_361)
);

FAx1_ASAP7_75t_SL g333 ( 
.A(n_306),
.B(n_23),
.CI(n_30),
.CON(n_333),
.SN(n_333)
);

NAND2xp5_ASAP7_75t_L g364 ( 
.A(n_333),
.B(n_343),
.Y(n_364)
);

NAND2xp5_ASAP7_75t_L g334 ( 
.A(n_304),
.B(n_120),
.Y(n_334)
);

INVx1_ASAP7_75t_L g356 ( 
.A(n_334),
.Y(n_356)
);

OAI22xp5_ASAP7_75t_SL g335 ( 
.A1(n_301),
.A2(n_180),
.B1(n_164),
.B2(n_124),
.Y(n_335)
);

INVx1_ASAP7_75t_L g336 ( 
.A(n_316),
.Y(n_336)
);

INVx1_ASAP7_75t_L g365 ( 
.A(n_336),
.Y(n_365)
);

MAJIxp5_ASAP7_75t_L g337 ( 
.A(n_297),
.B(n_120),
.C(n_90),
.Y(n_337)
);

MAJIxp5_ASAP7_75t_L g348 ( 
.A(n_337),
.B(n_298),
.C(n_307),
.Y(n_348)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_304),
.B(n_16),
.Y(n_339)
);

NOR2xp33_ASAP7_75t_L g349 ( 
.A(n_339),
.B(n_342),
.Y(n_349)
);

OAI21xp5_ASAP7_75t_SL g358 ( 
.A1(n_341),
.A2(n_340),
.B(n_328),
.Y(n_358)
);

NOR2xp33_ASAP7_75t_L g342 ( 
.A(n_308),
.B(n_16),
.Y(n_342)
);

INVx1_ASAP7_75t_L g343 ( 
.A(n_303),
.Y(n_343)
);

CKINVDCx20_ASAP7_75t_R g344 ( 
.A(n_303),
.Y(n_344)
);

NOR2xp33_ASAP7_75t_SL g351 ( 
.A(n_344),
.B(n_292),
.Y(n_351)
);

XOR2xp5_ASAP7_75t_L g345 ( 
.A(n_321),
.B(n_307),
.Y(n_345)
);

MAJIxp5_ASAP7_75t_L g371 ( 
.A(n_345),
.B(n_348),
.C(n_357),
.Y(n_371)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_329),
.A2(n_301),
.B1(n_295),
.B2(n_310),
.Y(n_346)
);

AOI22xp5_ASAP7_75t_L g377 ( 
.A1(n_346),
.A2(n_350),
.B1(n_355),
.B2(n_362),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g369 ( 
.A1(n_347),
.A2(n_326),
.B1(n_338),
.B2(n_320),
.Y(n_369)
);

INVx1_ASAP7_75t_L g386 ( 
.A(n_351),
.Y(n_386)
);

OAI22xp5_ASAP7_75t_SL g355 ( 
.A1(n_330),
.A2(n_299),
.B1(n_315),
.B2(n_313),
.Y(n_355)
);

MAJIxp5_ASAP7_75t_L g357 ( 
.A(n_321),
.B(n_299),
.C(n_296),
.Y(n_357)
);

NOR2xp33_ASAP7_75t_L g382 ( 
.A(n_358),
.B(n_365),
.Y(n_382)
);

OAI22xp5_ASAP7_75t_SL g362 ( 
.A1(n_324),
.A2(n_318),
.B1(n_300),
.B2(n_309),
.Y(n_362)
);

OAI22xp5_ASAP7_75t_SL g363 ( 
.A1(n_324),
.A2(n_69),
.B1(n_65),
.B2(n_61),
.Y(n_363)
);

AOI22xp5_ASAP7_75t_L g387 ( 
.A1(n_363),
.A2(n_366),
.B1(n_0),
.B2(n_1),
.Y(n_387)
);

OAI22xp5_ASAP7_75t_L g366 ( 
.A1(n_329),
.A2(n_59),
.B1(n_56),
.B2(n_49),
.Y(n_366)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_337),
.B(n_131),
.C(n_119),
.Y(n_367)
);

MAJIxp5_ASAP7_75t_L g372 ( 
.A(n_367),
.B(n_333),
.C(n_325),
.Y(n_372)
);

CKINVDCx20_ASAP7_75t_R g368 ( 
.A(n_349),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g388 ( 
.A(n_368),
.B(n_375),
.Y(n_388)
);

XNOR2xp5_ASAP7_75t_SL g389 ( 
.A(n_369),
.B(n_347),
.Y(n_389)
);

MAJIxp5_ASAP7_75t_L g370 ( 
.A(n_345),
.B(n_338),
.C(n_332),
.Y(n_370)
);

NAND2xp5_ASAP7_75t_SL g390 ( 
.A(n_370),
.B(n_376),
.Y(n_390)
);

XNOR2xp5_ASAP7_75t_L g396 ( 
.A(n_372),
.B(n_384),
.Y(n_396)
);

BUFx12_ASAP7_75t_L g373 ( 
.A(n_358),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_L g391 ( 
.A(n_373),
.B(n_381),
.Y(n_391)
);

A2O1A1O1Ixp25_ASAP7_75t_L g374 ( 
.A1(n_352),
.A2(n_320),
.B(n_334),
.C(n_323),
.D(n_333),
.Y(n_374)
);

INVx1_ASAP7_75t_L g402 ( 
.A(n_374),
.Y(n_402)
);

BUFx12f_ASAP7_75t_SL g375 ( 
.A(n_362),
.Y(n_375)
);

MAJIxp5_ASAP7_75t_L g376 ( 
.A(n_348),
.B(n_335),
.C(n_12),
.Y(n_376)
);

AND2x2_ASAP7_75t_L g378 ( 
.A(n_352),
.B(n_364),
.Y(n_378)
);

NAND2xp5_ASAP7_75t_L g401 ( 
.A(n_378),
.B(n_379),
.Y(n_401)
);

AO21x1_ASAP7_75t_L g379 ( 
.A1(n_353),
.A2(n_11),
.B(n_18),
.Y(n_379)
);

MAJIxp5_ASAP7_75t_L g380 ( 
.A(n_357),
.B(n_11),
.C(n_18),
.Y(n_380)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_380),
.B(n_359),
.C(n_364),
.Y(n_393)
);

CKINVDCx5p33_ASAP7_75t_R g381 ( 
.A(n_356),
.Y(n_381)
);

NOR2xp33_ASAP7_75t_SL g398 ( 
.A(n_382),
.B(n_385),
.Y(n_398)
);

MAJIxp5_ASAP7_75t_L g383 ( 
.A(n_354),
.B(n_23),
.C(n_31),
.Y(n_383)
);

MAJIxp5_ASAP7_75t_L g394 ( 
.A(n_383),
.B(n_367),
.C(n_355),
.Y(n_394)
);

HB1xp67_ASAP7_75t_L g384 ( 
.A(n_365),
.Y(n_384)
);

INVx2_ASAP7_75t_L g385 ( 
.A(n_360),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g395 ( 
.A1(n_387),
.A2(n_361),
.B1(n_356),
.B2(n_350),
.Y(n_395)
);

XOR2xp5_ASAP7_75t_L g407 ( 
.A(n_389),
.B(n_392),
.Y(n_407)
);

XOR2xp5_ASAP7_75t_L g392 ( 
.A(n_377),
.B(n_354),
.Y(n_392)
);

NAND2xp5_ASAP7_75t_L g409 ( 
.A(n_393),
.B(n_394),
.Y(n_409)
);

AOI22xp5_ASAP7_75t_L g408 ( 
.A1(n_395),
.A2(n_374),
.B1(n_379),
.B2(n_373),
.Y(n_408)
);

MAJIxp5_ASAP7_75t_L g397 ( 
.A(n_371),
.B(n_363),
.C(n_23),
.Y(n_397)
);

MAJIxp5_ASAP7_75t_L g406 ( 
.A(n_397),
.B(n_400),
.C(n_381),
.Y(n_406)
);

XNOR2xp5_ASAP7_75t_L g399 ( 
.A(n_371),
.B(n_11),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_L g412 ( 
.A(n_399),
.B(n_14),
.Y(n_412)
);

MAJIxp5_ASAP7_75t_L g400 ( 
.A(n_383),
.B(n_23),
.C(n_30),
.Y(n_400)
);

AOI21xp5_ASAP7_75t_SL g403 ( 
.A1(n_391),
.A2(n_375),
.B(n_378),
.Y(n_403)
);

CKINVDCx20_ASAP7_75t_R g419 ( 
.A(n_403),
.Y(n_419)
);

AOI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_402),
.A2(n_386),
.B1(n_373),
.B2(n_372),
.Y(n_404)
);

AND2x2_ASAP7_75t_L g425 ( 
.A(n_404),
.B(n_410),
.Y(n_425)
);

CKINVDCx20_ASAP7_75t_R g405 ( 
.A(n_388),
.Y(n_405)
);

NAND2xp5_ASAP7_75t_L g417 ( 
.A(n_405),
.B(n_406),
.Y(n_417)
);

INVx1_ASAP7_75t_L g424 ( 
.A(n_408),
.Y(n_424)
);

AOI22xp33_ASAP7_75t_SL g410 ( 
.A1(n_401),
.A2(n_30),
.B1(n_9),
.B2(n_12),
.Y(n_410)
);

MAJIxp5_ASAP7_75t_L g411 ( 
.A(n_392),
.B(n_23),
.C(n_9),
.Y(n_411)
);

NOR2xp33_ASAP7_75t_L g423 ( 
.A(n_411),
.B(n_412),
.Y(n_423)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_390),
.A2(n_8),
.B1(n_15),
.B2(n_14),
.Y(n_413)
);

NOR2xp33_ASAP7_75t_L g426 ( 
.A(n_413),
.B(n_415),
.Y(n_426)
);

NOR2xp33_ASAP7_75t_L g414 ( 
.A(n_398),
.B(n_14),
.Y(n_414)
);

NOR2xp33_ASAP7_75t_L g427 ( 
.A(n_414),
.B(n_13),
.Y(n_427)
);

NOR2xp33_ASAP7_75t_SL g415 ( 
.A(n_396),
.B(n_17),
.Y(n_415)
);

XNOR2x1_ASAP7_75t_L g416 ( 
.A(n_407),
.B(n_394),
.Y(n_416)
);

MAJIxp5_ASAP7_75t_L g432 ( 
.A(n_416),
.B(n_12),
.C(n_8),
.Y(n_432)
);

NOR2x1_ASAP7_75t_SL g418 ( 
.A(n_403),
.B(n_409),
.Y(n_418)
);

INVx1_ASAP7_75t_L g428 ( 
.A(n_418),
.Y(n_428)
);

XNOR2xp5_ASAP7_75t_SL g420 ( 
.A(n_407),
.B(n_389),
.Y(n_420)
);

NAND2xp5_ASAP7_75t_SL g431 ( 
.A(n_420),
.B(n_422),
.Y(n_431)
);

NOR2xp33_ASAP7_75t_SL g421 ( 
.A(n_406),
.B(n_397),
.Y(n_421)
);

INVx1_ASAP7_75t_L g436 ( 
.A(n_421),
.Y(n_436)
);

MAJIxp5_ASAP7_75t_L g422 ( 
.A(n_411),
.B(n_400),
.C(n_17),
.Y(n_422)
);

NAND2xp5_ASAP7_75t_L g430 ( 
.A(n_427),
.B(n_13),
.Y(n_430)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_419),
.B(n_410),
.Y(n_429)
);

INVx1_ASAP7_75t_L g440 ( 
.A(n_429),
.Y(n_440)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_430),
.Y(n_442)
);

NAND2xp5_ASAP7_75t_SL g441 ( 
.A(n_432),
.B(n_433),
.Y(n_441)
);

NAND2xp5_ASAP7_75t_SL g433 ( 
.A(n_417),
.B(n_424),
.Y(n_433)
);

NOR2xp33_ASAP7_75t_SL g434 ( 
.A(n_426),
.B(n_0),
.Y(n_434)
);

NOR2x1_ASAP7_75t_L g439 ( 
.A(n_434),
.B(n_431),
.Y(n_439)
);

OAI22xp5_ASAP7_75t_L g435 ( 
.A1(n_425),
.A2(n_6),
.B1(n_3),
.B2(n_4),
.Y(n_435)
);

AOI21xp5_ASAP7_75t_L g437 ( 
.A1(n_435),
.A2(n_427),
.B(n_426),
.Y(n_437)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_437),
.B(n_439),
.Y(n_443)
);

OAI21xp5_ASAP7_75t_SL g438 ( 
.A1(n_428),
.A2(n_423),
.B(n_3),
.Y(n_438)
);

XNOR2x2_ASAP7_75t_SL g446 ( 
.A(n_438),
.B(n_5),
.Y(n_446)
);

OAI22xp5_ASAP7_75t_L g444 ( 
.A1(n_440),
.A2(n_436),
.B1(n_429),
.B2(n_5),
.Y(n_444)
);

NAND2x1_ASAP7_75t_L g448 ( 
.A(n_444),
.B(n_445),
.Y(n_448)
);

OAI22xp5_ASAP7_75t_L g445 ( 
.A1(n_441),
.A2(n_2),
.B1(n_4),
.B2(n_5),
.Y(n_445)
);

CKINVDCx20_ASAP7_75t_R g447 ( 
.A(n_446),
.Y(n_447)
);

INVx1_ASAP7_75t_L g449 ( 
.A(n_448),
.Y(n_449)
);

CKINVDCx20_ASAP7_75t_R g450 ( 
.A(n_449),
.Y(n_450)
);

AOI21xp5_ASAP7_75t_L g451 ( 
.A1(n_450),
.A2(n_443),
.B(n_447),
.Y(n_451)
);

MAJIxp5_ASAP7_75t_L g452 ( 
.A(n_451),
.B(n_442),
.C(n_6),
.Y(n_452)
);


endmodule