module real_aes_5800_n_249 (n_17, n_28, n_226, n_76, n_202, n_149, n_56, n_113, n_34, n_98, n_121, n_120, n_125, n_187, n_190, n_90, n_216, n_82, n_238, n_65, n_47, n_74, n_106, n_58, n_185, n_134, n_32, n_30, n_230, n_165, n_51, n_195, n_246, n_248, n_176, n_27, n_163, n_222, n_61, n_29, n_20, n_52, n_221, n_174, n_156, n_57, n_64, n_66, n_18, n_207, n_104, n_21, n_31, n_8, n_183, n_205, n_220, n_211, n_10, n_177, n_83, n_181, n_197, n_124, n_22, n_173, n_191, n_209, n_3, n_41, n_140, n_234, n_153, n_75, n_178, n_219, n_19, n_71, n_180, n_40, n_49, n_212, n_210, n_239, n_126, n_91, n_100, n_43, n_103, n_166, n_200, n_224, n_151, n_115, n_96, n_110, n_130, n_54, n_112, n_35, n_42, n_147, n_150, n_99, n_15, n_9, n_23, n_72, n_132, n_119, n_160, n_95, n_131, n_144, n_164, n_231, n_169, n_242, n_44, n_102, n_188, n_152, n_198, n_201, n_122, n_7, n_228, n_196, n_141, n_128, n_172, n_111, n_158, n_4, n_232, n_167, n_123, n_80, n_179, n_6, n_12, n_68, n_129, n_162, n_79, n_193, n_214, n_69, n_46, n_109, n_59, n_25, n_203, n_236, n_73, n_77, n_218, n_81, n_133, n_48, n_204, n_37, n_117, n_208, n_97, n_215, n_135, n_186, n_70, n_138, n_50, n_114, n_89, n_170, n_26, n_235, n_86, n_93, n_182, n_154, n_127, n_199, n_245, n_161, n_189, n_13, n_24, n_217, n_2, n_142, n_55, n_168, n_175, n_241, n_145, n_62, n_105, n_223, n_84, n_227, n_67, n_92, n_33, n_206, n_148, n_88, n_14, n_159, n_11, n_85, n_108, n_194, n_137, n_225, n_16, n_116, n_94, n_229, n_39, n_5, n_45, n_60, n_233, n_240, n_247, n_38, n_155, n_243, n_118, n_143, n_139, n_244, n_192, n_213, n_136, n_87, n_171, n_0, n_157, n_78, n_101, n_63, n_1, n_146, n_237, n_107, n_184, n_53, n_36, n_249);
input n_17;
input n_28;
input n_226;
input n_76;
input n_202;
input n_149;
input n_56;
input n_113;
input n_34;
input n_98;
input n_121;
input n_120;
input n_125;
input n_187;
input n_190;
input n_90;
input n_216;
input n_82;
input n_238;
input n_65;
input n_47;
input n_74;
input n_106;
input n_58;
input n_185;
input n_134;
input n_32;
input n_30;
input n_230;
input n_165;
input n_51;
input n_195;
input n_246;
input n_248;
input n_176;
input n_27;
input n_163;
input n_222;
input n_61;
input n_29;
input n_20;
input n_52;
input n_221;
input n_174;
input n_156;
input n_57;
input n_64;
input n_66;
input n_18;
input n_207;
input n_104;
input n_21;
input n_31;
input n_8;
input n_183;
input n_205;
input n_220;
input n_211;
input n_10;
input n_177;
input n_83;
input n_181;
input n_197;
input n_124;
input n_22;
input n_173;
input n_191;
input n_209;
input n_3;
input n_41;
input n_140;
input n_234;
input n_153;
input n_75;
input n_178;
input n_219;
input n_19;
input n_71;
input n_180;
input n_40;
input n_49;
input n_212;
input n_210;
input n_239;
input n_126;
input n_91;
input n_100;
input n_43;
input n_103;
input n_166;
input n_200;
input n_224;
input n_151;
input n_115;
input n_96;
input n_110;
input n_130;
input n_54;
input n_112;
input n_35;
input n_42;
input n_147;
input n_150;
input n_99;
input n_15;
input n_9;
input n_23;
input n_72;
input n_132;
input n_119;
input n_160;
input n_95;
input n_131;
input n_144;
input n_164;
input n_231;
input n_169;
input n_242;
input n_44;
input n_102;
input n_188;
input n_152;
input n_198;
input n_201;
input n_122;
input n_7;
input n_228;
input n_196;
input n_141;
input n_128;
input n_172;
input n_111;
input n_158;
input n_4;
input n_232;
input n_167;
input n_123;
input n_80;
input n_179;
input n_6;
input n_12;
input n_68;
input n_129;
input n_162;
input n_79;
input n_193;
input n_214;
input n_69;
input n_46;
input n_109;
input n_59;
input n_25;
input n_203;
input n_236;
input n_73;
input n_77;
input n_218;
input n_81;
input n_133;
input n_48;
input n_204;
input n_37;
input n_117;
input n_208;
input n_97;
input n_215;
input n_135;
input n_186;
input n_70;
input n_138;
input n_50;
input n_114;
input n_89;
input n_170;
input n_26;
input n_235;
input n_86;
input n_93;
input n_182;
input n_154;
input n_127;
input n_199;
input n_245;
input n_161;
input n_189;
input n_13;
input n_24;
input n_217;
input n_2;
input n_142;
input n_55;
input n_168;
input n_175;
input n_241;
input n_145;
input n_62;
input n_105;
input n_223;
input n_84;
input n_227;
input n_67;
input n_92;
input n_33;
input n_206;
input n_148;
input n_88;
input n_14;
input n_159;
input n_11;
input n_85;
input n_108;
input n_194;
input n_137;
input n_225;
input n_16;
input n_116;
input n_94;
input n_229;
input n_39;
input n_5;
input n_45;
input n_60;
input n_233;
input n_240;
input n_247;
input n_38;
input n_155;
input n_243;
input n_118;
input n_143;
input n_139;
input n_244;
input n_192;
input n_213;
input n_136;
input n_87;
input n_171;
input n_0;
input n_157;
input n_78;
input n_101;
input n_63;
input n_1;
input n_146;
input n_237;
input n_107;
input n_184;
input n_53;
input n_36;
output n_249;
wire n_480;
wire n_476;
wire n_758;
wire n_599;
wire n_436;
wire n_887;
wire n_684;
wire n_257;
wire n_390;
wire n_821;
wire n_830;
wire n_285;
wire n_624;
wire n_618;
wire n_800;
wire n_778;
wire n_522;
wire n_838;
wire n_933;
wire n_485;
wire n_822;
wire n_846;
wire n_750;
wire n_631;
wire n_943;
wire n_357;
wire n_503;
wire n_635;
wire n_287;
wire n_386;
wire n_673;
wire n_905;
wire n_518;
wire n_254;
wire n_792;
wire n_878;
wire n_665;
wire n_667;
wire n_580;
wire n_577;
wire n_469;
wire n_362;
wire n_759;
wire n_445;
wire n_596;
wire n_592;
wire n_540;
wire n_657;
wire n_299;
wire n_322;
wire n_900;
wire n_328;
wire n_718;
wire n_318;
wire n_841;
wire n_355;
wire n_669;
wire n_423;
wire n_458;
wire n_444;
wire n_736;
wire n_761;
wire n_742;
wire n_319;
wire n_364;
wire n_421;
wire n_555;
wire n_329;
wire n_766;
wire n_852;
wire n_857;
wire n_919;
wire n_461;
wire n_908;
wire n_376;
wire n_549;
wire n_571;
wire n_694;
wire n_308;
wire n_491;
wire n_894;
wire n_923;
wire n_429;
wire n_752;
wire n_448;
wire n_545;
wire n_556;
wire n_341;
wire n_593;
wire n_460;
wire n_937;
wire n_773;
wire n_401;
wire n_538;
wire n_317;
wire n_353;
wire n_431;
wire n_321;
wire n_865;
wire n_551;
wire n_320;
wire n_537;
wire n_666;
wire n_884;
wire n_560;
wire n_260;
wire n_660;
wire n_814;
wire n_944;
wire n_886;
wire n_594;
wire n_856;
wire n_767;
wire n_696;
wire n_889;
wire n_704;
wire n_941;
wire n_453;
wire n_374;
wire n_379;
wire n_647;
wire n_932;
wire n_399;
wire n_948;
wire n_700;
wire n_677;
wire n_378;
wire n_591;
wire n_775;
wire n_763;
wire n_870;
wire n_271;
wire n_489;
wire n_548;
wire n_427;
wire n_678;
wire n_415;
wire n_572;
wire n_519;
wire n_564;
wire n_638;
wire n_815;
wire n_573;
wire n_510;
wire n_709;
wire n_330;
wire n_388;
wire n_786;
wire n_512;
wire n_395;
wire n_332;
wire n_795;
wire n_626;
wire n_292;
wire n_539;
wire n_400;
wire n_816;
wire n_625;
wire n_289;
wire n_462;
wire n_280;
wire n_615;
wire n_550;
wire n_333;
wire n_670;
wire n_818;
wire n_716;
wire n_918;
wire n_356;
wire n_478;
wire n_883;
wire n_584;
wire n_896;
wire n_408;
wire n_553;
wire n_372;
wire n_528;
wire n_578;
wire n_892;
wire n_495;
wire n_370;
wire n_384;
wire n_744;
wire n_938;
wire n_352;
wire n_935;
wire n_824;
wire n_467;
wire n_875;
wire n_327;
wire n_774;
wire n_813;
wire n_791;
wire n_466;
wire n_559;
wire n_636;
wire n_872;
wire n_906;
wire n_263;
wire n_477;
wire n_515;
wire n_680;
wire n_595;
wire n_301;
wire n_343;
wire n_369;
wire n_726;
wire n_517;
wire n_683;
wire n_780;
wire n_904;
wire n_840;
wire n_570;
wire n_675;
wire n_931;
wire n_920;
wire n_530;
wire n_835;
wire n_535;
wire n_732;
wire n_834;
wire n_882;
wire n_784;
wire n_281;
wire n_496;
wire n_693;
wire n_468;
wire n_746;
wire n_284;
wire n_316;
wire n_532;
wire n_656;
wire n_755;
wire n_409;
wire n_860;
wire n_748;
wire n_909;
wire n_298;
wire n_523;
wire n_781;
wire n_439;
wire n_576;
wire n_924;
wire n_506;
wire n_606;
wire n_513;
wire n_651;
wire n_796;
wire n_874;
wire n_297;
wire n_801;
wire n_383;
wire n_529;
wire n_310;
wire n_455;
wire n_504;
wire n_725;
wire n_671;
wire n_547;
wire n_659;
wire n_682;
wire n_634;
wire n_903;
wire n_454;
wire n_812;
wire n_782;
wire n_443;
wire n_565;
wire n_817;
wire n_760;
wire n_608;
wire n_925;
wire n_534;
wire n_708;
wire n_457;
wire n_345;
wire n_304;
wire n_885;
wire n_381;
wire n_493;
wire n_311;
wire n_324;
wire n_664;
wire n_278;
wire n_367;
wire n_819;
wire n_267;
wire n_737;
wire n_581;
wire n_610;
wire n_936;
wire n_620;
wire n_582;
wire n_641;
wire n_828;
wire n_808;
wire n_770;
wire n_940;
wire n_745;
wire n_722;
wire n_867;
wire n_339;
wire n_398;
wire n_688;
wire n_277;
wire n_609;
wire n_425;
wire n_879;
wire n_331;
wire n_363;
wire n_417;
wire n_449;
wire n_607;
wire n_754;
wire n_323;
wire n_690;
wire n_629;
wire n_499;
wire n_508;
wire n_350;
wire n_706;
wire n_901;
wire n_561;
wire n_947;
wire n_876;
wire n_437;
wire n_428;
wire n_405;
wire n_621;
wire n_368;
wire n_783;
wire n_655;
wire n_654;
wire n_527;
wire n_434;
wire n_502;
wire n_505;
wire n_769;
wire n_600;
wire n_731;
wire n_250;
wire n_605;
wire n_672;
wire n_567;
wire n_916;
wire n_406;
wire n_426;
wire n_602;
wire n_402;
wire n_552;
wire n_617;
wire n_733;
wire n_676;
wire n_658;
wire n_531;
wire n_616;
wire n_590;
wire n_451;
wire n_432;
wire n_880;
wire n_807;
wire n_255;
wire n_286;
wire n_416;
wire n_790;
wire n_895;
wire n_832;
wire n_410;
wire n_799;
wire n_805;
wire n_751;
wire n_490;
wire n_261;
wire n_913;
wire n_619;
wire n_391;
wire n_360;
wire n_859;
wire n_695;
wire n_685;
wire n_881;
wire n_917;
wire n_361;
wire n_632;
wire n_768;
wire n_412;
wire n_542;
wire n_645;
wire n_557;
wire n_714;
wire n_777;
wire n_501;
wire n_488;
wire n_910;
wire n_251;
wire n_642;
wire n_613;
wire n_387;
wire n_296;
wire n_702;
wire n_256;
wire n_912;
wire n_302;
wire n_464;
wire n_351;
wire n_945;
wire n_898;
wire n_604;
wire n_734;
wire n_848;
wire n_392;
wire n_562;
wire n_288;
wire n_404;
wire n_598;
wire n_713;
wire n_728;
wire n_735;
wire n_756;
wire n_334;
wire n_274;
wire n_303;
wire n_569;
wire n_563;
wire n_785;
wire n_891;
wire n_269;
wire n_430;
wire n_568;
wire n_413;
wire n_471;
wire n_902;
wire n_853;
wire n_810;
wire n_843;
wire n_306;
wire n_579;
wire n_699;
wire n_533;
wire n_366;
wire n_346;
wire n_727;
wire n_397;
wire n_293;
wire n_358;
wire n_385;
wire n_275;
wire n_649;
wire n_663;
wire n_749;
wire n_588;
wire n_536;
wire n_914;
wire n_707;
wire n_622;
wire n_915;
wire n_470;
wire n_851;
wire n_934;
wire n_494;
wire n_711;
wire n_864;
wire n_377;
wire n_273;
wire n_927;
wire n_723;
wire n_662;
wire n_276;
wire n_295;
wire n_382;
wire n_845;
wire n_850;
wire n_265;
wire n_354;
wire n_720;
wire n_435;
wire n_511;
wire n_484;
wire n_326;
wire n_893;
wire n_492;
wire n_509;
wire n_407;
wire n_419;
wire n_730;
wire n_643;
wire n_747;
wire n_486;
wire n_930;
wire n_411;
wire n_697;
wire n_291;
wire n_847;
wire n_907;
wire n_779;
wire n_481;
wire n_498;
wire n_691;
wire n_765;
wire n_826;
wire n_648;
wire n_373;
wire n_589;
wire n_628;
wire n_939;
wire n_487;
wire n_831;
wire n_290;
wire n_365;
wire n_899;
wire n_526;
wire n_637;
wire n_653;
wire n_928;
wire n_692;
wire n_544;
wire n_268;
wire n_789;
wire n_282;
wire n_389;
wire n_738;
wire n_701;
wire n_309;
wire n_344;
wire n_827;
wire n_809;
wire n_922;
wire n_520;
wire n_482;
wire n_633;
wire n_926;
wire n_679;
wire n_942;
wire n_472;
wire n_866;
wire n_452;
wire n_787;
wire n_262;
wire n_630;
wire n_806;
wire n_689;
wire n_820;
wire n_715;
wire n_946;
wire n_349;
wire n_336;
wire n_420;
wire n_612;
wire n_858;
wire n_873;
wire n_438;
wire n_764;
wire n_794;
wire n_300;
wire n_252;
wire n_283;
wire n_314;
wire n_753;
wire n_741;
wire n_623;
wire n_446;
wire n_721;
wire n_681;
wire n_359;
wire n_456;
wire n_717;
wire n_312;
wire n_266;
wire n_712;
wire n_433;
wire n_335;
wire n_516;
wire n_313;
wire n_627;
wire n_739;
wire n_418;
wire n_521;
wire n_422;
wire n_771;
wire n_524;
wire n_861;
wire n_705;
wire n_575;
wire n_325;
wire n_762;
wire n_338;
wire n_479;
wire n_442;
wire n_825;
wire n_698;
wire n_371;
wire n_740;
wire n_541;
wire n_839;
wire n_546;
wire n_587;
wire n_639;
wire n_811;
wire n_253;
wire n_459;
wire n_558;
wire n_863;
wire n_724;
wire n_440;
wire n_525;
wire n_644;
wire n_674;
wire n_888;
wire n_836;
wire n_793;
wire n_272;
wire n_583;
wire n_347;
wire n_315;
wire n_833;
wire n_414;
wire n_757;
wire n_929;
wire n_279;
wire n_686;
wire n_776;
wire n_803;
wire n_890;
wire n_543;
wire n_497;
wire n_514;
wire n_507;
wire n_270;
wire n_614;
wire n_305;
wire n_586;
wire n_911;
wire n_772;
wire n_450;
wire n_788;
wire n_441;
wire n_585;
wire n_465;
wire n_473;
wire n_719;
wire n_566;
wire n_837;
wire n_871;
wire n_474;
wire n_829;
wire n_921;
wire n_375;
wire n_597;
wire n_340;
wire n_640;
wire n_483;
wire n_611;
wire n_380;
wire n_394;
wire n_687;
wire n_729;
wire n_844;
wire n_646;
wire n_650;
wire n_710;
wire n_743;
wire n_823;
wire n_393;
wire n_294;
wire n_258;
wire n_652;
wire n_703;
wire n_500;
wire n_307;
wire n_601;
wire n_661;
wire n_463;
wire n_396;
wire n_804;
wire n_447;
wire n_342;
wire n_348;
wire n_603;
wire n_403;
wire n_854;
wire n_424;
wire n_877;
wire n_802;
wire n_868;
wire n_574;
wire n_337;
wire n_842;
wire n_259;
wire n_849;
wire n_475;
wire n_554;
wire n_897;
wire n_264;
wire n_855;
wire n_798;
wire n_668;
wire n_797;
wire n_862;
wire n_869;
INVx1_ASAP7_75t_SL g400 ( .A(n_0), .Y(n_400) );
AOI22xp33_ASAP7_75t_SL g691 ( .A1(n_0), .A2(n_39), .B1(n_684), .B2(n_685), .Y(n_691) );
HB1xp67_ASAP7_75t_L g643 ( .A(n_1), .Y(n_643) );
AND2x4_ASAP7_75t_L g647 ( .A(n_1), .B(n_648), .Y(n_647) );
AND2x4_ASAP7_75t_L g660 ( .A(n_1), .B(n_243), .Y(n_660) );
AOI22xp33_ASAP7_75t_L g608 ( .A1(n_2), .A2(n_93), .B1(n_327), .B2(n_333), .Y(n_608) );
AOI22xp33_ASAP7_75t_L g557 ( .A1(n_3), .A2(n_131), .B1(n_372), .B2(n_558), .Y(n_557) );
AOI22xp33_ASAP7_75t_L g571 ( .A1(n_4), .A2(n_49), .B1(n_507), .B2(n_558), .Y(n_571) );
AOI22xp33_ASAP7_75t_L g708 ( .A1(n_5), .A2(n_98), .B1(n_657), .B2(n_661), .Y(n_708) );
NAND2xp5_ASAP7_75t_L g526 ( .A(n_6), .B(n_527), .Y(n_526) );
AOI22xp33_ASAP7_75t_L g538 ( .A1(n_7), .A2(n_188), .B1(n_348), .B2(n_539), .Y(n_538) );
INVx1_ASAP7_75t_L g417 ( .A(n_8), .Y(n_417) );
AOI21xp5_ASAP7_75t_L g547 ( .A1(n_9), .A2(n_548), .B(n_549), .Y(n_547) );
AOI22xp5_ASAP7_75t_L g623 ( .A1(n_10), .A2(n_204), .B1(n_375), .B2(n_576), .Y(n_623) );
INVx1_ASAP7_75t_L g460 ( .A(n_11), .Y(n_460) );
AOI22xp5_ASAP7_75t_L g505 ( .A1(n_12), .A2(n_23), .B1(n_506), .B2(n_507), .Y(n_505) );
AOI22xp33_ASAP7_75t_L g447 ( .A1(n_13), .A2(n_110), .B1(n_365), .B2(n_448), .Y(n_447) );
AOI22xp33_ASAP7_75t_L g552 ( .A1(n_14), .A2(n_220), .B1(n_363), .B2(n_541), .Y(n_552) );
AOI22xp33_ASAP7_75t_L g578 ( .A1(n_15), .A2(n_150), .B1(n_579), .B2(n_580), .Y(n_578) );
AOI22xp5_ASAP7_75t_L g369 ( .A1(n_16), .A2(n_177), .B1(n_370), .B2(n_372), .Y(n_369) );
AOI22xp33_ASAP7_75t_L g385 ( .A1(n_17), .A2(n_190), .B1(n_386), .B2(n_388), .Y(n_385) );
AOI22xp33_ASAP7_75t_L g559 ( .A1(n_18), .A2(n_141), .B1(n_375), .B2(n_501), .Y(n_559) );
AOI22xp33_ASAP7_75t_L g875 ( .A1(n_19), .A2(n_103), .B1(n_580), .B2(n_876), .Y(n_875) );
AOI22xp5_ASAP7_75t_L g467 ( .A1(n_20), .A2(n_54), .B1(n_286), .B2(n_298), .Y(n_467) );
INVx1_ASAP7_75t_L g523 ( .A(n_21), .Y(n_523) );
AOI22xp33_ASAP7_75t_L g259 ( .A1(n_22), .A2(n_90), .B1(n_260), .B2(n_283), .Y(n_259) );
AOI22xp5_ASAP7_75t_L g690 ( .A1(n_24), .A2(n_95), .B1(n_680), .B2(n_682), .Y(n_690) );
INVx1_ASAP7_75t_L g767 ( .A(n_25), .Y(n_767) );
AOI222xp33_ASAP7_75t_L g863 ( .A1(n_25), .A2(n_864), .B1(n_900), .B2(n_903), .C1(n_906), .C2(n_946), .Y(n_863) );
AO22x2_ASAP7_75t_L g908 ( .A1(n_25), .A2(n_767), .B1(n_909), .B2(n_945), .Y(n_908) );
INVx1_ASAP7_75t_L g280 ( .A(n_26), .Y(n_280) );
INVxp67_ASAP7_75t_L g305 ( .A(n_26), .Y(n_305) );
NOR2xp33_ASAP7_75t_L g312 ( .A(n_26), .B(n_191), .Y(n_312) );
AOI22xp33_ASAP7_75t_L g534 ( .A1(n_27), .A2(n_111), .B1(n_372), .B2(n_506), .Y(n_534) );
AOI22xp33_ASAP7_75t_L g625 ( .A1(n_28), .A2(n_202), .B1(n_525), .B2(n_579), .Y(n_625) );
CKINVDCx5p33_ASAP7_75t_R g878 ( .A(n_29), .Y(n_878) );
AOI22xp33_ASAP7_75t_L g894 ( .A1(n_30), .A2(n_83), .B1(n_895), .B2(n_897), .Y(n_894) );
AOI21xp33_ASAP7_75t_SL g487 ( .A1(n_31), .A2(n_488), .B(n_489), .Y(n_487) );
AOI22xp5_ASAP7_75t_L g437 ( .A1(n_32), .A2(n_136), .B1(n_370), .B2(n_438), .Y(n_437) );
AOI22xp5_ASAP7_75t_L g683 ( .A1(n_33), .A2(n_174), .B1(n_684), .B2(n_685), .Y(n_683) );
AOI22xp33_ASAP7_75t_L g768 ( .A1(n_34), .A2(n_234), .B1(n_673), .B2(n_676), .Y(n_768) );
AOI221xp5_ASAP7_75t_L g599 ( .A1(n_35), .A2(n_63), .B1(n_260), .B2(n_283), .C(n_600), .Y(n_599) );
NAND2xp5_ASAP7_75t_L g584 ( .A(n_36), .B(n_585), .Y(n_584) );
AOI22xp5_ASAP7_75t_L g569 ( .A1(n_37), .A2(n_96), .B1(n_330), .B2(n_570), .Y(n_569) );
NAND2xp5_ASAP7_75t_SL g276 ( .A(n_38), .B(n_264), .Y(n_276) );
AOI22xp33_ASAP7_75t_L g356 ( .A1(n_40), .A2(n_237), .B1(n_357), .B2(n_359), .Y(n_356) );
OAI21x1_ASAP7_75t_L g591 ( .A1(n_41), .A2(n_592), .B(n_609), .Y(n_591) );
NAND4xp25_ASAP7_75t_L g609 ( .A(n_41), .B(n_593), .C(n_598), .D(n_605), .Y(n_609) );
AOI221xp5_ASAP7_75t_L g347 ( .A1(n_42), .A2(n_66), .B1(n_348), .B2(n_350), .C(n_353), .Y(n_347) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_43), .A2(n_225), .B1(n_363), .B2(n_365), .Y(n_362) );
AOI22xp5_ASAP7_75t_L g573 ( .A1(n_44), .A2(n_166), .B1(n_574), .B2(n_576), .Y(n_573) );
AOI22xp33_ASAP7_75t_L g285 ( .A1(n_45), .A2(n_77), .B1(n_286), .B2(n_288), .Y(n_285) );
AOI22xp33_ASAP7_75t_L g594 ( .A1(n_46), .A2(n_172), .B1(n_576), .B2(n_595), .Y(n_594) );
AOI22xp33_ASAP7_75t_L g656 ( .A1(n_47), .A2(n_107), .B1(n_657), .B2(n_661), .Y(n_656) );
NAND2xp33_ASAP7_75t_L g463 ( .A(n_48), .B(n_464), .Y(n_463) );
AOI22xp33_ASAP7_75t_L g535 ( .A1(n_50), .A2(n_152), .B1(n_509), .B2(n_536), .Y(n_535) );
AOI22xp33_ASAP7_75t_L g540 ( .A1(n_51), .A2(n_97), .B1(n_363), .B2(n_541), .Y(n_540) );
INVx2_ASAP7_75t_L g641 ( .A(n_52), .Y(n_641) );
XNOR2x1_ASAP7_75t_L g427 ( .A(n_53), .B(n_428), .Y(n_427) );
AOI22xp33_ASAP7_75t_L g494 ( .A1(n_55), .A2(n_200), .B1(n_357), .B2(n_359), .Y(n_494) );
AOI21xp33_ASAP7_75t_L g586 ( .A1(n_56), .A2(n_587), .B(n_588), .Y(n_586) );
AND2x4_ASAP7_75t_L g649 ( .A(n_57), .B(n_641), .Y(n_649) );
INVx1_ASAP7_75t_L g659 ( .A(n_57), .Y(n_659) );
INVx1_ASAP7_75t_SL g681 ( .A(n_57), .Y(n_681) );
INVx1_ASAP7_75t_L g422 ( .A(n_58), .Y(n_422) );
AOI22xp33_ASAP7_75t_L g334 ( .A1(n_59), .A2(n_197), .B1(n_335), .B2(n_336), .Y(n_334) );
AOI22xp5_ASAP7_75t_L g374 ( .A1(n_60), .A2(n_61), .B1(n_375), .B2(n_377), .Y(n_374) );
XNOR2x1_ASAP7_75t_L g544 ( .A(n_62), .B(n_545), .Y(n_544) );
AOI21xp5_ASAP7_75t_L g519 ( .A1(n_64), .A2(n_520), .B(n_522), .Y(n_519) );
AOI22xp33_ASAP7_75t_L g916 ( .A1(n_65), .A2(n_156), .B1(n_917), .B2(n_918), .Y(n_916) );
AOI22xp5_ASAP7_75t_L g606 ( .A1(n_67), .A2(n_147), .B1(n_558), .B2(n_607), .Y(n_606) );
BUFx6f_ASAP7_75t_L g264 ( .A(n_68), .Y(n_264) );
AOI22xp33_ASAP7_75t_SL g296 ( .A1(n_69), .A2(n_142), .B1(n_297), .B2(n_298), .Y(n_296) );
INVx1_ASAP7_75t_L g476 ( .A(n_70), .Y(n_476) );
AOI22xp33_ASAP7_75t_L g604 ( .A1(n_71), .A2(n_173), .B1(n_286), .B2(n_288), .Y(n_604) );
AOI22xp5_ASAP7_75t_L g465 ( .A1(n_72), .A2(n_182), .B1(n_297), .B2(n_466), .Y(n_465) );
AOI22xp5_ASAP7_75t_L g694 ( .A1(n_73), .A2(n_148), .B1(n_684), .B2(n_685), .Y(n_694) );
AOI22xp33_ASAP7_75t_L g603 ( .A1(n_74), .A2(n_167), .B1(n_297), .B2(n_298), .Y(n_603) );
AOI22xp5_ASAP7_75t_L g596 ( .A1(n_75), .A2(n_235), .B1(n_330), .B2(n_597), .Y(n_596) );
INVx1_ASAP7_75t_L g670 ( .A(n_76), .Y(n_670) );
AOI22xp5_ASAP7_75t_L g621 ( .A1(n_78), .A2(n_219), .B1(n_570), .B2(n_622), .Y(n_621) );
NAND2xp5_ASAP7_75t_L g424 ( .A(n_79), .B(n_298), .Y(n_424) );
AOI22xp33_ASAP7_75t_L g430 ( .A1(n_80), .A2(n_124), .B1(n_382), .B2(n_431), .Y(n_430) );
AOI22xp33_ASAP7_75t_L g450 ( .A1(n_81), .A2(n_114), .B1(n_451), .B2(n_453), .Y(n_450) );
AOI22xp5_ASAP7_75t_L g679 ( .A1(n_82), .A2(n_244), .B1(n_680), .B2(n_682), .Y(n_679) );
INVx1_ASAP7_75t_L g268 ( .A(n_84), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g302 ( .A(n_84), .B(n_189), .Y(n_302) );
AOI22xp33_ASAP7_75t_L g936 ( .A1(n_85), .A2(n_161), .B1(n_937), .B2(n_939), .Y(n_936) );
AOI22xp5_ASAP7_75t_L g700 ( .A1(n_86), .A2(n_92), .B1(n_680), .B2(n_682), .Y(n_700) );
AOI22xp33_ASAP7_75t_L g555 ( .A1(n_87), .A2(n_154), .B1(n_435), .B2(n_556), .Y(n_555) );
INVx1_ASAP7_75t_L g601 ( .A(n_88), .Y(n_601) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_89), .A2(n_94), .B1(n_386), .B2(n_503), .Y(n_502) );
INVx1_ASAP7_75t_L g589 ( .A(n_91), .Y(n_589) );
AOI22xp33_ASAP7_75t_L g407 ( .A1(n_99), .A2(n_170), .B1(n_318), .B2(n_332), .Y(n_407) );
INVx1_ASAP7_75t_L g766 ( .A(n_100), .Y(n_766) );
AOI22xp5_ASAP7_75t_L g326 ( .A1(n_101), .A2(n_238), .B1(n_327), .B2(n_330), .Y(n_326) );
NAND2xp5_ASAP7_75t_L g445 ( .A(n_102), .B(n_446), .Y(n_445) );
AOI22xp33_ASAP7_75t_L g699 ( .A1(n_104), .A2(n_194), .B1(n_676), .B2(n_684), .Y(n_699) );
CKINVDCx5p33_ASAP7_75t_R g871 ( .A(n_105), .Y(n_871) );
AOI22xp5_ASAP7_75t_L g581 ( .A1(n_106), .A2(n_201), .B1(n_582), .B2(n_583), .Y(n_581) );
INVxp33_ASAP7_75t_SL g677 ( .A(n_108), .Y(n_677) );
INVx1_ASAP7_75t_L g630 ( .A(n_109), .Y(n_630) );
XNOR2x1_ASAP7_75t_L g614 ( .A(n_112), .B(n_615), .Y(n_614) );
AOI22xp33_ASAP7_75t_L g867 ( .A1(n_113), .A2(n_119), .B1(n_868), .B2(n_869), .Y(n_867) );
AOI22xp33_ASAP7_75t_L g662 ( .A1(n_115), .A2(n_151), .B1(n_663), .B2(n_664), .Y(n_662) );
AOI22xp33_ASAP7_75t_L g911 ( .A1(n_116), .A2(n_133), .B1(n_375), .B2(n_912), .Y(n_911) );
CKINVDCx20_ASAP7_75t_R g542 ( .A(n_117), .Y(n_542) );
AOI22xp33_ASAP7_75t_L g560 ( .A1(n_118), .A2(n_240), .B1(n_386), .B2(n_438), .Y(n_560) );
AOI22xp33_ASAP7_75t_L g499 ( .A1(n_120), .A2(n_129), .B1(n_500), .B2(n_501), .Y(n_499) );
AOI22xp33_ASAP7_75t_L g531 ( .A1(n_121), .A2(n_171), .B1(n_377), .B2(n_500), .Y(n_531) );
AOI22xp33_ASAP7_75t_L g885 ( .A1(n_122), .A2(n_138), .B1(n_595), .B2(n_886), .Y(n_885) );
AOI22xp33_ASAP7_75t_L g331 ( .A1(n_123), .A2(n_217), .B1(n_332), .B2(n_333), .Y(n_331) );
AOI22xp5_ASAP7_75t_L g317 ( .A1(n_125), .A2(n_199), .B1(n_318), .B2(n_324), .Y(n_317) );
AOI22xp5_ASAP7_75t_L g470 ( .A1(n_126), .A2(n_196), .B1(n_327), .B2(n_333), .Y(n_470) );
AOI22xp33_ASAP7_75t_L g617 ( .A1(n_127), .A2(n_211), .B1(n_370), .B2(n_372), .Y(n_617) );
AOI22xp5_ASAP7_75t_L g379 ( .A1(n_128), .A2(n_213), .B1(n_380), .B2(n_382), .Y(n_379) );
AOI22xp33_ASAP7_75t_L g532 ( .A1(n_130), .A2(n_218), .B1(n_386), .B2(n_438), .Y(n_532) );
INVx1_ASAP7_75t_L g419 ( .A(n_132), .Y(n_419) );
AOI22xp33_ASAP7_75t_L g495 ( .A1(n_134), .A2(n_139), .B1(n_496), .B2(n_497), .Y(n_495) );
AOI22xp33_ASAP7_75t_L g890 ( .A1(n_135), .A2(n_245), .B1(n_891), .B2(n_893), .Y(n_890) );
AOI22xp33_ASAP7_75t_L g572 ( .A1(n_137), .A2(n_206), .B1(n_327), .B2(n_333), .Y(n_572) );
AOI22xp33_ASAP7_75t_SL g940 ( .A1(n_140), .A2(n_168), .B1(n_941), .B2(n_943), .Y(n_940) );
CKINVDCx5p33_ASAP7_75t_R g881 ( .A(n_143), .Y(n_881) );
AOI22xp5_ASAP7_75t_L g469 ( .A1(n_144), .A2(n_157), .B1(n_324), .B2(n_330), .Y(n_469) );
INVx1_ASAP7_75t_L g674 ( .A(n_145), .Y(n_674) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_146), .B(n_484), .Y(n_483) );
CKINVDCx14_ASAP7_75t_R g255 ( .A(n_148), .Y(n_255) );
AOI22xp33_ASAP7_75t_L g913 ( .A1(n_149), .A2(n_183), .B1(n_914), .B2(n_915), .Y(n_913) );
AOI22xp33_ASAP7_75t_L g432 ( .A1(n_153), .A2(n_223), .B1(n_433), .B2(n_435), .Y(n_432) );
NAND2xp5_ASAP7_75t_L g306 ( .A(n_155), .B(n_307), .Y(n_306) );
INVx1_ASAP7_75t_L g415 ( .A(n_158), .Y(n_415) );
AOI22xp5_ASAP7_75t_L g618 ( .A1(n_159), .A2(n_222), .B1(n_386), .B2(n_619), .Y(n_618) );
AOI221xp5_ASAP7_75t_L g627 ( .A1(n_160), .A2(n_207), .B1(n_448), .B2(n_628), .C(n_629), .Y(n_627) );
AOI22xp33_ASAP7_75t_L g408 ( .A1(n_162), .A2(n_229), .B1(n_327), .B2(n_333), .Y(n_408) );
INVx1_ASAP7_75t_L g443 ( .A(n_163), .Y(n_443) );
NAND2xp5_ASAP7_75t_L g551 ( .A(n_164), .B(n_527), .Y(n_551) );
OA22x2_ASAP7_75t_L g262 ( .A1(n_165), .A2(n_191), .B1(n_263), .B2(n_264), .Y(n_262) );
INVx1_ASAP7_75t_L g293 ( .A(n_165), .Y(n_293) );
AOI21xp5_ASAP7_75t_SL g413 ( .A1(n_169), .A2(n_260), .B(n_414), .Y(n_413) );
AOI22xp33_ASAP7_75t_L g707 ( .A1(n_175), .A2(n_242), .B1(n_663), .B2(n_664), .Y(n_707) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_176), .A2(n_192), .B1(n_335), .B2(n_336), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g436 ( .A1(n_178), .A2(n_239), .B1(n_375), .B2(n_377), .Y(n_436) );
AOI21xp5_ASAP7_75t_L g925 ( .A1(n_179), .A2(n_926), .B(n_929), .Y(n_925) );
INVx1_ASAP7_75t_L g935 ( .A(n_180), .Y(n_935) );
INVx1_ASAP7_75t_L g932 ( .A(n_181), .Y(n_932) );
INVx1_ASAP7_75t_L g490 ( .A(n_184), .Y(n_490) );
OAI22xp5_ASAP7_75t_L g864 ( .A1(n_185), .A2(n_865), .B1(n_898), .B2(n_899), .Y(n_864) );
CKINVDCx5p33_ASAP7_75t_R g898 ( .A(n_185), .Y(n_898) );
AOI22xp33_ASAP7_75t_L g508 ( .A1(n_186), .A2(n_214), .B1(n_435), .B2(n_509), .Y(n_508) );
AOI22xp33_ASAP7_75t_L g553 ( .A1(n_187), .A2(n_232), .B1(n_451), .B2(n_539), .Y(n_553) );
INVx1_ASAP7_75t_L g282 ( .A(n_189), .Y(n_282) );
NAND2xp5_ASAP7_75t_L g315 ( .A(n_189), .B(n_291), .Y(n_315) );
OAI21xp33_ASAP7_75t_L g294 ( .A1(n_191), .A2(n_210), .B(n_295), .Y(n_294) );
INVx1_ASAP7_75t_L g411 ( .A(n_193), .Y(n_411) );
CKINVDCx5p33_ASAP7_75t_R g344 ( .A(n_194), .Y(n_344) );
AOI22xp5_ASAP7_75t_L g405 ( .A1(n_195), .A2(n_230), .B1(n_324), .B2(n_330), .Y(n_405) );
AOI22xp5_ASAP7_75t_L g472 ( .A1(n_198), .A2(n_208), .B1(n_335), .B2(n_336), .Y(n_472) );
AOI22xp5_ASAP7_75t_L g693 ( .A1(n_203), .A2(n_216), .B1(n_680), .B2(n_682), .Y(n_693) );
INVx1_ASAP7_75t_L g480 ( .A(n_205), .Y(n_480) );
AOI22xp5_ASAP7_75t_L g473 ( .A1(n_209), .A2(n_247), .B1(n_318), .B2(n_332), .Y(n_473) );
INVx1_ASAP7_75t_L g270 ( .A(n_210), .Y(n_270) );
NOR2xp33_ASAP7_75t_L g313 ( .A(n_210), .B(n_236), .Y(n_313) );
CKINVDCx16_ASAP7_75t_R g550 ( .A(n_212), .Y(n_550) );
AOI22xp5_ASAP7_75t_L g626 ( .A1(n_215), .A2(n_224), .B1(n_582), .B2(n_583), .Y(n_626) );
AOI21xp5_ASAP7_75t_L g440 ( .A1(n_221), .A2(n_441), .B(n_442), .Y(n_440) );
INVx1_ASAP7_75t_L g566 ( .A(n_226), .Y(n_566) );
AOI22xp33_ASAP7_75t_L g887 ( .A1(n_227), .A2(n_248), .B1(n_619), .B2(n_888), .Y(n_887) );
AOI22xp33_ASAP7_75t_L g920 ( .A1(n_228), .A2(n_233), .B1(n_921), .B2(n_922), .Y(n_920) );
AOI21xp33_ASAP7_75t_SL g474 ( .A1(n_231), .A2(n_260), .B(n_475), .Y(n_474) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_236), .B(n_275), .Y(n_274) );
INVxp33_ASAP7_75t_L g669 ( .A(n_241), .Y(n_669) );
INVx1_ASAP7_75t_L g648 ( .A(n_243), .Y(n_648) );
CKINVDCx20_ASAP7_75t_R g354 ( .A(n_246), .Y(n_354) );
O2A1O1Ixp33_ASAP7_75t_SL g249 ( .A1(n_250), .A2(n_513), .B(n_635), .C(n_644), .Y(n_249) );
AOI21xp5_ASAP7_75t_L g635 ( .A1(n_250), .A2(n_513), .B(n_636), .Y(n_635) );
XNOR2xp5_ASAP7_75t_L g250 ( .A(n_251), .B(n_394), .Y(n_250) );
INVx2_ASAP7_75t_SL g251 ( .A(n_252), .Y(n_251) );
AO22x2_ASAP7_75t_L g252 ( .A1(n_253), .A2(n_340), .B1(n_391), .B2(n_393), .Y(n_252) );
INVx2_ASAP7_75t_L g393 ( .A(n_253), .Y(n_393) );
INVx2_ASAP7_75t_L g253 ( .A(n_254), .Y(n_253) );
OAI21x1_ASAP7_75t_L g254 ( .A1(n_255), .A2(n_256), .B(n_337), .Y(n_254) );
NAND3xp33_ASAP7_75t_SL g337 ( .A(n_255), .B(n_338), .C(n_339), .Y(n_337) );
INVx1_ASAP7_75t_L g256 ( .A(n_257), .Y(n_256) );
OR2x2_ASAP7_75t_L g257 ( .A(n_258), .B(n_316), .Y(n_257) );
INVx1_ASAP7_75t_L g339 ( .A(n_258), .Y(n_339) );
NAND4xp25_ASAP7_75t_L g258 ( .A(n_259), .B(n_285), .C(n_296), .D(n_306), .Y(n_258) );
AND2x2_ASAP7_75t_L g260 ( .A(n_261), .B(n_271), .Y(n_260) );
AND2x4_ASAP7_75t_L g286 ( .A(n_261), .B(n_287), .Y(n_286) );
AND2x4_ASAP7_75t_L g349 ( .A(n_261), .B(n_287), .Y(n_349) );
AND2x4_ASAP7_75t_L g364 ( .A(n_261), .B(n_271), .Y(n_364) );
AND2x2_ASAP7_75t_L g261 ( .A(n_262), .B(n_265), .Y(n_261) );
AND2x2_ASAP7_75t_L g284 ( .A(n_262), .B(n_266), .Y(n_284) );
AND2x2_ASAP7_75t_L g303 ( .A(n_262), .B(n_304), .Y(n_303) );
INVx1_ASAP7_75t_L g320 ( .A(n_262), .Y(n_320) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_263), .B(n_270), .Y(n_269) );
INVx2_ASAP7_75t_L g263 ( .A(n_264), .Y(n_263) );
NAND2xp33_ASAP7_75t_L g267 ( .A(n_264), .B(n_268), .Y(n_267) );
INVx3_ASAP7_75t_L g275 ( .A(n_264), .Y(n_275) );
NAND2xp33_ASAP7_75t_L g281 ( .A(n_264), .B(n_282), .Y(n_281) );
INVx1_ASAP7_75t_L g295 ( .A(n_264), .Y(n_295) );
HB1xp67_ASAP7_75t_L g301 ( .A(n_264), .Y(n_301) );
AND2x4_ASAP7_75t_L g319 ( .A(n_265), .B(n_320), .Y(n_319) );
INVx1_ASAP7_75t_L g265 ( .A(n_266), .Y(n_265) );
NAND2xp5_ASAP7_75t_L g266 ( .A(n_267), .B(n_269), .Y(n_266) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_268), .B(n_293), .Y(n_292) );
OAI21xp5_ASAP7_75t_L g304 ( .A1(n_270), .A2(n_295), .B(n_305), .Y(n_304) );
AND2x2_ASAP7_75t_L g283 ( .A(n_271), .B(n_284), .Y(n_283) );
AND2x4_ASAP7_75t_L g288 ( .A(n_271), .B(n_289), .Y(n_288) );
AND2x4_ASAP7_75t_L g336 ( .A(n_271), .B(n_319), .Y(n_336) );
AND2x2_ASAP7_75t_L g352 ( .A(n_271), .B(n_284), .Y(n_352) );
AND2x4_ASAP7_75t_L g367 ( .A(n_271), .B(n_289), .Y(n_367) );
AND2x2_ASAP7_75t_L g378 ( .A(n_271), .B(n_319), .Y(n_378) );
AND2x4_ASAP7_75t_L g271 ( .A(n_272), .B(n_277), .Y(n_271) );
INVx2_ASAP7_75t_L g272 ( .A(n_273), .Y(n_272) );
AND2x4_ASAP7_75t_L g287 ( .A(n_273), .B(n_277), .Y(n_287) );
AND2x2_ASAP7_75t_L g299 ( .A(n_273), .B(n_300), .Y(n_299) );
OR2x2_ASAP7_75t_L g322 ( .A(n_273), .B(n_323), .Y(n_322) );
AND2x4_ASAP7_75t_L g328 ( .A(n_273), .B(n_329), .Y(n_328) );
AND2x4_ASAP7_75t_L g273 ( .A(n_274), .B(n_276), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g279 ( .A(n_275), .B(n_280), .Y(n_279) );
INVxp67_ASAP7_75t_L g291 ( .A(n_275), .Y(n_291) );
NAND3xp33_ASAP7_75t_L g314 ( .A(n_276), .B(n_290), .C(n_315), .Y(n_314) );
INVx1_ASAP7_75t_L g277 ( .A(n_278), .Y(n_277) );
INVx1_ASAP7_75t_L g323 ( .A(n_278), .Y(n_323) );
AND2x2_ASAP7_75t_L g278 ( .A(n_279), .B(n_281), .Y(n_278) );
INVx2_ASAP7_75t_L g412 ( .A(n_283), .Y(n_412) );
HB1xp67_ASAP7_75t_L g464 ( .A(n_283), .Y(n_464) );
AND2x4_ASAP7_75t_L g297 ( .A(n_284), .B(n_287), .Y(n_297) );
AND2x4_ASAP7_75t_L g327 ( .A(n_284), .B(n_328), .Y(n_327) );
AND2x4_ASAP7_75t_L g330 ( .A(n_284), .B(n_325), .Y(n_330) );
AND2x2_ASAP7_75t_L g358 ( .A(n_284), .B(n_287), .Y(n_358) );
AND2x4_ASAP7_75t_L g381 ( .A(n_284), .B(n_321), .Y(n_381) );
AND2x2_ASAP7_75t_L g387 ( .A(n_284), .B(n_328), .Y(n_387) );
AND2x2_ASAP7_75t_L g434 ( .A(n_284), .B(n_328), .Y(n_434) );
INVx2_ASAP7_75t_L g418 ( .A(n_286), .Y(n_418) );
AND2x4_ASAP7_75t_L g335 ( .A(n_287), .B(n_319), .Y(n_335) );
AND2x4_ASAP7_75t_L g376 ( .A(n_287), .B(n_319), .Y(n_376) );
INVx2_ASAP7_75t_L g420 ( .A(n_288), .Y(n_420) );
AND2x4_ASAP7_75t_L g324 ( .A(n_289), .B(n_325), .Y(n_324) );
AND2x4_ASAP7_75t_L g333 ( .A(n_289), .B(n_328), .Y(n_333) );
AND2x4_ASAP7_75t_L g384 ( .A(n_289), .B(n_325), .Y(n_384) );
AND2x4_ASAP7_75t_L g390 ( .A(n_289), .B(n_328), .Y(n_390) );
AND2x2_ASAP7_75t_L g289 ( .A(n_290), .B(n_294), .Y(n_289) );
NAND2xp5_ASAP7_75t_L g290 ( .A(n_291), .B(n_292), .Y(n_290) );
INVx1_ASAP7_75t_L g423 ( .A(n_297), .Y(n_423) );
INVx4_ASAP7_75t_L g444 ( .A(n_298), .Y(n_444) );
AND2x4_ASAP7_75t_L g298 ( .A(n_299), .B(n_303), .Y(n_298) );
AND2x4_ASAP7_75t_L g361 ( .A(n_299), .B(n_303), .Y(n_361) );
NAND2xp5_ASAP7_75t_L g300 ( .A(n_301), .B(n_302), .Y(n_300) );
INVx1_ASAP7_75t_L g310 ( .A(n_301), .Y(n_310) );
INVx2_ASAP7_75t_SL g631 ( .A(n_307), .Y(n_631) );
INVx2_ASAP7_75t_SL g307 ( .A(n_308), .Y(n_307) );
BUFx6f_ASAP7_75t_L g355 ( .A(n_308), .Y(n_355) );
NOR2xp33_ASAP7_75t_L g414 ( .A(n_308), .B(n_415), .Y(n_414) );
INVx2_ASAP7_75t_L g492 ( .A(n_308), .Y(n_492) );
BUFx6f_ASAP7_75t_L g308 ( .A(n_309), .Y(n_308) );
INVx3_ASAP7_75t_L g529 ( .A(n_309), .Y(n_529) );
AO21x2_ASAP7_75t_L g309 ( .A1(n_310), .A2(n_311), .B(n_314), .Y(n_309) );
HB1xp67_ASAP7_75t_L g642 ( .A(n_311), .Y(n_642) );
NAND2xp5_ASAP7_75t_L g311 ( .A(n_312), .B(n_313), .Y(n_311) );
INVxp67_ASAP7_75t_L g338 ( .A(n_316), .Y(n_338) );
NAND4xp25_ASAP7_75t_L g316 ( .A(n_317), .B(n_326), .C(n_331), .D(n_334), .Y(n_316) );
AND2x4_ASAP7_75t_L g318 ( .A(n_319), .B(n_321), .Y(n_318) );
AND2x4_ASAP7_75t_L g332 ( .A(n_319), .B(n_328), .Y(n_332) );
AND2x4_ASAP7_75t_L g371 ( .A(n_319), .B(n_328), .Y(n_371) );
AND2x4_ASAP7_75t_L g373 ( .A(n_319), .B(n_325), .Y(n_373) );
INVx2_ASAP7_75t_L g321 ( .A(n_322), .Y(n_321) );
INVx2_ASAP7_75t_L g325 ( .A(n_322), .Y(n_325) );
INVx1_ASAP7_75t_L g329 ( .A(n_323), .Y(n_329) );
INVxp67_ASAP7_75t_SL g340 ( .A(n_341), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_342), .Y(n_341) );
INVx1_ASAP7_75t_L g342 ( .A(n_343), .Y(n_342) );
INVxp67_ASAP7_75t_SL g392 ( .A(n_343), .Y(n_392) );
XNOR2x1_ASAP7_75t_L g343 ( .A(n_344), .B(n_345), .Y(n_343) );
OR2x2_ASAP7_75t_L g345 ( .A(n_346), .B(n_368), .Y(n_345) );
NAND3xp33_ASAP7_75t_L g346 ( .A(n_347), .B(n_356), .C(n_362), .Y(n_346) );
BUFx6f_ASAP7_75t_L g348 ( .A(n_349), .Y(n_348) );
INVx1_ASAP7_75t_L g452 ( .A(n_349), .Y(n_452) );
BUFx3_ASAP7_75t_L g579 ( .A(n_349), .Y(n_579) );
BUFx3_ASAP7_75t_L g942 ( .A(n_349), .Y(n_942) );
INVx2_ASAP7_75t_L g521 ( .A(n_350), .Y(n_521) );
INVx2_ASAP7_75t_L g350 ( .A(n_351), .Y(n_350) );
INVx2_ASAP7_75t_L g441 ( .A(n_351), .Y(n_441) );
INVx2_ASAP7_75t_L g585 ( .A(n_351), .Y(n_585) );
INVx3_ASAP7_75t_L g351 ( .A(n_352), .Y(n_351) );
INVx2_ASAP7_75t_L g486 ( .A(n_352), .Y(n_486) );
BUFx3_ASAP7_75t_L g874 ( .A(n_352), .Y(n_874) );
NOR2xp33_ASAP7_75t_L g353 ( .A(n_354), .B(n_355), .Y(n_353) );
INVx2_ASAP7_75t_L g446 ( .A(n_355), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g475 ( .A(n_355), .B(n_476), .Y(n_475) );
INVx2_ASAP7_75t_L g944 ( .A(n_357), .Y(n_944) );
BUFx3_ASAP7_75t_L g357 ( .A(n_358), .Y(n_357) );
INVx2_ASAP7_75t_L g454 ( .A(n_358), .Y(n_454) );
BUFx6f_ASAP7_75t_L g539 ( .A(n_358), .Y(n_539) );
INVx2_ASAP7_75t_L g359 ( .A(n_360), .Y(n_359) );
INVx4_ASAP7_75t_L g525 ( .A(n_360), .Y(n_525) );
INVx2_ASAP7_75t_L g931 ( .A(n_360), .Y(n_931) );
INVx5_ASAP7_75t_L g360 ( .A(n_361), .Y(n_360) );
BUFx4f_ASAP7_75t_L g580 ( .A(n_361), .Y(n_580) );
BUFx3_ASAP7_75t_L g363 ( .A(n_364), .Y(n_363) );
INVx2_ASAP7_75t_L g449 ( .A(n_364), .Y(n_449) );
BUFx6f_ASAP7_75t_L g587 ( .A(n_364), .Y(n_587) );
INVx2_ASAP7_75t_L g896 ( .A(n_364), .Y(n_896) );
BUFx8_ASAP7_75t_SL g938 ( .A(n_364), .Y(n_938) );
INVx2_ASAP7_75t_L g365 ( .A(n_366), .Y(n_365) );
INVx3_ASAP7_75t_L g541 ( .A(n_366), .Y(n_541) );
INVx2_ASAP7_75t_L g897 ( .A(n_366), .Y(n_897) );
INVx3_ASAP7_75t_L g366 ( .A(n_367), .Y(n_366) );
BUFx6f_ASAP7_75t_L g497 ( .A(n_367), .Y(n_497) );
BUFx6f_ASAP7_75t_L g583 ( .A(n_367), .Y(n_583) );
NAND4xp25_ASAP7_75t_SL g368 ( .A(n_369), .B(n_374), .C(n_379), .D(n_385), .Y(n_368) );
BUFx2_ASAP7_75t_SL g917 ( .A(n_370), .Y(n_917) );
BUFx6f_ASAP7_75t_L g370 ( .A(n_371), .Y(n_370) );
BUFx6f_ASAP7_75t_L g506 ( .A(n_371), .Y(n_506) );
BUFx12f_ASAP7_75t_L g558 ( .A(n_371), .Y(n_558) );
BUFx3_ASAP7_75t_L g914 ( .A(n_372), .Y(n_914) );
BUFx6f_ASAP7_75t_L g372 ( .A(n_373), .Y(n_372) );
BUFx6f_ASAP7_75t_L g431 ( .A(n_373), .Y(n_431) );
BUFx6f_ASAP7_75t_L g507 ( .A(n_373), .Y(n_507) );
BUFx6f_ASAP7_75t_L g607 ( .A(n_373), .Y(n_607) );
BUFx12f_ASAP7_75t_L g375 ( .A(n_376), .Y(n_375) );
BUFx6f_ASAP7_75t_L g500 ( .A(n_376), .Y(n_500) );
INVx3_ASAP7_75t_L g575 ( .A(n_376), .Y(n_575) );
BUFx6f_ASAP7_75t_L g377 ( .A(n_378), .Y(n_377) );
BUFx5_ASAP7_75t_L g501 ( .A(n_378), .Y(n_501) );
BUFx3_ASAP7_75t_L g576 ( .A(n_378), .Y(n_576) );
BUFx6f_ASAP7_75t_L g380 ( .A(n_381), .Y(n_380) );
BUFx6f_ASAP7_75t_L g435 ( .A(n_381), .Y(n_435) );
BUFx3_ASAP7_75t_L g536 ( .A(n_381), .Y(n_536) );
BUFx6f_ASAP7_75t_L g622 ( .A(n_381), .Y(n_622) );
BUFx12f_ASAP7_75t_L g923 ( .A(n_381), .Y(n_923) );
INVx2_ASAP7_75t_L g382 ( .A(n_383), .Y(n_382) );
INVx5_ASAP7_75t_L g556 ( .A(n_383), .Y(n_556) );
INVx2_ASAP7_75t_L g570 ( .A(n_383), .Y(n_570) );
INVx3_ASAP7_75t_L g597 ( .A(n_383), .Y(n_597) );
INVx6_ASAP7_75t_L g383 ( .A(n_384), .Y(n_383) );
BUFx12f_ASAP7_75t_L g509 ( .A(n_384), .Y(n_509) );
BUFx3_ASAP7_75t_L g921 ( .A(n_386), .Y(n_921) );
BUFx6f_ASAP7_75t_L g386 ( .A(n_387), .Y(n_386) );
BUFx8_ASAP7_75t_L g888 ( .A(n_387), .Y(n_888) );
INVx4_ASAP7_75t_L g388 ( .A(n_389), .Y(n_388) );
INVx4_ASAP7_75t_L g438 ( .A(n_389), .Y(n_438) );
INVx2_ASAP7_75t_L g503 ( .A(n_389), .Y(n_503) );
INVx4_ASAP7_75t_L g619 ( .A(n_389), .Y(n_619) );
INVx2_ASAP7_75t_L g919 ( .A(n_389), .Y(n_919) );
INVx8_ASAP7_75t_L g389 ( .A(n_390), .Y(n_389) );
INVx1_ASAP7_75t_L g391 ( .A(n_392), .Y(n_391) );
AOI22xp5_ASAP7_75t_L g394 ( .A1(n_395), .A2(n_457), .B1(n_511), .B2(n_512), .Y(n_394) );
INVx1_ASAP7_75t_L g511 ( .A(n_395), .Y(n_511) );
OAI22xp5_ASAP7_75t_L g395 ( .A1(n_396), .A2(n_425), .B1(n_426), .B2(n_455), .Y(n_395) );
INVx1_ASAP7_75t_L g396 ( .A(n_397), .Y(n_396) );
INVx1_ASAP7_75t_L g456 ( .A(n_397), .Y(n_456) );
INVx1_ASAP7_75t_L g397 ( .A(n_398), .Y(n_397) );
INVx1_ASAP7_75t_L g398 ( .A(n_399), .Y(n_398) );
XNOR2x1_ASAP7_75t_L g399 ( .A(n_400), .B(n_401), .Y(n_399) );
AND2x2_ASAP7_75t_L g401 ( .A(n_402), .B(n_409), .Y(n_401) );
NOR2xp33_ASAP7_75t_L g402 ( .A(n_403), .B(n_406), .Y(n_402) );
NAND2xp5_ASAP7_75t_L g403 ( .A(n_404), .B(n_405), .Y(n_403) );
NAND2xp5_ASAP7_75t_L g406 ( .A(n_407), .B(n_408), .Y(n_406) );
NOR3xp33_ASAP7_75t_L g409 ( .A(n_410), .B(n_416), .C(n_421), .Y(n_409) );
OAI21xp33_ASAP7_75t_L g410 ( .A1(n_411), .A2(n_412), .B(n_413), .Y(n_410) );
INVx2_ASAP7_75t_L g628 ( .A(n_412), .Y(n_628) );
OAI22xp33_ASAP7_75t_L g416 ( .A1(n_417), .A2(n_418), .B1(n_419), .B2(n_420), .Y(n_416) );
INVxp67_ASAP7_75t_L g466 ( .A(n_420), .Y(n_466) );
OAI21xp5_ASAP7_75t_SL g421 ( .A1(n_422), .A2(n_423), .B(n_424), .Y(n_421) );
INVx2_ASAP7_75t_L g425 ( .A(n_426), .Y(n_425) );
INVx1_ASAP7_75t_L g426 ( .A(n_427), .Y(n_426) );
OR2x2_ASAP7_75t_L g428 ( .A(n_429), .B(n_439), .Y(n_428) );
NAND4xp25_ASAP7_75t_L g429 ( .A(n_430), .B(n_432), .C(n_436), .D(n_437), .Y(n_429) );
HB1xp67_ASAP7_75t_L g880 ( .A(n_431), .Y(n_880) );
BUFx4f_ASAP7_75t_L g433 ( .A(n_434), .Y(n_433) );
NAND3xp33_ASAP7_75t_SL g439 ( .A(n_440), .B(n_447), .C(n_450), .Y(n_439) );
OAI21xp5_ASAP7_75t_L g442 ( .A1(n_443), .A2(n_444), .B(n_445), .Y(n_442) );
OAI21xp5_ASAP7_75t_L g549 ( .A1(n_444), .A2(n_550), .B(n_551), .Y(n_549) );
INVx2_ASAP7_75t_SL g448 ( .A(n_449), .Y(n_448) );
INVx2_ASAP7_75t_SL g496 ( .A(n_449), .Y(n_496) );
INVx2_ASAP7_75t_L g451 ( .A(n_452), .Y(n_451) );
INVx2_ASAP7_75t_L g488 ( .A(n_452), .Y(n_488) );
INVx1_ASAP7_75t_L g453 ( .A(n_454), .Y(n_453) );
INVx2_ASAP7_75t_L g582 ( .A(n_454), .Y(n_582) );
INVx1_ASAP7_75t_L g455 ( .A(n_456), .Y(n_455) );
INVx1_ASAP7_75t_L g512 ( .A(n_457), .Y(n_512) );
OA22x2_ASAP7_75t_L g457 ( .A1(n_458), .A2(n_477), .B1(n_478), .B2(n_510), .Y(n_457) );
INVx2_ASAP7_75t_SL g510 ( .A(n_458), .Y(n_510) );
INVx3_ASAP7_75t_SL g458 ( .A(n_459), .Y(n_458) );
XNOR2x1_ASAP7_75t_L g459 ( .A(n_460), .B(n_461), .Y(n_459) );
NOR2x1_ASAP7_75t_L g461 ( .A(n_462), .B(n_468), .Y(n_461) );
NAND3xp33_ASAP7_75t_L g462 ( .A(n_463), .B(n_465), .C(n_467), .Y(n_462) );
NAND4xp25_ASAP7_75t_SL g468 ( .A(n_469), .B(n_470), .C(n_471), .D(n_474), .Y(n_468) );
AND2x2_ASAP7_75t_L g471 ( .A(n_472), .B(n_473), .Y(n_471) );
INVx1_ASAP7_75t_L g477 ( .A(n_478), .Y(n_477) );
INVx2_ASAP7_75t_SL g478 ( .A(n_479), .Y(n_478) );
XNOR2x1_ASAP7_75t_L g479 ( .A(n_480), .B(n_481), .Y(n_479) );
NOR4xp75_ASAP7_75t_L g481 ( .A(n_482), .B(n_493), .C(n_498), .D(n_504), .Y(n_481) );
NAND2xp5_ASAP7_75t_L g482 ( .A(n_483), .B(n_487), .Y(n_482) );
INVx2_ASAP7_75t_L g484 ( .A(n_485), .Y(n_484) );
INVx2_ASAP7_75t_L g548 ( .A(n_485), .Y(n_548) );
INVx2_ASAP7_75t_L g928 ( .A(n_485), .Y(n_928) );
BUFx6f_ASAP7_75t_L g485 ( .A(n_486), .Y(n_485) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_490), .B(n_491), .Y(n_489) );
INVx3_ASAP7_75t_L g491 ( .A(n_492), .Y(n_491) );
NAND2xp5_ASAP7_75t_L g493 ( .A(n_494), .B(n_495), .Y(n_493) );
BUFx3_ASAP7_75t_L g939 ( .A(n_497), .Y(n_939) );
NAND2xp5_ASAP7_75t_SL g498 ( .A(n_499), .B(n_502), .Y(n_498) );
BUFx3_ASAP7_75t_L g912 ( .A(n_501), .Y(n_912) );
NAND2xp5_ASAP7_75t_SL g504 ( .A(n_505), .B(n_508), .Y(n_504) );
BUFx3_ASAP7_75t_L g915 ( .A(n_509), .Y(n_915) );
XNOR2xp5_ASAP7_75t_L g513 ( .A(n_514), .B(n_562), .Y(n_513) );
OAI22xp33_ASAP7_75t_SL g514 ( .A1(n_515), .A2(n_516), .B1(n_543), .B2(n_561), .Y(n_514) );
INVx2_ASAP7_75t_SL g515 ( .A(n_516), .Y(n_515) );
INVx1_ASAP7_75t_L g516 ( .A(n_517), .Y(n_516) );
XNOR2x1_ASAP7_75t_L g517 ( .A(n_518), .B(n_542), .Y(n_517) );
NAND4xp75_ASAP7_75t_L g518 ( .A(n_519), .B(n_530), .C(n_533), .D(n_537), .Y(n_518) );
INVx1_ASAP7_75t_L g520 ( .A(n_521), .Y(n_520) );
OAI21xp5_ASAP7_75t_L g522 ( .A1(n_523), .A2(n_524), .B(n_526), .Y(n_522) );
INVx2_ASAP7_75t_L g524 ( .A(n_525), .Y(n_524) );
INVx4_ASAP7_75t_L g527 ( .A(n_528), .Y(n_527) );
INVx1_ASAP7_75t_L g876 ( .A(n_528), .Y(n_876) );
INVx4_ASAP7_75t_L g528 ( .A(n_529), .Y(n_528) );
INVx3_ASAP7_75t_L g590 ( .A(n_529), .Y(n_590) );
AND2x2_ASAP7_75t_L g530 ( .A(n_531), .B(n_532), .Y(n_530) );
AND2x2_ASAP7_75t_L g533 ( .A(n_534), .B(n_535), .Y(n_533) );
AND2x2_ASAP7_75t_L g537 ( .A(n_538), .B(n_540), .Y(n_537) );
BUFx3_ASAP7_75t_L g893 ( .A(n_539), .Y(n_893) );
INVx1_ASAP7_75t_L g561 ( .A(n_543), .Y(n_561) );
INVx1_ASAP7_75t_L g543 ( .A(n_544), .Y(n_543) );
OR2x2_ASAP7_75t_L g545 ( .A(n_546), .B(n_554), .Y(n_545) );
NAND3xp33_ASAP7_75t_L g546 ( .A(n_547), .B(n_552), .C(n_553), .Y(n_546) );
NAND4xp25_ASAP7_75t_SL g554 ( .A(n_555), .B(n_557), .C(n_559), .D(n_560), .Y(n_554) );
BUFx6f_ASAP7_75t_L g883 ( .A(n_558), .Y(n_883) );
AO22x2_ASAP7_75t_L g562 ( .A1(n_563), .A2(n_611), .B1(n_632), .B2(n_634), .Y(n_562) );
INVx1_ASAP7_75t_L g634 ( .A(n_563), .Y(n_634) );
AO22x2_ASAP7_75t_L g563 ( .A1(n_564), .A2(n_565), .B1(n_591), .B2(n_610), .Y(n_563) );
INVx2_ASAP7_75t_L g564 ( .A(n_565), .Y(n_564) );
XNOR2x1_ASAP7_75t_L g565 ( .A(n_566), .B(n_567), .Y(n_565) );
NOR2x1_ASAP7_75t_L g567 ( .A(n_568), .B(n_577), .Y(n_567) );
NAND4xp25_ASAP7_75t_L g568 ( .A(n_569), .B(n_571), .C(n_572), .D(n_573), .Y(n_568) );
HB1xp67_ASAP7_75t_L g869 ( .A(n_570), .Y(n_869) );
INVx2_ASAP7_75t_L g574 ( .A(n_575), .Y(n_574) );
INVx1_ASAP7_75t_L g595 ( .A(n_575), .Y(n_595) );
BUFx2_ASAP7_75t_L g886 ( .A(n_576), .Y(n_886) );
NAND4xp25_ASAP7_75t_L g577 ( .A(n_578), .B(n_581), .C(n_584), .D(n_586), .Y(n_577) );
INVx2_ASAP7_75t_L g892 ( .A(n_579), .Y(n_892) );
NOR2xp33_ASAP7_75t_L g588 ( .A(n_589), .B(n_590), .Y(n_588) );
NOR2xp33_ASAP7_75t_L g600 ( .A(n_590), .B(n_601), .Y(n_600) );
INVx4_ASAP7_75t_L g934 ( .A(n_590), .Y(n_934) );
INVx2_ASAP7_75t_L g610 ( .A(n_591), .Y(n_610) );
AND3x1_ASAP7_75t_L g592 ( .A(n_593), .B(n_598), .C(n_605), .Y(n_592) );
AND2x2_ASAP7_75t_L g593 ( .A(n_594), .B(n_596), .Y(n_593) );
AND2x2_ASAP7_75t_L g598 ( .A(n_599), .B(n_602), .Y(n_598) );
AND2x2_ASAP7_75t_L g602 ( .A(n_603), .B(n_604), .Y(n_602) );
AND2x2_ASAP7_75t_L g605 ( .A(n_606), .B(n_608), .Y(n_605) );
INVx1_ASAP7_75t_L g611 ( .A(n_612), .Y(n_611) );
HB1xp67_ASAP7_75t_L g612 ( .A(n_613), .Y(n_612) );
INVx1_ASAP7_75t_L g633 ( .A(n_613), .Y(n_633) );
INVx1_ASAP7_75t_L g613 ( .A(n_614), .Y(n_613) );
NAND4xp75_ASAP7_75t_L g615 ( .A(n_616), .B(n_620), .C(n_624), .D(n_627), .Y(n_615) );
AND2x2_ASAP7_75t_L g616 ( .A(n_617), .B(n_618), .Y(n_616) );
AND2x2_ASAP7_75t_L g620 ( .A(n_621), .B(n_623), .Y(n_620) );
BUFx3_ASAP7_75t_L g868 ( .A(n_622), .Y(n_868) );
AND2x2_ASAP7_75t_L g624 ( .A(n_625), .B(n_626), .Y(n_624) );
NOR2xp33_ASAP7_75t_L g629 ( .A(n_630), .B(n_631), .Y(n_629) );
INVxp67_ASAP7_75t_L g632 ( .A(n_633), .Y(n_632) );
BUFx10_ASAP7_75t_L g636 ( .A(n_637), .Y(n_636) );
HB1xp67_ASAP7_75t_L g637 ( .A(n_638), .Y(n_637) );
NAND3xp33_ASAP7_75t_L g638 ( .A(n_639), .B(n_642), .C(n_643), .Y(n_638) );
AND2x2_ASAP7_75t_L g901 ( .A(n_639), .B(n_902), .Y(n_901) );
AND2x2_ASAP7_75t_L g947 ( .A(n_639), .B(n_948), .Y(n_947) );
INVx1_ASAP7_75t_L g639 ( .A(n_640), .Y(n_639) );
OA21x2_ASAP7_75t_L g904 ( .A1(n_640), .A2(n_681), .B(n_905), .Y(n_904) );
HB1xp67_ASAP7_75t_L g640 ( .A(n_641), .Y(n_640) );
AND2x2_ASAP7_75t_L g658 ( .A(n_641), .B(n_659), .Y(n_658) );
AND3x4_ASAP7_75t_L g680 ( .A(n_641), .B(n_647), .C(n_681), .Y(n_680) );
NOR2xp33_ASAP7_75t_L g948 ( .A(n_642), .B(n_902), .Y(n_948) );
INVx1_ASAP7_75t_L g902 ( .A(n_643), .Y(n_902) );
OAI21xp5_ASAP7_75t_L g644 ( .A1(n_645), .A2(n_650), .B(n_863), .Y(n_644) );
BUFx2_ASAP7_75t_L g645 ( .A(n_646), .Y(n_645) );
OAI22xp5_ASAP7_75t_L g667 ( .A1(n_646), .A2(n_668), .B1(n_669), .B2(n_670), .Y(n_667) );
OAI221xp5_ASAP7_75t_L g765 ( .A1(n_646), .A2(n_668), .B1(n_766), .B2(n_767), .C(n_768), .Y(n_765) );
NAND2xp5_ASAP7_75t_L g646 ( .A(n_647), .B(n_649), .Y(n_646) );
AND2x4_ASAP7_75t_L g663 ( .A(n_647), .B(n_658), .Y(n_663) );
AND2x4_ASAP7_75t_L g664 ( .A(n_647), .B(n_649), .Y(n_664) );
AND2x4_ASAP7_75t_L g682 ( .A(n_647), .B(n_649), .Y(n_682) );
CKINVDCx5p33_ASAP7_75t_R g905 ( .A(n_647), .Y(n_905) );
AND2x2_ASAP7_75t_L g661 ( .A(n_649), .B(n_660), .Y(n_661) );
AND2x4_ASAP7_75t_L g676 ( .A(n_649), .B(n_660), .Y(n_676) );
AND2x2_ASAP7_75t_L g685 ( .A(n_649), .B(n_660), .Y(n_685) );
AOI211x1_ASAP7_75t_L g650 ( .A1(n_651), .A2(n_763), .B(n_769), .C(n_844), .Y(n_650) );
NAND5xp2_ASAP7_75t_L g651 ( .A(n_652), .B(n_721), .C(n_739), .D(n_749), .E(n_754), .Y(n_651) );
AOI332xp33_ASAP7_75t_L g652 ( .A1(n_653), .A2(n_686), .A3(n_696), .B1(n_697), .B2(n_701), .B3(n_710), .C1(n_711), .C2(n_715), .Y(n_652) );
NOR2xp33_ASAP7_75t_L g653 ( .A(n_654), .B(n_665), .Y(n_653) );
INVx2_ASAP7_75t_L g709 ( .A(n_654), .Y(n_709) );
BUFx3_ASAP7_75t_L g782 ( .A(n_654), .Y(n_782) );
NOR2xp33_ASAP7_75t_L g789 ( .A(n_654), .B(n_705), .Y(n_789) );
INVx1_ASAP7_75t_L g654 ( .A(n_655), .Y(n_654) );
INVx1_ASAP7_75t_L g719 ( .A(n_655), .Y(n_719) );
OR2x2_ASAP7_75t_L g816 ( .A(n_655), .B(n_678), .Y(n_816) );
NAND2xp5_ASAP7_75t_L g655 ( .A(n_656), .B(n_662), .Y(n_655) );
AND2x2_ASAP7_75t_L g657 ( .A(n_658), .B(n_660), .Y(n_657) );
AND2x4_ASAP7_75t_L g673 ( .A(n_658), .B(n_660), .Y(n_673) );
AND2x2_ASAP7_75t_L g684 ( .A(n_658), .B(n_660), .Y(n_684) );
INVx3_ASAP7_75t_L g668 ( .A(n_663), .Y(n_668) );
INVx1_ASAP7_75t_L g779 ( .A(n_665), .Y(n_779) );
NOR2xp33_ASAP7_75t_L g828 ( .A(n_665), .B(n_829), .Y(n_828) );
OR2x2_ASAP7_75t_L g665 ( .A(n_666), .B(n_678), .Y(n_665) );
INVx1_ASAP7_75t_L g704 ( .A(n_666), .Y(n_704) );
INVx2_ASAP7_75t_L g742 ( .A(n_666), .Y(n_742) );
AND2x2_ASAP7_75t_L g750 ( .A(n_666), .B(n_751), .Y(n_750) );
AND2x2_ASAP7_75t_L g758 ( .A(n_666), .B(n_678), .Y(n_758) );
AND2x2_ASAP7_75t_L g761 ( .A(n_666), .B(n_705), .Y(n_761) );
AND2x2_ASAP7_75t_L g811 ( .A(n_666), .B(n_706), .Y(n_811) );
OR2x2_ASAP7_75t_L g666 ( .A(n_667), .B(n_671), .Y(n_666) );
OAI22xp5_ASAP7_75t_L g671 ( .A1(n_672), .A2(n_674), .B1(n_675), .B2(n_677), .Y(n_671) );
INVx3_ASAP7_75t_L g672 ( .A(n_673), .Y(n_672) );
INVx2_ASAP7_75t_L g675 ( .A(n_676), .Y(n_675) );
HB1xp67_ASAP7_75t_L g710 ( .A(n_678), .Y(n_710) );
INVx2_ASAP7_75t_L g729 ( .A(n_678), .Y(n_729) );
OR2x2_ASAP7_75t_L g738 ( .A(n_678), .B(n_719), .Y(n_738) );
AND2x2_ASAP7_75t_L g751 ( .A(n_678), .B(n_719), .Y(n_751) );
AND2x2_ASAP7_75t_L g771 ( .A(n_678), .B(n_718), .Y(n_771) );
OR2x2_ASAP7_75t_L g800 ( .A(n_678), .B(n_742), .Y(n_800) );
AND2x2_ASAP7_75t_L g834 ( .A(n_678), .B(n_742), .Y(n_834) );
AND2x2_ASAP7_75t_L g678 ( .A(n_679), .B(n_683), .Y(n_678) );
INVxp67_ASAP7_75t_SL g686 ( .A(n_687), .Y(n_686) );
NAND2xp5_ASAP7_75t_L g687 ( .A(n_688), .B(n_695), .Y(n_687) );
INVx1_ASAP7_75t_L g714 ( .A(n_688), .Y(n_714) );
OR2x2_ASAP7_75t_L g748 ( .A(n_688), .B(n_698), .Y(n_748) );
OAI32xp33_ASAP7_75t_L g853 ( .A1(n_688), .A2(n_753), .A3(n_770), .B1(n_829), .B2(n_849), .Y(n_853) );
NOR2xp33_ASAP7_75t_L g862 ( .A(n_688), .B(n_746), .Y(n_862) );
OR2x2_ASAP7_75t_L g688 ( .A(n_689), .B(n_692), .Y(n_688) );
AND2x2_ASAP7_75t_L g696 ( .A(n_689), .B(n_692), .Y(n_696) );
INVx1_ASAP7_75t_L g726 ( .A(n_689), .Y(n_726) );
NAND2xp5_ASAP7_75t_L g737 ( .A(n_689), .B(n_697), .Y(n_737) );
AND2x2_ASAP7_75t_L g689 ( .A(n_690), .B(n_691), .Y(n_689) );
OR2x2_ASAP7_75t_L g725 ( .A(n_692), .B(n_726), .Y(n_725) );
INVx1_ASAP7_75t_L g744 ( .A(n_692), .Y(n_744) );
AND2x2_ASAP7_75t_L g762 ( .A(n_692), .B(n_712), .Y(n_762) );
AND2x2_ASAP7_75t_L g777 ( .A(n_692), .B(n_726), .Y(n_777) );
NAND2xp5_ASAP7_75t_L g788 ( .A(n_692), .B(n_697), .Y(n_788) );
AOI211xp5_ASAP7_75t_SL g856 ( .A1(n_692), .A2(n_857), .B(n_858), .C(n_859), .Y(n_856) );
AND2x2_ASAP7_75t_L g692 ( .A(n_693), .B(n_694), .Y(n_692) );
INVx1_ASAP7_75t_L g695 ( .A(n_696), .Y(n_695) );
AND2x2_ASAP7_75t_L g732 ( .A(n_696), .B(n_712), .Y(n_732) );
NAND2xp5_ASAP7_75t_L g796 ( .A(n_696), .B(n_797), .Y(n_796) );
AND2x2_ASAP7_75t_L g822 ( .A(n_696), .B(n_697), .Y(n_822) );
NOR2x1_ASAP7_75t_R g722 ( .A(n_697), .B(n_723), .Y(n_722) );
AND2x2_ASAP7_75t_L g743 ( .A(n_697), .B(n_744), .Y(n_743) );
AND2x2_ASAP7_75t_L g785 ( .A(n_697), .B(n_777), .Y(n_785) );
INVx1_ASAP7_75t_L g697 ( .A(n_698), .Y(n_697) );
INVx1_ASAP7_75t_SL g713 ( .A(n_698), .Y(n_713) );
OR2x2_ASAP7_75t_L g753 ( .A(n_698), .B(n_725), .Y(n_753) );
NAND2xp5_ASAP7_75t_L g794 ( .A(n_698), .B(n_724), .Y(n_794) );
AND2x2_ASAP7_75t_L g818 ( .A(n_698), .B(n_744), .Y(n_818) );
AND2x2_ASAP7_75t_L g698 ( .A(n_699), .B(n_700), .Y(n_698) );
INVx1_ASAP7_75t_L g701 ( .A(n_702), .Y(n_701) );
NAND2xp5_ASAP7_75t_L g702 ( .A(n_703), .B(n_709), .Y(n_702) );
AOI221xp5_ASAP7_75t_L g772 ( .A1(n_703), .A2(n_711), .B1(n_740), .B2(n_747), .C(n_773), .Y(n_772) );
AND2x2_ASAP7_75t_L g703 ( .A(n_704), .B(n_705), .Y(n_703) );
INVx2_ASAP7_75t_L g720 ( .A(n_704), .Y(n_720) );
NAND2xp5_ASAP7_75t_L g842 ( .A(n_704), .B(n_843), .Y(n_842) );
NAND2xp5_ASAP7_75t_SL g723 ( .A(n_705), .B(n_724), .Y(n_723) );
BUFx6f_ASAP7_75t_L g735 ( .A(n_705), .Y(n_735) );
INVx2_ASAP7_75t_L g746 ( .A(n_705), .Y(n_746) );
INVx2_ASAP7_75t_L g757 ( .A(n_705), .Y(n_757) );
NAND2xp5_ASAP7_75t_L g806 ( .A(n_705), .B(n_743), .Y(n_806) );
AND2x2_ASAP7_75t_L g817 ( .A(n_705), .B(n_818), .Y(n_817) );
INVx1_ASAP7_75t_L g829 ( .A(n_705), .Y(n_829) );
NAND2xp5_ASAP7_75t_SL g860 ( .A(n_705), .B(n_736), .Y(n_860) );
INVx4_ASAP7_75t_L g705 ( .A(n_706), .Y(n_705) );
NAND2xp5_ASAP7_75t_L g741 ( .A(n_706), .B(n_742), .Y(n_741) );
OR2x2_ASAP7_75t_L g798 ( .A(n_706), .B(n_712), .Y(n_798) );
AND2x2_ASAP7_75t_L g706 ( .A(n_707), .B(n_708), .Y(n_706) );
A2O1A1Ixp33_ASAP7_75t_L g739 ( .A1(n_709), .A2(n_740), .B(n_743), .C(n_745), .Y(n_739) );
NAND2xp5_ASAP7_75t_L g760 ( .A(n_709), .B(n_761), .Y(n_760) );
INVx1_ASAP7_75t_L g792 ( .A(n_709), .Y(n_792) );
NOR2xp33_ASAP7_75t_L g855 ( .A(n_709), .B(n_845), .Y(n_855) );
OAI221xp5_ASAP7_75t_L g859 ( .A1(n_710), .A2(n_725), .B1(n_800), .B2(n_860), .C(n_861), .Y(n_859) );
OAI21xp33_ASAP7_75t_L g786 ( .A1(n_711), .A2(n_787), .B(n_789), .Y(n_786) );
AND2x2_ASAP7_75t_L g843 ( .A(n_711), .B(n_746), .Y(n_843) );
A2O1A1O1Ixp25_ASAP7_75t_L g846 ( .A1(n_711), .A2(n_785), .B(n_834), .C(n_847), .D(n_848), .Y(n_846) );
INVx2_ASAP7_75t_SL g852 ( .A(n_711), .Y(n_852) );
AND2x4_ASAP7_75t_L g711 ( .A(n_712), .B(n_714), .Y(n_711) );
AND2x2_ASAP7_75t_L g776 ( .A(n_712), .B(n_777), .Y(n_776) );
INVx1_ASAP7_75t_L g712 ( .A(n_713), .Y(n_712) );
AOI221xp5_ASAP7_75t_L g804 ( .A1(n_715), .A2(n_758), .B1(n_805), .B2(n_807), .C(n_809), .Y(n_804) );
INVx1_ASAP7_75t_L g715 ( .A(n_716), .Y(n_715) );
NAND2xp5_ASAP7_75t_L g716 ( .A(n_717), .B(n_720), .Y(n_716) );
INVx1_ASAP7_75t_SL g847 ( .A(n_717), .Y(n_847) );
INVx1_ASAP7_75t_L g717 ( .A(n_718), .Y(n_717) );
INVx1_ASAP7_75t_L g718 ( .A(n_719), .Y(n_718) );
NAND2xp5_ASAP7_75t_L g823 ( .A(n_720), .B(n_771), .Y(n_823) );
NOR2xp33_ASAP7_75t_L g858 ( .A(n_720), .B(n_838), .Y(n_858) );
AOI21xp5_ASAP7_75t_L g721 ( .A1(n_722), .A2(n_727), .B(n_730), .Y(n_721) );
NAND2xp5_ASAP7_75t_L g808 ( .A(n_724), .B(n_797), .Y(n_808) );
INVx3_ASAP7_75t_SL g724 ( .A(n_725), .Y(n_724) );
NAND2xp5_ASAP7_75t_L g810 ( .A(n_726), .B(n_811), .Y(n_810) );
AOI221xp5_ASAP7_75t_L g861 ( .A1(n_726), .A2(n_747), .B1(n_761), .B2(n_774), .C(n_862), .Y(n_861) );
CKINVDCx14_ASAP7_75t_R g727 ( .A(n_728), .Y(n_727) );
CKINVDCx14_ASAP7_75t_R g728 ( .A(n_729), .Y(n_728) );
AND2x2_ASAP7_75t_L g826 ( .A(n_729), .B(n_811), .Y(n_826) );
AOI21xp33_ASAP7_75t_SL g730 ( .A1(n_731), .A2(n_733), .B(n_738), .Y(n_730) );
INVx1_ASAP7_75t_L g731 ( .A(n_732), .Y(n_731) );
NOR2xp33_ASAP7_75t_L g824 ( .A(n_732), .B(n_747), .Y(n_824) );
NAND2xp5_ASAP7_75t_L g838 ( .A(n_732), .B(n_839), .Y(n_838) );
NAND2xp5_ASAP7_75t_L g733 ( .A(n_734), .B(n_736), .Y(n_733) );
AND2x2_ASAP7_75t_L g821 ( .A(n_734), .B(n_822), .Y(n_821) );
NAND2xp5_ASAP7_75t_L g833 ( .A(n_734), .B(n_834), .Y(n_833) );
INVx2_ASAP7_75t_L g734 ( .A(n_735), .Y(n_734) );
NAND2xp5_ASAP7_75t_L g836 ( .A(n_735), .B(n_744), .Y(n_836) );
INVx1_ASAP7_75t_L g736 ( .A(n_737), .Y(n_736) );
A2O1A1Ixp33_ASAP7_75t_L g848 ( .A1(n_737), .A2(n_823), .B(n_849), .C(n_850), .Y(n_848) );
INVx1_ASAP7_75t_L g813 ( .A(n_738), .Y(n_813) );
NOR2xp33_ASAP7_75t_L g837 ( .A(n_738), .B(n_838), .Y(n_837) );
INVx1_ASAP7_75t_L g740 ( .A(n_741), .Y(n_740) );
INVx2_ASAP7_75t_L g774 ( .A(n_742), .Y(n_774) );
AND2x2_ASAP7_75t_L g745 ( .A(n_746), .B(n_747), .Y(n_745) );
NAND2xp5_ASAP7_75t_L g784 ( .A(n_746), .B(n_785), .Y(n_784) );
NOR2xp33_ASAP7_75t_L g803 ( .A(n_746), .B(n_748), .Y(n_803) );
INVx1_ASAP7_75t_L g839 ( .A(n_746), .Y(n_839) );
INVx1_ASAP7_75t_L g747 ( .A(n_748), .Y(n_747) );
NAND2xp5_ASAP7_75t_L g749 ( .A(n_750), .B(n_752), .Y(n_749) );
OAI21xp5_ASAP7_75t_L g801 ( .A1(n_751), .A2(n_802), .B(n_803), .Y(n_801) );
INVx1_ASAP7_75t_L g841 ( .A(n_751), .Y(n_841) );
INVx1_ASAP7_75t_L g752 ( .A(n_753), .Y(n_752) );
OAI21xp33_ASAP7_75t_L g754 ( .A1(n_755), .A2(n_759), .B(n_762), .Y(n_754) );
INVx1_ASAP7_75t_L g755 ( .A(n_756), .Y(n_755) );
NAND2xp5_ASAP7_75t_L g756 ( .A(n_757), .B(n_758), .Y(n_756) );
NAND2xp67_ASAP7_75t_L g775 ( .A(n_757), .B(n_776), .Y(n_775) );
INVx1_ASAP7_75t_L g835 ( .A(n_758), .Y(n_835) );
INVxp67_ASAP7_75t_SL g759 ( .A(n_760), .Y(n_759) );
INVx1_ASAP7_75t_L g849 ( .A(n_761), .Y(n_849) );
NAND2xp5_ASAP7_75t_L g827 ( .A(n_762), .B(n_828), .Y(n_827) );
INVx1_ASAP7_75t_L g832 ( .A(n_762), .Y(n_832) );
INVx2_ASAP7_75t_L g763 ( .A(n_764), .Y(n_763) );
AOI211xp5_ASAP7_75t_SL g830 ( .A1(n_764), .A2(n_831), .B(n_837), .C(n_840), .Y(n_830) );
HB1xp67_ASAP7_75t_L g764 ( .A(n_765), .Y(n_764) );
NAND2xp5_ASAP7_75t_L g812 ( .A(n_765), .B(n_813), .Y(n_812) );
INVx2_ASAP7_75t_L g845 ( .A(n_765), .Y(n_845) );
OAI211xp5_ASAP7_75t_L g769 ( .A1(n_770), .A2(n_772), .B(n_778), .C(n_830), .Y(n_769) );
INVx1_ASAP7_75t_L g770 ( .A(n_771), .Y(n_770) );
NOR2xp67_ASAP7_75t_SL g773 ( .A(n_774), .B(n_775), .Y(n_773) );
NOR2xp33_ASAP7_75t_L g851 ( .A(n_774), .B(n_852), .Y(n_851) );
INVx1_ASAP7_75t_L g783 ( .A(n_776), .Y(n_783) );
AOI211xp5_ASAP7_75t_L g778 ( .A1(n_779), .A2(n_780), .B(n_790), .C(n_819), .Y(n_778) );
OAI211xp5_ASAP7_75t_SL g780 ( .A1(n_781), .A2(n_783), .B(n_784), .C(n_786), .Y(n_780) );
INVx2_ASAP7_75t_L g781 ( .A(n_782), .Y(n_781) );
INVx1_ASAP7_75t_L g802 ( .A(n_784), .Y(n_802) );
INVx1_ASAP7_75t_L g787 ( .A(n_788), .Y(n_787) );
NAND3xp33_ASAP7_75t_SL g790 ( .A(n_791), .B(n_801), .C(n_804), .Y(n_790) );
A2O1A1Ixp33_ASAP7_75t_SL g791 ( .A1(n_792), .A2(n_793), .B(n_795), .C(n_799), .Y(n_791) );
INVx1_ASAP7_75t_L g793 ( .A(n_794), .Y(n_793) );
INVx1_ASAP7_75t_L g795 ( .A(n_796), .Y(n_795) );
INVx1_ASAP7_75t_L g797 ( .A(n_798), .Y(n_797) );
INVx1_ASAP7_75t_L g799 ( .A(n_800), .Y(n_799) );
INVx1_ASAP7_75t_L g805 ( .A(n_806), .Y(n_805) );
INVx1_ASAP7_75t_L g807 ( .A(n_808), .Y(n_807) );
OAI21xp33_ASAP7_75t_L g809 ( .A1(n_810), .A2(n_812), .B(n_814), .Y(n_809) );
NAND2xp5_ASAP7_75t_L g814 ( .A(n_815), .B(n_817), .Y(n_814) );
INVx1_ASAP7_75t_L g815 ( .A(n_816), .Y(n_815) );
OAI221xp5_ASAP7_75t_L g819 ( .A1(n_820), .A2(n_823), .B1(n_824), .B2(n_825), .C(n_827), .Y(n_819) );
INVx1_ASAP7_75t_L g820 ( .A(n_821), .Y(n_820) );
INVx1_ASAP7_75t_L g825 ( .A(n_826), .Y(n_825) );
OAI22xp5_ASAP7_75t_L g831 ( .A1(n_832), .A2(n_833), .B1(n_835), .B2(n_836), .Y(n_831) );
INVx1_ASAP7_75t_L g857 ( .A(n_833), .Y(n_857) );
NOR2xp33_ASAP7_75t_L g840 ( .A(n_841), .B(n_842), .Y(n_840) );
OAI22xp33_ASAP7_75t_L g844 ( .A1(n_845), .A2(n_846), .B1(n_854), .B2(n_856), .Y(n_844) );
NOR2xp33_ASAP7_75t_SL g850 ( .A(n_851), .B(n_853), .Y(n_850) );
INVx1_ASAP7_75t_L g854 ( .A(n_855), .Y(n_854) );
INVx1_ASAP7_75t_L g899 ( .A(n_865), .Y(n_899) );
OR4x1_ASAP7_75t_L g865 ( .A(n_866), .B(n_877), .C(n_884), .D(n_889), .Y(n_865) );
NAND2x1_ASAP7_75t_L g866 ( .A(n_867), .B(n_870), .Y(n_866) );
OA21x2_ASAP7_75t_L g870 ( .A1(n_871), .A2(n_872), .B(n_875), .Y(n_870) );
INVx1_ASAP7_75t_SL g872 ( .A(n_873), .Y(n_872) );
BUFx3_ASAP7_75t_L g873 ( .A(n_874), .Y(n_873) );
OAI22xp5_ASAP7_75t_L g877 ( .A1(n_878), .A2(n_879), .B1(n_881), .B2(n_882), .Y(n_877) );
INVx1_ASAP7_75t_L g879 ( .A(n_880), .Y(n_879) );
INVx1_ASAP7_75t_L g882 ( .A(n_883), .Y(n_882) );
NAND2xp5_ASAP7_75t_SL g884 ( .A(n_885), .B(n_887), .Y(n_884) );
NAND2xp5_ASAP7_75t_L g889 ( .A(n_890), .B(n_894), .Y(n_889) );
INVx2_ASAP7_75t_L g891 ( .A(n_892), .Y(n_891) );
INVx2_ASAP7_75t_L g895 ( .A(n_896), .Y(n_895) );
BUFx2_ASAP7_75t_SL g900 ( .A(n_901), .Y(n_900) );
HB1xp67_ASAP7_75t_L g903 ( .A(n_904), .Y(n_903) );
INVx1_ASAP7_75t_L g906 ( .A(n_907), .Y(n_906) );
INVx4_ASAP7_75t_L g907 ( .A(n_908), .Y(n_907) );
INVx1_ASAP7_75t_L g945 ( .A(n_909), .Y(n_945) );
NOR2x1_ASAP7_75t_L g909 ( .A(n_910), .B(n_924), .Y(n_909) );
NAND4xp25_ASAP7_75t_L g910 ( .A(n_911), .B(n_913), .C(n_916), .D(n_920), .Y(n_910) );
BUFx2_ASAP7_75t_SL g918 ( .A(n_919), .Y(n_918) );
BUFx3_ASAP7_75t_L g922 ( .A(n_923), .Y(n_922) );
NAND3xp33_ASAP7_75t_L g924 ( .A(n_925), .B(n_936), .C(n_940), .Y(n_924) );
INVx2_ASAP7_75t_SL g926 ( .A(n_927), .Y(n_926) );
INVx2_ASAP7_75t_L g927 ( .A(n_928), .Y(n_927) );
OAI22xp5_ASAP7_75t_L g929 ( .A1(n_930), .A2(n_932), .B1(n_933), .B2(n_935), .Y(n_929) );
INVx1_ASAP7_75t_L g930 ( .A(n_931), .Y(n_930) );
INVx1_ASAP7_75t_L g933 ( .A(n_934), .Y(n_933) );
HB1xp67_ASAP7_75t_L g937 ( .A(n_938), .Y(n_937) );
BUFx2_ASAP7_75t_L g941 ( .A(n_942), .Y(n_941) );
INVx2_ASAP7_75t_L g943 ( .A(n_944), .Y(n_943) );
HB1xp67_ASAP7_75t_L g946 ( .A(n_947), .Y(n_946) );
endmodule