module fake_aes_2071_n_583 (n_53, n_67, n_45, n_20, n_2, n_38, n_44, n_64, n_54, n_62, n_36, n_47, n_37, n_69, n_34, n_5, n_23, n_8, n_28, n_31, n_22, n_46, n_48, n_58, n_57, n_11, n_25, n_16, n_26, n_13, n_30, n_33, n_50, n_52, n_49, n_59, n_73, n_3, n_18, n_60, n_66, n_32, n_0, n_41, n_1, n_35, n_55, n_65, n_12, n_9, n_70, n_17, n_63, n_14, n_10, n_15, n_56, n_71, n_42, n_24, n_19, n_61, n_21, n_6, n_4, n_72, n_51, n_29, n_43, n_7, n_68, n_40, n_27, n_39, n_583);
input n_53;
input n_67;
input n_45;
input n_20;
input n_2;
input n_38;
input n_44;
input n_64;
input n_54;
input n_62;
input n_36;
input n_47;
input n_37;
input n_69;
input n_34;
input n_5;
input n_23;
input n_8;
input n_28;
input n_31;
input n_22;
input n_46;
input n_48;
input n_58;
input n_57;
input n_11;
input n_25;
input n_16;
input n_26;
input n_13;
input n_30;
input n_33;
input n_50;
input n_52;
input n_49;
input n_59;
input n_73;
input n_3;
input n_18;
input n_60;
input n_66;
input n_32;
input n_0;
input n_41;
input n_1;
input n_35;
input n_55;
input n_65;
input n_12;
input n_9;
input n_70;
input n_17;
input n_63;
input n_14;
input n_10;
input n_15;
input n_56;
input n_71;
input n_42;
input n_24;
input n_19;
input n_61;
input n_21;
input n_6;
input n_4;
input n_72;
input n_51;
input n_29;
input n_43;
input n_7;
input n_68;
input n_40;
input n_27;
input n_39;
output n_583;
wire n_117;
wire n_361;
wire n_513;
wire n_185;
wire n_407;
wire n_284;
wire n_278;
wire n_500;
wire n_114;
wire n_94;
wire n_125;
wire n_431;
wire n_484;
wire n_161;
wire n_496;
wire n_177;
wire n_130;
wire n_189;
wire n_311;
wire n_292;
wire n_309;
wire n_160;
wire n_154;
wire n_328;
wire n_468;
wire n_523;
wire n_229;
wire n_336;
wire n_464;
wire n_448;
wire n_348;
wire n_252;
wire n_152;
wire n_113;
wire n_353;
wire n_564;
wire n_528;
wire n_206;
wire n_383;
wire n_288;
wire n_532;
wire n_544;
wire n_400;
wire n_296;
wire n_157;
wire n_79;
wire n_202;
wire n_386;
wire n_432;
wire n_142;
wire n_232;
wire n_462;
wire n_316;
wire n_545;
wire n_211;
wire n_334;
wire n_389;
wire n_548;
wire n_436;
wire n_275;
wire n_463;
wire n_131;
wire n_112;
wire n_205;
wire n_330;
wire n_162;
wire n_387;
wire n_163;
wire n_434;
wire n_105;
wire n_227;
wire n_384;
wire n_476;
wire n_231;
wire n_452;
wire n_518;
wire n_547;
wire n_298;
wire n_411;
wire n_144;
wire n_183;
wire n_489;
wire n_199;
wire n_351;
wire n_83;
wire n_401;
wire n_100;
wire n_305;
wire n_461;
wire n_228;
wire n_360;
wire n_345;
wire n_236;
wire n_340;
wire n_481;
wire n_443;
wire n_150;
wire n_373;
wire n_576;
wire n_301;
wire n_222;
wire n_234;
wire n_465;
wire n_366;
wire n_286;
wire n_190;
wire n_246;
wire n_321;
wire n_572;
wire n_324;
wire n_392;
wire n_279;
wire n_303;
wire n_437;
wire n_512;
wire n_326;
wire n_289;
wire n_333;
wire n_249;
wire n_244;
wire n_540;
wire n_563;
wire n_119;
wire n_141;
wire n_517;
wire n_560;
wire n_479;
wire n_97;
wire n_167;
wire n_554;
wire n_447;
wire n_171;
wire n_567;
wire n_196;
wire n_580;
wire n_192;
wire n_502;
wire n_543;
wire n_312;
wire n_455;
wire n_529;
wire n_137;
wire n_511;
wire n_277;
wire n_467;
wire n_367;
wire n_85;
wire n_250;
wire n_314;
wire n_237;
wire n_181;
wire n_101;
wire n_255;
wire n_426;
wire n_91;
wire n_108;
wire n_116;
wire n_230;
wire n_209;
wire n_274;
wire n_282;
wire n_319;
wire n_499;
wire n_417;
wire n_241;
wire n_575;
wire n_95;
wire n_238;
wire n_318;
wire n_471;
wire n_293;
wire n_506;
wire n_533;
wire n_135;
wire n_393;
wire n_247;
wire n_490;
wire n_381;
wire n_550;
wire n_304;
wire n_399;
wire n_571;
wire n_294;
wire n_459;
wire n_313;
wire n_210;
wire n_184;
wire n_322;
wire n_310;
wire n_191;
wire n_307;
wire n_474;
wire n_354;
wire n_402;
wire n_413;
wire n_391;
wire n_427;
wire n_460;
wire n_478;
wire n_243;
wire n_415;
wire n_482;
wire n_394;
wire n_235;
wire n_442;
wire n_331;
wire n_485;
wire n_352;
wire n_268;
wire n_174;
wire n_501;
wire n_248;
wire n_299;
wire n_89;
wire n_338;
wire n_519;
wire n_256;
wire n_77;
wire n_551;
wire n_404;
wire n_369;
wire n_509;
wire n_172;
wire n_329;
wire n_251;
wire n_525;
wire n_218;
wire n_507;
wire n_271;
wire n_302;
wire n_466;
wire n_270;
wire n_362;
wire n_153;
wire n_259;
wire n_308;
wire n_546;
wire n_93;
wire n_412;
wire n_140;
wire n_207;
wire n_565;
wire n_224;
wire n_96;
wire n_219;
wire n_475;
wire n_578;
wire n_133;
wire n_149;
wire n_542;
wire n_81;
wire n_537;
wire n_214;
wire n_204;
wire n_430;
wire n_88;
wire n_450;
wire n_579;
wire n_107;
wire n_403;
wire n_557;
wire n_516;
wire n_254;
wire n_549;
wire n_262;
wire n_556;
wire n_239;
wire n_439;
wire n_87;
wire n_379;
wire n_527;
wire n_98;
wire n_526;
wire n_276;
wire n_320;
wire n_285;
wire n_195;
wire n_165;
wire n_446;
wire n_423;
wire n_342;
wire n_420;
wire n_370;
wire n_574;
wire n_217;
wire n_139;
wire n_388;
wire n_454;
wire n_193;
wire n_273;
wire n_505;
wire n_390;
wire n_120;
wire n_514;
wire n_486;
wire n_568;
wire n_245;
wire n_357;
wire n_90;
wire n_260;
wire n_78;
wire n_539;
wire n_197;
wire n_201;
wire n_317;
wire n_416;
wire n_374;
wire n_111;
wire n_536;
wire n_265;
wire n_264;
wire n_522;
wire n_208;
wire n_200;
wire n_573;
wire n_126;
wire n_178;
wire n_118;
wire n_365;
wire n_541;
wire n_179;
wire n_315;
wire n_363;
wire n_409;
wire n_86;
wire n_143;
wire n_295;
wire n_263;
wire n_166;
wire n_495;
wire n_186;
wire n_364;
wire n_428;
wire n_566;
wire n_75;
wire n_376;
wire n_552;
wire n_344;
wire n_136;
wire n_503;
wire n_283;
wire n_76;
wire n_520;
wire n_435;
wire n_216;
wire n_577;
wire n_147;
wire n_148;
wire n_212;
wire n_472;
wire n_92;
wire n_419;
wire n_396;
wire n_168;
wire n_477;
wire n_508;
wire n_570;
wire n_398;
wire n_445;
wire n_438;
wire n_134;
wire n_429;
wire n_488;
wire n_233;
wire n_82;
wire n_106;
wire n_440;
wire n_553;
wire n_173;
wire n_422;
wire n_327;
wire n_325;
wire n_349;
wire n_498;
wire n_225;
wire n_535;
wire n_530;
wire n_220;
wire n_358;
wire n_267;
wire n_221;
wire n_456;
wire n_203;
wire n_102;
wire n_449;
wire n_115;
wire n_80;
wire n_300;
wire n_158;
wire n_524;
wire n_121;
wire n_497;
wire n_339;
wire n_240;
wire n_378;
wire n_582;
wire n_359;
wire n_346;
wire n_103;
wire n_180;
wire n_441;
wire n_104;
wire n_74;
wire n_561;
wire n_335;
wire n_272;
wire n_534;
wire n_531;
wire n_146;
wire n_397;
wire n_306;
wire n_215;
wire n_242;
wire n_155;
wire n_198;
wire n_169;
wire n_424;
wire n_156;
wire n_124;
wire n_569;
wire n_297;
wire n_128;
wire n_129;
wire n_410;
wire n_188;
wire n_377;
wire n_510;
wire n_343;
wire n_127;
wire n_291;
wire n_170;
wire n_504;
wire n_458;
wire n_581;
wire n_418;
wire n_493;
wire n_555;
wire n_380;
wire n_356;
wire n_281;
wire n_341;
wire n_470;
wire n_122;
wire n_187;
wire n_375;
wire n_138;
wire n_487;
wire n_451;
wire n_371;
wire n_323;
wire n_473;
wire n_347;
wire n_558;
wire n_258;
wire n_253;
wire n_515;
wire n_84;
wire n_266;
wire n_213;
wire n_538;
wire n_182;
wire n_492;
wire n_368;
wire n_355;
wire n_226;
wire n_382;
wire n_159;
wire n_337;
wire n_444;
wire n_176;
wire n_521;
wire n_469;
wire n_123;
wire n_457;
wire n_223;
wire n_494;
wire n_559;
wire n_480;
wire n_372;
wire n_453;
wire n_194;
wire n_287;
wire n_110;
wire n_261;
wire n_425;
wire n_332;
wire n_414;
wire n_562;
wire n_350;
wire n_433;
wire n_164;
wire n_421;
wire n_175;
wire n_145;
wire n_483;
wire n_408;
wire n_290;
wire n_405;
wire n_280;
wire n_99;
wire n_109;
wire n_132;
wire n_395;
wire n_406;
wire n_491;
wire n_151;
wire n_385;
wire n_257;
wire n_269;
BUFx3_ASAP7_75t_L g74 ( .A(n_34), .Y(n_74) );
INVx1_ASAP7_75t_L g75 ( .A(n_23), .Y(n_75) );
BUFx2_ASAP7_75t_L g76 ( .A(n_66), .Y(n_76) );
INVx1_ASAP7_75t_L g77 ( .A(n_65), .Y(n_77) );
INVx1_ASAP7_75t_L g78 ( .A(n_21), .Y(n_78) );
INVx1_ASAP7_75t_L g79 ( .A(n_73), .Y(n_79) );
INVx1_ASAP7_75t_L g80 ( .A(n_67), .Y(n_80) );
INVxp33_ASAP7_75t_L g81 ( .A(n_52), .Y(n_81) );
CKINVDCx5p33_ASAP7_75t_R g82 ( .A(n_19), .Y(n_82) );
INVx1_ASAP7_75t_L g83 ( .A(n_21), .Y(n_83) );
INVx1_ASAP7_75t_L g84 ( .A(n_27), .Y(n_84) );
INVx1_ASAP7_75t_L g85 ( .A(n_15), .Y(n_85) );
INVx1_ASAP7_75t_L g86 ( .A(n_43), .Y(n_86) );
INVx1_ASAP7_75t_L g87 ( .A(n_53), .Y(n_87) );
HB1xp67_ASAP7_75t_L g88 ( .A(n_22), .Y(n_88) );
INVx1_ASAP7_75t_L g89 ( .A(n_22), .Y(n_89) );
CKINVDCx5p33_ASAP7_75t_R g90 ( .A(n_4), .Y(n_90) );
INVx1_ASAP7_75t_L g91 ( .A(n_36), .Y(n_91) );
CKINVDCx20_ASAP7_75t_R g92 ( .A(n_56), .Y(n_92) );
INVxp33_ASAP7_75t_SL g93 ( .A(n_59), .Y(n_93) );
INVx1_ASAP7_75t_L g94 ( .A(n_37), .Y(n_94) );
INVx1_ASAP7_75t_L g95 ( .A(n_8), .Y(n_95) );
INVxp67_ASAP7_75t_SL g96 ( .A(n_68), .Y(n_96) );
INVxp67_ASAP7_75t_SL g97 ( .A(n_5), .Y(n_97) );
INVx1_ASAP7_75t_L g98 ( .A(n_11), .Y(n_98) );
CKINVDCx5p33_ASAP7_75t_R g99 ( .A(n_24), .Y(n_99) );
INVx1_ASAP7_75t_L g100 ( .A(n_32), .Y(n_100) );
CKINVDCx20_ASAP7_75t_R g101 ( .A(n_46), .Y(n_101) );
INVxp67_ASAP7_75t_SL g102 ( .A(n_2), .Y(n_102) );
INVx1_ASAP7_75t_L g103 ( .A(n_29), .Y(n_103) );
INVx1_ASAP7_75t_L g104 ( .A(n_41), .Y(n_104) );
INVx1_ASAP7_75t_L g105 ( .A(n_60), .Y(n_105) );
INVx2_ASAP7_75t_L g106 ( .A(n_28), .Y(n_106) );
INVx1_ASAP7_75t_L g107 ( .A(n_38), .Y(n_107) );
INVx1_ASAP7_75t_L g108 ( .A(n_58), .Y(n_108) );
INVx1_ASAP7_75t_L g109 ( .A(n_17), .Y(n_109) );
INVx1_ASAP7_75t_L g110 ( .A(n_7), .Y(n_110) );
INVx1_ASAP7_75t_L g111 ( .A(n_15), .Y(n_111) );
CKINVDCx5p33_ASAP7_75t_R g112 ( .A(n_57), .Y(n_112) );
INVx1_ASAP7_75t_L g113 ( .A(n_42), .Y(n_113) );
INVx1_ASAP7_75t_L g114 ( .A(n_0), .Y(n_114) );
CKINVDCx5p33_ASAP7_75t_R g115 ( .A(n_63), .Y(n_115) );
INVxp33_ASAP7_75t_SL g116 ( .A(n_54), .Y(n_116) );
INVx2_ASAP7_75t_L g117 ( .A(n_69), .Y(n_117) );
INVx1_ASAP7_75t_L g118 ( .A(n_39), .Y(n_118) );
INVx1_ASAP7_75t_L g119 ( .A(n_0), .Y(n_119) );
INVx1_ASAP7_75t_L g120 ( .A(n_7), .Y(n_120) );
INVx1_ASAP7_75t_L g121 ( .A(n_77), .Y(n_121) );
INVx1_ASAP7_75t_L g122 ( .A(n_77), .Y(n_122) );
HB1xp67_ASAP7_75t_L g123 ( .A(n_88), .Y(n_123) );
INVx1_ASAP7_75t_L g124 ( .A(n_79), .Y(n_124) );
NOR2xp33_ASAP7_75t_L g125 ( .A(n_76), .B(n_1), .Y(n_125) );
CKINVDCx5p33_ASAP7_75t_R g126 ( .A(n_92), .Y(n_126) );
INVx1_ASAP7_75t_L g127 ( .A(n_79), .Y(n_127) );
NAND2xp5_ASAP7_75t_SL g128 ( .A(n_76), .B(n_1), .Y(n_128) );
INVx1_ASAP7_75t_L g129 ( .A(n_80), .Y(n_129) );
CKINVDCx5p33_ASAP7_75t_R g130 ( .A(n_101), .Y(n_130) );
INVx1_ASAP7_75t_L g131 ( .A(n_80), .Y(n_131) );
NAND2xp33_ASAP7_75t_R g132 ( .A(n_93), .B(n_26), .Y(n_132) );
INVx2_ASAP7_75t_L g133 ( .A(n_106), .Y(n_133) );
INVx1_ASAP7_75t_L g134 ( .A(n_84), .Y(n_134) );
INVx1_ASAP7_75t_L g135 ( .A(n_84), .Y(n_135) );
HB1xp67_ASAP7_75t_L g136 ( .A(n_82), .Y(n_136) );
INVx1_ASAP7_75t_L g137 ( .A(n_86), .Y(n_137) );
INVx5_ASAP7_75t_L g138 ( .A(n_74), .Y(n_138) );
INVx1_ASAP7_75t_L g139 ( .A(n_86), .Y(n_139) );
INVx1_ASAP7_75t_L g140 ( .A(n_87), .Y(n_140) );
NAND2xp5_ASAP7_75t_L g141 ( .A(n_106), .B(n_2), .Y(n_141) );
CKINVDCx20_ASAP7_75t_R g142 ( .A(n_90), .Y(n_142) );
CKINVDCx5p33_ASAP7_75t_R g143 ( .A(n_99), .Y(n_143) );
BUFx6f_ASAP7_75t_L g144 ( .A(n_74), .Y(n_144) );
CKINVDCx5p33_ASAP7_75t_R g145 ( .A(n_116), .Y(n_145) );
AND2x4_ASAP7_75t_L g146 ( .A(n_74), .B(n_3), .Y(n_146) );
INVx2_ASAP7_75t_L g147 ( .A(n_117), .Y(n_147) );
NAND2xp33_ASAP7_75t_R g148 ( .A(n_112), .B(n_30), .Y(n_148) );
CKINVDCx20_ASAP7_75t_R g149 ( .A(n_75), .Y(n_149) );
INVx3_ASAP7_75t_L g150 ( .A(n_87), .Y(n_150) );
BUFx3_ASAP7_75t_L g151 ( .A(n_117), .Y(n_151) );
NOR2xp33_ASAP7_75t_L g152 ( .A(n_91), .B(n_3), .Y(n_152) );
INVx1_ASAP7_75t_SL g153 ( .A(n_81), .Y(n_153) );
CKINVDCx20_ASAP7_75t_R g154 ( .A(n_75), .Y(n_154) );
INVx2_ASAP7_75t_L g155 ( .A(n_91), .Y(n_155) );
NAND2xp5_ASAP7_75t_L g156 ( .A(n_94), .B(n_4), .Y(n_156) );
CKINVDCx5p33_ASAP7_75t_R g157 ( .A(n_115), .Y(n_157) );
NOR2xp33_ASAP7_75t_R g158 ( .A(n_94), .B(n_100), .Y(n_158) );
OAI22xp5_ASAP7_75t_L g159 ( .A1(n_78), .A2(n_5), .B1(n_6), .B2(n_8), .Y(n_159) );
CKINVDCx20_ASAP7_75t_R g160 ( .A(n_78), .Y(n_160) );
INVx1_ASAP7_75t_L g161 ( .A(n_100), .Y(n_161) );
NAND2xp5_ASAP7_75t_L g162 ( .A(n_153), .B(n_105), .Y(n_162) );
INVx2_ASAP7_75t_L g163 ( .A(n_144), .Y(n_163) );
NAND2x1_ASAP7_75t_L g164 ( .A(n_146), .B(n_105), .Y(n_164) );
AND3x1_ASAP7_75t_L g165 ( .A(n_125), .B(n_120), .C(n_119), .Y(n_165) );
NAND2x1p5_ASAP7_75t_L g166 ( .A(n_146), .B(n_104), .Y(n_166) );
INVx2_ASAP7_75t_L g167 ( .A(n_144), .Y(n_167) );
NAND2x1p5_ASAP7_75t_L g168 ( .A(n_146), .B(n_104), .Y(n_168) );
INVx3_ASAP7_75t_L g169 ( .A(n_146), .Y(n_169) );
INVx1_ASAP7_75t_L g170 ( .A(n_150), .Y(n_170) );
INVx4_ASAP7_75t_L g171 ( .A(n_138), .Y(n_171) );
CKINVDCx5p33_ASAP7_75t_R g172 ( .A(n_142), .Y(n_172) );
OAI22xp5_ASAP7_75t_L g173 ( .A1(n_123), .A2(n_120), .B1(n_119), .B2(n_85), .Y(n_173) );
NAND2xp5_ASAP7_75t_L g174 ( .A(n_121), .B(n_118), .Y(n_174) );
NOR2xp33_ASAP7_75t_L g175 ( .A(n_145), .B(n_118), .Y(n_175) );
BUFx6f_ASAP7_75t_L g176 ( .A(n_144), .Y(n_176) );
OR2x2_ASAP7_75t_SL g177 ( .A(n_136), .B(n_114), .Y(n_177) );
INVx1_ASAP7_75t_L g178 ( .A(n_155), .Y(n_178) );
NOR2xp33_ASAP7_75t_L g179 ( .A(n_157), .B(n_113), .Y(n_179) );
AND2x2_ASAP7_75t_L g180 ( .A(n_121), .B(n_114), .Y(n_180) );
BUFx6f_ASAP7_75t_L g181 ( .A(n_144), .Y(n_181) );
OAI221xp5_ASAP7_75t_L g182 ( .A1(n_122), .A2(n_83), .B1(n_111), .B2(n_110), .C(n_109), .Y(n_182) );
NAND2x1p5_ASAP7_75t_L g183 ( .A(n_150), .B(n_113), .Y(n_183) );
INVx2_ASAP7_75t_L g184 ( .A(n_144), .Y(n_184) );
INVx3_ASAP7_75t_L g185 ( .A(n_151), .Y(n_185) );
INVx3_ASAP7_75t_L g186 ( .A(n_151), .Y(n_186) );
AO22x2_ASAP7_75t_L g187 ( .A1(n_159), .A2(n_103), .B1(n_107), .B2(n_108), .Y(n_187) );
AOI22xp5_ASAP7_75t_L g188 ( .A1(n_149), .A2(n_111), .B1(n_110), .B2(n_109), .Y(n_188) );
NOR2xp33_ASAP7_75t_L g189 ( .A(n_143), .B(n_108), .Y(n_189) );
AND2x2_ASAP7_75t_L g190 ( .A(n_122), .B(n_124), .Y(n_190) );
INVx1_ASAP7_75t_L g191 ( .A(n_155), .Y(n_191) );
BUFx6f_ASAP7_75t_L g192 ( .A(n_144), .Y(n_192) );
INVx1_ASAP7_75t_L g193 ( .A(n_150), .Y(n_193) );
NAND2xp5_ASAP7_75t_SL g194 ( .A(n_158), .B(n_124), .Y(n_194) );
NAND2xp5_ASAP7_75t_SL g195 ( .A(n_127), .B(n_107), .Y(n_195) );
AND2x2_ASAP7_75t_L g196 ( .A(n_127), .B(n_83), .Y(n_196) );
BUFx6f_ASAP7_75t_L g197 ( .A(n_138), .Y(n_197) );
INVx2_ASAP7_75t_L g198 ( .A(n_133), .Y(n_198) );
AO22x2_ASAP7_75t_L g199 ( .A1(n_129), .A2(n_103), .B1(n_85), .B2(n_98), .Y(n_199) );
HB1xp67_ASAP7_75t_L g200 ( .A(n_126), .Y(n_200) );
AO22x2_ASAP7_75t_L g201 ( .A1(n_129), .A2(n_98), .B1(n_95), .B2(n_89), .Y(n_201) );
BUFx3_ASAP7_75t_L g202 ( .A(n_138), .Y(n_202) );
INVx1_ASAP7_75t_SL g203 ( .A(n_154), .Y(n_203) );
NAND2xp5_ASAP7_75t_L g204 ( .A(n_131), .B(n_95), .Y(n_204) );
INVx1_ASAP7_75t_L g205 ( .A(n_155), .Y(n_205) );
INVx1_ASAP7_75t_L g206 ( .A(n_150), .Y(n_206) );
AND2x2_ASAP7_75t_L g207 ( .A(n_131), .B(n_89), .Y(n_207) );
CKINVDCx5p33_ASAP7_75t_R g208 ( .A(n_130), .Y(n_208) );
AOI22xp5_ASAP7_75t_L g209 ( .A1(n_160), .A2(n_102), .B1(n_97), .B2(n_96), .Y(n_209) );
NOR2xp33_ASAP7_75t_L g210 ( .A(n_134), .B(n_35), .Y(n_210) );
NAND2xp5_ASAP7_75t_L g211 ( .A(n_134), .B(n_6), .Y(n_211) );
BUFx2_ASAP7_75t_L g212 ( .A(n_135), .Y(n_212) );
INVx1_ASAP7_75t_L g213 ( .A(n_133), .Y(n_213) );
CKINVDCx5p33_ASAP7_75t_R g214 ( .A(n_132), .Y(n_214) );
INVx3_ASAP7_75t_L g215 ( .A(n_151), .Y(n_215) );
NAND3x1_ASAP7_75t_L g216 ( .A(n_156), .B(n_9), .C(n_10), .Y(n_216) );
NAND2xp5_ASAP7_75t_L g217 ( .A(n_135), .B(n_9), .Y(n_217) );
INVx2_ASAP7_75t_SL g218 ( .A(n_138), .Y(n_218) );
HB1xp67_ASAP7_75t_L g219 ( .A(n_137), .Y(n_219) );
NOR3xp33_ASAP7_75t_SL g220 ( .A(n_208), .B(n_128), .C(n_152), .Y(n_220) );
BUFx3_ASAP7_75t_L g221 ( .A(n_185), .Y(n_221) );
NAND2xp5_ASAP7_75t_L g222 ( .A(n_212), .B(n_161), .Y(n_222) );
INVx4_ASAP7_75t_L g223 ( .A(n_166), .Y(n_223) );
INVxp67_ASAP7_75t_SL g224 ( .A(n_166), .Y(n_224) );
BUFx6f_ASAP7_75t_L g225 ( .A(n_183), .Y(n_225) );
NOR3xp33_ASAP7_75t_SL g226 ( .A(n_208), .B(n_148), .C(n_141), .Y(n_226) );
AO22x1_ASAP7_75t_L g227 ( .A1(n_214), .A2(n_161), .B1(n_140), .B2(n_139), .Y(n_227) );
INVx2_ASAP7_75t_L g228 ( .A(n_178), .Y(n_228) );
AND2x2_ASAP7_75t_L g229 ( .A(n_212), .B(n_140), .Y(n_229) );
BUFx4f_ASAP7_75t_L g230 ( .A(n_166), .Y(n_230) );
INVx2_ASAP7_75t_L g231 ( .A(n_178), .Y(n_231) );
INVx1_ASAP7_75t_L g232 ( .A(n_191), .Y(n_232) );
BUFx6f_ASAP7_75t_L g233 ( .A(n_183), .Y(n_233) );
AND2x2_ASAP7_75t_L g234 ( .A(n_219), .B(n_139), .Y(n_234) );
INVx5_ASAP7_75t_L g235 ( .A(n_197), .Y(n_235) );
AND2x2_ASAP7_75t_L g236 ( .A(n_190), .B(n_137), .Y(n_236) );
OR2x6_ASAP7_75t_L g237 ( .A(n_168), .B(n_147), .Y(n_237) );
INVx2_ASAP7_75t_L g238 ( .A(n_191), .Y(n_238) );
INVx2_ASAP7_75t_L g239 ( .A(n_205), .Y(n_239) );
AND3x1_ASAP7_75t_L g240 ( .A(n_209), .B(n_147), .C(n_133), .Y(n_240) );
INVx1_ASAP7_75t_L g241 ( .A(n_205), .Y(n_241) );
NAND2xp5_ASAP7_75t_L g242 ( .A(n_190), .B(n_138), .Y(n_242) );
CKINVDCx20_ASAP7_75t_R g243 ( .A(n_172), .Y(n_243) );
NAND2xp5_ASAP7_75t_L g244 ( .A(n_162), .B(n_138), .Y(n_244) );
INVx1_ASAP7_75t_L g245 ( .A(n_206), .Y(n_245) );
OR2x2_ASAP7_75t_L g246 ( .A(n_203), .B(n_147), .Y(n_246) );
INVx2_ASAP7_75t_L g247 ( .A(n_206), .Y(n_247) );
NOR2xp33_ASAP7_75t_L g248 ( .A(n_175), .B(n_40), .Y(n_248) );
INVx3_ASAP7_75t_L g249 ( .A(n_185), .Y(n_249) );
BUFx3_ASAP7_75t_L g250 ( .A(n_185), .Y(n_250) );
INVx1_ASAP7_75t_L g251 ( .A(n_170), .Y(n_251) );
INVx2_ASAP7_75t_L g252 ( .A(n_193), .Y(n_252) );
NOR3xp33_ASAP7_75t_SL g253 ( .A(n_172), .B(n_10), .C(n_11), .Y(n_253) );
NOR2xp33_ASAP7_75t_SL g254 ( .A(n_168), .B(n_45), .Y(n_254) );
INVx3_ASAP7_75t_L g255 ( .A(n_186), .Y(n_255) );
AND2x4_ASAP7_75t_L g256 ( .A(n_180), .B(n_12), .Y(n_256) );
OR2x2_ASAP7_75t_SL g257 ( .A(n_200), .B(n_12), .Y(n_257) );
BUFx2_ASAP7_75t_L g258 ( .A(n_201), .Y(n_258) );
INVx1_ASAP7_75t_L g259 ( .A(n_213), .Y(n_259) );
INVx1_ASAP7_75t_L g260 ( .A(n_213), .Y(n_260) );
NOR3xp33_ASAP7_75t_SL g261 ( .A(n_182), .B(n_13), .C(n_14), .Y(n_261) );
NAND2xp5_ASAP7_75t_L g262 ( .A(n_180), .B(n_13), .Y(n_262) );
INVx1_ASAP7_75t_L g263 ( .A(n_169), .Y(n_263) );
OR2x4_ASAP7_75t_L g264 ( .A(n_189), .B(n_179), .Y(n_264) );
NAND2xp5_ASAP7_75t_L g265 ( .A(n_196), .B(n_14), .Y(n_265) );
INVx4_ASAP7_75t_L g266 ( .A(n_168), .Y(n_266) );
CKINVDCx11_ASAP7_75t_R g267 ( .A(n_173), .Y(n_267) );
AND2x6_ASAP7_75t_L g268 ( .A(n_169), .B(n_48), .Y(n_268) );
NAND2xp5_ASAP7_75t_L g269 ( .A(n_196), .B(n_16), .Y(n_269) );
INVx3_ASAP7_75t_L g270 ( .A(n_186), .Y(n_270) );
INVx2_ASAP7_75t_SL g271 ( .A(n_183), .Y(n_271) );
NAND2xp33_ASAP7_75t_SL g272 ( .A(n_214), .B(n_16), .Y(n_272) );
INVx2_ASAP7_75t_SL g273 ( .A(n_164), .Y(n_273) );
NAND2xp5_ASAP7_75t_L g274 ( .A(n_207), .B(n_17), .Y(n_274) );
INVx1_ASAP7_75t_L g275 ( .A(n_169), .Y(n_275) );
NAND2xp5_ASAP7_75t_L g276 ( .A(n_207), .B(n_18), .Y(n_276) );
NAND2xp5_ASAP7_75t_L g277 ( .A(n_186), .B(n_18), .Y(n_277) );
INVx5_ASAP7_75t_L g278 ( .A(n_197), .Y(n_278) );
BUFx6f_ASAP7_75t_L g279 ( .A(n_176), .Y(n_279) );
INVx2_ASAP7_75t_SL g280 ( .A(n_164), .Y(n_280) );
INVx2_ASAP7_75t_L g281 ( .A(n_247), .Y(n_281) );
AOI22xp5_ASAP7_75t_L g282 ( .A1(n_224), .A2(n_165), .B1(n_194), .B2(n_187), .Y(n_282) );
INVx1_ASAP7_75t_L g283 ( .A(n_236), .Y(n_283) );
OR2x6_ASAP7_75t_L g284 ( .A(n_223), .B(n_187), .Y(n_284) );
NAND2xp5_ASAP7_75t_L g285 ( .A(n_229), .B(n_215), .Y(n_285) );
OR2x6_ASAP7_75t_L g286 ( .A(n_223), .B(n_187), .Y(n_286) );
INVx1_ASAP7_75t_L g287 ( .A(n_236), .Y(n_287) );
BUFx3_ASAP7_75t_L g288 ( .A(n_225), .Y(n_288) );
CKINVDCx20_ASAP7_75t_R g289 ( .A(n_243), .Y(n_289) );
AOI22xp33_ASAP7_75t_L g290 ( .A1(n_258), .A2(n_199), .B1(n_201), .B2(n_187), .Y(n_290) );
NAND3xp33_ASAP7_75t_SL g291 ( .A(n_253), .B(n_188), .C(n_217), .Y(n_291) );
NAND2xp5_ASAP7_75t_L g292 ( .A(n_229), .B(n_215), .Y(n_292) );
BUFx3_ASAP7_75t_L g293 ( .A(n_225), .Y(n_293) );
BUFx6f_ASAP7_75t_L g294 ( .A(n_225), .Y(n_294) );
CKINVDCx5p33_ASAP7_75t_R g295 ( .A(n_267), .Y(n_295) );
BUFx2_ASAP7_75t_L g296 ( .A(n_258), .Y(n_296) );
INVx1_ASAP7_75t_L g297 ( .A(n_256), .Y(n_297) );
NOR2xp33_ASAP7_75t_L g298 ( .A(n_264), .B(n_177), .Y(n_298) );
BUFx4f_ASAP7_75t_SL g299 ( .A(n_223), .Y(n_299) );
OR2x6_ASAP7_75t_L g300 ( .A(n_266), .B(n_201), .Y(n_300) );
OR2x2_ASAP7_75t_L g301 ( .A(n_246), .B(n_177), .Y(n_301) );
OR2x2_ASAP7_75t_L g302 ( .A(n_246), .B(n_204), .Y(n_302) );
INVx1_ASAP7_75t_L g303 ( .A(n_256), .Y(n_303) );
INVx2_ASAP7_75t_SL g304 ( .A(n_230), .Y(n_304) );
NAND2xp5_ASAP7_75t_L g305 ( .A(n_234), .B(n_215), .Y(n_305) );
AND2x4_ASAP7_75t_L g306 ( .A(n_266), .B(n_195), .Y(n_306) );
NAND2xp5_ASAP7_75t_L g307 ( .A(n_234), .B(n_201), .Y(n_307) );
NOR2x1_ASAP7_75t_SL g308 ( .A(n_237), .B(n_174), .Y(n_308) );
INVx1_ASAP7_75t_L g309 ( .A(n_256), .Y(n_309) );
BUFx3_ASAP7_75t_L g310 ( .A(n_225), .Y(n_310) );
NOR2xp67_ASAP7_75t_L g311 ( .A(n_266), .B(n_211), .Y(n_311) );
AOI21xp5_ASAP7_75t_L g312 ( .A1(n_245), .A2(n_218), .B(n_199), .Y(n_312) );
OR2x6_ASAP7_75t_L g313 ( .A(n_237), .B(n_199), .Y(n_313) );
AOI21xp5_ASAP7_75t_L g314 ( .A1(n_245), .A2(n_218), .B(n_199), .Y(n_314) );
NOR2xp33_ASAP7_75t_L g315 ( .A(n_264), .B(n_210), .Y(n_315) );
AOI22xp33_ASAP7_75t_SL g316 ( .A1(n_230), .A2(n_216), .B1(n_198), .B2(n_171), .Y(n_316) );
OR2x6_ASAP7_75t_L g317 ( .A(n_237), .B(n_216), .Y(n_317) );
BUFx12f_ASAP7_75t_L g318 ( .A(n_257), .Y(n_318) );
INVx2_ASAP7_75t_L g319 ( .A(n_247), .Y(n_319) );
INVx2_ASAP7_75t_L g320 ( .A(n_228), .Y(n_320) );
AOI222xp33_ASAP7_75t_L g321 ( .A1(n_256), .A2(n_198), .B1(n_163), .B2(n_167), .C1(n_184), .C2(n_181), .Y(n_321) );
CKINVDCx5p33_ASAP7_75t_R g322 ( .A(n_226), .Y(n_322) );
OAI22xp33_ASAP7_75t_SL g323 ( .A1(n_230), .A2(n_19), .B1(n_20), .B2(n_23), .Y(n_323) );
BUFx2_ASAP7_75t_L g324 ( .A(n_237), .Y(n_324) );
OAI22xp5_ASAP7_75t_L g325 ( .A1(n_237), .A2(n_171), .B1(n_167), .B2(n_163), .Y(n_325) );
AOI221xp5_ASAP7_75t_L g326 ( .A1(n_240), .A2(n_171), .B1(n_184), .B2(n_192), .C(n_181), .Y(n_326) );
INVx3_ASAP7_75t_L g327 ( .A(n_225), .Y(n_327) );
NAND2xp5_ASAP7_75t_L g328 ( .A(n_222), .B(n_202), .Y(n_328) );
NAND2xp5_ASAP7_75t_L g329 ( .A(n_302), .B(n_227), .Y(n_329) );
NAND2xp5_ASAP7_75t_SL g330 ( .A(n_294), .B(n_233), .Y(n_330) );
INVx1_ASAP7_75t_L g331 ( .A(n_320), .Y(n_331) );
A2O1A1Ixp33_ASAP7_75t_L g332 ( .A1(n_315), .A2(n_312), .B(n_314), .C(n_290), .Y(n_332) );
CKINVDCx6p67_ASAP7_75t_R g333 ( .A(n_313), .Y(n_333) );
CKINVDCx5p33_ASAP7_75t_R g334 ( .A(n_289), .Y(n_334) );
BUFx3_ASAP7_75t_L g335 ( .A(n_299), .Y(n_335) );
INVx4_ASAP7_75t_L g336 ( .A(n_313), .Y(n_336) );
OAI21xp33_ASAP7_75t_SL g337 ( .A1(n_313), .A2(n_271), .B(n_241), .Y(n_337) );
OR2x2_ASAP7_75t_L g338 ( .A(n_300), .B(n_227), .Y(n_338) );
INVx2_ASAP7_75t_L g339 ( .A(n_320), .Y(n_339) );
AOI21xp5_ASAP7_75t_L g340 ( .A1(n_315), .A2(n_242), .B(n_244), .Y(n_340) );
INVx1_ASAP7_75t_L g341 ( .A(n_281), .Y(n_341) );
BUFx6f_ASAP7_75t_L g342 ( .A(n_294), .Y(n_342) );
BUFx3_ASAP7_75t_L g343 ( .A(n_299), .Y(n_343) );
OR2x2_ASAP7_75t_L g344 ( .A(n_300), .B(n_262), .Y(n_344) );
NAND2x1_ASAP7_75t_L g345 ( .A(n_294), .B(n_233), .Y(n_345) );
OAI22xp5_ASAP7_75t_L g346 ( .A1(n_300), .A2(n_271), .B1(n_233), .B2(n_241), .Y(n_346) );
AND2x2_ASAP7_75t_L g347 ( .A(n_283), .B(n_228), .Y(n_347) );
INVx1_ASAP7_75t_L g348 ( .A(n_281), .Y(n_348) );
AOI22xp33_ASAP7_75t_SL g349 ( .A1(n_318), .A2(n_254), .B1(n_257), .B2(n_268), .Y(n_349) );
AND2x2_ASAP7_75t_L g350 ( .A(n_287), .B(n_231), .Y(n_350) );
INVx3_ASAP7_75t_L g351 ( .A(n_294), .Y(n_351) );
INVx2_ASAP7_75t_L g352 ( .A(n_319), .Y(n_352) );
AO21x2_ASAP7_75t_L g353 ( .A1(n_291), .A2(n_277), .B(n_261), .Y(n_353) );
OAI21x1_ASAP7_75t_L g354 ( .A1(n_327), .A2(n_274), .B(n_265), .Y(n_354) );
AO21x2_ASAP7_75t_L g355 ( .A1(n_297), .A2(n_276), .B(n_269), .Y(n_355) );
AOI22xp5_ASAP7_75t_L g356 ( .A1(n_290), .A2(n_240), .B1(n_272), .B2(n_254), .Y(n_356) );
HB1xp67_ASAP7_75t_L g357 ( .A(n_324), .Y(n_357) );
NAND2xp5_ASAP7_75t_L g358 ( .A(n_307), .B(n_259), .Y(n_358) );
AND2x2_ASAP7_75t_L g359 ( .A(n_347), .B(n_350), .Y(n_359) );
AOI22xp33_ASAP7_75t_L g360 ( .A1(n_349), .A2(n_318), .B1(n_284), .B2(n_286), .Y(n_360) );
BUFx2_ASAP7_75t_L g361 ( .A(n_337), .Y(n_361) );
AOI22xp33_ASAP7_75t_L g362 ( .A1(n_349), .A2(n_286), .B1(n_284), .B2(n_298), .Y(n_362) );
INVx1_ASAP7_75t_L g363 ( .A(n_331), .Y(n_363) );
OAI21x1_ASAP7_75t_L g364 ( .A1(n_354), .A2(n_327), .B(n_325), .Y(n_364) );
AOI22xp33_ASAP7_75t_L g365 ( .A1(n_353), .A2(n_286), .B1(n_284), .B2(n_298), .Y(n_365) );
OAI21x1_ASAP7_75t_L g366 ( .A1(n_354), .A2(n_319), .B(n_326), .Y(n_366) );
OAI22xp5_ASAP7_75t_L g367 ( .A1(n_333), .A2(n_338), .B1(n_356), .B2(n_336), .Y(n_367) );
OAI221xp5_ASAP7_75t_L g368 ( .A1(n_356), .A2(n_301), .B1(n_220), .B2(n_282), .C(n_316), .Y(n_368) );
AOI21xp5_ASAP7_75t_L g369 ( .A1(n_340), .A2(n_233), .B(n_303), .Y(n_369) );
INVx2_ASAP7_75t_L g370 ( .A(n_339), .Y(n_370) );
OAI22xp33_ASAP7_75t_L g371 ( .A1(n_333), .A2(n_317), .B1(n_295), .B2(n_296), .Y(n_371) );
OAI22xp5_ASAP7_75t_SL g372 ( .A1(n_334), .A2(n_295), .B1(n_317), .B2(n_264), .Y(n_372) );
AOI22xp33_ASAP7_75t_L g373 ( .A1(n_353), .A2(n_317), .B1(n_322), .B2(n_309), .Y(n_373) );
AOI221xp5_ASAP7_75t_L g374 ( .A1(n_329), .A2(n_305), .B1(n_292), .B2(n_285), .C(n_323), .Y(n_374) );
AND2x2_ASAP7_75t_L g375 ( .A(n_347), .B(n_308), .Y(n_375) );
NAND2x1_ASAP7_75t_L g376 ( .A(n_339), .B(n_268), .Y(n_376) );
AOI221xp5_ASAP7_75t_L g377 ( .A1(n_329), .A2(n_232), .B1(n_259), .B2(n_260), .C(n_263), .Y(n_377) );
OAI22xp33_ASAP7_75t_L g378 ( .A1(n_333), .A2(n_304), .B1(n_233), .B2(n_311), .Y(n_378) );
OAI22xp5_ASAP7_75t_L g379 ( .A1(n_338), .A2(n_260), .B1(n_232), .B2(n_231), .Y(n_379) );
OAI22xp5_ASAP7_75t_L g380 ( .A1(n_338), .A2(n_239), .B1(n_238), .B2(n_310), .Y(n_380) );
INVx4_ASAP7_75t_SL g381 ( .A(n_335), .Y(n_381) );
AO21x2_ASAP7_75t_L g382 ( .A1(n_332), .A2(n_248), .B(n_328), .Y(n_382) );
INVx1_ASAP7_75t_L g383 ( .A(n_331), .Y(n_383) );
INVx1_ASAP7_75t_L g384 ( .A(n_341), .Y(n_384) );
AOI22xp5_ASAP7_75t_L g385 ( .A1(n_368), .A2(n_337), .B1(n_353), .B2(n_336), .Y(n_385) );
OR2x2_ASAP7_75t_L g386 ( .A(n_359), .B(n_336), .Y(n_386) );
AND2x2_ASAP7_75t_L g387 ( .A(n_359), .B(n_341), .Y(n_387) );
OAI221xp5_ASAP7_75t_L g388 ( .A1(n_374), .A2(n_332), .B1(n_344), .B2(n_357), .C(n_340), .Y(n_388) );
NAND2xp5_ASAP7_75t_L g389 ( .A(n_363), .B(n_350), .Y(n_389) );
INVx1_ASAP7_75t_L g390 ( .A(n_363), .Y(n_390) );
INVx2_ASAP7_75t_L g391 ( .A(n_370), .Y(n_391) );
OAI22xp33_ASAP7_75t_L g392 ( .A1(n_379), .A2(n_336), .B1(n_346), .B2(n_335), .Y(n_392) );
INVx1_ASAP7_75t_L g393 ( .A(n_383), .Y(n_393) );
NAND2xp5_ASAP7_75t_L g394 ( .A(n_383), .B(n_350), .Y(n_394) );
AOI222xp33_ASAP7_75t_L g395 ( .A1(n_372), .A2(n_336), .B1(n_358), .B2(n_346), .C1(n_343), .C2(n_335), .Y(n_395) );
AND2x2_ASAP7_75t_L g396 ( .A(n_375), .B(n_348), .Y(n_396) );
AND2x2_ASAP7_75t_L g397 ( .A(n_375), .B(n_348), .Y(n_397) );
OAI21xp33_ASAP7_75t_L g398 ( .A1(n_360), .A2(n_339), .B(n_352), .Y(n_398) );
INVx1_ASAP7_75t_L g399 ( .A(n_384), .Y(n_399) );
BUFx2_ASAP7_75t_L g400 ( .A(n_361), .Y(n_400) );
OAI221xp5_ASAP7_75t_L g401 ( .A1(n_372), .A2(n_344), .B1(n_357), .B2(n_358), .C(n_343), .Y(n_401) );
INVx1_ASAP7_75t_L g402 ( .A(n_384), .Y(n_402) );
AND2x2_ASAP7_75t_L g403 ( .A(n_370), .B(n_352), .Y(n_403) );
AOI22xp33_ASAP7_75t_L g404 ( .A1(n_362), .A2(n_353), .B1(n_344), .B2(n_343), .Y(n_404) );
AOI22xp33_ASAP7_75t_L g405 ( .A1(n_367), .A2(n_353), .B1(n_268), .B2(n_355), .Y(n_405) );
AOI21xp5_ASAP7_75t_L g406 ( .A1(n_376), .A2(n_330), .B(n_345), .Y(n_406) );
HB1xp67_ASAP7_75t_L g407 ( .A(n_370), .Y(n_407) );
OAI211xp5_ASAP7_75t_SL g408 ( .A1(n_365), .A2(n_321), .B(n_330), .C(n_280), .Y(n_408) );
INVx1_ASAP7_75t_L g409 ( .A(n_366), .Y(n_409) );
HB1xp67_ASAP7_75t_L g410 ( .A(n_381), .Y(n_410) );
NOR4xp25_ASAP7_75t_SL g411 ( .A(n_381), .B(n_268), .C(n_345), .D(n_354), .Y(n_411) );
OAI22xp5_ASAP7_75t_L g412 ( .A1(n_379), .A2(n_293), .B1(n_310), .B2(n_288), .Y(n_412) );
AOI22xp33_ASAP7_75t_L g413 ( .A1(n_367), .A2(n_268), .B1(n_355), .B2(n_306), .Y(n_413) );
INVx3_ASAP7_75t_L g414 ( .A(n_376), .Y(n_414) );
AND2x4_ASAP7_75t_SL g415 ( .A(n_373), .B(n_351), .Y(n_415) );
INVx1_ASAP7_75t_L g416 ( .A(n_366), .Y(n_416) );
AND2x2_ASAP7_75t_L g417 ( .A(n_391), .B(n_382), .Y(n_417) );
AOI22xp33_ASAP7_75t_L g418 ( .A1(n_395), .A2(n_371), .B1(n_382), .B2(n_380), .Y(n_418) );
INVxp67_ASAP7_75t_SL g419 ( .A(n_407), .Y(n_419) );
OR2x2_ASAP7_75t_L g420 ( .A(n_390), .B(n_382), .Y(n_420) );
INVxp67_ASAP7_75t_SL g421 ( .A(n_391), .Y(n_421) );
NAND2xp5_ASAP7_75t_L g422 ( .A(n_393), .B(n_380), .Y(n_422) );
INVx1_ASAP7_75t_L g423 ( .A(n_393), .Y(n_423) );
AO31x2_ASAP7_75t_L g424 ( .A1(n_416), .A2(n_369), .A3(n_238), .B(n_239), .Y(n_424) );
AND2x2_ASAP7_75t_L g425 ( .A(n_391), .B(n_364), .Y(n_425) );
AND2x2_ASAP7_75t_L g426 ( .A(n_403), .B(n_364), .Y(n_426) );
AND2x2_ASAP7_75t_L g427 ( .A(n_403), .B(n_355), .Y(n_427) );
AND2x2_ASAP7_75t_L g428 ( .A(n_400), .B(n_355), .Y(n_428) );
AND2x2_ASAP7_75t_L g429 ( .A(n_400), .B(n_351), .Y(n_429) );
INVxp67_ASAP7_75t_L g430 ( .A(n_399), .Y(n_430) );
AND2x2_ASAP7_75t_L g431 ( .A(n_399), .B(n_351), .Y(n_431) );
AND2x2_ASAP7_75t_L g432 ( .A(n_402), .B(n_351), .Y(n_432) );
AND2x2_ASAP7_75t_SL g433 ( .A(n_413), .B(n_342), .Y(n_433) );
OAI221xp5_ASAP7_75t_SL g434 ( .A1(n_395), .A2(n_378), .B1(n_377), .B2(n_381), .C(n_280), .Y(n_434) );
NOR2xp33_ASAP7_75t_L g435 ( .A(n_401), .B(n_306), .Y(n_435) );
NOR2xp67_ASAP7_75t_SL g436 ( .A(n_410), .B(n_342), .Y(n_436) );
INVx1_ASAP7_75t_L g437 ( .A(n_402), .Y(n_437) );
AND2x2_ASAP7_75t_L g438 ( .A(n_396), .B(n_351), .Y(n_438) );
INVx2_ASAP7_75t_L g439 ( .A(n_409), .Y(n_439) );
INVx1_ASAP7_75t_L g440 ( .A(n_409), .Y(n_440) );
BUFx3_ASAP7_75t_L g441 ( .A(n_396), .Y(n_441) );
INVx2_ASAP7_75t_L g442 ( .A(n_414), .Y(n_442) );
NOR2xp33_ASAP7_75t_L g443 ( .A(n_386), .B(n_20), .Y(n_443) );
AND2x2_ASAP7_75t_L g444 ( .A(n_397), .B(n_342), .Y(n_444) );
INVx2_ASAP7_75t_L g445 ( .A(n_414), .Y(n_445) );
INVx3_ASAP7_75t_L g446 ( .A(n_414), .Y(n_446) );
NOR2xp33_ASAP7_75t_L g447 ( .A(n_386), .B(n_24), .Y(n_447) );
INVx2_ASAP7_75t_SL g448 ( .A(n_415), .Y(n_448) );
AOI221xp5_ASAP7_75t_L g449 ( .A1(n_388), .A2(n_263), .B1(n_275), .B2(n_251), .C(n_273), .Y(n_449) );
NOR2xp33_ASAP7_75t_L g450 ( .A(n_387), .B(n_273), .Y(n_450) );
NOR4xp75_ASAP7_75t_L g451 ( .A(n_398), .B(n_381), .C(n_268), .D(n_31), .Y(n_451) );
AND2x2_ASAP7_75t_L g452 ( .A(n_397), .B(n_342), .Y(n_452) );
OR2x2_ASAP7_75t_L g453 ( .A(n_404), .B(n_342), .Y(n_453) );
INVx2_ASAP7_75t_L g454 ( .A(n_414), .Y(n_454) );
INVx1_ASAP7_75t_SL g455 ( .A(n_415), .Y(n_455) );
INVx2_ASAP7_75t_L g456 ( .A(n_415), .Y(n_456) );
AOI211xp5_ASAP7_75t_SL g457 ( .A1(n_392), .A2(n_381), .B(n_268), .C(n_255), .Y(n_457) );
NAND2x1p5_ASAP7_75t_L g458 ( .A(n_385), .B(n_342), .Y(n_458) );
AND2x2_ASAP7_75t_L g459 ( .A(n_405), .B(n_342), .Y(n_459) );
OR2x2_ASAP7_75t_L g460 ( .A(n_385), .B(n_293), .Y(n_460) );
NAND4xp25_ASAP7_75t_L g461 ( .A(n_418), .B(n_398), .C(n_408), .D(n_389), .Y(n_461) );
AND2x2_ASAP7_75t_L g462 ( .A(n_441), .B(n_394), .Y(n_462) );
AND2x4_ASAP7_75t_L g463 ( .A(n_441), .B(n_406), .Y(n_463) );
OAI31xp33_ASAP7_75t_SL g464 ( .A1(n_443), .A2(n_412), .A3(n_411), .B(n_33), .Y(n_464) );
INVx1_ASAP7_75t_L g465 ( .A(n_423), .Y(n_465) );
INVx2_ASAP7_75t_L g466 ( .A(n_439), .Y(n_466) );
NAND2xp5_ASAP7_75t_L g467 ( .A(n_441), .B(n_288), .Y(n_467) );
AOI22xp33_ASAP7_75t_L g468 ( .A1(n_418), .A2(n_270), .B1(n_255), .B2(n_249), .Y(n_468) );
AND2x2_ASAP7_75t_L g469 ( .A(n_438), .B(n_25), .Y(n_469) );
INVx1_ASAP7_75t_SL g470 ( .A(n_444), .Y(n_470) );
BUFx8_ASAP7_75t_L g471 ( .A(n_438), .Y(n_471) );
INVx1_ASAP7_75t_L g472 ( .A(n_423), .Y(n_472) );
OR2x2_ASAP7_75t_L g473 ( .A(n_419), .B(n_270), .Y(n_473) );
NAND2xp5_ASAP7_75t_L g474 ( .A(n_437), .B(n_251), .Y(n_474) );
INVx1_ASAP7_75t_L g475 ( .A(n_437), .Y(n_475) );
OR2x2_ASAP7_75t_L g476 ( .A(n_419), .B(n_270), .Y(n_476) );
NAND2xp5_ASAP7_75t_L g477 ( .A(n_430), .B(n_275), .Y(n_477) );
NOR2xp33_ASAP7_75t_L g478 ( .A(n_443), .B(n_447), .Y(n_478) );
OR2x2_ASAP7_75t_L g479 ( .A(n_427), .B(n_255), .Y(n_479) );
INVx1_ASAP7_75t_L g480 ( .A(n_431), .Y(n_480) );
INVx1_ASAP7_75t_L g481 ( .A(n_431), .Y(n_481) );
OR2x2_ASAP7_75t_L g482 ( .A(n_427), .B(n_249), .Y(n_482) );
NAND2xp5_ASAP7_75t_L g483 ( .A(n_447), .B(n_252), .Y(n_483) );
AOI21xp33_ASAP7_75t_SL g484 ( .A1(n_434), .A2(n_44), .B(n_47), .Y(n_484) );
INVx2_ASAP7_75t_L g485 ( .A(n_439), .Y(n_485) );
HB1xp67_ASAP7_75t_L g486 ( .A(n_421), .Y(n_486) );
AND2x2_ASAP7_75t_L g487 ( .A(n_438), .B(n_49), .Y(n_487) );
NOR2xp33_ASAP7_75t_R g488 ( .A(n_433), .B(n_50), .Y(n_488) );
NOR2xp33_ASAP7_75t_L g489 ( .A(n_435), .B(n_434), .Y(n_489) );
OR2x2_ASAP7_75t_L g490 ( .A(n_421), .B(n_249), .Y(n_490) );
INVx2_ASAP7_75t_L g491 ( .A(n_440), .Y(n_491) );
AOI31xp67_ASAP7_75t_SL g492 ( .A1(n_457), .A2(n_51), .A3(n_55), .B(n_61), .Y(n_492) );
NOR2xp33_ASAP7_75t_R g493 ( .A(n_433), .B(n_62), .Y(n_493) );
OR2x2_ASAP7_75t_L g494 ( .A(n_444), .B(n_192), .Y(n_494) );
NAND2xp33_ASAP7_75t_SL g495 ( .A(n_448), .B(n_192), .Y(n_495) );
INVx1_ASAP7_75t_L g496 ( .A(n_432), .Y(n_496) );
INVx1_ASAP7_75t_L g497 ( .A(n_440), .Y(n_497) );
OR2x6_ASAP7_75t_L g498 ( .A(n_448), .B(n_192), .Y(n_498) );
NAND2xp5_ASAP7_75t_SL g499 ( .A(n_446), .B(n_278), .Y(n_499) );
NAND2xp5_ASAP7_75t_L g500 ( .A(n_428), .B(n_252), .Y(n_500) );
AND2x2_ASAP7_75t_L g501 ( .A(n_452), .B(n_64), .Y(n_501) );
AOI22xp33_ASAP7_75t_L g502 ( .A1(n_489), .A2(n_433), .B1(n_435), .B2(n_448), .Y(n_502) );
INVxp67_ASAP7_75t_L g503 ( .A(n_486), .Y(n_503) );
INVx1_ASAP7_75t_L g504 ( .A(n_465), .Y(n_504) );
INVx1_ASAP7_75t_L g505 ( .A(n_472), .Y(n_505) );
INVx1_ASAP7_75t_L g506 ( .A(n_475), .Y(n_506) );
NAND2xp5_ASAP7_75t_L g507 ( .A(n_462), .B(n_428), .Y(n_507) );
NAND2xp5_ASAP7_75t_L g508 ( .A(n_480), .B(n_422), .Y(n_508) );
O2A1O1Ixp33_ASAP7_75t_L g509 ( .A1(n_484), .A2(n_450), .B(n_449), .C(n_420), .Y(n_509) );
NAND2xp33_ASAP7_75t_SL g510 ( .A(n_488), .B(n_436), .Y(n_510) );
INVxp67_ASAP7_75t_L g511 ( .A(n_486), .Y(n_511) );
OAI22xp33_ASAP7_75t_L g512 ( .A1(n_461), .A2(n_478), .B1(n_455), .B2(n_498), .Y(n_512) );
NOR2xp33_ASAP7_75t_L g513 ( .A(n_478), .B(n_450), .Y(n_513) );
NAND2xp5_ASAP7_75t_L g514 ( .A(n_481), .B(n_417), .Y(n_514) );
OAI21xp33_ASAP7_75t_L g515 ( .A1(n_464), .A2(n_420), .B(n_458), .Y(n_515) );
AOI222xp33_ASAP7_75t_L g516 ( .A1(n_483), .A2(n_433), .B1(n_455), .B2(n_426), .C1(n_417), .C2(n_456), .Y(n_516) );
AOI322xp5_ASAP7_75t_L g517 ( .A1(n_468), .A2(n_456), .A3(n_429), .B1(n_426), .B2(n_452), .C1(n_459), .C2(n_425), .Y(n_517) );
INVx1_ASAP7_75t_L g518 ( .A(n_497), .Y(n_518) );
AOI21x1_ASAP7_75t_L g519 ( .A1(n_499), .A2(n_498), .B(n_487), .Y(n_519) );
INVxp67_ASAP7_75t_L g520 ( .A(n_495), .Y(n_520) );
NAND2x1_ASAP7_75t_L g521 ( .A(n_498), .B(n_446), .Y(n_521) );
NAND2xp5_ASAP7_75t_L g522 ( .A(n_496), .B(n_425), .Y(n_522) );
AOI22xp33_ASAP7_75t_L g523 ( .A1(n_468), .A2(n_458), .B1(n_460), .B2(n_459), .Y(n_523) );
HB1xp67_ASAP7_75t_L g524 ( .A(n_466), .Y(n_524) );
NAND2x1_ASAP7_75t_L g525 ( .A(n_463), .B(n_446), .Y(n_525) );
INVx1_ASAP7_75t_L g526 ( .A(n_491), .Y(n_526) );
AOI221xp5_ASAP7_75t_L g527 ( .A1(n_470), .A2(n_454), .B1(n_445), .B2(n_442), .C(n_192), .Y(n_527) );
OAI32xp33_ASAP7_75t_L g528 ( .A1(n_492), .A2(n_453), .A3(n_445), .B1(n_442), .B2(n_451), .Y(n_528) );
OAI22xp33_ASAP7_75t_L g529 ( .A1(n_477), .A2(n_424), .B1(n_250), .B2(n_221), .Y(n_529) );
AND2x4_ASAP7_75t_L g530 ( .A(n_463), .B(n_424), .Y(n_530) );
NAND3xp33_ASAP7_75t_SL g531 ( .A(n_509), .B(n_493), .C(n_488), .Y(n_531) );
NAND2xp5_ASAP7_75t_SL g532 ( .A(n_510), .B(n_471), .Y(n_532) );
XNOR2xp5_ASAP7_75t_L g533 ( .A(n_507), .B(n_469), .Y(n_533) );
O2A1O1Ixp5_ASAP7_75t_L g534 ( .A1(n_512), .A2(n_467), .B(n_500), .C(n_501), .Y(n_534) );
INVx4_ASAP7_75t_L g535 ( .A(n_530), .Y(n_535) );
OAI21xp33_ASAP7_75t_L g536 ( .A1(n_517), .A2(n_494), .B(n_485), .Y(n_536) );
O2A1O1Ixp33_ASAP7_75t_SL g537 ( .A1(n_512), .A2(n_476), .B(n_473), .C(n_474), .Y(n_537) );
INVx1_ASAP7_75t_L g538 ( .A(n_504), .Y(n_538) );
INVx1_ASAP7_75t_L g539 ( .A(n_505), .Y(n_539) );
AOI221xp5_ASAP7_75t_L g540 ( .A1(n_513), .A2(n_482), .B1(n_479), .B2(n_490), .C(n_181), .Y(n_540) );
INVx1_ASAP7_75t_L g541 ( .A(n_506), .Y(n_541) );
INVx1_ASAP7_75t_L g542 ( .A(n_518), .Y(n_542) );
INVx1_ASAP7_75t_SL g543 ( .A(n_521), .Y(n_543) );
INVx2_ASAP7_75t_L g544 ( .A(n_524), .Y(n_544) );
INVx1_ASAP7_75t_L g545 ( .A(n_526), .Y(n_545) );
BUFx3_ASAP7_75t_L g546 ( .A(n_525), .Y(n_546) );
NAND2xp5_ASAP7_75t_L g547 ( .A(n_508), .B(n_424), .Y(n_547) );
INVx1_ASAP7_75t_L g548 ( .A(n_503), .Y(n_548) );
NOR2xp33_ASAP7_75t_R g549 ( .A(n_519), .B(n_70), .Y(n_549) );
OAI32xp33_ASAP7_75t_L g550 ( .A1(n_520), .A2(n_250), .A3(n_221), .B1(n_71), .B2(n_72), .Y(n_550) );
OR2x2_ASAP7_75t_L g551 ( .A(n_522), .B(n_176), .Y(n_551) );
OAI21xp5_ASAP7_75t_SL g552 ( .A1(n_532), .A2(n_531), .B(n_543), .Y(n_552) );
CKINVDCx20_ASAP7_75t_R g553 ( .A(n_533), .Y(n_553) );
NOR2x1_ASAP7_75t_L g554 ( .A(n_532), .B(n_509), .Y(n_554) );
AOI322xp5_ASAP7_75t_L g555 ( .A1(n_536), .A2(n_502), .A3(n_515), .B1(n_511), .B2(n_523), .C1(n_520), .C2(n_530), .Y(n_555) );
NAND4xp25_ASAP7_75t_L g556 ( .A(n_534), .B(n_516), .C(n_528), .D(n_527), .Y(n_556) );
NAND3xp33_ASAP7_75t_L g557 ( .A(n_548), .B(n_529), .C(n_514), .Y(n_557) );
INVx2_ASAP7_75t_SL g558 ( .A(n_535), .Y(n_558) );
AOI32xp33_ASAP7_75t_L g559 ( .A1(n_546), .A2(n_235), .A3(n_278), .B1(n_279), .B2(n_197), .Y(n_559) );
NOR2xp33_ASAP7_75t_L g560 ( .A(n_553), .B(n_542), .Y(n_560) );
BUFx2_ASAP7_75t_L g561 ( .A(n_558), .Y(n_561) );
AOI21xp5_ASAP7_75t_L g562 ( .A1(n_552), .A2(n_537), .B(n_550), .Y(n_562) );
AND2x4_ASAP7_75t_L g563 ( .A(n_554), .B(n_541), .Y(n_563) );
NAND2xp5_ASAP7_75t_L g564 ( .A(n_555), .B(n_538), .Y(n_564) );
AOI21xp5_ASAP7_75t_L g565 ( .A1(n_552), .A2(n_537), .B(n_547), .Y(n_565) );
NOR2x1_ASAP7_75t_SL g566 ( .A(n_557), .B(n_544), .Y(n_566) );
AOI221xp5_ASAP7_75t_L g567 ( .A1(n_556), .A2(n_539), .B1(n_540), .B2(n_545), .C(n_544), .Y(n_567) );
AOI221xp5_ASAP7_75t_SL g568 ( .A1(n_556), .A2(n_551), .B1(n_549), .B2(n_279), .C(n_197), .Y(n_568) );
AOI211xp5_ASAP7_75t_L g569 ( .A1(n_559), .A2(n_235), .B(n_552), .C(n_556), .Y(n_569) );
OA22x2_ASAP7_75t_L g570 ( .A1(n_552), .A2(n_558), .B1(n_532), .B2(n_535), .Y(n_570) );
O2A1O1Ixp33_ASAP7_75t_L g571 ( .A1(n_552), .A2(n_554), .B(n_556), .C(n_537), .Y(n_571) );
NOR2x1p5_ASAP7_75t_L g572 ( .A(n_564), .B(n_570), .Y(n_572) );
NOR3xp33_ASAP7_75t_L g573 ( .A(n_571), .B(n_569), .C(n_568), .Y(n_573) );
INVx1_ASAP7_75t_SL g574 ( .A(n_561), .Y(n_574) );
NOR3xp33_ASAP7_75t_SL g575 ( .A(n_562), .B(n_564), .C(n_565), .Y(n_575) );
HB1xp67_ASAP7_75t_L g576 ( .A(n_574), .Y(n_576) );
NAND2xp5_ASAP7_75t_L g577 ( .A(n_575), .B(n_567), .Y(n_577) );
NOR2x1_ASAP7_75t_L g578 ( .A(n_572), .B(n_563), .Y(n_578) );
INVx1_ASAP7_75t_SL g579 ( .A(n_576), .Y(n_579) );
NAND2xp5_ASAP7_75t_L g580 ( .A(n_577), .B(n_573), .Y(n_580) );
INVx1_ASAP7_75t_L g581 ( .A(n_579), .Y(n_581) );
AOI22xp5_ASAP7_75t_SL g582 ( .A1(n_581), .A2(n_580), .B1(n_563), .B2(n_560), .Y(n_582) );
AOI21xp5_ASAP7_75t_L g583 ( .A1(n_582), .A2(n_578), .B(n_566), .Y(n_583) );
endmodule