module fake_jpeg_1090_n_615 (n_13, n_1, n_10, n_6, n_14, n_18, n_4, n_16, n_3, n_0, n_9, n_5, n_11, n_17, n_2, n_12, n_8, n_15, n_7, n_615);

input n_13;
input n_1;
input n_10;
input n_6;
input n_14;
input n_18;
input n_4;
input n_16;
input n_3;
input n_0;
input n_9;
input n_5;
input n_11;
input n_17;
input n_2;
input n_12;
input n_8;
input n_15;
input n_7;

output n_615;

wire n_529;
wire n_595;
wire n_390;
wire n_552;
wire n_253;
wire n_330;
wire n_369;
wire n_158;
wire n_73;
wire n_152;
wire n_252;
wire n_19;
wire n_182;
wire n_525;
wire n_385;
wire n_464;
wire n_228;
wire n_134;
wire n_428;
wire n_127;
wire n_502;
wire n_295;
wire n_28;
wire n_38;
wire n_293;
wire n_432;
wire n_340;
wire n_381;
wire n_466;
wire n_586;
wire n_377;
wire n_291;
wire n_236;
wire n_483;
wire n_394;
wire n_392;
wire n_141;
wire n_331;
wire n_175;
wire n_284;
wire n_171;
wire n_263;
wire n_336;
wire n_27;
wire n_365;
wire n_179;
wire n_185;
wire n_338;
wire n_129;
wire n_451;
wire n_148;
wire n_434;
wire n_324;
wire n_611;
wire n_44;
wire n_355;
wire n_519;
wire n_276;
wire n_143;
wire n_431;
wire n_102;
wire n_549;
wire n_196;
wire n_66;
wire n_374;
wire n_566;
wire n_142;
wire n_362;
wire n_417;
wire n_470;
wire n_597;
wire n_172;
wire n_547;
wire n_345;
wire n_591;
wire n_78;
wire n_241;
wire n_359;
wire n_214;
wire n_461;
wire n_304;
wire n_60;
wire n_513;
wire n_283;
wire n_107;
wire n_490;
wire n_517;
wire n_479;
wire n_415;
wire n_543;
wire n_357;
wire n_89;
wire n_131;
wire n_607;
wire n_294;
wire n_230;
wire n_170;
wire n_602;
wire n_313;
wire n_542;
wire n_574;
wire n_264;
wire n_437;
wire n_93;
wire n_227;
wire n_559;
wire n_48;
wire n_465;
wire n_200;
wire n_582;
wire n_192;
wire n_265;
wire n_115;
wire n_270;
wire n_387;
wire n_579;
wire n_416;
wire n_221;
wire n_256;
wire n_454;
wire n_540;
wire n_213;
wire n_292;
wire n_135;
wire n_435;
wire n_189;
wire n_370;
wire n_410;
wire n_571;
wire n_82;
wire n_155;
wire n_508;
wire n_309;
wire n_286;
wire n_427;
wire n_225;
wire n_105;
wire n_401;
wire n_493;
wire n_326;
wire n_51;
wire n_59;
wire n_84;
wire n_606;
wire n_496;
wire n_166;
wire n_65;
wire n_191;
wire n_193;
wire n_487;
wire n_42;
wire n_49;
wire n_569;
wire n_596;
wire n_400;
wire n_319;
wire n_116;
wire n_126;
wire n_220;
wire n_74;
wire n_137;
wire n_455;
wire n_544;
wire n_31;
wire n_277;
wire n_255;
wire n_605;
wire n_601;
wire n_406;
wire n_124;
wire n_447;
wire n_223;
wire n_288;
wire n_21;
wire n_349;
wire n_393;
wire n_234;
wire n_530;
wire n_23;
wire n_69;
wire n_195;
wire n_450;
wire n_557;
wire n_408;
wire n_80;
wire n_562;
wire n_204;
wire n_306;
wire n_429;
wire n_497;
wire n_368;
wire n_298;
wire n_106;
wire n_545;
wire n_386;
wire n_418;
wire n_327;
wire n_75;
wire n_122;
wire n_246;
wire n_233;
wire n_99;
wire n_130;
wire n_70;
wire n_458;
wire n_423;
wire n_85;
wire n_163;
wire n_136;
wire n_448;
wire n_139;
wire n_584;
wire n_254;
wire n_608;
wire n_323;
wire n_165;
wire n_108;
wire n_68;
wire n_52;
wire n_388;
wire n_94;
wire n_206;
wire n_463;
wire n_92;
wire n_332;
wire n_310;
wire n_346;
wire n_34;
wire n_425;
wire n_39;
wire n_371;
wire n_164;
wire n_505;
wire n_474;
wire n_539;
wire n_261;
wire n_146;
wire n_104;
wire n_285;
wire n_300;
wire n_299;
wire n_442;
wire n_211;
wire n_79;
wire n_162;
wire n_67;
wire n_271;
wire n_575;
wire n_268;
wire n_404;
wire n_91;
wire n_511;
wire n_486;
wire n_305;
wire n_161;
wire n_441;
wire n_555;
wire n_342;
wire n_101;
wire n_226;
wire n_509;
wire n_149;
wire n_87;
wire n_46;
wire n_578;
wire n_589;
wire n_176;
wire n_315;
wire n_222;
wire n_353;
wire n_614;
wire n_97;
wire n_573;
wire n_498;
wire n_382;
wire n_460;
wire n_237;
wire n_188;
wire n_610;
wire n_174;
wire n_198;
wire n_422;
wire n_560;
wire n_190;
wire n_510;
wire n_32;
wire n_100;
wire n_258;
wire n_128;
wire n_366;
wire n_536;
wire n_289;
wire n_316;
wire n_229;
wire n_144;
wire n_64;
wire n_180;
wire n_245;
wire n_414;
wire n_178;
wire n_231;
wire n_203;
wire n_537;
wire n_110;
wire n_594;
wire n_590;
wire n_531;
wire n_76;
wire n_278;
wire n_343;
wire n_577;
wire n_26;
wire n_88;
wire n_397;
wire n_592;
wire n_363;
wire n_570;
wire n_238;
wire n_598;
wire n_29;
wire n_103;
wire n_150;
wire n_350;
wire n_352;
wire n_488;
wire n_367;
wire n_383;
wire n_187;
wire n_272;
wire n_280;
wire n_554;
wire n_301;
wire n_609;
wire n_201;
wire n_420;
wire n_321;
wire n_40;
wire n_250;
wire n_71;
wire n_456;
wire n_501;
wire n_389;
wire n_457;
wire n_523;
wire n_339;
wire n_109;
wire n_267;
wire n_480;
wire n_533;
wire n_612;
wire n_296;
wire n_384;
wire n_588;
wire n_168;
wire n_459;
wire n_274;
wire n_485;
wire n_585;
wire n_491;
wire n_24;
wire n_526;
wire n_467;
wire n_269;
wire n_572;
wire n_546;
wire n_287;
wire n_219;
wire n_452;
wire n_433;
wire n_77;
wire n_473;
wire n_45;
wire n_520;
wire n_476;
wire n_337;
wire n_317;
wire n_20;
wire n_145;
wire n_360;
wire n_407;
wire n_303;
wire n_259;
wire n_399;
wire n_90;
wire n_328;
wire n_344;
wire n_218;
wire n_63;
wire n_599;
wire n_239;
wire n_243;
wire n_481;
wire n_348;
wire n_587;
wire n_439;
wire n_262;
wire n_240;
wire n_398;
wire n_56;
wire n_583;
wire n_522;
wire n_333;
wire n_518;
wire n_132;
wire n_133;
wire n_378;
wire n_419;
wire n_565;
wire n_302;
wire n_216;
wire n_528;
wire n_184;
wire n_311;
wire n_329;
wire n_314;
wire n_208;
wire n_308;
wire n_421;
wire n_297;
wire n_320;
wire n_210;
wire n_35;
wire n_123;
wire n_453;
wire n_500;
wire n_260;
wire n_199;
wire n_550;
wire n_413;
wire n_275;
wire n_494;
wire n_604;
wire n_169;
wire n_153;
wire n_411;
wire n_322;
wire n_551;
wire n_36;
wire n_62;
wire n_600;
wire n_492;
wire n_603;
wire n_478;
wire n_118;
wire n_140;
wire n_361;
wire n_567;
wire n_318;
wire n_96;
wire n_159;
wire n_117;
wire n_354;
wire n_515;
wire n_347;
wire n_521;
wire n_424;
wire n_55;
wire n_312;
wire n_358;
wire n_47;
wire n_538;
wire n_147;
wire n_449;
wire n_98;
wire n_251;
wire n_534;
wire n_472;
wire n_279;
wire n_593;
wire n_154;
wire n_495;
wire n_205;
wire n_507;
wire n_379;
wire n_503;
wire n_114;
wire n_444;
wire n_499;
wire n_281;
wire n_376;
wire n_207;
wire n_235;
wire n_50;
wire n_160;
wire n_194;
wire n_506;
wire n_57;
wire n_405;
wire n_356;
wire n_119;
wire n_484;
wire n_568;
wire n_83;
wire n_395;
wire n_125;
wire n_81;
wire n_224;
wire n_403;
wire n_113;
wire n_248;
wire n_380;
wire n_30;
wire n_307;
wire n_446;
wire n_576;
wire n_469;
wire n_111;
wire n_197;
wire n_375;
wire n_396;
wire n_186;
wire n_440;
wire n_202;
wire n_430;
wire n_25;
wire n_436;
wire n_37;
wire n_121;
wire n_334;
wire n_177;
wire n_364;
wire n_553;
wire n_257;
wire n_61;
wire n_173;
wire n_561;
wire n_244;
wire n_232;
wire n_527;
wire n_482;
wire n_58;
wire n_41;
wire n_613;
wire n_266;
wire n_548;
wire n_72;
wire n_512;
wire n_445;
wire n_443;
wire n_215;
wire n_212;
wire n_516;
wire n_183;
wire n_409;
wire n_532;
wire n_249;
wire n_412;
wire n_581;
wire n_217;
wire n_471;
wire n_580;
wire n_541;
wire n_53;
wire n_372;
wire n_558;
wire n_33;
wire n_54;
wire n_477;
wire n_391;
wire n_535;
wire n_489;
wire n_209;
wire n_22;
wire n_138;
wire n_556;
wire n_524;
wire n_402;
wire n_563;
wire n_504;
wire n_438;
wire n_475;
wire n_157;
wire n_247;
wire n_273;
wire n_86;
wire n_156;
wire n_373;
wire n_112;
wire n_95;
wire n_341;
wire n_151;
wire n_426;
wire n_290;
wire n_242;
wire n_514;
wire n_564;
wire n_351;
wire n_325;
wire n_462;
wire n_167;
wire n_335;
wire n_120;
wire n_43;
wire n_468;
wire n_282;
wire n_181;

INVxp67_ASAP7_75t_L g19 ( 
.A(n_14),
.Y(n_19)
);

BUFx12f_ASAP7_75t_L g20 ( 
.A(n_11),
.Y(n_20)
);

CKINVDCx20_ASAP7_75t_R g21 ( 
.A(n_16),
.Y(n_21)
);

BUFx3_ASAP7_75t_L g22 ( 
.A(n_5),
.Y(n_22)
);

BUFx12f_ASAP7_75t_L g23 ( 
.A(n_12),
.Y(n_23)
);

BUFx12f_ASAP7_75t_L g24 ( 
.A(n_16),
.Y(n_24)
);

CKINVDCx20_ASAP7_75t_R g25 ( 
.A(n_15),
.Y(n_25)
);

BUFx6f_ASAP7_75t_L g26 ( 
.A(n_0),
.Y(n_26)
);

INVx2_ASAP7_75t_L g27 ( 
.A(n_8),
.Y(n_27)
);

BUFx6f_ASAP7_75t_L g28 ( 
.A(n_13),
.Y(n_28)
);

INVx1_ASAP7_75t_L g29 ( 
.A(n_14),
.Y(n_29)
);

BUFx3_ASAP7_75t_L g30 ( 
.A(n_6),
.Y(n_30)
);

BUFx6f_ASAP7_75t_L g31 ( 
.A(n_17),
.Y(n_31)
);

INVx3_ASAP7_75t_L g32 ( 
.A(n_1),
.Y(n_32)
);

BUFx12f_ASAP7_75t_L g33 ( 
.A(n_14),
.Y(n_33)
);

NOR2xp33_ASAP7_75t_L g34 ( 
.A(n_2),
.B(n_14),
.Y(n_34)
);

CKINVDCx20_ASAP7_75t_R g35 ( 
.A(n_18),
.Y(n_35)
);

BUFx5_ASAP7_75t_L g36 ( 
.A(n_7),
.Y(n_36)
);

CKINVDCx16_ASAP7_75t_R g37 ( 
.A(n_12),
.Y(n_37)
);

BUFx12f_ASAP7_75t_L g38 ( 
.A(n_11),
.Y(n_38)
);

BUFx16f_ASAP7_75t_L g39 ( 
.A(n_10),
.Y(n_39)
);

BUFx6f_ASAP7_75t_L g40 ( 
.A(n_6),
.Y(n_40)
);

CKINVDCx20_ASAP7_75t_R g41 ( 
.A(n_0),
.Y(n_41)
);

BUFx2_ASAP7_75t_L g42 ( 
.A(n_16),
.Y(n_42)
);

CKINVDCx20_ASAP7_75t_R g43 ( 
.A(n_9),
.Y(n_43)
);

INVx3_ASAP7_75t_L g44 ( 
.A(n_6),
.Y(n_44)
);

INVx13_ASAP7_75t_L g45 ( 
.A(n_12),
.Y(n_45)
);

CKINVDCx20_ASAP7_75t_R g46 ( 
.A(n_6),
.Y(n_46)
);

INVx1_ASAP7_75t_L g47 ( 
.A(n_9),
.Y(n_47)
);

INVx1_ASAP7_75t_L g48 ( 
.A(n_13),
.Y(n_48)
);

CKINVDCx20_ASAP7_75t_R g49 ( 
.A(n_13),
.Y(n_49)
);

CKINVDCx20_ASAP7_75t_R g50 ( 
.A(n_9),
.Y(n_50)
);

INVx2_ASAP7_75t_L g51 ( 
.A(n_12),
.Y(n_51)
);

BUFx6f_ASAP7_75t_L g52 ( 
.A(n_7),
.Y(n_52)
);

BUFx5_ASAP7_75t_L g53 ( 
.A(n_7),
.Y(n_53)
);

BUFx8_ASAP7_75t_L g54 ( 
.A(n_18),
.Y(n_54)
);

BUFx12_ASAP7_75t_L g55 ( 
.A(n_10),
.Y(n_55)
);

INVx3_ASAP7_75t_L g56 ( 
.A(n_17),
.Y(n_56)
);

INVx1_ASAP7_75t_L g57 ( 
.A(n_10),
.Y(n_57)
);

INVx1_ASAP7_75t_L g58 ( 
.A(n_29),
.Y(n_58)
);

INVx1_ASAP7_75t_L g193 ( 
.A(n_58),
.Y(n_193)
);

INVx1_ASAP7_75t_L g59 ( 
.A(n_29),
.Y(n_59)
);

INVx1_ASAP7_75t_L g205 ( 
.A(n_59),
.Y(n_205)
);

INVx2_ASAP7_75t_L g60 ( 
.A(n_27),
.Y(n_60)
);

INVx2_ASAP7_75t_L g140 ( 
.A(n_60),
.Y(n_140)
);

CKINVDCx20_ASAP7_75t_R g61 ( 
.A(n_42),
.Y(n_61)
);

NOR2xp33_ASAP7_75t_L g130 ( 
.A(n_61),
.B(n_70),
.Y(n_130)
);

INVx4_ASAP7_75t_L g62 ( 
.A(n_36),
.Y(n_62)
);

INVx2_ASAP7_75t_SL g185 ( 
.A(n_62),
.Y(n_185)
);

BUFx6f_ASAP7_75t_L g63 ( 
.A(n_40),
.Y(n_63)
);

BUFx6f_ASAP7_75t_L g135 ( 
.A(n_63),
.Y(n_135)
);

INVx3_ASAP7_75t_L g64 ( 
.A(n_54),
.Y(n_64)
);

INVx4_ASAP7_75t_SL g217 ( 
.A(n_64),
.Y(n_217)
);

BUFx6f_ASAP7_75t_L g65 ( 
.A(n_40),
.Y(n_65)
);

BUFx6f_ASAP7_75t_L g154 ( 
.A(n_65),
.Y(n_154)
);

INVx2_ASAP7_75t_L g66 ( 
.A(n_27),
.Y(n_66)
);

INVx2_ASAP7_75t_L g143 ( 
.A(n_66),
.Y(n_143)
);

BUFx6f_ASAP7_75t_L g67 ( 
.A(n_40),
.Y(n_67)
);

BUFx6f_ASAP7_75t_L g171 ( 
.A(n_67),
.Y(n_171)
);

INVx8_ASAP7_75t_L g68 ( 
.A(n_39),
.Y(n_68)
);

BUFx2_ASAP7_75t_L g129 ( 
.A(n_68),
.Y(n_129)
);

INVx4_ASAP7_75t_SL g69 ( 
.A(n_54),
.Y(n_69)
);

BUFx3_ASAP7_75t_L g138 ( 
.A(n_69),
.Y(n_138)
);

CKINVDCx20_ASAP7_75t_R g70 ( 
.A(n_42),
.Y(n_70)
);

OR2x2_ASAP7_75t_L g71 ( 
.A(n_34),
.B(n_18),
.Y(n_71)
);

NAND2xp33_ASAP7_75t_SL g215 ( 
.A(n_71),
.B(n_91),
.Y(n_215)
);

BUFx12f_ASAP7_75t_L g72 ( 
.A(n_54),
.Y(n_72)
);

INVx5_ASAP7_75t_L g146 ( 
.A(n_72),
.Y(n_146)
);

INVx4_ASAP7_75t_L g73 ( 
.A(n_39),
.Y(n_73)
);

INVx3_ASAP7_75t_L g153 ( 
.A(n_73),
.Y(n_153)
);

INVx6_ASAP7_75t_L g74 ( 
.A(n_26),
.Y(n_74)
);

BUFx6f_ASAP7_75t_L g173 ( 
.A(n_74),
.Y(n_173)
);

INVx2_ASAP7_75t_L g75 ( 
.A(n_51),
.Y(n_75)
);

INVx2_ASAP7_75t_L g152 ( 
.A(n_75),
.Y(n_152)
);

BUFx10_ASAP7_75t_L g76 ( 
.A(n_39),
.Y(n_76)
);

BUFx2_ASAP7_75t_L g142 ( 
.A(n_76),
.Y(n_142)
);

NAND2xp5_ASAP7_75t_L g77 ( 
.A(n_51),
.B(n_17),
.Y(n_77)
);

NAND2xp5_ASAP7_75t_L g128 ( 
.A(n_77),
.B(n_99),
.Y(n_128)
);

INVx3_ASAP7_75t_L g78 ( 
.A(n_54),
.Y(n_78)
);

INVx3_ASAP7_75t_L g160 ( 
.A(n_78),
.Y(n_160)
);

INVx2_ASAP7_75t_L g79 ( 
.A(n_32),
.Y(n_79)
);

INVx2_ASAP7_75t_L g158 ( 
.A(n_79),
.Y(n_158)
);

INVx13_ASAP7_75t_L g80 ( 
.A(n_45),
.Y(n_80)
);

BUFx16f_ASAP7_75t_L g149 ( 
.A(n_80),
.Y(n_149)
);

INVx2_ASAP7_75t_L g81 ( 
.A(n_32),
.Y(n_81)
);

INVx2_ASAP7_75t_L g167 ( 
.A(n_81),
.Y(n_167)
);

BUFx6f_ASAP7_75t_L g82 ( 
.A(n_26),
.Y(n_82)
);

BUFx6f_ASAP7_75t_L g177 ( 
.A(n_82),
.Y(n_177)
);

BUFx8_ASAP7_75t_L g83 ( 
.A(n_37),
.Y(n_83)
);

BUFx12f_ASAP7_75t_L g131 ( 
.A(n_83),
.Y(n_131)
);

INVx1_ASAP7_75t_L g84 ( 
.A(n_47),
.Y(n_84)
);

NOR2xp33_ASAP7_75t_L g150 ( 
.A(n_84),
.B(n_92),
.Y(n_150)
);

BUFx3_ASAP7_75t_L g85 ( 
.A(n_22),
.Y(n_85)
);

BUFx2_ASAP7_75t_L g169 ( 
.A(n_85),
.Y(n_169)
);

BUFx3_ASAP7_75t_L g86 ( 
.A(n_22),
.Y(n_86)
);

INVx5_ASAP7_75t_L g166 ( 
.A(n_86),
.Y(n_166)
);

BUFx24_ASAP7_75t_L g87 ( 
.A(n_45),
.Y(n_87)
);

INVx11_ASAP7_75t_L g207 ( 
.A(n_87),
.Y(n_207)
);

INVx11_ASAP7_75t_L g88 ( 
.A(n_20),
.Y(n_88)
);

INVx11_ASAP7_75t_L g137 ( 
.A(n_88),
.Y(n_137)
);

INVx3_ASAP7_75t_L g89 ( 
.A(n_24),
.Y(n_89)
);

INVx3_ASAP7_75t_L g161 ( 
.A(n_89),
.Y(n_161)
);

INVx11_ASAP7_75t_L g90 ( 
.A(n_20),
.Y(n_90)
);

INVx11_ASAP7_75t_L g147 ( 
.A(n_90),
.Y(n_147)
);

INVx1_ASAP7_75t_SL g91 ( 
.A(n_20),
.Y(n_91)
);

INVx1_ASAP7_75t_L g92 ( 
.A(n_47),
.Y(n_92)
);

BUFx6f_ASAP7_75t_L g93 ( 
.A(n_28),
.Y(n_93)
);

BUFx6f_ASAP7_75t_L g178 ( 
.A(n_93),
.Y(n_178)
);

CKINVDCx20_ASAP7_75t_R g94 ( 
.A(n_42),
.Y(n_94)
);

NOR2xp33_ASAP7_75t_L g176 ( 
.A(n_94),
.B(n_96),
.Y(n_176)
);

BUFx6f_ASAP7_75t_L g95 ( 
.A(n_28),
.Y(n_95)
);

BUFx6f_ASAP7_75t_L g182 ( 
.A(n_95),
.Y(n_182)
);

CKINVDCx20_ASAP7_75t_R g96 ( 
.A(n_31),
.Y(n_96)
);

BUFx10_ASAP7_75t_L g97 ( 
.A(n_20),
.Y(n_97)
);

BUFx12f_ASAP7_75t_L g132 ( 
.A(n_97),
.Y(n_132)
);

INVx3_ASAP7_75t_L g98 ( 
.A(n_24),
.Y(n_98)
);

INVx3_ASAP7_75t_L g162 ( 
.A(n_98),
.Y(n_162)
);

NAND2xp5_ASAP7_75t_L g99 ( 
.A(n_21),
.B(n_15),
.Y(n_99)
);

INVx8_ASAP7_75t_L g100 ( 
.A(n_23),
.Y(n_100)
);

INVx5_ASAP7_75t_L g194 ( 
.A(n_100),
.Y(n_194)
);

CKINVDCx20_ASAP7_75t_R g101 ( 
.A(n_31),
.Y(n_101)
);

NOR2xp33_ASAP7_75t_L g197 ( 
.A(n_101),
.B(n_112),
.Y(n_197)
);

BUFx6f_ASAP7_75t_L g102 ( 
.A(n_52),
.Y(n_102)
);

BUFx6f_ASAP7_75t_L g188 ( 
.A(n_102),
.Y(n_188)
);

INVx2_ASAP7_75t_L g103 ( 
.A(n_44),
.Y(n_103)
);

INVx2_ASAP7_75t_L g168 ( 
.A(n_103),
.Y(n_168)
);

INVx6_ASAP7_75t_L g104 ( 
.A(n_52),
.Y(n_104)
);

BUFx6f_ASAP7_75t_L g199 ( 
.A(n_104),
.Y(n_199)
);

BUFx16f_ASAP7_75t_L g105 ( 
.A(n_19),
.Y(n_105)
);

BUFx12f_ASAP7_75t_L g202 ( 
.A(n_105),
.Y(n_202)
);

BUFx24_ASAP7_75t_L g106 ( 
.A(n_19),
.Y(n_106)
);

CKINVDCx16_ASAP7_75t_R g201 ( 
.A(n_106),
.Y(n_201)
);

NOR2xp33_ASAP7_75t_L g107 ( 
.A(n_21),
.B(n_15),
.Y(n_107)
);

NOR2xp33_ASAP7_75t_SL g148 ( 
.A(n_107),
.B(n_35),
.Y(n_148)
);

BUFx5_ASAP7_75t_L g108 ( 
.A(n_36),
.Y(n_108)
);

INVx4_ASAP7_75t_L g218 ( 
.A(n_108),
.Y(n_218)
);

BUFx6f_ASAP7_75t_L g109 ( 
.A(n_30),
.Y(n_109)
);

BUFx6f_ASAP7_75t_L g204 ( 
.A(n_109),
.Y(n_204)
);

BUFx3_ASAP7_75t_L g110 ( 
.A(n_30),
.Y(n_110)
);

INVx5_ASAP7_75t_L g208 ( 
.A(n_110),
.Y(n_208)
);

INVx3_ASAP7_75t_L g111 ( 
.A(n_24),
.Y(n_111)
);

HB1xp67_ASAP7_75t_L g220 ( 
.A(n_111),
.Y(n_220)
);

CKINVDCx16_ASAP7_75t_R g112 ( 
.A(n_24),
.Y(n_112)
);

BUFx12_ASAP7_75t_L g113 ( 
.A(n_56),
.Y(n_113)
);

CKINVDCx16_ASAP7_75t_R g211 ( 
.A(n_113),
.Y(n_211)
);

CKINVDCx20_ASAP7_75t_R g114 ( 
.A(n_25),
.Y(n_114)
);

NOR2xp33_ASAP7_75t_L g209 ( 
.A(n_114),
.B(n_115),
.Y(n_209)
);

CKINVDCx20_ASAP7_75t_R g115 ( 
.A(n_25),
.Y(n_115)
);

BUFx6f_ASAP7_75t_L g116 ( 
.A(n_23),
.Y(n_116)
);

BUFx6f_ASAP7_75t_L g210 ( 
.A(n_116),
.Y(n_210)
);

BUFx6f_ASAP7_75t_L g117 ( 
.A(n_23),
.Y(n_117)
);

INVx6_ASAP7_75t_L g151 ( 
.A(n_117),
.Y(n_151)
);

INVx1_ASAP7_75t_L g118 ( 
.A(n_48),
.Y(n_118)
);

INVx2_ASAP7_75t_L g184 ( 
.A(n_118),
.Y(n_184)
);

INVx2_ASAP7_75t_L g119 ( 
.A(n_44),
.Y(n_119)
);

INVx2_ASAP7_75t_L g186 ( 
.A(n_119),
.Y(n_186)
);

AND2x4_ASAP7_75t_L g120 ( 
.A(n_56),
.B(n_0),
.Y(n_120)
);

NAND2x1_ASAP7_75t_SL g200 ( 
.A(n_120),
.B(n_0),
.Y(n_200)
);

BUFx6f_ASAP7_75t_L g121 ( 
.A(n_23),
.Y(n_121)
);

INVx6_ASAP7_75t_L g164 ( 
.A(n_121),
.Y(n_164)
);

BUFx6f_ASAP7_75t_L g122 ( 
.A(n_33),
.Y(n_122)
);

INVx8_ASAP7_75t_L g139 ( 
.A(n_122),
.Y(n_139)
);

BUFx6f_ASAP7_75t_L g123 ( 
.A(n_33),
.Y(n_123)
);

INVx8_ASAP7_75t_L g180 ( 
.A(n_123),
.Y(n_180)
);

INVx4_ASAP7_75t_L g124 ( 
.A(n_53),
.Y(n_124)
);

INVx4_ASAP7_75t_L g136 ( 
.A(n_124),
.Y(n_136)
);

INVx8_ASAP7_75t_L g125 ( 
.A(n_33),
.Y(n_125)
);

INVx4_ASAP7_75t_L g145 ( 
.A(n_125),
.Y(n_145)
);

INVx6_ASAP7_75t_L g126 ( 
.A(n_33),
.Y(n_126)
);

INVx2_ASAP7_75t_L g189 ( 
.A(n_126),
.Y(n_189)
);

INVx4_ASAP7_75t_L g127 ( 
.A(n_53),
.Y(n_127)
);

INVx4_ASAP7_75t_L g155 ( 
.A(n_127),
.Y(n_155)
);

NAND2xp5_ASAP7_75t_SL g133 ( 
.A(n_71),
.B(n_107),
.Y(n_133)
);

NOR2xp33_ASAP7_75t_SL g225 ( 
.A(n_133),
.B(n_141),
.Y(n_225)
);

AOI22xp33_ASAP7_75t_SL g134 ( 
.A1(n_72),
.A2(n_38),
.B1(n_35),
.B2(n_57),
.Y(n_134)
);

AOI22xp33_ASAP7_75t_SL g227 ( 
.A1(n_134),
.A2(n_214),
.B1(n_125),
.B2(n_80),
.Y(n_227)
);

CKINVDCx20_ASAP7_75t_R g141 ( 
.A(n_105),
.Y(n_141)
);

CKINVDCx20_ASAP7_75t_R g144 ( 
.A(n_83),
.Y(n_144)
);

NOR2xp33_ASAP7_75t_L g222 ( 
.A(n_144),
.B(n_148),
.Y(n_222)
);

NOR2xp33_ASAP7_75t_SL g156 ( 
.A(n_73),
.B(n_50),
.Y(n_156)
);

NOR2xp33_ASAP7_75t_L g265 ( 
.A(n_156),
.B(n_163),
.Y(n_265)
);

OR2x2_ASAP7_75t_L g157 ( 
.A(n_69),
.B(n_57),
.Y(n_157)
);

NAND2x1_ASAP7_75t_SL g226 ( 
.A(n_157),
.B(n_200),
.Y(n_226)
);

INVx4_ASAP7_75t_L g159 ( 
.A(n_68),
.Y(n_159)
);

INVx4_ASAP7_75t_L g279 ( 
.A(n_159),
.Y(n_279)
);

NOR2xp33_ASAP7_75t_SL g163 ( 
.A(n_85),
.B(n_50),
.Y(n_163)
);

INVx11_ASAP7_75t_L g165 ( 
.A(n_72),
.Y(n_165)
);

INVx4_ASAP7_75t_L g257 ( 
.A(n_165),
.Y(n_257)
);

CKINVDCx20_ASAP7_75t_R g170 ( 
.A(n_126),
.Y(n_170)
);

NOR2xp33_ASAP7_75t_L g271 ( 
.A(n_170),
.B(n_191),
.Y(n_271)
);

NAND2xp5_ASAP7_75t_SL g172 ( 
.A(n_86),
.B(n_48),
.Y(n_172)
);

NAND2xp5_ASAP7_75t_L g223 ( 
.A(n_172),
.B(n_174),
.Y(n_223)
);

NAND2xp5_ASAP7_75t_L g174 ( 
.A(n_120),
.B(n_49),
.Y(n_174)
);

INVx4_ASAP7_75t_L g175 ( 
.A(n_88),
.Y(n_175)
);

INVx4_ASAP7_75t_L g259 ( 
.A(n_175),
.Y(n_259)
);

NAND2xp5_ASAP7_75t_L g179 ( 
.A(n_120),
.B(n_49),
.Y(n_179)
);

NAND2xp5_ASAP7_75t_L g224 ( 
.A(n_179),
.B(n_181),
.Y(n_224)
);

NAND2xp5_ASAP7_75t_L g181 ( 
.A(n_63),
.B(n_46),
.Y(n_181)
);

INVx11_ASAP7_75t_L g183 ( 
.A(n_87),
.Y(n_183)
);

INVx4_ASAP7_75t_L g293 ( 
.A(n_183),
.Y(n_293)
);

AOI22xp5_ASAP7_75t_L g187 ( 
.A1(n_82),
.A2(n_46),
.B1(n_43),
.B2(n_41),
.Y(n_187)
);

OAI22xp5_ASAP7_75t_L g229 ( 
.A1(n_187),
.A2(n_219),
.B1(n_123),
.B2(n_97),
.Y(n_229)
);

NAND2xp5_ASAP7_75t_L g190 ( 
.A(n_65),
.B(n_43),
.Y(n_190)
);

NAND2xp5_ASAP7_75t_L g233 ( 
.A(n_190),
.B(n_192),
.Y(n_233)
);

CKINVDCx20_ASAP7_75t_R g191 ( 
.A(n_116),
.Y(n_191)
);

NAND2xp5_ASAP7_75t_SL g192 ( 
.A(n_110),
.B(n_41),
.Y(n_192)
);

NAND2xp5_ASAP7_75t_SL g195 ( 
.A(n_109),
.B(n_38),
.Y(n_195)
);

NAND2xp5_ASAP7_75t_L g248 ( 
.A(n_195),
.B(n_212),
.Y(n_248)
);

INVx4_ASAP7_75t_L g196 ( 
.A(n_90),
.Y(n_196)
);

INVx3_ASAP7_75t_L g240 ( 
.A(n_196),
.Y(n_240)
);

INVx2_ASAP7_75t_L g198 ( 
.A(n_74),
.Y(n_198)
);

INVx2_ASAP7_75t_L g230 ( 
.A(n_198),
.Y(n_230)
);

INVx4_ASAP7_75t_L g203 ( 
.A(n_100),
.Y(n_203)
);

INVx3_ASAP7_75t_L g262 ( 
.A(n_203),
.Y(n_262)
);

CKINVDCx20_ASAP7_75t_R g206 ( 
.A(n_117),
.Y(n_206)
);

NOR2xp33_ASAP7_75t_L g276 ( 
.A(n_206),
.B(n_11),
.Y(n_276)
);

NAND2xp5_ASAP7_75t_L g212 ( 
.A(n_67),
.B(n_38),
.Y(n_212)
);

INVx2_ASAP7_75t_L g213 ( 
.A(n_104),
.Y(n_213)
);

INVx2_ASAP7_75t_L g243 ( 
.A(n_213),
.Y(n_243)
);

AOI22xp33_ASAP7_75t_SL g214 ( 
.A1(n_127),
.A2(n_38),
.B1(n_55),
.B2(n_3),
.Y(n_214)
);

NAND2xp5_ASAP7_75t_L g216 ( 
.A(n_121),
.B(n_1),
.Y(n_216)
);

NAND2xp5_ASAP7_75t_L g282 ( 
.A(n_216),
.B(n_4),
.Y(n_282)
);

AOI22xp33_ASAP7_75t_L g219 ( 
.A1(n_93),
.A2(n_102),
.B1(n_95),
.B2(n_122),
.Y(n_219)
);

BUFx4f_ASAP7_75t_SL g221 ( 
.A(n_202),
.Y(n_221)
);

CKINVDCx16_ASAP7_75t_R g300 ( 
.A(n_221),
.Y(n_300)
);

INVxp67_ASAP7_75t_L g323 ( 
.A(n_227),
.Y(n_323)
);

INVx1_ASAP7_75t_L g228 ( 
.A(n_193),
.Y(n_228)
);

HB1xp67_ASAP7_75t_L g332 ( 
.A(n_228),
.Y(n_332)
);

AOI22xp33_ASAP7_75t_SL g303 ( 
.A1(n_229),
.A2(n_232),
.B1(n_245),
.B2(n_246),
.Y(n_303)
);

INVx1_ASAP7_75t_L g231 ( 
.A(n_205),
.Y(n_231)
);

HB1xp67_ASAP7_75t_L g334 ( 
.A(n_231),
.Y(n_334)
);

AOI22xp33_ASAP7_75t_SL g232 ( 
.A1(n_218),
.A2(n_76),
.B1(n_97),
.B2(n_113),
.Y(n_232)
);

XNOR2xp5_ASAP7_75t_SL g234 ( 
.A(n_128),
.B(n_150),
.Y(n_234)
);

MAJx2_ASAP7_75t_L g317 ( 
.A(n_234),
.B(n_211),
.C(n_201),
.Y(n_317)
);

INVx1_ASAP7_75t_L g235 ( 
.A(n_176),
.Y(n_235)
);

INVx1_ASAP7_75t_L g307 ( 
.A(n_235),
.Y(n_307)
);

AND2x2_ASAP7_75t_SL g236 ( 
.A(n_200),
.B(n_76),
.Y(n_236)
);

CKINVDCx16_ASAP7_75t_R g320 ( 
.A(n_236),
.Y(n_320)
);

INVx8_ASAP7_75t_L g237 ( 
.A(n_132),
.Y(n_237)
);

BUFx2_ASAP7_75t_L g338 ( 
.A(n_237),
.Y(n_338)
);

AND2x2_ASAP7_75t_L g238 ( 
.A(n_215),
.B(n_106),
.Y(n_238)
);

NOR2xp33_ASAP7_75t_SL g339 ( 
.A(n_238),
.B(n_254),
.Y(n_339)
);

OAI22xp5_ASAP7_75t_SL g239 ( 
.A1(n_219),
.A2(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_239)
);

AOI22xp5_ASAP7_75t_L g313 ( 
.A1(n_239),
.A2(n_266),
.B1(n_171),
.B2(n_154),
.Y(n_313)
);

INVx1_ASAP7_75t_L g241 ( 
.A(n_130),
.Y(n_241)
);

INVx1_ASAP7_75t_L g328 ( 
.A(n_241),
.Y(n_328)
);

INVx1_ASAP7_75t_L g242 ( 
.A(n_184),
.Y(n_242)
);

INVx1_ASAP7_75t_L g353 ( 
.A(n_242),
.Y(n_353)
);

INVx6_ASAP7_75t_L g244 ( 
.A(n_177),
.Y(n_244)
);

BUFx6f_ASAP7_75t_L g337 ( 
.A(n_244),
.Y(n_337)
);

AOI22xp33_ASAP7_75t_SL g245 ( 
.A1(n_169),
.A2(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_245)
);

AOI22xp33_ASAP7_75t_SL g246 ( 
.A1(n_169),
.A2(n_55),
.B1(n_2),
.B2(n_3),
.Y(n_246)
);

INVx6_ASAP7_75t_L g247 ( 
.A(n_177),
.Y(n_247)
);

BUFx6f_ASAP7_75t_L g344 ( 
.A(n_247),
.Y(n_344)
);

BUFx3_ASAP7_75t_L g249 ( 
.A(n_142),
.Y(n_249)
);

BUFx3_ASAP7_75t_L g308 ( 
.A(n_249),
.Y(n_308)
);

OAI21xp33_ASAP7_75t_L g250 ( 
.A1(n_157),
.A2(n_13),
.B(n_4),
.Y(n_250)
);

AND2x2_ASAP7_75t_L g304 ( 
.A(n_250),
.B(n_272),
.Y(n_304)
);

INVx1_ASAP7_75t_L g251 ( 
.A(n_197),
.Y(n_251)
);

INVx1_ASAP7_75t_L g355 ( 
.A(n_251),
.Y(n_355)
);

INVx2_ASAP7_75t_L g252 ( 
.A(n_189),
.Y(n_252)
);

INVx2_ASAP7_75t_L g347 ( 
.A(n_252),
.Y(n_347)
);

INVx13_ASAP7_75t_L g253 ( 
.A(n_149),
.Y(n_253)
);

CKINVDCx16_ASAP7_75t_R g335 ( 
.A(n_253),
.Y(n_335)
);

AND2x2_ASAP7_75t_L g254 ( 
.A(n_140),
.B(n_152),
.Y(n_254)
);

INVx2_ASAP7_75t_L g255 ( 
.A(n_161),
.Y(n_255)
);

INVx2_ASAP7_75t_L g351 ( 
.A(n_255),
.Y(n_351)
);

INVx1_ASAP7_75t_L g256 ( 
.A(n_220),
.Y(n_256)
);

INVx2_ASAP7_75t_L g352 ( 
.A(n_256),
.Y(n_352)
);

BUFx6f_ASAP7_75t_L g258 ( 
.A(n_178),
.Y(n_258)
);

INVx5_ASAP7_75t_L g299 ( 
.A(n_258),
.Y(n_299)
);

INVx2_ASAP7_75t_L g260 ( 
.A(n_162),
.Y(n_260)
);

INVx4_ASAP7_75t_L g326 ( 
.A(n_260),
.Y(n_326)
);

BUFx12f_ASAP7_75t_L g261 ( 
.A(n_149),
.Y(n_261)
);

INVx5_ASAP7_75t_L g340 ( 
.A(n_261),
.Y(n_340)
);

INVx13_ASAP7_75t_L g263 ( 
.A(n_202),
.Y(n_263)
);

INVxp33_ASAP7_75t_L g309 ( 
.A(n_263),
.Y(n_309)
);

INVx3_ASAP7_75t_L g264 ( 
.A(n_138),
.Y(n_264)
);

INVx4_ASAP7_75t_L g333 ( 
.A(n_264),
.Y(n_333)
);

OAI22xp5_ASAP7_75t_SL g266 ( 
.A1(n_173),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_266)
);

CKINVDCx14_ASAP7_75t_R g267 ( 
.A(n_142),
.Y(n_267)
);

NAND2xp33_ASAP7_75t_SL g310 ( 
.A(n_267),
.B(n_294),
.Y(n_310)
);

CKINVDCx20_ASAP7_75t_R g268 ( 
.A(n_209),
.Y(n_268)
);

NAND2xp5_ASAP7_75t_SL g314 ( 
.A(n_268),
.B(n_282),
.Y(n_314)
);

INVx1_ASAP7_75t_L g269 ( 
.A(n_220),
.Y(n_269)
);

INVxp67_ASAP7_75t_L g354 ( 
.A(n_269),
.Y(n_354)
);

AOI22xp33_ASAP7_75t_L g270 ( 
.A1(n_158),
.A2(n_1),
.B1(n_4),
.B2(n_5),
.Y(n_270)
);

OAI22xp5_ASAP7_75t_L g330 ( 
.A1(n_270),
.A2(n_165),
.B1(n_137),
.B2(n_147),
.Y(n_330)
);

INVx3_ASAP7_75t_L g272 ( 
.A(n_138),
.Y(n_272)
);

BUFx6f_ASAP7_75t_L g273 ( 
.A(n_178),
.Y(n_273)
);

CKINVDCx20_ASAP7_75t_R g302 ( 
.A(n_273),
.Y(n_302)
);

INVx2_ASAP7_75t_L g274 ( 
.A(n_167),
.Y(n_274)
);

AND2x2_ASAP7_75t_L g318 ( 
.A(n_274),
.B(n_277),
.Y(n_318)
);

INVx1_ASAP7_75t_L g275 ( 
.A(n_168),
.Y(n_275)
);

NOR2xp33_ASAP7_75t_L g301 ( 
.A(n_275),
.B(n_276),
.Y(n_301)
);

INVx3_ASAP7_75t_L g277 ( 
.A(n_159),
.Y(n_277)
);

INVx3_ASAP7_75t_L g278 ( 
.A(n_145),
.Y(n_278)
);

AND2x2_ASAP7_75t_L g331 ( 
.A(n_278),
.B(n_284),
.Y(n_331)
);

INVx1_ASAP7_75t_L g280 ( 
.A(n_186),
.Y(n_280)
);

NOR2xp33_ASAP7_75t_L g319 ( 
.A(n_280),
.B(n_287),
.Y(n_319)
);

INVx6_ASAP7_75t_L g281 ( 
.A(n_182),
.Y(n_281)
);

CKINVDCx20_ASAP7_75t_R g336 ( 
.A(n_281),
.Y(n_336)
);

BUFx6f_ASAP7_75t_L g283 ( 
.A(n_182),
.Y(n_283)
);

CKINVDCx20_ASAP7_75t_R g343 ( 
.A(n_283),
.Y(n_343)
);

INVx2_ASAP7_75t_L g284 ( 
.A(n_143),
.Y(n_284)
);

INVx2_ASAP7_75t_L g285 ( 
.A(n_173),
.Y(n_285)
);

AND2x2_ASAP7_75t_L g349 ( 
.A(n_285),
.B(n_286),
.Y(n_349)
);

AND2x2_ASAP7_75t_L g286 ( 
.A(n_153),
.B(n_5),
.Y(n_286)
);

INVxp67_ASAP7_75t_L g287 ( 
.A(n_185),
.Y(n_287)
);

CKINVDCx16_ASAP7_75t_R g288 ( 
.A(n_129),
.Y(n_288)
);

NAND2xp5_ASAP7_75t_SL g342 ( 
.A(n_288),
.B(n_289),
.Y(n_342)
);

NAND2xp5_ASAP7_75t_L g289 ( 
.A(n_185),
.B(n_7),
.Y(n_289)
);

NAND2xp5_ASAP7_75t_L g290 ( 
.A(n_217),
.B(n_8),
.Y(n_290)
);

NOR2xp33_ASAP7_75t_SL g311 ( 
.A(n_290),
.B(n_8),
.Y(n_311)
);

INVx3_ASAP7_75t_L g291 ( 
.A(n_145),
.Y(n_291)
);

NOR2xp33_ASAP7_75t_L g345 ( 
.A(n_291),
.B(n_292),
.Y(n_345)
);

BUFx3_ASAP7_75t_L g292 ( 
.A(n_146),
.Y(n_292)
);

INVx8_ASAP7_75t_L g294 ( 
.A(n_132),
.Y(n_294)
);

INVx2_ASAP7_75t_SL g295 ( 
.A(n_129),
.Y(n_295)
);

NAND2xp5_ASAP7_75t_L g312 ( 
.A(n_295),
.B(n_296),
.Y(n_312)
);

INVx2_ASAP7_75t_L g296 ( 
.A(n_199),
.Y(n_296)
);

INVx4_ASAP7_75t_SL g297 ( 
.A(n_131),
.Y(n_297)
);

NAND2xp5_ASAP7_75t_L g315 ( 
.A(n_297),
.B(n_298),
.Y(n_315)
);

BUFx6f_ASAP7_75t_L g298 ( 
.A(n_188),
.Y(n_298)
);

OAI22xp33_ASAP7_75t_L g305 ( 
.A1(n_227),
.A2(n_134),
.B1(n_214),
.B2(n_204),
.Y(n_305)
);

OAI22xp5_ASAP7_75t_L g359 ( 
.A1(n_305),
.A2(n_306),
.B1(n_313),
.B2(n_325),
.Y(n_359)
);

AOI22xp33_ASAP7_75t_L g306 ( 
.A1(n_250),
.A2(n_160),
.B1(n_188),
.B2(n_217),
.Y(n_306)
);

NAND2xp5_ASAP7_75t_SL g385 ( 
.A(n_311),
.B(n_321),
.Y(n_385)
);

OAI22xp5_ASAP7_75t_SL g316 ( 
.A1(n_248),
.A2(n_199),
.B1(n_204),
.B2(n_154),
.Y(n_316)
);

AOI22xp5_ASAP7_75t_SL g376 ( 
.A1(n_316),
.A2(n_322),
.B1(n_298),
.B2(n_258),
.Y(n_376)
);

XNOR2xp5_ASAP7_75t_L g373 ( 
.A(n_317),
.B(n_232),
.Y(n_373)
);

NOR2xp33_ASAP7_75t_SL g321 ( 
.A(n_265),
.B(n_136),
.Y(n_321)
);

OAI22xp5_ASAP7_75t_SL g322 ( 
.A1(n_233),
.A2(n_135),
.B1(n_171),
.B2(n_155),
.Y(n_322)
);

NAND2xp5_ASAP7_75t_L g324 ( 
.A(n_224),
.B(n_155),
.Y(n_324)
);

NAND2xp5_ASAP7_75t_L g357 ( 
.A(n_324),
.B(n_350),
.Y(n_357)
);

AOI22xp5_ASAP7_75t_L g325 ( 
.A1(n_223),
.A2(n_135),
.B1(n_136),
.B2(n_210),
.Y(n_325)
);

NOR2xp33_ASAP7_75t_SL g327 ( 
.A(n_222),
.B(n_166),
.Y(n_327)
);

NAND2xp5_ASAP7_75t_SL g397 ( 
.A(n_327),
.B(n_202),
.Y(n_397)
);

AOI22xp5_ASAP7_75t_SL g329 ( 
.A1(n_238),
.A2(n_208),
.B1(n_194),
.B2(n_203),
.Y(n_329)
);

OAI21xp5_ASAP7_75t_SL g377 ( 
.A1(n_329),
.A2(n_246),
.B(n_245),
.Y(n_377)
);

OAI22xp5_ASAP7_75t_L g391 ( 
.A1(n_330),
.A2(n_341),
.B1(n_346),
.B2(n_348),
.Y(n_391)
);

OAI22xp5_ASAP7_75t_L g341 ( 
.A1(n_270),
.A2(n_151),
.B1(n_164),
.B2(n_210),
.Y(n_341)
);

OAI22xp5_ASAP7_75t_L g346 ( 
.A1(n_271),
.A2(n_164),
.B1(n_151),
.B2(n_139),
.Y(n_346)
);

OAI22xp5_ASAP7_75t_L g348 ( 
.A1(n_286),
.A2(n_139),
.B1(n_180),
.B2(n_147),
.Y(n_348)
);

NAND2xp5_ASAP7_75t_L g350 ( 
.A(n_236),
.B(n_196),
.Y(n_350)
);

AOI22xp5_ASAP7_75t_L g356 ( 
.A1(n_254),
.A2(n_180),
.B1(n_175),
.B2(n_137),
.Y(n_356)
);

NAND2xp5_ASAP7_75t_L g360 ( 
.A(n_356),
.B(n_267),
.Y(n_360)
);

INVx1_ASAP7_75t_L g358 ( 
.A(n_312),
.Y(n_358)
);

INVx1_ASAP7_75t_L g421 ( 
.A(n_358),
.Y(n_421)
);

AND2x2_ASAP7_75t_L g403 ( 
.A(n_360),
.B(n_376),
.Y(n_403)
);

BUFx3_ASAP7_75t_L g361 ( 
.A(n_340),
.Y(n_361)
);

INVx4_ASAP7_75t_L g411 ( 
.A(n_361),
.Y(n_411)
);

INVx1_ASAP7_75t_L g362 ( 
.A(n_312),
.Y(n_362)
);

INVx1_ASAP7_75t_L g435 ( 
.A(n_362),
.Y(n_435)
);

NOR2xp33_ASAP7_75t_L g363 ( 
.A(n_307),
.B(n_328),
.Y(n_363)
);

CKINVDCx14_ASAP7_75t_R g408 ( 
.A(n_363),
.Y(n_408)
);

CKINVDCx16_ASAP7_75t_R g364 ( 
.A(n_318),
.Y(n_364)
);

NOR2xp33_ASAP7_75t_L g410 ( 
.A(n_364),
.B(n_371),
.Y(n_410)
);

AND2x6_ASAP7_75t_L g365 ( 
.A(n_317),
.B(n_225),
.Y(n_365)
);

NOR2xp33_ASAP7_75t_L g429 ( 
.A(n_365),
.B(n_379),
.Y(n_429)
);

AOI22xp33_ASAP7_75t_SL g366 ( 
.A1(n_323),
.A2(n_262),
.B1(n_295),
.B2(n_279),
.Y(n_366)
);

AOI22xp33_ASAP7_75t_SL g405 ( 
.A1(n_366),
.A2(n_368),
.B1(n_370),
.B2(n_372),
.Y(n_405)
);

MAJIxp5_ASAP7_75t_L g367 ( 
.A(n_320),
.B(n_226),
.C(n_243),
.Y(n_367)
);

XNOR2xp5_ASAP7_75t_L g437 ( 
.A(n_367),
.B(n_373),
.Y(n_437)
);

AOI22xp33_ASAP7_75t_SL g368 ( 
.A1(n_323),
.A2(n_302),
.B1(n_343),
.B2(n_304),
.Y(n_368)
);

NAND2xp5_ASAP7_75t_L g369 ( 
.A(n_324),
.B(n_226),
.Y(n_369)
);

NAND2xp5_ASAP7_75t_L g407 ( 
.A(n_369),
.B(n_374),
.Y(n_407)
);

AOI22xp33_ASAP7_75t_SL g370 ( 
.A1(n_302),
.A2(n_292),
.B1(n_131),
.B2(n_297),
.Y(n_370)
);

INVxp33_ASAP7_75t_SL g371 ( 
.A(n_329),
.Y(n_371)
);

INVx13_ASAP7_75t_L g372 ( 
.A(n_335),
.Y(n_372)
);

NAND2xp5_ASAP7_75t_L g374 ( 
.A(n_301),
.B(n_230),
.Y(n_374)
);

NOR2xp33_ASAP7_75t_SL g375 ( 
.A(n_314),
.B(n_240),
.Y(n_375)
);

NOR2xp33_ASAP7_75t_SL g427 ( 
.A(n_375),
.B(n_386),
.Y(n_427)
);

INVxp67_ASAP7_75t_L g418 ( 
.A(n_377),
.Y(n_418)
);

XNOR2xp5_ASAP7_75t_L g378 ( 
.A(n_339),
.B(n_287),
.Y(n_378)
);

XOR2xp5_ASAP7_75t_L g412 ( 
.A(n_378),
.B(n_387),
.Y(n_412)
);

AND2x6_ASAP7_75t_L g379 ( 
.A(n_350),
.B(n_131),
.Y(n_379)
);

CKINVDCx20_ASAP7_75t_R g380 ( 
.A(n_332),
.Y(n_380)
);

NOR2xp33_ASAP7_75t_L g419 ( 
.A(n_380),
.B(n_388),
.Y(n_419)
);

INVx1_ASAP7_75t_L g381 ( 
.A(n_352),
.Y(n_381)
);

INVx1_ASAP7_75t_L g438 ( 
.A(n_381),
.Y(n_438)
);

INVx1_ASAP7_75t_L g382 ( 
.A(n_352),
.Y(n_382)
);

INVx2_ASAP7_75t_L g430 ( 
.A(n_382),
.Y(n_430)
);

BUFx6f_ASAP7_75t_L g383 ( 
.A(n_337),
.Y(n_383)
);

INVxp67_ASAP7_75t_L g426 ( 
.A(n_383),
.Y(n_426)
);

A2O1A1Ixp33_ASAP7_75t_L g384 ( 
.A1(n_304),
.A2(n_342),
.B(n_349),
.C(n_339),
.Y(n_384)
);

NAND2xp5_ASAP7_75t_SL g402 ( 
.A(n_384),
.B(n_389),
.Y(n_402)
);

MAJIxp5_ASAP7_75t_SL g386 ( 
.A(n_304),
.B(n_183),
.C(n_294),
.Y(n_386)
);

MAJIxp5_ASAP7_75t_L g387 ( 
.A(n_355),
.B(n_259),
.C(n_249),
.Y(n_387)
);

INVx1_ASAP7_75t_L g388 ( 
.A(n_353),
.Y(n_388)
);

NOR2xp33_ASAP7_75t_L g389 ( 
.A(n_307),
.B(n_328),
.Y(n_389)
);

INVx1_ASAP7_75t_SL g390 ( 
.A(n_310),
.Y(n_390)
);

NAND2xp5_ASAP7_75t_L g415 ( 
.A(n_390),
.B(n_396),
.Y(n_415)
);

INVx13_ASAP7_75t_L g392 ( 
.A(n_309),
.Y(n_392)
);

CKINVDCx20_ASAP7_75t_R g414 ( 
.A(n_392),
.Y(n_414)
);

MAJIxp5_ASAP7_75t_L g393 ( 
.A(n_355),
.B(n_259),
.C(n_257),
.Y(n_393)
);

XOR2xp5_ASAP7_75t_L g416 ( 
.A(n_393),
.B(n_310),
.Y(n_416)
);

INVx13_ASAP7_75t_L g394 ( 
.A(n_309),
.Y(n_394)
);

CKINVDCx20_ASAP7_75t_R g417 ( 
.A(n_394),
.Y(n_417)
);

AOI22xp33_ASAP7_75t_SL g395 ( 
.A1(n_343),
.A2(n_257),
.B1(n_132),
.B2(n_207),
.Y(n_395)
);

OAI21xp5_ASAP7_75t_L g428 ( 
.A1(n_395),
.A2(n_300),
.B(n_293),
.Y(n_428)
);

INVx2_ASAP7_75t_L g396 ( 
.A(n_337),
.Y(n_396)
);

NAND2xp5_ASAP7_75t_SL g406 ( 
.A(n_397),
.B(n_398),
.Y(n_406)
);

NOR2xp33_ASAP7_75t_L g398 ( 
.A(n_334),
.B(n_221),
.Y(n_398)
);

INVx1_ASAP7_75t_L g399 ( 
.A(n_353),
.Y(n_399)
);

NAND2xp5_ASAP7_75t_SL g425 ( 
.A(n_399),
.B(n_400),
.Y(n_425)
);

INVx1_ASAP7_75t_L g400 ( 
.A(n_318),
.Y(n_400)
);

INVx3_ASAP7_75t_L g401 ( 
.A(n_299),
.Y(n_401)
);

NAND2xp5_ASAP7_75t_L g420 ( 
.A(n_401),
.B(n_336),
.Y(n_420)
);

OAI22xp5_ASAP7_75t_SL g404 ( 
.A1(n_358),
.A2(n_313),
.B1(n_303),
.B2(n_325),
.Y(n_404)
);

AOI22xp5_ASAP7_75t_L g441 ( 
.A1(n_404),
.A2(n_409),
.B1(n_413),
.B2(n_422),
.Y(n_441)
);

OAI22xp5_ASAP7_75t_L g409 ( 
.A1(n_362),
.A2(n_305),
.B1(n_349),
.B2(n_315),
.Y(n_409)
);

OAI22xp5_ASAP7_75t_SL g413 ( 
.A1(n_376),
.A2(n_349),
.B1(n_336),
.B2(n_316),
.Y(n_413)
);

MAJIxp5_ASAP7_75t_L g457 ( 
.A(n_416),
.B(n_331),
.C(n_333),
.Y(n_457)
);

INVx1_ASAP7_75t_L g442 ( 
.A(n_420),
.Y(n_442)
);

OAI22xp5_ASAP7_75t_SL g422 ( 
.A1(n_357),
.A2(n_315),
.B1(n_322),
.B2(n_356),
.Y(n_422)
);

CKINVDCx20_ASAP7_75t_R g423 ( 
.A(n_374),
.Y(n_423)
);

NOR2xp33_ASAP7_75t_L g455 ( 
.A(n_423),
.B(n_381),
.Y(n_455)
);

AOI22xp5_ASAP7_75t_L g424 ( 
.A1(n_359),
.A2(n_345),
.B1(n_344),
.B2(n_299),
.Y(n_424)
);

OAI22xp5_ASAP7_75t_SL g461 ( 
.A1(n_424),
.A2(n_436),
.B1(n_383),
.B2(n_361),
.Y(n_461)
);

OAI21xp5_ASAP7_75t_SL g440 ( 
.A1(n_428),
.A2(n_433),
.B(n_400),
.Y(n_440)
);

OAI22xp5_ASAP7_75t_SL g431 ( 
.A1(n_357),
.A2(n_244),
.B1(n_281),
.B2(n_247),
.Y(n_431)
);

AOI22xp5_ASAP7_75t_L g470 ( 
.A1(n_431),
.A2(n_354),
.B1(n_347),
.B2(n_326),
.Y(n_470)
);

NAND2xp5_ASAP7_75t_L g432 ( 
.A(n_369),
.B(n_319),
.Y(n_432)
);

NAND2xp5_ASAP7_75t_L g443 ( 
.A(n_432),
.B(n_434),
.Y(n_443)
);

AOI21xp5_ASAP7_75t_L g433 ( 
.A1(n_390),
.A2(n_377),
.B(n_373),
.Y(n_433)
);

OA21x2_ASAP7_75t_L g434 ( 
.A1(n_360),
.A2(n_331),
.B(n_318),
.Y(n_434)
);

AOI22xp5_ASAP7_75t_L g436 ( 
.A1(n_391),
.A2(n_344),
.B1(n_331),
.B2(n_333),
.Y(n_436)
);

OAI21xp5_ASAP7_75t_L g439 ( 
.A1(n_433),
.A2(n_384),
.B(n_378),
.Y(n_439)
);

OAI21xp5_ASAP7_75t_SL g489 ( 
.A1(n_439),
.A2(n_440),
.B(n_447),
.Y(n_489)
);

OR2x2_ASAP7_75t_L g444 ( 
.A(n_402),
.B(n_386),
.Y(n_444)
);

CKINVDCx20_ASAP7_75t_R g486 ( 
.A(n_444),
.Y(n_486)
);

NAND3xp33_ASAP7_75t_L g445 ( 
.A(n_402),
.B(n_367),
.C(n_375),
.Y(n_445)
);

NOR2xp33_ASAP7_75t_L g475 ( 
.A(n_445),
.B(n_466),
.Y(n_475)
);

CKINVDCx10_ASAP7_75t_R g446 ( 
.A(n_405),
.Y(n_446)
);

CKINVDCx20_ASAP7_75t_R g497 ( 
.A(n_446),
.Y(n_497)
);

AOI22xp5_ASAP7_75t_SL g447 ( 
.A1(n_418),
.A2(n_379),
.B1(n_380),
.B2(n_385),
.Y(n_447)
);

CKINVDCx20_ASAP7_75t_R g448 ( 
.A(n_408),
.Y(n_448)
);

NAND2xp5_ASAP7_75t_L g476 ( 
.A(n_448),
.B(n_454),
.Y(n_476)
);

NAND2xp5_ASAP7_75t_L g449 ( 
.A(n_423),
.B(n_388),
.Y(n_449)
);

INVx1_ASAP7_75t_L g482 ( 
.A(n_449),
.Y(n_482)
);

NOR2xp33_ASAP7_75t_SL g450 ( 
.A(n_406),
.B(n_387),
.Y(n_450)
);

NOR2xp33_ASAP7_75t_SL g490 ( 
.A(n_450),
.B(n_451),
.Y(n_490)
);

NAND2xp5_ASAP7_75t_SL g451 ( 
.A(n_421),
.B(n_399),
.Y(n_451)
);

NAND2xp5_ASAP7_75t_L g452 ( 
.A(n_425),
.B(n_382),
.Y(n_452)
);

INVx1_ASAP7_75t_L g484 ( 
.A(n_452),
.Y(n_484)
);

CKINVDCx16_ASAP7_75t_R g453 ( 
.A(n_419),
.Y(n_453)
);

INVx1_ASAP7_75t_L g488 ( 
.A(n_453),
.Y(n_488)
);

CKINVDCx20_ASAP7_75t_R g454 ( 
.A(n_419),
.Y(n_454)
);

INVx1_ASAP7_75t_L g492 ( 
.A(n_455),
.Y(n_492)
);

NOR2xp33_ASAP7_75t_L g456 ( 
.A(n_414),
.B(n_393),
.Y(n_456)
);

NAND2xp5_ASAP7_75t_SL g499 ( 
.A(n_456),
.B(n_458),
.Y(n_499)
);

MAJIxp5_ASAP7_75t_L g477 ( 
.A(n_457),
.B(n_412),
.C(n_416),
.Y(n_477)
);

NOR2xp33_ASAP7_75t_L g458 ( 
.A(n_414),
.B(n_401),
.Y(n_458)
);

INVx1_ASAP7_75t_L g459 ( 
.A(n_438),
.Y(n_459)
);

INVx1_ASAP7_75t_L g503 ( 
.A(n_459),
.Y(n_503)
);

NAND2xp5_ASAP7_75t_L g460 ( 
.A(n_425),
.B(n_396),
.Y(n_460)
);

NAND2xp5_ASAP7_75t_L g498 ( 
.A(n_460),
.B(n_464),
.Y(n_498)
);

AOI22xp5_ASAP7_75t_SL g494 ( 
.A1(n_461),
.A2(n_471),
.B1(n_446),
.B2(n_409),
.Y(n_494)
);

OAI22xp5_ASAP7_75t_SL g462 ( 
.A1(n_421),
.A2(n_365),
.B1(n_273),
.B2(n_283),
.Y(n_462)
);

AOI22xp5_ASAP7_75t_L g485 ( 
.A1(n_462),
.A2(n_463),
.B1(n_470),
.B2(n_413),
.Y(n_485)
);

OAI22xp5_ASAP7_75t_SL g463 ( 
.A1(n_435),
.A2(n_338),
.B1(n_326),
.B2(n_351),
.Y(n_463)
);

CKINVDCx14_ASAP7_75t_R g464 ( 
.A(n_406),
.Y(n_464)
);

CKINVDCx20_ASAP7_75t_R g465 ( 
.A(n_420),
.Y(n_465)
);

CKINVDCx20_ASAP7_75t_R g500 ( 
.A(n_465),
.Y(n_500)
);

NAND2xp5_ASAP7_75t_L g466 ( 
.A(n_435),
.B(n_347),
.Y(n_466)
);

NOR2xp33_ASAP7_75t_L g467 ( 
.A(n_417),
.B(n_351),
.Y(n_467)
);

NOR2xp33_ASAP7_75t_L g480 ( 
.A(n_467),
.B(n_468),
.Y(n_480)
);

INVx1_ASAP7_75t_L g468 ( 
.A(n_438),
.Y(n_468)
);

CKINVDCx20_ASAP7_75t_R g469 ( 
.A(n_434),
.Y(n_469)
);

NOR2xp33_ASAP7_75t_L g493 ( 
.A(n_469),
.B(n_472),
.Y(n_493)
);

AOI22xp5_ASAP7_75t_SL g471 ( 
.A1(n_403),
.A2(n_338),
.B1(n_372),
.B2(n_340),
.Y(n_471)
);

AOI32xp33_ASAP7_75t_L g472 ( 
.A1(n_429),
.A2(n_392),
.A3(n_394),
.B1(n_293),
.B2(n_354),
.Y(n_472)
);

AOI21xp5_ASAP7_75t_L g473 ( 
.A1(n_440),
.A2(n_410),
.B(n_403),
.Y(n_473)
);

OAI21xp5_ASAP7_75t_SL g515 ( 
.A1(n_473),
.A2(n_478),
.B(n_494),
.Y(n_515)
);

XNOR2xp5_ASAP7_75t_SL g474 ( 
.A(n_439),
.B(n_437),
.Y(n_474)
);

XNOR2xp5_ASAP7_75t_SL g516 ( 
.A(n_474),
.B(n_441),
.Y(n_516)
);

MAJIxp5_ASAP7_75t_L g505 ( 
.A(n_477),
.B(n_479),
.C(n_496),
.Y(n_505)
);

AOI21xp5_ASAP7_75t_L g478 ( 
.A1(n_469),
.A2(n_410),
.B(n_403),
.Y(n_478)
);

MAJIxp5_ASAP7_75t_L g479 ( 
.A(n_457),
.B(n_437),
.C(n_412),
.Y(n_479)
);

XNOR2xp5_ASAP7_75t_L g481 ( 
.A(n_457),
.B(n_432),
.Y(n_481)
);

XNOR2xp5_ASAP7_75t_L g506 ( 
.A(n_481),
.B(n_483),
.Y(n_506)
);

XNOR2xp5_ASAP7_75t_L g483 ( 
.A(n_443),
.B(n_407),
.Y(n_483)
);

OAI22xp5_ASAP7_75t_L g522 ( 
.A1(n_485),
.A2(n_460),
.B1(n_434),
.B2(n_470),
.Y(n_522)
);

BUFx24_ASAP7_75t_SL g487 ( 
.A(n_448),
.Y(n_487)
);

NOR2xp33_ASAP7_75t_SL g510 ( 
.A(n_487),
.B(n_495),
.Y(n_510)
);

FAx1_ASAP7_75t_SL g491 ( 
.A(n_444),
.B(n_407),
.CI(n_427),
.CON(n_491),
.SN(n_491)
);

OAI31xp33_ASAP7_75t_SL g509 ( 
.A1(n_491),
.A2(n_445),
.A3(n_444),
.B(n_449),
.Y(n_509)
);

NOR2xp33_ASAP7_75t_L g495 ( 
.A(n_450),
.B(n_464),
.Y(n_495)
);

XOR2xp5_ASAP7_75t_L g496 ( 
.A(n_443),
.B(n_427),
.Y(n_496)
);

OAI22xp5_ASAP7_75t_SL g501 ( 
.A1(n_441),
.A2(n_424),
.B1(n_436),
.B2(n_415),
.Y(n_501)
);

AOI22xp5_ASAP7_75t_L g525 ( 
.A1(n_501),
.A2(n_404),
.B1(n_461),
.B2(n_422),
.Y(n_525)
);

NOR2xp33_ASAP7_75t_L g502 ( 
.A(n_454),
.B(n_411),
.Y(n_502)
);

NAND2xp5_ASAP7_75t_L g526 ( 
.A(n_502),
.B(n_458),
.Y(n_526)
);

NAND2xp5_ASAP7_75t_L g504 ( 
.A(n_476),
.B(n_451),
.Y(n_504)
);

INVx1_ASAP7_75t_L g532 ( 
.A(n_504),
.Y(n_532)
);

INVx1_ASAP7_75t_L g507 ( 
.A(n_476),
.Y(n_507)
);

INVx1_ASAP7_75t_L g541 ( 
.A(n_507),
.Y(n_541)
);

INVx1_ASAP7_75t_L g508 ( 
.A(n_492),
.Y(n_508)
);

NAND2xp5_ASAP7_75t_L g534 ( 
.A(n_508),
.B(n_514),
.Y(n_534)
);

XNOR2xp5_ASAP7_75t_L g533 ( 
.A(n_509),
.B(n_517),
.Y(n_533)
);

MAJIxp5_ASAP7_75t_L g511 ( 
.A(n_479),
.B(n_456),
.C(n_442),
.Y(n_511)
);

MAJIxp5_ASAP7_75t_L g538 ( 
.A(n_511),
.B(n_512),
.C(n_513),
.Y(n_538)
);

MAJIxp5_ASAP7_75t_L g512 ( 
.A(n_477),
.B(n_442),
.C(n_447),
.Y(n_512)
);

MAJIxp5_ASAP7_75t_L g513 ( 
.A(n_474),
.B(n_453),
.C(n_452),
.Y(n_513)
);

NOR2xp33_ASAP7_75t_L g514 ( 
.A(n_490),
.B(n_475),
.Y(n_514)
);

XNOR2xp5_ASAP7_75t_SL g536 ( 
.A(n_516),
.B(n_489),
.Y(n_536)
);

XNOR2xp5_ASAP7_75t_L g517 ( 
.A(n_481),
.B(n_455),
.Y(n_517)
);

INVx1_ASAP7_75t_L g518 ( 
.A(n_492),
.Y(n_518)
);

HB1xp67_ASAP7_75t_L g542 ( 
.A(n_518),
.Y(n_542)
);

INVx1_ASAP7_75t_L g519 ( 
.A(n_498),
.Y(n_519)
);

INVxp33_ASAP7_75t_L g545 ( 
.A(n_519),
.Y(n_545)
);

NAND2xp5_ASAP7_75t_SL g520 ( 
.A(n_490),
.B(n_462),
.Y(n_520)
);

OAI22xp5_ASAP7_75t_L g539 ( 
.A1(n_520),
.A2(n_522),
.B1(n_523),
.B2(n_525),
.Y(n_539)
);

OAI21xp5_ASAP7_75t_SL g521 ( 
.A1(n_493),
.A2(n_465),
.B(n_471),
.Y(n_521)
);

OAI21xp5_ASAP7_75t_L g531 ( 
.A1(n_521),
.A2(n_473),
.B(n_478),
.Y(n_531)
);

NOR2xp33_ASAP7_75t_L g523 ( 
.A(n_496),
.B(n_411),
.Y(n_523)
);

MAJIxp5_ASAP7_75t_L g524 ( 
.A(n_499),
.B(n_415),
.C(n_468),
.Y(n_524)
);

MAJIxp5_ASAP7_75t_L g540 ( 
.A(n_524),
.B(n_488),
.C(n_482),
.Y(n_540)
);

OAI22xp5_ASAP7_75t_SL g537 ( 
.A1(n_526),
.A2(n_528),
.B1(n_529),
.B2(n_530),
.Y(n_537)
);

XNOR2xp5_ASAP7_75t_L g527 ( 
.A(n_499),
.B(n_466),
.Y(n_527)
);

XNOR2xp5_ASAP7_75t_L g544 ( 
.A(n_527),
.B(n_498),
.Y(n_544)
);

AOI22xp5_ASAP7_75t_L g528 ( 
.A1(n_500),
.A2(n_434),
.B1(n_431),
.B2(n_459),
.Y(n_528)
);

AOI22xp5_ASAP7_75t_L g529 ( 
.A1(n_500),
.A2(n_472),
.B1(n_467),
.B2(n_463),
.Y(n_529)
);

NOR2xp33_ASAP7_75t_L g530 ( 
.A(n_483),
.B(n_417),
.Y(n_530)
);

OAI21xp5_ASAP7_75t_SL g556 ( 
.A1(n_531),
.A2(n_550),
.B(n_491),
.Y(n_556)
);

XOR2xp5_ASAP7_75t_L g535 ( 
.A(n_505),
.B(n_511),
.Y(n_535)
);

XOR2xp5_ASAP7_75t_L g565 ( 
.A(n_535),
.B(n_536),
.Y(n_565)
);

NAND2xp5_ASAP7_75t_SL g558 ( 
.A(n_540),
.B(n_546),
.Y(n_558)
);

XNOR2x1_ASAP7_75t_L g543 ( 
.A(n_516),
.B(n_494),
.Y(n_543)
);

XNOR2xp5_ASAP7_75t_L g562 ( 
.A(n_543),
.B(n_501),
.Y(n_562)
);

NAND2xp5_ASAP7_75t_L g554 ( 
.A(n_544),
.B(n_524),
.Y(n_554)
);

MAJIxp5_ASAP7_75t_L g546 ( 
.A(n_505),
.B(n_512),
.C(n_506),
.Y(n_546)
);

MAJIxp5_ASAP7_75t_L g547 ( 
.A(n_506),
.B(n_489),
.C(n_488),
.Y(n_547)
);

NAND2xp5_ASAP7_75t_SL g560 ( 
.A(n_547),
.B(n_527),
.Y(n_560)
);

OAI22xp5_ASAP7_75t_SL g548 ( 
.A1(n_525),
.A2(n_482),
.B1(n_484),
.B2(n_486),
.Y(n_548)
);

AOI22xp5_ASAP7_75t_L g563 ( 
.A1(n_548),
.A2(n_549),
.B1(n_503),
.B2(n_497),
.Y(n_563)
);

OAI22xp5_ASAP7_75t_SL g549 ( 
.A1(n_529),
.A2(n_484),
.B1(n_486),
.B2(n_485),
.Y(n_549)
);

OAI21xp5_ASAP7_75t_L g550 ( 
.A1(n_515),
.A2(n_491),
.B(n_480),
.Y(n_550)
);

MAJIxp5_ASAP7_75t_L g551 ( 
.A(n_535),
.B(n_513),
.C(n_515),
.Y(n_551)
);

NAND2xp5_ASAP7_75t_L g569 ( 
.A(n_551),
.B(n_553),
.Y(n_569)
);

OAI22xp5_ASAP7_75t_SL g552 ( 
.A1(n_532),
.A2(n_528),
.B1(n_504),
.B2(n_509),
.Y(n_552)
);

AOI22xp5_ASAP7_75t_L g579 ( 
.A1(n_552),
.A2(n_559),
.B1(n_566),
.B2(n_548),
.Y(n_579)
);

MAJIxp5_ASAP7_75t_L g553 ( 
.A(n_546),
.B(n_517),
.C(n_521),
.Y(n_553)
);

INVxp67_ASAP7_75t_L g572 ( 
.A(n_554),
.Y(n_572)
);

INVx1_ASAP7_75t_L g555 ( 
.A(n_534),
.Y(n_555)
);

INVx1_ASAP7_75t_L g574 ( 
.A(n_555),
.Y(n_574)
);

OAI21xp5_ASAP7_75t_L g575 ( 
.A1(n_556),
.A2(n_533),
.B(n_545),
.Y(n_575)
);

INVx1_ASAP7_75t_L g557 ( 
.A(n_542),
.Y(n_557)
);

INVx1_ASAP7_75t_L g578 ( 
.A(n_557),
.Y(n_578)
);

INVx1_ASAP7_75t_L g559 ( 
.A(n_544),
.Y(n_559)
);

XNOR2xp5_ASAP7_75t_L g576 ( 
.A(n_560),
.B(n_562),
.Y(n_576)
);

CKINVDCx20_ASAP7_75t_R g561 ( 
.A(n_550),
.Y(n_561)
);

NOR2xp33_ASAP7_75t_SL g577 ( 
.A(n_561),
.B(n_556),
.Y(n_577)
);

OAI22xp5_ASAP7_75t_SL g570 ( 
.A1(n_563),
.A2(n_545),
.B1(n_541),
.B2(n_531),
.Y(n_570)
);

MAJIxp5_ASAP7_75t_L g564 ( 
.A(n_538),
.B(n_503),
.C(n_497),
.Y(n_564)
);

MAJIxp5_ASAP7_75t_L g571 ( 
.A(n_564),
.B(n_567),
.C(n_558),
.Y(n_571)
);

INVx1_ASAP7_75t_L g566 ( 
.A(n_540),
.Y(n_566)
);

MAJIxp5_ASAP7_75t_L g567 ( 
.A(n_538),
.B(n_430),
.C(n_426),
.Y(n_567)
);

AOI22xp5_ASAP7_75t_L g568 ( 
.A1(n_552),
.A2(n_549),
.B1(n_537),
.B2(n_539),
.Y(n_568)
);

OAI22xp5_ASAP7_75t_L g588 ( 
.A1(n_568),
.A2(n_577),
.B1(n_564),
.B2(n_576),
.Y(n_588)
);

INVx1_ASAP7_75t_L g590 ( 
.A(n_570),
.Y(n_590)
);

XNOR2xp5_ASAP7_75t_L g582 ( 
.A(n_571),
.B(n_575),
.Y(n_582)
);

MAJIxp5_ASAP7_75t_L g573 ( 
.A(n_567),
.B(n_547),
.C(n_533),
.Y(n_573)
);

NAND2xp5_ASAP7_75t_SL g587 ( 
.A(n_573),
.B(n_580),
.Y(n_587)
);

INVx1_ASAP7_75t_L g591 ( 
.A(n_579),
.Y(n_591)
);

MAJIxp5_ASAP7_75t_L g580 ( 
.A(n_551),
.B(n_543),
.C(n_536),
.Y(n_580)
);

MAJIxp5_ASAP7_75t_L g581 ( 
.A(n_553),
.B(n_430),
.C(n_428),
.Y(n_581)
);

MAJIxp5_ASAP7_75t_L g592 ( 
.A(n_581),
.B(n_565),
.C(n_562),
.Y(n_592)
);

CKINVDCx20_ASAP7_75t_R g583 ( 
.A(n_575),
.Y(n_583)
);

NOR2xp33_ASAP7_75t_L g595 ( 
.A(n_583),
.B(n_589),
.Y(n_595)
);

OAI22xp33_ASAP7_75t_SL g584 ( 
.A1(n_574),
.A2(n_563),
.B1(n_557),
.B2(n_559),
.Y(n_584)
);

INVx1_ASAP7_75t_L g597 ( 
.A(n_584),
.Y(n_597)
);

NOR2xp33_ASAP7_75t_L g585 ( 
.A(n_571),
.B(n_510),
.Y(n_585)
);

NOR2xp33_ASAP7_75t_L g600 ( 
.A(n_585),
.B(n_588),
.Y(n_600)
);

XOR2xp5_ASAP7_75t_L g586 ( 
.A(n_576),
.B(n_554),
.Y(n_586)
);

MAJIxp5_ASAP7_75t_L g593 ( 
.A(n_586),
.B(n_592),
.C(n_587),
.Y(n_593)
);

NOR2xp33_ASAP7_75t_SL g589 ( 
.A(n_569),
.B(n_565),
.Y(n_589)
);

NAND2xp5_ASAP7_75t_L g605 ( 
.A(n_593),
.B(n_594),
.Y(n_605)
);

MAJIxp5_ASAP7_75t_L g594 ( 
.A(n_582),
.B(n_572),
.C(n_573),
.Y(n_594)
);

AOI21x1_ASAP7_75t_SL g596 ( 
.A1(n_590),
.A2(n_572),
.B(n_568),
.Y(n_596)
);

OAI21xp5_ASAP7_75t_L g604 ( 
.A1(n_596),
.A2(n_591),
.B(n_237),
.Y(n_604)
);

MAJIxp5_ASAP7_75t_L g598 ( 
.A(n_582),
.B(n_578),
.C(n_580),
.Y(n_598)
);

NOR2xp33_ASAP7_75t_SL g603 ( 
.A(n_598),
.B(n_592),
.Y(n_603)
);

OAI21xp5_ASAP7_75t_SL g599 ( 
.A1(n_590),
.A2(n_581),
.B(n_263),
.Y(n_599)
);

OAI21xp5_ASAP7_75t_SL g602 ( 
.A1(n_599),
.A2(n_591),
.B(n_253),
.Y(n_602)
);

MAJIxp5_ASAP7_75t_L g601 ( 
.A(n_600),
.B(n_595),
.C(n_586),
.Y(n_601)
);

NOR2xp33_ASAP7_75t_SL g607 ( 
.A(n_601),
.B(n_602),
.Y(n_607)
);

NOR2x1_ASAP7_75t_L g608 ( 
.A(n_603),
.B(n_604),
.Y(n_608)
);

OAI21xp5_ASAP7_75t_SL g606 ( 
.A1(n_605),
.A2(n_600),
.B(n_597),
.Y(n_606)
);

NOR2xp33_ASAP7_75t_L g609 ( 
.A(n_606),
.B(n_308),
.Y(n_609)
);

INVx1_ASAP7_75t_L g611 ( 
.A(n_609),
.Y(n_611)
);

NOR2xp33_ASAP7_75t_L g610 ( 
.A(n_607),
.B(n_308),
.Y(n_610)
);

AOI322xp5_ASAP7_75t_L g612 ( 
.A1(n_611),
.A2(n_610),
.A3(n_608),
.B1(n_261),
.B2(n_11),
.C1(n_10),
.C2(n_9),
.Y(n_612)
);

NAND2xp5_ASAP7_75t_L g613 ( 
.A(n_612),
.B(n_8),
.Y(n_613)
);

BUFx24_ASAP7_75t_SL g614 ( 
.A(n_613),
.Y(n_614)
);

NAND2xp5_ASAP7_75t_L g615 ( 
.A(n_614),
.B(n_261),
.Y(n_615)
);


endmodule